module basic_3000_30000_3500_15_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2836,In_1688);
nor U1 (N_1,In_1994,In_2884);
xor U2 (N_2,In_1320,In_2384);
xnor U3 (N_3,In_2854,In_918);
nand U4 (N_4,In_1500,In_1765);
or U5 (N_5,In_2831,In_1394);
xnor U6 (N_6,In_1223,In_1849);
nand U7 (N_7,In_498,In_1083);
nand U8 (N_8,In_1966,In_166);
and U9 (N_9,In_1786,In_1101);
nor U10 (N_10,In_2839,In_1766);
or U11 (N_11,In_336,In_1593);
nor U12 (N_12,In_816,In_1597);
nor U13 (N_13,In_433,In_947);
or U14 (N_14,In_2353,In_2638);
and U15 (N_15,In_223,In_2050);
or U16 (N_16,In_2263,In_2182);
or U17 (N_17,In_1465,In_2357);
nor U18 (N_18,In_1276,In_868);
or U19 (N_19,In_293,In_751);
nand U20 (N_20,In_296,In_1353);
nand U21 (N_21,In_1438,In_1654);
nand U22 (N_22,In_1960,In_829);
xor U23 (N_23,In_1344,In_1508);
xnor U24 (N_24,In_567,In_1722);
and U25 (N_25,In_922,In_365);
or U26 (N_26,In_131,In_1801);
nor U27 (N_27,In_1651,In_2790);
or U28 (N_28,In_2968,In_1697);
or U29 (N_29,In_2589,In_2150);
nor U30 (N_30,In_2605,In_1436);
and U31 (N_31,In_2480,In_1947);
xnor U32 (N_32,In_1481,In_2147);
xnor U33 (N_33,In_1279,In_1264);
nand U34 (N_34,In_1477,In_2786);
nand U35 (N_35,In_51,In_1628);
or U36 (N_36,In_1044,In_1602);
nor U37 (N_37,In_688,In_2917);
or U38 (N_38,In_1708,In_833);
and U39 (N_39,In_2334,In_198);
and U40 (N_40,In_1024,In_360);
xor U41 (N_41,In_1975,In_169);
and U42 (N_42,In_771,In_427);
and U43 (N_43,In_2751,In_853);
xor U44 (N_44,In_204,In_732);
xor U45 (N_45,In_1090,In_1814);
and U46 (N_46,In_2979,In_1634);
nand U47 (N_47,In_2984,In_136);
nor U48 (N_48,In_620,In_1625);
xnor U49 (N_49,In_202,In_1990);
or U50 (N_50,In_2468,In_2097);
nand U51 (N_51,In_1555,In_420);
nand U52 (N_52,In_2170,In_2032);
xnor U53 (N_53,In_236,In_395);
nand U54 (N_54,In_1586,In_141);
nor U55 (N_55,In_2485,In_2642);
and U56 (N_56,In_389,In_1749);
nand U57 (N_57,In_605,In_2525);
nor U58 (N_58,In_2828,In_1168);
nor U59 (N_59,In_888,In_1452);
nor U60 (N_60,In_1346,In_504);
and U61 (N_61,In_2875,In_1203);
nand U62 (N_62,In_2542,In_1497);
and U63 (N_63,In_2207,In_2973);
and U64 (N_64,In_487,In_683);
nand U65 (N_65,In_2154,In_938);
xor U66 (N_66,In_1466,In_1871);
or U67 (N_67,In_2346,In_304);
nor U68 (N_68,In_272,In_1630);
and U69 (N_69,In_68,In_1948);
nand U70 (N_70,In_1608,In_2634);
xnor U71 (N_71,In_2023,In_2081);
or U72 (N_72,In_2721,In_2418);
nand U73 (N_73,In_2570,In_475);
and U74 (N_74,In_737,In_1140);
nand U75 (N_75,In_762,In_989);
or U76 (N_76,In_254,In_875);
and U77 (N_77,In_539,In_640);
or U78 (N_78,In_1425,In_1207);
nor U79 (N_79,In_2530,In_676);
xnor U80 (N_80,In_2964,In_1810);
nor U81 (N_81,In_2131,In_285);
nand U82 (N_82,In_2407,In_787);
nand U83 (N_83,In_2408,In_1231);
nor U84 (N_84,In_1850,In_1301);
nor U85 (N_85,In_220,In_2319);
nor U86 (N_86,In_2993,In_2393);
and U87 (N_87,In_1443,In_581);
or U88 (N_88,In_1284,In_2083);
and U89 (N_89,In_2300,In_1288);
and U90 (N_90,In_986,In_744);
and U91 (N_91,In_2791,In_748);
nor U92 (N_92,In_1569,In_2004);
xnor U93 (N_93,In_1208,In_1351);
and U94 (N_94,In_2261,In_2227);
nor U95 (N_95,In_1306,In_378);
nand U96 (N_96,In_1173,In_2178);
nor U97 (N_97,In_2168,In_1897);
nor U98 (N_98,In_177,In_760);
nor U99 (N_99,In_982,In_2116);
and U100 (N_100,In_521,In_1028);
nand U101 (N_101,In_1777,In_2996);
and U102 (N_102,In_1085,In_459);
xor U103 (N_103,In_380,In_207);
and U104 (N_104,In_2354,In_1403);
and U105 (N_105,In_428,In_1050);
xor U106 (N_106,In_1987,In_412);
or U107 (N_107,In_2515,In_2539);
or U108 (N_108,In_1717,In_759);
xor U109 (N_109,In_677,In_526);
xor U110 (N_110,In_1266,In_2636);
nand U111 (N_111,In_595,In_438);
or U112 (N_112,In_2342,In_308);
and U113 (N_113,In_2748,In_1951);
and U114 (N_114,In_2484,In_2286);
xnor U115 (N_115,In_2419,In_2936);
and U116 (N_116,In_2882,In_2630);
and U117 (N_117,In_2703,In_1632);
nor U118 (N_118,In_2406,In_1084);
nand U119 (N_119,In_933,In_1241);
nand U120 (N_120,In_2585,In_1635);
xor U121 (N_121,In_2362,In_507);
nand U122 (N_122,In_256,In_1535);
nor U123 (N_123,In_2104,In_1304);
nor U124 (N_124,In_1931,In_2678);
and U125 (N_125,In_15,In_739);
and U126 (N_126,In_1996,In_715);
nand U127 (N_127,In_667,In_297);
xor U128 (N_128,In_2404,In_2205);
and U129 (N_129,In_2315,In_276);
xnor U130 (N_130,In_2604,In_1369);
xor U131 (N_131,In_2329,In_435);
and U132 (N_132,In_92,In_1354);
xnor U133 (N_133,In_446,In_550);
nand U134 (N_134,In_1549,In_1311);
and U135 (N_135,In_2091,In_1411);
nand U136 (N_136,In_956,In_181);
nand U137 (N_137,In_520,In_154);
xnor U138 (N_138,In_1903,In_2185);
xnor U139 (N_139,In_1778,In_1845);
nor U140 (N_140,In_634,In_2820);
or U141 (N_141,In_1169,In_554);
xnor U142 (N_142,In_416,In_2251);
or U143 (N_143,In_1864,In_578);
nor U144 (N_144,In_1904,In_1912);
nor U145 (N_145,In_437,In_2567);
or U146 (N_146,In_1326,In_990);
xor U147 (N_147,In_2618,In_883);
xor U148 (N_148,In_1859,In_2487);
nor U149 (N_149,In_1531,In_2632);
and U150 (N_150,In_1695,In_1468);
nand U151 (N_151,In_16,In_1771);
nor U152 (N_152,In_294,In_37);
nand U153 (N_153,In_167,In_472);
nor U154 (N_154,In_134,In_2305);
nand U155 (N_155,In_2193,In_1398);
nor U156 (N_156,In_2297,In_2211);
nand U157 (N_157,In_1141,In_1890);
nand U158 (N_158,In_1045,In_94);
nand U159 (N_159,In_2559,In_2568);
and U160 (N_160,In_2864,In_1123);
nor U161 (N_161,In_2947,In_2220);
and U162 (N_162,In_801,In_224);
nor U163 (N_163,In_2612,In_175);
nand U164 (N_164,In_1748,In_1236);
or U165 (N_165,In_925,In_2490);
and U166 (N_166,In_1730,In_1544);
or U167 (N_167,In_383,In_1488);
xnor U168 (N_168,In_1509,In_1170);
or U169 (N_169,In_2201,In_2990);
nand U170 (N_170,In_841,In_2218);
nor U171 (N_171,In_840,In_2714);
and U172 (N_172,In_586,In_785);
nand U173 (N_173,In_1056,In_2675);
or U174 (N_174,In_115,In_2078);
xor U175 (N_175,In_1661,In_2537);
nor U176 (N_176,In_235,In_2119);
and U177 (N_177,In_479,In_1027);
nand U178 (N_178,In_2765,In_2086);
xnor U179 (N_179,In_1572,In_1536);
xnor U180 (N_180,In_1454,In_592);
and U181 (N_181,In_636,In_2026);
nor U182 (N_182,In_1338,In_670);
and U183 (N_183,In_939,In_2093);
nand U184 (N_184,In_1830,In_2551);
and U185 (N_185,In_2761,In_2173);
or U186 (N_186,In_1482,In_924);
nand U187 (N_187,In_302,In_2586);
and U188 (N_188,In_2064,In_2992);
or U189 (N_189,In_2111,In_1435);
xor U190 (N_190,In_1191,In_1940);
nor U191 (N_191,In_2662,In_2972);
and U192 (N_192,In_680,In_2728);
nand U193 (N_193,In_1787,In_2123);
and U194 (N_194,In_805,In_1718);
nor U195 (N_195,In_1147,In_2505);
or U196 (N_196,In_242,In_1092);
nand U197 (N_197,In_1225,In_877);
and U198 (N_198,In_971,In_1327);
or U199 (N_199,In_1906,In_642);
nand U200 (N_200,In_1390,In_80);
nor U201 (N_201,In_2210,In_1568);
or U202 (N_202,In_746,In_1333);
or U203 (N_203,In_2654,In_1737);
nor U204 (N_204,In_240,In_1965);
or U205 (N_205,In_2325,In_2360);
nand U206 (N_206,In_2293,In_1253);
xor U207 (N_207,In_1023,In_541);
nor U208 (N_208,In_2517,In_547);
or U209 (N_209,In_2045,In_2219);
or U210 (N_210,In_1348,In_371);
or U211 (N_211,In_78,In_1725);
nand U212 (N_212,In_2596,In_2049);
nor U213 (N_213,In_1703,In_691);
nand U214 (N_214,In_2228,In_2750);
nor U215 (N_215,In_260,In_2035);
nor U216 (N_216,In_1218,In_241);
nor U217 (N_217,In_514,In_497);
xnor U218 (N_218,In_28,In_1026);
nor U219 (N_219,In_2158,In_1901);
or U220 (N_220,In_2274,In_1973);
and U221 (N_221,In_222,In_1972);
nand U222 (N_222,In_865,In_716);
nand U223 (N_223,In_2680,In_4);
and U224 (N_224,In_1564,In_156);
and U225 (N_225,In_1504,In_1583);
or U226 (N_226,In_2981,In_2617);
and U227 (N_227,In_1215,In_1899);
and U228 (N_228,In_2132,In_2808);
and U229 (N_229,In_923,In_1721);
xor U230 (N_230,In_2094,In_976);
nand U231 (N_231,In_2633,In_2373);
and U232 (N_232,In_824,In_2595);
nand U233 (N_233,In_54,In_1616);
nand U234 (N_234,In_1122,In_267);
or U235 (N_235,In_406,In_1066);
nand U236 (N_236,In_1683,In_82);
nand U237 (N_237,In_2143,In_2526);
or U238 (N_238,In_891,In_89);
xor U239 (N_239,In_1924,In_1910);
xnor U240 (N_240,In_1278,In_1345);
xnor U241 (N_241,In_1809,In_2673);
xnor U242 (N_242,In_413,In_896);
or U243 (N_243,In_1734,In_1374);
or U244 (N_244,In_1007,In_2768);
or U245 (N_245,In_218,In_2098);
nand U246 (N_246,In_2987,In_615);
and U247 (N_247,In_692,In_71);
nor U248 (N_248,In_571,In_621);
or U249 (N_249,In_2108,In_2496);
or U250 (N_250,In_2090,In_1493);
and U251 (N_251,In_2212,In_121);
or U252 (N_252,In_2804,In_1395);
and U253 (N_253,In_1352,In_1197);
xor U254 (N_254,In_261,In_894);
nand U255 (N_255,In_577,In_1756);
and U256 (N_256,In_2802,In_2783);
xor U257 (N_257,In_1793,In_2477);
nor U258 (N_258,In_2381,In_119);
or U259 (N_259,In_1356,In_210);
nand U260 (N_260,In_2061,In_2065);
or U261 (N_261,In_125,In_1794);
xor U262 (N_262,In_596,In_2348);
nand U263 (N_263,In_103,In_2054);
nor U264 (N_264,In_1214,In_1724);
and U265 (N_265,In_1047,In_216);
xor U266 (N_266,In_644,In_1112);
nand U267 (N_267,In_1815,In_2590);
or U268 (N_268,In_1260,In_1652);
nand U269 (N_269,In_1001,In_2088);
nand U270 (N_270,In_2421,In_247);
and U271 (N_271,In_1323,In_1257);
or U272 (N_272,In_1510,In_1726);
and U273 (N_273,In_36,In_2195);
nand U274 (N_274,In_1707,In_286);
nor U275 (N_275,In_1785,In_1711);
and U276 (N_276,In_3,In_2247);
nand U277 (N_277,In_1020,In_1470);
nand U278 (N_278,In_75,In_139);
nand U279 (N_279,In_1545,In_985);
nand U280 (N_280,In_1689,In_2025);
nand U281 (N_281,In_602,In_850);
or U282 (N_282,In_363,In_1773);
or U283 (N_283,In_280,In_803);
nor U284 (N_284,In_1506,In_738);
or U285 (N_285,In_1919,In_1762);
and U286 (N_286,In_834,In_2647);
nand U287 (N_287,In_2503,In_344);
xnor U288 (N_288,In_49,In_1177);
or U289 (N_289,In_698,In_432);
nand U290 (N_290,In_98,In_1881);
nand U291 (N_291,In_1701,In_2506);
nor U292 (N_292,In_742,In_1513);
nand U293 (N_293,In_1832,In_763);
nor U294 (N_294,In_2403,In_869);
nor U295 (N_295,In_2848,In_2606);
xnor U296 (N_296,In_910,In_1249);
or U297 (N_297,In_1402,In_1124);
xor U298 (N_298,In_2695,In_1639);
nand U299 (N_299,In_2914,In_2311);
xor U300 (N_300,In_2600,In_1275);
and U301 (N_301,In_251,In_1532);
or U302 (N_302,In_600,In_1592);
nor U303 (N_303,In_93,In_2370);
xor U304 (N_304,In_1811,In_560);
xnor U305 (N_305,In_2508,In_1552);
xor U306 (N_306,In_467,In_2137);
xor U307 (N_307,In_164,In_1546);
nand U308 (N_308,In_2256,In_1512);
nor U309 (N_309,In_2157,In_2152);
or U310 (N_310,In_2242,In_1846);
or U311 (N_311,In_2085,In_1959);
nand U312 (N_312,In_2394,In_702);
and U313 (N_313,In_2336,In_2609);
nor U314 (N_314,In_2744,In_2805);
nand U315 (N_315,In_303,In_484);
nand U316 (N_316,In_84,In_2577);
and U317 (N_317,In_2361,In_627);
nor U318 (N_318,In_2717,In_1999);
or U319 (N_319,In_2060,In_2007);
xor U320 (N_320,In_2611,In_2892);
xnor U321 (N_321,In_320,In_516);
nor U322 (N_322,In_209,In_2328);
or U323 (N_323,In_706,In_1378);
xor U324 (N_324,In_1033,In_1464);
xor U325 (N_325,In_1322,In_1097);
nand U326 (N_326,In_245,In_1799);
and U327 (N_327,In_384,In_1219);
or U328 (N_328,In_843,In_2041);
nand U329 (N_329,In_150,In_291);
nor U330 (N_330,In_1181,In_1984);
nor U331 (N_331,In_1991,In_1364);
xnor U332 (N_332,In_2658,In_1538);
or U333 (N_333,In_1942,In_1054);
nand U334 (N_334,In_2012,In_2204);
or U335 (N_335,In_2890,In_466);
or U336 (N_336,In_1331,In_1918);
nand U337 (N_337,In_262,In_259);
nand U338 (N_338,In_2430,In_515);
and U339 (N_339,In_2115,In_788);
nand U340 (N_340,In_268,In_2493);
nand U341 (N_341,In_1473,In_2146);
and U342 (N_342,In_332,In_1911);
and U343 (N_343,In_2509,In_208);
and U344 (N_344,In_2375,In_2928);
nand U345 (N_345,In_312,In_783);
nand U346 (N_346,In_1507,In_2067);
nor U347 (N_347,In_1647,In_159);
and U348 (N_348,In_87,In_2033);
and U349 (N_349,In_1343,In_1167);
and U350 (N_350,In_270,In_1824);
nor U351 (N_351,In_2202,In_781);
or U352 (N_352,In_431,In_21);
nand U353 (N_353,In_2613,In_2135);
and U354 (N_354,In_1710,In_2314);
and U355 (N_355,In_2646,In_2891);
nand U356 (N_356,In_810,In_2667);
xnor U357 (N_357,In_1818,In_2747);
nand U358 (N_358,In_534,In_864);
xor U359 (N_359,In_229,In_1666);
or U360 (N_360,In_61,In_1246);
and U361 (N_361,In_518,In_306);
xor U362 (N_362,In_2557,In_884);
nand U363 (N_363,In_2639,In_2075);
nand U364 (N_364,In_1530,In_393);
xor U365 (N_365,In_2925,In_1080);
or U366 (N_366,In_1606,In_2316);
and U367 (N_367,In_2465,In_915);
or U368 (N_368,In_2056,In_2870);
or U369 (N_369,In_618,In_2701);
or U370 (N_370,In_1212,In_2295);
and U371 (N_371,In_2462,In_2196);
or U372 (N_372,In_1895,In_2929);
or U373 (N_373,In_1952,In_1983);
and U374 (N_374,In_2840,In_1727);
and U375 (N_375,In_419,In_246);
nand U376 (N_376,In_775,In_2597);
xor U377 (N_377,In_2977,In_1086);
and U378 (N_378,In_860,In_1759);
nand U379 (N_379,In_774,In_1735);
and U380 (N_380,In_1025,In_2034);
nand U381 (N_381,In_1637,In_2058);
nor U382 (N_382,In_172,In_163);
nor U383 (N_383,In_1034,In_352);
and U384 (N_384,In_1143,In_2440);
nand U385 (N_385,In_2005,In_2766);
xor U386 (N_386,In_381,In_663);
and U387 (N_387,In_287,In_890);
or U388 (N_388,In_2089,In_1837);
nand U389 (N_389,In_1106,In_658);
nor U390 (N_390,In_606,In_83);
or U391 (N_391,In_1315,In_1360);
xnor U392 (N_392,In_122,In_528);
and U393 (N_393,In_1957,In_1584);
nand U394 (N_394,In_1865,In_391);
nand U395 (N_395,In_31,In_705);
nor U396 (N_396,In_2941,In_1277);
nand U397 (N_397,In_948,In_356);
and U398 (N_398,In_58,In_490);
and U399 (N_399,In_1758,In_2299);
nand U400 (N_400,In_2935,In_32);
nand U401 (N_401,In_2663,In_24);
nand U402 (N_402,In_2415,In_127);
nand U403 (N_403,In_480,In_2223);
and U404 (N_404,In_1969,In_2006);
xnor U405 (N_405,In_1457,In_442);
xor U406 (N_406,In_1082,In_2507);
or U407 (N_407,In_2413,In_2704);
and U408 (N_408,In_2079,In_1303);
nor U409 (N_409,In_2520,In_2326);
nand U410 (N_410,In_2866,In_650);
nand U411 (N_411,In_111,In_2934);
nor U412 (N_412,In_885,In_696);
xnor U413 (N_413,In_279,In_1998);
or U414 (N_414,In_2792,In_2958);
nand U415 (N_415,In_1359,In_1292);
nor U416 (N_416,In_1077,In_2930);
and U417 (N_417,In_1062,In_1676);
xor U418 (N_418,In_1800,In_1294);
xor U419 (N_419,In_2163,In_1105);
or U420 (N_420,In_2306,In_2057);
nand U421 (N_421,In_1646,In_1888);
xor U422 (N_422,In_2851,In_929);
and U423 (N_423,In_81,In_2429);
and U424 (N_424,In_559,In_2533);
or U425 (N_425,In_1560,In_858);
and U426 (N_426,In_1529,In_2923);
xnor U427 (N_427,In_2082,In_1185);
and U428 (N_428,In_275,In_2450);
and U429 (N_429,In_1607,In_996);
and U430 (N_430,In_2153,In_2277);
or U431 (N_431,In_257,In_2573);
xnor U432 (N_432,In_2463,In_1188);
nand U433 (N_433,In_196,In_1366);
nor U434 (N_434,In_2754,In_1650);
and U435 (N_435,In_2491,In_2814);
and U436 (N_436,In_1937,In_394);
nor U437 (N_437,In_2829,In_811);
nor U438 (N_438,In_2736,In_2409);
nand U439 (N_439,In_1989,In_1685);
xor U440 (N_440,In_1199,In_1131);
xor U441 (N_441,In_187,In_2347);
and U442 (N_442,In_368,In_2340);
nor U443 (N_443,In_1004,In_1605);
nand U444 (N_444,In_2248,In_1829);
or U445 (N_445,In_1067,In_2124);
xor U446 (N_446,In_1856,In_597);
and U447 (N_447,In_1967,In_2234);
nor U448 (N_448,In_1934,In_2113);
and U449 (N_449,In_2339,In_687);
nand U450 (N_450,In_784,In_1005);
and U451 (N_451,In_2017,In_1515);
and U452 (N_452,In_2458,In_2010);
nand U453 (N_453,In_2742,In_460);
nand U454 (N_454,In_1298,In_881);
and U455 (N_455,In_1019,In_1165);
nor U456 (N_456,In_1180,In_17);
or U457 (N_457,In_1979,In_2363);
and U458 (N_458,In_1035,In_2666);
nand U459 (N_459,In_1553,In_817);
nand U460 (N_460,In_1491,In_1626);
xnor U461 (N_461,In_2187,In_1295);
nor U462 (N_462,In_1687,In_2232);
xnor U463 (N_463,In_1598,In_1776);
and U464 (N_464,In_2259,In_2881);
nor U465 (N_465,In_1614,In_1096);
nand U466 (N_466,In_1933,In_1636);
or U467 (N_467,In_362,In_2402);
and U468 (N_468,In_1833,In_2694);
or U469 (N_469,In_733,In_128);
xor U470 (N_470,In_2907,In_1358);
and U471 (N_471,In_1006,In_2267);
and U472 (N_472,In_837,In_157);
nor U473 (N_473,In_779,In_1878);
nand U474 (N_474,In_999,In_1060);
or U475 (N_475,In_2599,In_1094);
xor U476 (N_476,In_1828,In_1949);
or U477 (N_477,In_1342,In_673);
xnor U478 (N_478,In_1977,In_463);
nor U479 (N_479,In_2386,In_2343);
xor U480 (N_480,In_792,In_1715);
and U481 (N_481,In_188,In_85);
or U482 (N_482,In_1115,In_1521);
nor U483 (N_483,In_887,In_2757);
nand U484 (N_484,In_1015,In_57);
xnor U485 (N_485,In_324,In_269);
and U486 (N_486,In_1479,In_682);
or U487 (N_487,In_2591,In_1254);
or U488 (N_488,In_132,In_2823);
nand U489 (N_489,In_836,In_1953);
or U490 (N_490,In_2240,In_2784);
nor U491 (N_491,In_1770,In_1677);
xnor U492 (N_492,In_2063,In_594);
nand U493 (N_493,In_2653,In_1523);
xnor U494 (N_494,In_2184,In_1875);
or U495 (N_495,In_102,In_1618);
nand U496 (N_496,In_2615,In_1179);
nor U497 (N_497,In_2344,In_866);
nand U498 (N_498,In_2674,In_239);
or U499 (N_499,In_822,In_1672);
nand U500 (N_500,In_2700,In_2983);
or U501 (N_501,In_1806,In_1961);
and U502 (N_502,In_761,In_243);
nor U503 (N_503,In_1698,In_1270);
and U504 (N_504,In_815,In_277);
xnor U505 (N_505,In_2976,In_2576);
or U506 (N_506,In_2015,In_1855);
or U507 (N_507,In_1763,In_609);
xnor U508 (N_508,In_1950,In_2812);
and U509 (N_509,In_2560,In_46);
nor U510 (N_510,In_138,In_2873);
nand U511 (N_511,In_2745,In_964);
xnor U512 (N_512,In_174,In_233);
xor U513 (N_513,In_2366,In_1091);
nor U514 (N_514,In_1423,In_622);
nor U515 (N_515,In_109,In_2356);
and U516 (N_516,In_713,In_940);
nand U517 (N_517,In_2036,In_537);
nor U518 (N_518,In_347,In_2691);
nand U519 (N_519,In_255,In_2974);
and U520 (N_520,In_2352,In_2955);
xor U521 (N_521,In_728,In_142);
or U522 (N_522,In_852,In_2416);
or U523 (N_523,In_2250,In_6);
and U524 (N_524,In_1095,In_2109);
and U525 (N_525,In_1641,In_1980);
nand U526 (N_526,In_357,In_1825);
xor U527 (N_527,In_443,In_2452);
xor U528 (N_528,In_1995,In_2358);
nor U529 (N_529,In_1736,In_906);
nand U530 (N_530,In_1603,In_1838);
nor U531 (N_531,In_2817,In_1932);
nor U532 (N_532,In_1391,In_2351);
nand U533 (N_533,In_513,In_1843);
nor U534 (N_534,In_2948,In_576);
nor U535 (N_535,In_2852,In_1458);
xor U536 (N_536,In_662,In_1709);
nor U537 (N_537,In_1410,In_1892);
and U538 (N_538,In_2203,In_646);
xor U539 (N_539,In_720,In_2475);
and U540 (N_540,In_1242,In_1853);
xnor U541 (N_541,In_2535,In_2149);
or U542 (N_542,In_153,In_703);
xnor U543 (N_543,In_2298,In_1923);
or U544 (N_544,In_2661,In_2371);
nor U545 (N_545,In_2579,In_2669);
xor U546 (N_546,In_660,In_1363);
nand U547 (N_547,In_1139,In_629);
or U548 (N_548,In_2534,In_1289);
or U549 (N_549,In_1699,In_582);
xor U550 (N_550,In_2279,In_2698);
and U551 (N_551,In_1857,In_430);
and U552 (N_552,In_2114,In_264);
xor U553 (N_553,In_114,In_830);
xor U554 (N_554,In_1820,In_2846);
nor U555 (N_555,In_2994,In_838);
or U556 (N_556,In_2956,In_397);
nor U557 (N_557,In_1335,In_619);
nor U558 (N_558,In_694,In_1399);
and U559 (N_559,In_182,In_135);
and U560 (N_560,In_29,In_2231);
xor U561 (N_561,In_1002,In_2690);
xnor U562 (N_562,In_2194,In_2702);
xnor U563 (N_563,In_1981,In_828);
and U564 (N_564,In_53,In_1213);
xnor U565 (N_565,In_701,In_334);
or U566 (N_566,In_1908,In_2697);
nor U567 (N_567,In_399,In_876);
nor U568 (N_568,In_2338,In_2550);
xor U569 (N_569,In_955,In_2206);
and U570 (N_570,In_140,In_2922);
or U571 (N_571,In_1051,In_2376);
nand U572 (N_572,In_1831,In_2320);
or U573 (N_573,In_2810,In_1587);
nand U574 (N_574,In_1944,In_664);
or U575 (N_575,In_411,In_1472);
nand U576 (N_576,In_700,In_1319);
nand U577 (N_577,In_711,In_2377);
or U578 (N_578,In_2624,In_2582);
and U579 (N_579,In_1621,In_1245);
and U580 (N_580,In_2179,In_203);
or U581 (N_581,In_486,In_1424);
nor U582 (N_582,In_1642,In_1779);
nor U583 (N_583,In_358,In_1471);
xor U584 (N_584,In_1362,In_952);
nand U585 (N_585,In_2683,In_2889);
nor U586 (N_586,In_512,In_1702);
or U587 (N_587,In_2029,In_2159);
or U588 (N_588,In_2637,In_983);
nand U589 (N_589,In_1873,In_2723);
or U590 (N_590,In_1964,In_808);
or U591 (N_591,In_1017,In_386);
and U592 (N_592,In_1003,In_1381);
xnor U593 (N_593,In_2906,In_2896);
xor U594 (N_594,In_2969,In_481);
xnor U595 (N_595,In_1373,In_2221);
or U596 (N_596,In_2608,In_227);
nor U597 (N_597,In_1663,In_1669);
nor U598 (N_598,In_2838,In_1633);
and U599 (N_599,In_2975,In_1891);
nor U600 (N_600,In_2729,In_743);
or U601 (N_601,In_1135,In_1445);
and U602 (N_602,In_252,In_10);
nand U603 (N_603,In_278,In_695);
and U604 (N_604,In_1437,In_1262);
and U605 (N_605,In_143,In_2488);
nor U606 (N_606,In_1414,In_86);
nand U607 (N_607,In_548,In_1372);
xor U608 (N_608,In_1772,In_2688);
and U609 (N_609,In_1041,In_1063);
and U610 (N_610,In_659,In_2562);
xor U611 (N_611,In_942,In_856);
or U612 (N_612,In_734,In_2815);
or U613 (N_613,In_1922,In_2913);
or U614 (N_614,In_2322,In_2909);
nor U615 (N_615,In_2249,In_2492);
and U616 (N_616,In_517,In_11);
and U617 (N_617,In_1451,In_1098);
and U618 (N_618,In_714,In_1406);
nand U619 (N_619,In_1255,In_1909);
nor U620 (N_620,In_770,In_2368);
or U621 (N_621,In_1137,In_2200);
nor U622 (N_622,In_2933,In_2470);
nor U623 (N_623,In_2937,In_524);
and U624 (N_624,In_45,In_1556);
nor U625 (N_625,In_1533,In_1740);
nand U626 (N_626,In_2013,In_1591);
nand U627 (N_627,In_2502,In_2382);
and U628 (N_628,In_1588,In_950);
nor U629 (N_629,In_2997,In_1201);
nor U630 (N_630,In_1182,In_570);
xnor U631 (N_631,In_1671,In_1037);
xor U632 (N_632,In_772,In_2481);
nand U633 (N_633,In_66,In_2213);
or U634 (N_634,In_1744,In_2827);
or U635 (N_635,In_1171,In_892);
xnor U636 (N_636,In_392,In_2885);
or U637 (N_637,In_1797,In_2656);
nand U638 (N_638,In_797,In_1622);
or U639 (N_639,In_2785,In_452);
xnor U640 (N_640,In_9,In_2944);
nor U641 (N_641,In_1039,In_2243);
nand U642 (N_642,In_390,In_1397);
xor U643 (N_643,In_2603,In_1145);
or U644 (N_644,In_2799,In_335);
or U645 (N_645,In_2857,In_2304);
or U646 (N_646,In_1935,In_1417);
nor U647 (N_647,In_2169,In_1049);
xnor U648 (N_648,In_1839,In_1580);
nand U649 (N_649,In_1519,In_2048);
and U650 (N_650,In_2862,In_1259);
xor U651 (N_651,In_2952,In_2264);
and U652 (N_652,In_920,In_2616);
and U653 (N_653,In_2631,In_1539);
xor U654 (N_654,In_2924,In_2388);
and U655 (N_655,In_684,In_1387);
or U656 (N_656,In_2869,In_1184);
xor U657 (N_657,In_2764,In_2425);
and U658 (N_658,In_2074,In_2448);
nand U659 (N_659,In_2883,In_451);
and U660 (N_660,In_1475,In_165);
nor U661 (N_661,In_2781,In_2133);
nand U662 (N_662,In_1609,In_1681);
nand U663 (N_663,In_2853,In_458);
xnor U664 (N_664,In_758,In_1574);
xnor U665 (N_665,In_2174,In_2392);
xnor U666 (N_666,In_2457,In_861);
or U667 (N_667,In_1601,In_160);
or U668 (N_668,In_305,In_152);
and U669 (N_669,In_1914,In_967);
xor U670 (N_670,In_2456,In_1594);
or U671 (N_671,In_2028,In_1927);
nor U672 (N_672,In_2001,In_1404);
and U673 (N_673,In_1655,In_201);
or U674 (N_674,In_2125,In_2252);
or U675 (N_675,In_193,In_1496);
nand U676 (N_676,In_2192,In_879);
or U677 (N_677,In_941,In_67);
or U678 (N_678,In_250,In_2165);
nand U679 (N_679,In_1528,In_1713);
or U680 (N_680,In_1930,In_464);
and U681 (N_681,In_806,In_1227);
and U682 (N_682,In_200,In_807);
nor U683 (N_683,In_2332,In_848);
xor U684 (N_684,In_563,In_666);
xor U685 (N_685,In_14,In_1469);
xor U686 (N_686,In_1870,In_1194);
xnor U687 (N_687,In_2294,In_1876);
xor U688 (N_688,In_913,In_2733);
nor U689 (N_689,In_2209,In_2878);
nor U690 (N_690,In_529,In_921);
nor U691 (N_691,In_773,In_2003);
or U692 (N_692,In_2980,In_2712);
or U693 (N_693,In_519,In_1526);
nor U694 (N_694,In_2426,In_2540);
or U695 (N_695,In_905,In_1291);
or U696 (N_696,In_2767,In_2197);
nand U697 (N_697,In_1453,In_2437);
and U698 (N_698,In_2302,In_281);
or U699 (N_699,In_1840,In_2743);
xor U700 (N_700,In_721,In_316);
and U701 (N_701,In_1172,In_2105);
or U702 (N_702,In_1819,In_2389);
nand U703 (N_703,In_693,In_987);
and U704 (N_704,In_1585,In_558);
xor U705 (N_705,In_1883,In_2385);
xor U706 (N_706,In_813,In_2436);
nor U707 (N_707,In_74,In_1929);
xor U708 (N_708,In_1841,In_979);
or U709 (N_709,In_1244,In_1673);
or U710 (N_710,In_553,In_648);
xor U711 (N_711,In_791,In_2886);
and U712 (N_712,In_2333,In_2651);
and U713 (N_713,In_2161,In_980);
nand U714 (N_714,In_1383,In_1450);
xor U715 (N_715,In_1520,In_1134);
nand U716 (N_716,In_2833,In_1440);
and U717 (N_717,In_863,In_2879);
or U718 (N_718,In_1071,In_1578);
nor U719 (N_719,In_1290,In_1679);
or U720 (N_720,In_1768,In_2850);
nor U721 (N_721,In_1729,In_862);
or U722 (N_722,In_1222,In_2275);
or U723 (N_723,In_1456,In_2208);
and U724 (N_724,In_2798,In_1272);
nor U725 (N_725,In_786,In_2705);
and U726 (N_726,In_2970,In_1382);
nor U727 (N_727,In_1619,In_489);
or U728 (N_728,In_1745,In_1130);
and U729 (N_729,In_552,In_1032);
nand U730 (N_730,In_722,In_314);
and U731 (N_731,In_556,In_2739);
xor U732 (N_732,In_1221,In_1146);
xnor U733 (N_733,In_333,In_930);
nand U734 (N_734,In_421,In_1396);
or U735 (N_735,In_909,In_678);
nand U736 (N_736,In_96,In_690);
nand U737 (N_737,In_2037,In_372);
nor U738 (N_738,In_2059,In_2069);
and U739 (N_739,In_1128,In_1334);
and U740 (N_740,In_1065,In_1835);
and U741 (N_741,In_1175,In_1110);
and U742 (N_742,In_2527,In_1321);
nor U743 (N_743,In_282,In_2272);
xnor U744 (N_744,In_1653,In_408);
or U745 (N_745,In_1014,In_1732);
or U746 (N_746,In_2610,In_557);
nand U747 (N_747,In_448,In_361);
nor U748 (N_748,In_2672,In_655);
nand U749 (N_749,In_217,In_1848);
xor U750 (N_750,In_1079,In_2134);
or U751 (N_751,In_2002,In_2623);
and U752 (N_752,In_19,In_2245);
and U753 (N_753,In_1662,In_1107);
nand U754 (N_754,In_2856,In_1059);
nor U755 (N_755,In_436,In_2156);
nor U756 (N_756,In_2660,In_226);
xnor U757 (N_757,In_2350,In_709);
nor U758 (N_758,In_936,In_377);
xor U759 (N_759,In_59,In_2991);
nor U760 (N_760,In_133,In_723);
or U761 (N_761,In_661,In_645);
or U762 (N_762,In_1746,In_477);
or U763 (N_763,In_1088,In_340);
or U764 (N_764,In_587,In_1144);
nor U765 (N_765,In_373,In_886);
nor U766 (N_766,In_162,In_185);
nor U767 (N_767,In_1741,In_984);
nand U768 (N_768,In_1668,In_161);
and U769 (N_769,In_2420,In_1596);
nor U770 (N_770,In_2355,In_1480);
nand U771 (N_771,In_1325,In_1483);
and U772 (N_772,In_1629,In_56);
nor U773 (N_773,In_2071,In_972);
nand U774 (N_774,In_2581,In_710);
nand U775 (N_775,In_2391,In_2988);
xor U776 (N_776,In_2166,In_1103);
xnor U777 (N_777,In_2148,In_2614);
xnor U778 (N_778,In_1649,In_355);
nor U779 (N_779,In_898,In_1237);
nand U780 (N_780,In_818,In_1238);
nor U781 (N_781,In_2793,In_981);
or U782 (N_782,In_345,In_726);
and U783 (N_783,In_2021,In_43);
or U784 (N_784,In_1534,In_1386);
xnor U785 (N_785,In_963,In_1738);
and U786 (N_786,In_542,In_1422);
nand U787 (N_787,In_1189,In_441);
nand U788 (N_788,In_105,In_769);
nand U789 (N_789,In_248,In_2051);
xnor U790 (N_790,In_376,In_2769);
nand U791 (N_791,In_604,In_2268);
or U792 (N_792,In_809,In_844);
xor U793 (N_793,In_1670,In_403);
and U794 (N_794,In_2432,In_614);
and U795 (N_795,In_584,In_1783);
or U796 (N_796,In_2536,In_842);
nand U797 (N_797,In_2730,In_2327);
xor U798 (N_798,In_2276,In_1600);
and U799 (N_799,In_1499,In_2224);
nor U800 (N_800,In_1656,In_831);
and U801 (N_801,In_1309,In_1114);
nand U802 (N_802,In_1297,In_106);
nand U803 (N_803,In_551,In_342);
nand U804 (N_804,In_253,In_2910);
nor U805 (N_805,In_1341,In_99);
and U806 (N_806,In_1567,In_847);
or U807 (N_807,In_1658,In_186);
xor U808 (N_808,In_2825,In_35);
and U809 (N_809,In_2861,In_343);
nand U810 (N_810,In_908,In_995);
or U811 (N_811,In_353,In_1118);
nor U812 (N_812,In_1243,In_2244);
nor U813 (N_813,In_318,In_1657);
or U814 (N_814,In_1016,In_426);
xnor U815 (N_815,In_1376,In_1176);
or U816 (N_816,In_2424,In_369);
nand U817 (N_817,In_1070,In_1862);
xnor U818 (N_818,In_2395,In_704);
nand U819 (N_819,In_263,In_1036);
or U820 (N_820,In_641,In_2172);
nor U821 (N_821,In_346,In_2076);
xor U822 (N_822,In_2464,In_630);
xor U823 (N_823,In_1367,In_2038);
nor U824 (N_824,In_2966,In_2953);
or U825 (N_825,In_991,In_632);
xor U826 (N_826,In_1064,In_2313);
nand U827 (N_827,In_1154,In_540);
xor U828 (N_828,In_800,In_2096);
or U829 (N_829,In_2397,In_2710);
and U830 (N_830,In_2241,In_2258);
xnor U831 (N_831,In_1743,In_536);
nand U832 (N_832,In_1566,In_2707);
or U833 (N_833,In_904,In_1575);
nand U834 (N_834,In_1645,In_396);
and U835 (N_835,In_1009,In_1099);
xnor U836 (N_836,In_1885,In_2685);
nand U837 (N_837,In_1102,In_2122);
nor U838 (N_838,In_1789,In_1211);
and U839 (N_839,In_1571,In_1719);
xnor U840 (N_840,In_1731,In_2020);
nor U841 (N_841,In_832,In_502);
nand U842 (N_842,In_1694,In_2398);
and U843 (N_843,In_1429,In_1807);
xor U844 (N_844,In_1187,In_410);
nor U845 (N_845,In_2471,In_1161);
xor U846 (N_846,In_2659,In_41);
nor U847 (N_847,In_2405,In_1527);
or U848 (N_848,In_1256,In_2734);
and U849 (N_849,In_1705,In_483);
nor U850 (N_850,In_2920,In_1573);
or U851 (N_851,In_1186,In_501);
or U852 (N_852,In_1487,In_2900);
xor U853 (N_853,In_2281,In_900);
xor U854 (N_854,In_736,In_565);
nand U855 (N_855,In_1867,In_814);
xnor U856 (N_856,In_1674,In_2901);
nor U857 (N_857,In_1728,In_2867);
xnor U858 (N_858,In_1224,In_2578);
or U859 (N_859,In_364,In_2335);
nand U860 (N_860,In_2140,In_2040);
nor U861 (N_861,In_2588,In_1781);
xnor U862 (N_862,In_199,In_2811);
or U863 (N_863,In_2543,In_969);
or U864 (N_864,In_1784,In_1976);
and U865 (N_865,In_348,In_1877);
or U866 (N_866,In_561,In_190);
and U867 (N_867,In_638,In_1804);
nand U868 (N_868,In_798,In_825);
nand U869 (N_869,In_1792,In_2621);
and U870 (N_870,In_2842,In_1565);
nor U871 (N_871,In_766,In_2649);
nand U872 (N_872,In_2569,In_0);
or U873 (N_873,In_735,In_1613);
nor U874 (N_874,In_994,In_2417);
or U875 (N_875,In_2459,In_184);
nor U876 (N_876,In_2167,In_932);
and U877 (N_877,In_992,In_951);
xnor U878 (N_878,In_1505,In_60);
nand U879 (N_879,In_323,In_1985);
and U880 (N_880,In_2926,In_2776);
xor U881 (N_881,In_2565,In_764);
xor U882 (N_882,In_2773,In_2584);
nand U883 (N_883,In_151,In_2819);
or U884 (N_884,In_2323,In_2451);
or U885 (N_885,In_754,In_79);
nor U886 (N_886,In_665,In_1305);
nand U887 (N_887,In_1251,In_48);
nand U888 (N_888,In_740,In_1502);
and U889 (N_889,In_1882,In_1489);
xnor U890 (N_890,In_2479,In_2899);
or U891 (N_891,In_385,In_2439);
nand U892 (N_892,In_2387,In_2238);
and U893 (N_893,In_1282,In_730);
xnor U894 (N_894,In_1089,In_1328);
xnor U895 (N_895,In_1936,In_2444);
nor U896 (N_896,In_2859,In_2715);
nor U897 (N_897,In_1299,In_643);
nor U898 (N_898,In_522,In_2824);
xnor U899 (N_899,In_482,In_455);
nor U900 (N_900,In_1913,In_1153);
and U901 (N_901,In_2217,In_1116);
nor U902 (N_902,In_1537,In_1774);
and U903 (N_903,In_1310,In_2215);
xnor U904 (N_904,In_1577,In_1956);
xor U905 (N_905,In_966,In_2627);
nand U906 (N_906,In_2999,In_1893);
and U907 (N_907,In_767,In_76);
and U908 (N_908,In_2894,In_284);
nor U909 (N_909,In_1193,In_1413);
nand U910 (N_910,In_1155,In_2843);
nand U911 (N_911,In_2927,In_2982);
and U912 (N_912,In_753,In_749);
and U913 (N_913,In_1057,In_1816);
nor U914 (N_914,In_2310,In_2273);
nor U915 (N_915,In_1233,In_1754);
nor U916 (N_916,In_2778,In_2500);
nor U917 (N_917,In_1263,In_2548);
and U918 (N_918,In_1678,In_1008);
xor U919 (N_919,In_719,In_757);
nor U920 (N_920,In_1692,In_2874);
nor U921 (N_921,In_1667,In_588);
or U922 (N_922,In_2138,In_1132);
or U923 (N_923,In_1716,In_902);
nand U924 (N_924,In_1720,In_27);
or U925 (N_925,In_1285,In_1195);
nor U926 (N_926,In_2962,In_566);
nand U927 (N_927,In_699,In_1013);
nand U928 (N_928,In_2772,In_2971);
nor U929 (N_929,In_598,In_912);
xnor U930 (N_930,In_322,In_1970);
and U931 (N_931,In_2620,In_493);
nand U932 (N_932,In_33,In_1190);
or U933 (N_933,In_544,In_112);
and U934 (N_934,In_569,In_2681);
nor U935 (N_935,In_2070,In_2942);
xor U936 (N_936,In_1239,In_409);
nor U937 (N_937,In_819,In_789);
nand U938 (N_938,In_1220,In_485);
xor U939 (N_939,In_2303,In_1235);
and U940 (N_940,In_494,In_2832);
or U941 (N_941,In_1337,In_593);
nand U942 (N_942,In_799,In_2722);
and U943 (N_943,In_23,In_1992);
or U944 (N_944,In_439,In_1557);
nand U945 (N_945,In_415,In_2180);
nor U946 (N_946,In_1069,In_2102);
nand U947 (N_947,In_1946,In_123);
xnor U948 (N_948,In_607,In_2803);
or U949 (N_949,In_2511,In_2478);
or U950 (N_950,In_708,In_2236);
xnor U951 (N_951,In_2435,In_1550);
or U952 (N_952,In_315,In_1795);
and U953 (N_953,In_1813,In_2198);
nand U954 (N_954,In_1905,In_2253);
and U955 (N_955,In_2725,In_341);
or U956 (N_956,In_616,In_1675);
xnor U957 (N_957,In_2278,In_231);
or U958 (N_958,In_2472,In_1631);
or U959 (N_959,In_367,In_626);
or U960 (N_960,In_674,In_2741);
and U961 (N_961,In_1928,In_750);
and U962 (N_962,In_2246,In_974);
and U963 (N_963,In_313,In_2237);
or U964 (N_964,In_2752,In_2018);
nor U965 (N_965,In_2504,In_1162);
or U966 (N_966,In_295,In_1460);
xor U967 (N_967,In_2190,In_1462);
nor U968 (N_968,In_2822,In_2438);
nand U969 (N_969,In_1844,In_1022);
or U970 (N_970,In_531,In_729);
nor U971 (N_971,In_1271,In_1485);
nor U972 (N_972,In_1455,In_1660);
nor U973 (N_973,In_1812,In_1120);
nor U974 (N_974,In_2737,In_2547);
and U975 (N_975,In_2112,In_583);
or U976 (N_976,In_2538,In_1336);
and U977 (N_977,In_2188,In_532);
and U978 (N_978,In_72,In_1926);
nand U979 (N_979,In_589,In_454);
nand U980 (N_980,In_398,In_2270);
or U981 (N_981,In_1700,In_1159);
xnor U982 (N_982,In_564,In_1151);
nand U983 (N_983,In_2657,In_471);
or U984 (N_984,In_654,In_2476);
nand U985 (N_985,In_2746,In_1075);
nand U986 (N_986,In_1370,In_1503);
nand U987 (N_987,In_585,In_148);
or U988 (N_988,In_234,In_2898);
xnor U989 (N_989,In_290,In_2410);
nand U990 (N_990,In_2308,In_2142);
nor U991 (N_991,In_931,In_1582);
nand U992 (N_992,In_899,In_1907);
xnor U993 (N_993,In_2607,In_274);
nor U994 (N_994,In_2324,In_2524);
or U995 (N_995,In_155,In_2644);
nand U996 (N_996,In_755,In_1293);
nand U997 (N_997,In_2186,In_855);
or U998 (N_998,In_2068,In_1511);
nor U999 (N_999,In_474,In_2931);
or U1000 (N_1000,In_1548,In_1886);
nor U1001 (N_1001,In_1836,In_1081);
xnor U1002 (N_1002,In_2374,In_1494);
or U1003 (N_1003,In_2740,In_2959);
nor U1004 (N_1004,In_1042,In_1093);
nand U1005 (N_1005,In_953,In_2285);
and U1006 (N_1006,In_903,In_2062);
nand U1007 (N_1007,In_194,In_2235);
nand U1008 (N_1008,In_2495,In_100);
and U1009 (N_1009,In_2000,In_707);
and U1010 (N_1010,In_1712,In_960);
nand U1011 (N_1011,In_573,In_349);
and U1012 (N_1012,In_2189,In_2225);
or U1013 (N_1013,In_2687,In_311);
nor U1014 (N_1014,In_158,In_1248);
and U1015 (N_1015,In_2447,In_2307);
xnor U1016 (N_1016,In_823,In_2482);
or U1017 (N_1017,In_1076,In_2961);
and U1018 (N_1018,In_1955,In_1887);
nor U1019 (N_1019,In_685,In_469);
nor U1020 (N_1020,In_1704,In_1230);
nand U1021 (N_1021,In_1287,In_2321);
xnor U1022 (N_1022,In_1682,In_2260);
or U1023 (N_1023,In_2443,In_1226);
nand U1024 (N_1024,In_171,In_321);
nand U1025 (N_1025,In_1068,In_244);
nand U1026 (N_1026,In_1788,In_2794);
nand U1027 (N_1027,In_653,In_1866);
or U1028 (N_1028,In_2379,In_129);
nand U1029 (N_1029,In_962,In_2863);
or U1030 (N_1030,In_2486,In_301);
nand U1031 (N_1031,In_2497,In_2713);
xor U1032 (N_1032,In_689,In_70);
xor U1033 (N_1033,In_2554,In_1418);
and U1034 (N_1034,In_197,In_2289);
nand U1035 (N_1035,In_401,In_943);
nor U1036 (N_1036,In_69,In_1126);
or U1037 (N_1037,In_1680,In_2473);
nand U1038 (N_1038,In_851,In_1775);
xor U1039 (N_1039,In_1441,In_1296);
xnor U1040 (N_1040,In_288,In_429);
and U1041 (N_1041,In_2872,In_2871);
nand U1042 (N_1042,In_1474,In_724);
nor U1043 (N_1043,In_2510,In_874);
xor U1044 (N_1044,In_1884,In_213);
or U1045 (N_1045,In_2183,In_2139);
nor U1046 (N_1046,In_2466,In_2445);
and U1047 (N_1047,In_1149,In_2126);
nand U1048 (N_1048,In_1563,In_2796);
nand U1049 (N_1049,In_1595,In_2309);
xnor U1050 (N_1050,In_2380,In_1412);
and U1051 (N_1051,In_846,In_2708);
or U1052 (N_1052,In_1316,In_1780);
or U1053 (N_1053,In_776,In_1385);
nor U1054 (N_1054,In_2575,In_747);
xor U1055 (N_1055,In_1939,In_2181);
or U1056 (N_1056,In_1617,In_1751);
xnor U1057 (N_1057,In_1317,In_997);
xor U1058 (N_1058,In_1228,In_2893);
and U1059 (N_1059,In_2528,In_2055);
nor U1060 (N_1060,In_1380,In_2571);
nor U1061 (N_1061,In_2269,In_2758);
or U1062 (N_1062,In_73,In_2066);
and U1063 (N_1063,In_2330,In_628);
and U1064 (N_1064,In_1400,In_2629);
nor U1065 (N_1065,In_120,In_2199);
xor U1066 (N_1066,In_2908,In_434);
or U1067 (N_1067,In_2519,In_782);
xnor U1068 (N_1068,In_1300,In_476);
and U1069 (N_1069,In_417,In_2106);
and U1070 (N_1070,In_1659,In_1620);
nand U1071 (N_1071,In_414,In_444);
nand U1072 (N_1072,In_2911,In_2921);
or U1073 (N_1073,In_2222,In_1590);
xnor U1074 (N_1074,In_1261,In_298);
and U1075 (N_1075,In_2868,In_2684);
and U1076 (N_1076,In_2727,In_1318);
nor U1077 (N_1077,In_2151,In_1377);
nor U1078 (N_1078,In_258,In_101);
nor U1079 (N_1079,In_2731,In_1486);
xnor U1080 (N_1080,In_104,In_652);
xnor U1081 (N_1081,In_2233,In_1796);
and U1082 (N_1082,In_1823,In_1852);
xor U1083 (N_1083,In_2441,In_1686);
and U1084 (N_1084,In_211,In_1365);
and U1085 (N_1085,In_2383,In_1915);
and U1086 (N_1086,In_1073,In_2706);
xnor U1087 (N_1087,In_2905,In_2960);
nor U1088 (N_1088,In_25,In_379);
and U1089 (N_1089,In_145,In_2813);
or U1090 (N_1090,In_2762,In_2043);
nand U1091 (N_1091,In_1894,In_574);
or U1092 (N_1092,In_1558,In_2732);
nor U1093 (N_1093,In_2622,In_2749);
nor U1094 (N_1094,In_2696,In_2655);
or U1095 (N_1095,In_1962,In_914);
nand U1096 (N_1096,In_1802,In_1133);
or U1097 (N_1097,In_168,In_465);
or U1098 (N_1098,In_331,In_2523);
xor U1099 (N_1099,In_2835,In_826);
nand U1100 (N_1100,In_1324,In_2312);
and U1101 (N_1101,In_1900,In_624);
and U1102 (N_1102,In_1046,In_1880);
nand U1103 (N_1103,In_2101,In_1229);
xnor U1104 (N_1104,In_176,In_271);
nand U1105 (N_1105,In_1158,In_2978);
nor U1106 (N_1106,In_1896,In_77);
nor U1107 (N_1107,In_1525,In_2103);
nand U1108 (N_1108,In_2719,In_639);
xnor U1109 (N_1109,In_1954,In_2483);
nor U1110 (N_1110,In_2118,In_1274);
or U1111 (N_1111,In_872,In_1847);
and U1112 (N_1112,In_2428,In_1517);
xnor U1113 (N_1113,In_2720,In_2128);
or U1114 (N_1114,In_2014,In_2809);
and U1115 (N_1115,In_1043,In_1803);
and U1116 (N_1116,In_2022,In_1827);
nand U1117 (N_1117,In_2558,In_878);
and U1118 (N_1118,In_1072,In_611);
nor U1119 (N_1119,In_2372,In_820);
nand U1120 (N_1120,In_2177,In_2593);
nor U1121 (N_1121,In_215,In_2643);
xor U1122 (N_1122,In_1627,In_327);
or U1123 (N_1123,In_13,In_1808);
xnor U1124 (N_1124,In_1430,In_656);
or U1125 (N_1125,In_1834,In_2841);
xor U1126 (N_1126,In_1340,In_62);
nor U1127 (N_1127,In_40,In_1113);
xnor U1128 (N_1128,In_108,In_468);
and U1129 (N_1129,In_1769,In_1917);
or U1130 (N_1130,In_1148,In_2214);
nor U1131 (N_1131,In_2665,In_2271);
or U1132 (N_1132,In_2830,In_1302);
nand U1133 (N_1133,In_973,In_1968);
xor U1134 (N_1134,In_591,In_2939);
nor U1135 (N_1135,In_1307,In_752);
and U1136 (N_1136,In_2865,In_2938);
and U1137 (N_1137,In_63,In_1061);
nand U1138 (N_1138,In_2009,In_511);
or U1139 (N_1139,In_2399,In_170);
nor U1140 (N_1140,In_2738,In_2532);
xor U1141 (N_1141,In_1611,In_538);
or U1142 (N_1142,In_488,In_2292);
xor U1143 (N_1143,In_1157,In_2801);
nor U1144 (N_1144,In_2916,In_1421);
nor U1145 (N_1145,In_893,In_657);
nand U1146 (N_1146,In_1286,In_1514);
nor U1147 (N_1147,In_608,In_2943);
xnor U1148 (N_1148,In_549,In_2396);
and U1149 (N_1149,In_1868,In_2628);
or U1150 (N_1150,In_2652,In_1916);
nand U1151 (N_1151,In_857,In_946);
and U1152 (N_1152,In_2008,In_1313);
and U1153 (N_1153,In_926,In_1192);
and U1154 (N_1154,In_1426,In_2880);
xnor U1155 (N_1155,In_1696,In_1127);
nand U1156 (N_1156,In_802,In_1031);
or U1157 (N_1157,In_450,In_2423);
nand U1158 (N_1158,In_651,In_500);
nand U1159 (N_1159,In_1379,In_672);
and U1160 (N_1160,In_2164,In_351);
nor U1161 (N_1161,In_1869,In_1142);
or U1162 (N_1162,In_509,In_1416);
and U1163 (N_1163,In_423,In_631);
nor U1164 (N_1164,In_777,In_2141);
xnor U1165 (N_1165,In_2521,In_649);
and U1166 (N_1166,In_2601,In_1854);
xnor U1167 (N_1167,In_1863,In_1119);
and U1168 (N_1168,In_2807,In_601);
nand U1169 (N_1169,In_1200,In_214);
nand U1170 (N_1170,In_1401,In_328);
nand U1171 (N_1171,In_2489,In_725);
nand U1172 (N_1172,In_2592,In_1210);
xor U1173 (N_1173,In_499,In_2024);
or U1174 (N_1174,In_1432,In_1053);
and U1175 (N_1175,In_107,In_1183);
and U1176 (N_1176,In_1052,In_147);
nand U1177 (N_1177,In_2561,In_2341);
xnor U1178 (N_1178,In_2718,In_1842);
and U1179 (N_1179,In_90,In_1693);
or U1180 (N_1180,In_575,In_2378);
nor U1181 (N_1181,In_473,In_1384);
or U1182 (N_1182,In_2677,In_1492);
nor U1183 (N_1183,In_2682,In_1393);
or U1184 (N_1184,In_533,In_827);
nand U1185 (N_1185,In_388,In_1943);
and U1186 (N_1186,In_1478,In_633);
and U1187 (N_1187,In_523,In_2284);
nand U1188 (N_1188,In_1561,In_113);
xnor U1189 (N_1189,In_1428,In_1357);
and U1190 (N_1190,In_492,In_970);
and U1191 (N_1191,In_206,In_1516);
xnor U1192 (N_1192,In_205,In_130);
nor U1193 (N_1193,In_1038,In_2296);
xor U1194 (N_1194,In_1021,In_835);
nand U1195 (N_1195,In_339,In_1982);
and U1196 (N_1196,In_993,In_2467);
or U1197 (N_1197,In_1389,In_859);
xnor U1198 (N_1198,In_225,In_2501);
nor U1199 (N_1199,In_191,In_712);
xnor U1200 (N_1200,In_527,In_2845);
nand U1201 (N_1201,In_731,In_2711);
nor U1202 (N_1202,In_2262,In_179);
or U1203 (N_1203,In_2780,In_2770);
or U1204 (N_1204,In_2145,In_965);
xnor U1205 (N_1205,In_555,In_617);
nand U1206 (N_1206,In_1753,In_1347);
nor U1207 (N_1207,In_1559,In_1442);
or U1208 (N_1208,In_1925,In_2693);
and U1209 (N_1209,In_2016,In_212);
xor U1210 (N_1210,In_1216,In_1551);
nor U1211 (N_1211,In_1986,In_299);
nand U1212 (N_1212,In_2556,In_1997);
xor U1213 (N_1213,In_283,In_337);
nand U1214 (N_1214,In_470,In_2092);
nand U1215 (N_1215,In_1206,In_2171);
and U1216 (N_1216,In_1767,In_681);
or U1217 (N_1217,In_2779,In_2760);
xnor U1218 (N_1218,In_2453,In_382);
nor U1219 (N_1219,In_768,In_2775);
nand U1220 (N_1220,In_496,In_266);
nand U1221 (N_1221,In_957,In_2162);
xor U1222 (N_1222,In_2541,In_623);
and U1223 (N_1223,In_2902,In_1805);
and U1224 (N_1224,In_2120,In_2849);
xnor U1225 (N_1225,In_2897,In_562);
and U1226 (N_1226,In_954,In_2844);
and U1227 (N_1227,In_1439,In_697);
or U1228 (N_1228,In_2155,In_2668);
nor U1229 (N_1229,In_945,In_2265);
and U1230 (N_1230,In_2455,In_1448);
or U1231 (N_1231,In_1570,In_2099);
and U1232 (N_1232,In_1643,In_1408);
and U1233 (N_1233,In_1791,In_2671);
xor U1234 (N_1234,In_1109,In_2110);
or U1235 (N_1235,In_1166,In_1858);
or U1236 (N_1236,In_422,In_1000);
xnor U1237 (N_1237,In_2073,In_1498);
or U1238 (N_1238,In_2774,In_1879);
nand U1239 (N_1239,In_610,In_1117);
and U1240 (N_1240,In_765,In_1074);
nor U1241 (N_1241,In_1217,In_2699);
or U1242 (N_1242,In_2788,In_978);
nor U1243 (N_1243,In_2985,In_1125);
or U1244 (N_1244,In_2512,In_2789);
or U1245 (N_1245,In_1055,In_1283);
and U1246 (N_1246,In_2454,In_445);
or U1247 (N_1247,In_668,In_1623);
nand U1248 (N_1248,In_2257,In_2755);
nand U1249 (N_1249,In_1375,In_1640);
nand U1250 (N_1250,In_2782,In_2046);
nand U1251 (N_1251,In_65,In_2529);
nor U1252 (N_1252,In_2,In_124);
nor U1253 (N_1253,In_1258,In_2422);
nor U1254 (N_1254,In_1898,In_793);
nor U1255 (N_1255,In_1202,In_2689);
nor U1256 (N_1256,In_2400,In_2641);
or U1257 (N_1257,In_2771,In_1459);
and U1258 (N_1258,In_2912,In_2107);
or U1259 (N_1259,In_1314,In_934);
nand U1260 (N_1260,In_796,In_927);
or U1261 (N_1261,In_97,In_2564);
or U1262 (N_1262,In_1714,In_1554);
xor U1263 (N_1263,In_1581,In_2640);
and U1264 (N_1264,In_2087,In_2301);
nor U1265 (N_1265,In_310,In_178);
nand U1266 (N_1266,In_2756,In_1);
or U1267 (N_1267,In_2084,In_1644);
or U1268 (N_1268,In_612,In_375);
or U1269 (N_1269,In_2860,In_2753);
and U1270 (N_1270,In_2679,In_1542);
nand U1271 (N_1271,In_2821,In_2549);
or U1272 (N_1272,In_2442,In_2635);
or U1273 (N_1273,In_1129,In_330);
xor U1274 (N_1274,In_1433,In_1111);
and U1275 (N_1275,In_2230,In_2763);
nand U1276 (N_1276,In_1495,In_1874);
or U1277 (N_1277,In_1339,In_2583);
and U1278 (N_1278,In_456,In_1543);
nand U1279 (N_1279,In_1449,In_2555);
nand U1280 (N_1280,In_1547,In_2291);
nand U1281 (N_1281,In_146,In_545);
nand U1282 (N_1282,In_370,In_407);
nand U1283 (N_1283,In_637,In_2011);
and U1284 (N_1284,In_230,In_232);
or U1285 (N_1285,In_1501,In_580);
and U1286 (N_1286,In_1160,In_1739);
xor U1287 (N_1287,In_30,In_647);
or U1288 (N_1288,In_26,In_1540);
or U1289 (N_1289,In_2287,In_2390);
nand U1290 (N_1290,In_1589,In_2806);
and U1291 (N_1291,In_2431,In_546);
nor U1292 (N_1292,In_1247,In_425);
nor U1293 (N_1293,In_568,In_2858);
or U1294 (N_1294,In_1963,In_1860);
nand U1295 (N_1295,In_2572,In_1945);
and U1296 (N_1296,In_1010,In_192);
nor U1297 (N_1297,In_1579,In_2787);
nand U1298 (N_1298,In_1624,In_2411);
or U1299 (N_1299,In_2563,In_1752);
or U1300 (N_1300,In_144,In_2136);
and U1301 (N_1301,In_1958,In_2676);
xor U1302 (N_1302,In_968,In_1250);
or U1303 (N_1303,In_1100,In_2280);
nor U1304 (N_1304,In_1163,In_1447);
nor U1305 (N_1305,In_599,In_916);
xor U1306 (N_1306,In_2795,In_2957);
and U1307 (N_1307,In_1446,In_2919);
or U1308 (N_1308,In_870,In_2522);
or U1309 (N_1309,In_2544,In_1790);
and U1310 (N_1310,In_1415,In_508);
xor U1311 (N_1311,In_1821,In_91);
or U1312 (N_1312,In_745,In_2877);
nand U1313 (N_1313,In_38,In_2759);
xor U1314 (N_1314,In_845,In_889);
nor U1315 (N_1315,In_2349,In_2989);
nor U1316 (N_1316,In_2837,In_2469);
and U1317 (N_1317,In_1164,In_958);
and U1318 (N_1318,In_173,In_300);
and U1319 (N_1319,In_289,In_686);
nand U1320 (N_1320,In_2460,In_2318);
and U1321 (N_1321,In_20,In_1204);
or U1322 (N_1322,In_2895,In_1750);
and U1323 (N_1323,In_64,In_2963);
nor U1324 (N_1324,In_5,In_928);
xor U1325 (N_1325,In_1690,In_1861);
xnor U1326 (N_1326,In_1691,In_2494);
xnor U1327 (N_1327,In_2282,In_2288);
nor U1328 (N_1328,In_2816,In_505);
nand U1329 (N_1329,In_1312,In_2077);
or U1330 (N_1330,In_2229,In_988);
nand U1331 (N_1331,In_2531,In_977);
nor U1332 (N_1332,In_1757,In_1269);
nor U1333 (N_1333,In_1273,In_7);
nor U1334 (N_1334,In_1150,In_2255);
or U1335 (N_1335,In_55,In_2735);
and U1336 (N_1336,In_1329,In_1371);
and U1337 (N_1337,In_1889,In_195);
nand U1338 (N_1338,In_8,In_440);
nor U1339 (N_1339,In_22,In_2986);
or U1340 (N_1340,In_447,In_2160);
xnor U1341 (N_1341,In_839,In_907);
and U1342 (N_1342,In_1541,In_510);
or U1343 (N_1343,In_1388,In_1988);
or U1344 (N_1344,In_1664,In_118);
nor U1345 (N_1345,In_1938,In_1030);
or U1346 (N_1346,In_2645,In_2461);
xnor U1347 (N_1347,In_1240,In_1764);
nor U1348 (N_1348,In_1108,In_1029);
and U1349 (N_1349,In_219,In_2580);
xnor U1350 (N_1350,In_2954,In_727);
xnor U1351 (N_1351,In_1174,In_2724);
xnor U1352 (N_1352,In_2367,In_880);
xnor U1353 (N_1353,In_2052,In_2144);
xnor U1354 (N_1354,In_794,In_2047);
or U1355 (N_1355,In_1522,In_2664);
xor U1356 (N_1356,In_1484,In_1040);
and U1357 (N_1357,In_2226,In_1361);
or U1358 (N_1358,In_998,In_1723);
and U1359 (N_1359,In_12,In_675);
xor U1360 (N_1360,In_1747,In_307);
xnor U1361 (N_1361,In_935,In_2915);
and U1362 (N_1362,In_506,In_2998);
or U1363 (N_1363,In_149,In_871);
nor U1364 (N_1364,In_572,In_2216);
nand U1365 (N_1365,In_1665,In_2412);
nor U1366 (N_1366,In_1971,In_2499);
nor U1367 (N_1367,In_2650,In_329);
nand U1368 (N_1368,In_503,In_2290);
xor U1369 (N_1369,In_2474,In_238);
xor U1370 (N_1370,In_1078,In_1974);
or U1371 (N_1371,In_449,In_1476);
nor U1372 (N_1372,In_402,In_2648);
xnor U1373 (N_1373,In_1902,In_461);
nand U1374 (N_1374,In_2726,In_18);
nand U1375 (N_1375,In_1232,In_959);
nor U1376 (N_1376,In_221,In_625);
nor U1377 (N_1377,In_2566,In_183);
nand U1378 (N_1378,In_400,In_919);
or U1379 (N_1379,In_1978,In_1684);
or U1380 (N_1380,In_1461,In_1308);
nand U1381 (N_1381,In_2345,In_1872);
nor U1382 (N_1382,In_2826,In_273);
or U1383 (N_1383,In_2716,In_882);
nand U1384 (N_1384,In_1993,In_1196);
nand U1385 (N_1385,In_2876,In_1941);
and U1386 (N_1386,In_453,In_1349);
nand U1387 (N_1387,In_1782,In_2446);
or U1388 (N_1388,In_1612,In_1755);
nand U1389 (N_1389,In_2433,In_47);
and U1390 (N_1390,In_1610,In_854);
and U1391 (N_1391,In_2516,In_2019);
nor U1392 (N_1392,In_1524,In_2619);
or U1393 (N_1393,In_2117,In_867);
xnor U1394 (N_1394,In_1138,In_975);
nand U1395 (N_1395,In_718,In_937);
xor U1396 (N_1396,In_613,In_2176);
and U1397 (N_1397,In_354,In_2887);
or U1398 (N_1398,In_404,In_2053);
nor U1399 (N_1399,In_405,In_1431);
nor U1400 (N_1400,In_1760,In_2031);
nor U1401 (N_1401,In_2546,In_2449);
nand U1402 (N_1402,In_50,In_778);
and U1403 (N_1403,In_387,In_495);
xnor U1404 (N_1404,In_679,In_2995);
nand U1405 (N_1405,In_2364,In_491);
nand U1406 (N_1406,In_1121,In_2039);
and U1407 (N_1407,In_1518,In_1018);
nand U1408 (N_1408,In_338,In_603);
xnor U1409 (N_1409,In_543,In_2625);
nor U1410 (N_1410,In_1434,In_2777);
or U1411 (N_1411,In_2834,In_2239);
and U1412 (N_1412,In_1706,In_1205);
nand U1413 (N_1413,In_2692,In_2191);
nand U1414 (N_1414,In_350,In_95);
nor U1415 (N_1415,In_917,In_1058);
nand U1416 (N_1416,In_1234,In_1562);
nand U1417 (N_1417,In_2498,In_821);
and U1418 (N_1418,In_2574,In_2709);
xor U1419 (N_1419,In_944,In_1330);
xnor U1420 (N_1420,In_2553,In_2030);
or U1421 (N_1421,In_790,In_2518);
xor U1422 (N_1422,In_2626,In_2317);
xor U1423 (N_1423,In_2847,In_804);
nand U1424 (N_1424,In_478,In_457);
nand U1425 (N_1425,In_2594,In_2129);
and U1426 (N_1426,In_359,In_2080);
and U1427 (N_1427,In_1444,In_525);
nor U1428 (N_1428,In_366,In_374);
and U1429 (N_1429,In_1087,In_237);
and U1430 (N_1430,In_2951,In_2359);
nor U1431 (N_1431,In_897,In_2127);
or U1432 (N_1432,In_1419,In_1604);
xor U1433 (N_1433,In_717,In_1427);
and U1434 (N_1434,In_1463,In_961);
and U1435 (N_1435,In_1822,In_2945);
nor U1436 (N_1436,In_2903,In_2514);
or U1437 (N_1437,In_265,In_741);
and U1438 (N_1438,In_2602,In_1152);
and U1439 (N_1439,In_1209,In_2095);
nand U1440 (N_1440,In_590,In_895);
nor U1441 (N_1441,In_1368,In_1817);
xor U1442 (N_1442,In_780,In_2949);
and U1443 (N_1443,In_1798,In_795);
and U1444 (N_1444,In_2042,In_1136);
nor U1445 (N_1445,In_1576,In_137);
xor U1446 (N_1446,In_2130,In_42);
nor U1447 (N_1447,In_2027,In_812);
nand U1448 (N_1448,In_1156,In_39);
nor U1449 (N_1449,In_1280,In_180);
or U1450 (N_1450,In_1407,In_1011);
xor U1451 (N_1451,In_535,In_2946);
nand U1452 (N_1452,In_2904,In_2800);
or U1453 (N_1453,In_1392,In_1467);
xnor U1454 (N_1454,In_34,In_2414);
nand U1455 (N_1455,In_2175,In_2888);
xor U1456 (N_1456,In_1048,In_2266);
or U1457 (N_1457,In_462,In_1265);
xor U1458 (N_1458,In_1648,In_116);
nand U1459 (N_1459,In_2797,In_2365);
or U1460 (N_1460,In_1012,In_1104);
nand U1461 (N_1461,In_2670,In_1761);
and U1462 (N_1462,In_949,In_2283);
nor U1463 (N_1463,In_873,In_635);
nand U1464 (N_1464,In_2121,In_2100);
or U1465 (N_1465,In_424,In_911);
nor U1466 (N_1466,In_2855,In_756);
and U1467 (N_1467,In_292,In_1350);
or U1468 (N_1468,In_2072,In_1178);
or U1469 (N_1469,In_2686,In_901);
nor U1470 (N_1470,In_117,In_2967);
and U1471 (N_1471,In_2369,In_1268);
and U1472 (N_1472,In_1490,In_326);
nor U1473 (N_1473,In_2337,In_2950);
xor U1474 (N_1474,In_2427,In_1405);
and U1475 (N_1475,In_1638,In_1921);
and U1476 (N_1476,In_2598,In_1267);
xnor U1477 (N_1477,In_110,In_2587);
nand U1478 (N_1478,In_2932,In_319);
or U1479 (N_1479,In_2044,In_317);
xor U1480 (N_1480,In_1920,In_249);
nor U1481 (N_1481,In_671,In_88);
nand U1482 (N_1482,In_849,In_418);
xor U1483 (N_1483,In_228,In_1733);
nand U1484 (N_1484,In_52,In_1599);
or U1485 (N_1485,In_1742,In_1615);
nor U1486 (N_1486,In_1420,In_309);
nand U1487 (N_1487,In_2513,In_2965);
xnor U1488 (N_1488,In_1826,In_2552);
and U1489 (N_1489,In_2818,In_2918);
or U1490 (N_1490,In_669,In_2434);
xnor U1491 (N_1491,In_530,In_1355);
xor U1492 (N_1492,In_1198,In_1851);
nor U1493 (N_1493,In_1252,In_1281);
nor U1494 (N_1494,In_325,In_2545);
and U1495 (N_1495,In_126,In_2401);
or U1496 (N_1496,In_2331,In_1332);
nor U1497 (N_1497,In_2254,In_1409);
nand U1498 (N_1498,In_2940,In_189);
nand U1499 (N_1499,In_44,In_579);
nand U1500 (N_1500,In_1262,In_786);
nand U1501 (N_1501,In_953,In_548);
nor U1502 (N_1502,In_994,In_2267);
and U1503 (N_1503,In_2226,In_1349);
or U1504 (N_1504,In_2968,In_1579);
xnor U1505 (N_1505,In_1562,In_1838);
or U1506 (N_1506,In_347,In_2927);
or U1507 (N_1507,In_1819,In_355);
and U1508 (N_1508,In_2013,In_581);
or U1509 (N_1509,In_1529,In_1300);
nand U1510 (N_1510,In_672,In_895);
xnor U1511 (N_1511,In_1392,In_5);
or U1512 (N_1512,In_1541,In_1625);
and U1513 (N_1513,In_2326,In_395);
nand U1514 (N_1514,In_2875,In_1655);
nor U1515 (N_1515,In_1620,In_1035);
or U1516 (N_1516,In_870,In_1385);
xor U1517 (N_1517,In_2168,In_850);
or U1518 (N_1518,In_2010,In_55);
xor U1519 (N_1519,In_746,In_1176);
nor U1520 (N_1520,In_951,In_590);
nor U1521 (N_1521,In_2775,In_230);
xnor U1522 (N_1522,In_972,In_2181);
and U1523 (N_1523,In_2136,In_2318);
or U1524 (N_1524,In_2683,In_123);
nor U1525 (N_1525,In_1851,In_2438);
and U1526 (N_1526,In_2478,In_1089);
xnor U1527 (N_1527,In_1848,In_421);
xnor U1528 (N_1528,In_895,In_600);
xor U1529 (N_1529,In_1680,In_1537);
or U1530 (N_1530,In_153,In_2592);
nor U1531 (N_1531,In_2284,In_526);
nand U1532 (N_1532,In_41,In_1941);
nand U1533 (N_1533,In_544,In_2953);
nor U1534 (N_1534,In_781,In_673);
nand U1535 (N_1535,In_1443,In_2019);
and U1536 (N_1536,In_809,In_1758);
nor U1537 (N_1537,In_1849,In_2339);
and U1538 (N_1538,In_2252,In_934);
or U1539 (N_1539,In_1421,In_1803);
nand U1540 (N_1540,In_99,In_1518);
xnor U1541 (N_1541,In_2698,In_1479);
or U1542 (N_1542,In_1010,In_181);
nand U1543 (N_1543,In_1149,In_368);
nand U1544 (N_1544,In_2481,In_104);
and U1545 (N_1545,In_2321,In_359);
xor U1546 (N_1546,In_2922,In_869);
or U1547 (N_1547,In_2434,In_1571);
nor U1548 (N_1548,In_1276,In_84);
nor U1549 (N_1549,In_1465,In_1989);
xnor U1550 (N_1550,In_758,In_2458);
xor U1551 (N_1551,In_2103,In_2248);
and U1552 (N_1552,In_1201,In_771);
nor U1553 (N_1553,In_1751,In_721);
nor U1554 (N_1554,In_2044,In_1043);
nor U1555 (N_1555,In_2794,In_1832);
and U1556 (N_1556,In_298,In_2758);
and U1557 (N_1557,In_2597,In_1979);
nand U1558 (N_1558,In_1720,In_1234);
or U1559 (N_1559,In_701,In_223);
and U1560 (N_1560,In_2254,In_2771);
xnor U1561 (N_1561,In_1080,In_2393);
nand U1562 (N_1562,In_136,In_1787);
xor U1563 (N_1563,In_2012,In_802);
nor U1564 (N_1564,In_67,In_295);
nand U1565 (N_1565,In_1937,In_2531);
xor U1566 (N_1566,In_382,In_1704);
xor U1567 (N_1567,In_1651,In_2477);
xnor U1568 (N_1568,In_1102,In_2400);
nor U1569 (N_1569,In_240,In_372);
and U1570 (N_1570,In_2847,In_811);
and U1571 (N_1571,In_1541,In_1803);
xor U1572 (N_1572,In_404,In_2450);
nand U1573 (N_1573,In_1162,In_662);
and U1574 (N_1574,In_1963,In_1659);
or U1575 (N_1575,In_92,In_1589);
nor U1576 (N_1576,In_2021,In_2116);
xor U1577 (N_1577,In_179,In_1168);
nand U1578 (N_1578,In_1497,In_295);
and U1579 (N_1579,In_472,In_1325);
nor U1580 (N_1580,In_2606,In_1058);
and U1581 (N_1581,In_2779,In_1254);
and U1582 (N_1582,In_455,In_2600);
nand U1583 (N_1583,In_2068,In_2448);
nor U1584 (N_1584,In_2710,In_1058);
nand U1585 (N_1585,In_1719,In_878);
nand U1586 (N_1586,In_1100,In_29);
xor U1587 (N_1587,In_2083,In_1599);
nand U1588 (N_1588,In_2570,In_2758);
nand U1589 (N_1589,In_2134,In_2720);
nor U1590 (N_1590,In_2525,In_370);
xnor U1591 (N_1591,In_1884,In_2308);
and U1592 (N_1592,In_2272,In_848);
or U1593 (N_1593,In_1013,In_1586);
nand U1594 (N_1594,In_147,In_2789);
or U1595 (N_1595,In_1329,In_18);
or U1596 (N_1596,In_1551,In_2306);
nand U1597 (N_1597,In_1062,In_727);
xor U1598 (N_1598,In_2309,In_641);
or U1599 (N_1599,In_2302,In_2057);
nand U1600 (N_1600,In_661,In_159);
xnor U1601 (N_1601,In_2626,In_676);
and U1602 (N_1602,In_2292,In_2367);
nand U1603 (N_1603,In_666,In_2598);
and U1604 (N_1604,In_2632,In_864);
nand U1605 (N_1605,In_399,In_1940);
and U1606 (N_1606,In_10,In_1550);
nor U1607 (N_1607,In_2346,In_2626);
nand U1608 (N_1608,In_1484,In_1257);
xor U1609 (N_1609,In_1015,In_1038);
nand U1610 (N_1610,In_2159,In_1558);
xnor U1611 (N_1611,In_743,In_573);
nand U1612 (N_1612,In_245,In_698);
and U1613 (N_1613,In_658,In_2710);
xor U1614 (N_1614,In_2391,In_1691);
nand U1615 (N_1615,In_196,In_2762);
or U1616 (N_1616,In_1059,In_58);
or U1617 (N_1617,In_2272,In_448);
or U1618 (N_1618,In_727,In_604);
or U1619 (N_1619,In_1337,In_949);
nor U1620 (N_1620,In_679,In_2587);
nand U1621 (N_1621,In_67,In_958);
nand U1622 (N_1622,In_2643,In_31);
or U1623 (N_1623,In_111,In_1929);
nor U1624 (N_1624,In_891,In_272);
nand U1625 (N_1625,In_2334,In_2781);
nor U1626 (N_1626,In_989,In_2261);
xnor U1627 (N_1627,In_2570,In_769);
nor U1628 (N_1628,In_793,In_2207);
or U1629 (N_1629,In_1137,In_2013);
xor U1630 (N_1630,In_1155,In_787);
and U1631 (N_1631,In_1484,In_781);
nor U1632 (N_1632,In_430,In_1574);
nand U1633 (N_1633,In_1566,In_312);
nand U1634 (N_1634,In_1986,In_2844);
nand U1635 (N_1635,In_1301,In_1916);
nor U1636 (N_1636,In_1045,In_1696);
and U1637 (N_1637,In_2702,In_1750);
xnor U1638 (N_1638,In_2120,In_100);
and U1639 (N_1639,In_1034,In_2805);
or U1640 (N_1640,In_1170,In_731);
nand U1641 (N_1641,In_803,In_2994);
or U1642 (N_1642,In_770,In_344);
xor U1643 (N_1643,In_1489,In_1981);
and U1644 (N_1644,In_2085,In_923);
nand U1645 (N_1645,In_1202,In_787);
and U1646 (N_1646,In_1822,In_2674);
and U1647 (N_1647,In_537,In_180);
nand U1648 (N_1648,In_1357,In_2501);
xnor U1649 (N_1649,In_2036,In_695);
or U1650 (N_1650,In_42,In_2309);
and U1651 (N_1651,In_1948,In_2423);
nor U1652 (N_1652,In_367,In_2950);
nor U1653 (N_1653,In_727,In_1415);
xor U1654 (N_1654,In_828,In_1545);
nand U1655 (N_1655,In_2677,In_2934);
or U1656 (N_1656,In_798,In_2546);
nor U1657 (N_1657,In_988,In_1090);
or U1658 (N_1658,In_484,In_2201);
and U1659 (N_1659,In_1835,In_420);
nor U1660 (N_1660,In_696,In_2161);
and U1661 (N_1661,In_446,In_496);
nand U1662 (N_1662,In_1993,In_1661);
nor U1663 (N_1663,In_393,In_1302);
and U1664 (N_1664,In_1921,In_1474);
nand U1665 (N_1665,In_2365,In_2417);
nor U1666 (N_1666,In_2354,In_2478);
nand U1667 (N_1667,In_2521,In_2227);
or U1668 (N_1668,In_1770,In_2101);
nand U1669 (N_1669,In_2838,In_692);
nand U1670 (N_1670,In_2693,In_2051);
nand U1671 (N_1671,In_2752,In_867);
nand U1672 (N_1672,In_2669,In_1832);
xnor U1673 (N_1673,In_1631,In_1632);
and U1674 (N_1674,In_659,In_1018);
xnor U1675 (N_1675,In_2139,In_1890);
and U1676 (N_1676,In_148,In_744);
nor U1677 (N_1677,In_2302,In_1128);
and U1678 (N_1678,In_1364,In_1284);
or U1679 (N_1679,In_2955,In_191);
xor U1680 (N_1680,In_1403,In_2947);
or U1681 (N_1681,In_2651,In_394);
nand U1682 (N_1682,In_1257,In_820);
nand U1683 (N_1683,In_2058,In_2326);
nor U1684 (N_1684,In_1933,In_213);
xor U1685 (N_1685,In_578,In_297);
nor U1686 (N_1686,In_671,In_2115);
nor U1687 (N_1687,In_1524,In_2204);
or U1688 (N_1688,In_772,In_2193);
and U1689 (N_1689,In_811,In_1460);
and U1690 (N_1690,In_1709,In_1716);
and U1691 (N_1691,In_1240,In_222);
nor U1692 (N_1692,In_2614,In_2493);
and U1693 (N_1693,In_1130,In_590);
xnor U1694 (N_1694,In_850,In_1358);
and U1695 (N_1695,In_1161,In_2248);
nand U1696 (N_1696,In_984,In_1062);
nand U1697 (N_1697,In_1177,In_1332);
nand U1698 (N_1698,In_2330,In_2999);
xor U1699 (N_1699,In_2305,In_2595);
and U1700 (N_1700,In_1596,In_183);
nand U1701 (N_1701,In_261,In_1073);
nand U1702 (N_1702,In_1838,In_1313);
xnor U1703 (N_1703,In_2557,In_723);
and U1704 (N_1704,In_59,In_1094);
nor U1705 (N_1705,In_375,In_2107);
nand U1706 (N_1706,In_2281,In_2726);
nand U1707 (N_1707,In_2747,In_2783);
xnor U1708 (N_1708,In_1175,In_1051);
or U1709 (N_1709,In_979,In_2202);
nand U1710 (N_1710,In_2122,In_1942);
xor U1711 (N_1711,In_463,In_40);
and U1712 (N_1712,In_1175,In_2568);
and U1713 (N_1713,In_266,In_1625);
and U1714 (N_1714,In_1071,In_1979);
xor U1715 (N_1715,In_23,In_2896);
nor U1716 (N_1716,In_1866,In_2641);
nand U1717 (N_1717,In_48,In_2578);
and U1718 (N_1718,In_2145,In_1865);
nor U1719 (N_1719,In_792,In_1871);
xor U1720 (N_1720,In_1103,In_683);
or U1721 (N_1721,In_2498,In_681);
and U1722 (N_1722,In_1999,In_642);
xnor U1723 (N_1723,In_2929,In_705);
nand U1724 (N_1724,In_1425,In_2705);
xnor U1725 (N_1725,In_1352,In_1307);
nand U1726 (N_1726,In_1472,In_257);
or U1727 (N_1727,In_2868,In_2788);
and U1728 (N_1728,In_184,In_2950);
nor U1729 (N_1729,In_513,In_2608);
and U1730 (N_1730,In_452,In_1451);
nor U1731 (N_1731,In_2193,In_2553);
or U1732 (N_1732,In_799,In_2046);
nor U1733 (N_1733,In_1085,In_1221);
nand U1734 (N_1734,In_2081,In_1518);
nor U1735 (N_1735,In_148,In_2598);
nand U1736 (N_1736,In_1492,In_1383);
xor U1737 (N_1737,In_465,In_1851);
xor U1738 (N_1738,In_255,In_150);
or U1739 (N_1739,In_1444,In_2870);
or U1740 (N_1740,In_611,In_1649);
nand U1741 (N_1741,In_2087,In_2985);
nor U1742 (N_1742,In_2470,In_2883);
xor U1743 (N_1743,In_175,In_2099);
nor U1744 (N_1744,In_634,In_819);
and U1745 (N_1745,In_540,In_1204);
nand U1746 (N_1746,In_1637,In_352);
or U1747 (N_1747,In_1607,In_1115);
nand U1748 (N_1748,In_451,In_734);
and U1749 (N_1749,In_693,In_1057);
nand U1750 (N_1750,In_1791,In_1047);
nand U1751 (N_1751,In_2825,In_2195);
nor U1752 (N_1752,In_1793,In_436);
nand U1753 (N_1753,In_237,In_828);
or U1754 (N_1754,In_2545,In_118);
nor U1755 (N_1755,In_1195,In_2855);
or U1756 (N_1756,In_368,In_126);
or U1757 (N_1757,In_2095,In_2109);
or U1758 (N_1758,In_1843,In_2858);
or U1759 (N_1759,In_2415,In_751);
xor U1760 (N_1760,In_635,In_2615);
nor U1761 (N_1761,In_808,In_458);
and U1762 (N_1762,In_2985,In_1176);
nor U1763 (N_1763,In_1609,In_2587);
nand U1764 (N_1764,In_1808,In_193);
xor U1765 (N_1765,In_1673,In_2431);
or U1766 (N_1766,In_2431,In_2253);
nand U1767 (N_1767,In_1087,In_949);
xnor U1768 (N_1768,In_2933,In_1855);
and U1769 (N_1769,In_459,In_465);
xnor U1770 (N_1770,In_1941,In_780);
xnor U1771 (N_1771,In_191,In_1582);
nor U1772 (N_1772,In_2033,In_482);
and U1773 (N_1773,In_2482,In_240);
nor U1774 (N_1774,In_2358,In_0);
xor U1775 (N_1775,In_530,In_1958);
xor U1776 (N_1776,In_978,In_2696);
or U1777 (N_1777,In_2986,In_1434);
nand U1778 (N_1778,In_2139,In_2246);
or U1779 (N_1779,In_2114,In_2770);
nor U1780 (N_1780,In_2072,In_1172);
xor U1781 (N_1781,In_2023,In_2003);
nor U1782 (N_1782,In_1869,In_78);
nor U1783 (N_1783,In_2600,In_1032);
and U1784 (N_1784,In_1695,In_2993);
or U1785 (N_1785,In_1535,In_2179);
or U1786 (N_1786,In_1080,In_2154);
and U1787 (N_1787,In_2150,In_1240);
nor U1788 (N_1788,In_2949,In_1360);
nand U1789 (N_1789,In_732,In_2163);
and U1790 (N_1790,In_272,In_829);
or U1791 (N_1791,In_1272,In_1945);
and U1792 (N_1792,In_513,In_2534);
nand U1793 (N_1793,In_1306,In_2621);
nand U1794 (N_1794,In_865,In_1140);
xnor U1795 (N_1795,In_2057,In_698);
nor U1796 (N_1796,In_660,In_1003);
xnor U1797 (N_1797,In_2260,In_2721);
or U1798 (N_1798,In_2396,In_2722);
nand U1799 (N_1799,In_1803,In_82);
nor U1800 (N_1800,In_2173,In_1896);
nor U1801 (N_1801,In_2991,In_2775);
nand U1802 (N_1802,In_1021,In_1132);
xor U1803 (N_1803,In_2821,In_420);
and U1804 (N_1804,In_543,In_987);
xnor U1805 (N_1805,In_2026,In_884);
or U1806 (N_1806,In_1510,In_122);
xnor U1807 (N_1807,In_103,In_2354);
and U1808 (N_1808,In_1177,In_548);
nor U1809 (N_1809,In_343,In_379);
nand U1810 (N_1810,In_151,In_2271);
and U1811 (N_1811,In_2281,In_379);
or U1812 (N_1812,In_1906,In_2824);
nor U1813 (N_1813,In_2643,In_867);
and U1814 (N_1814,In_602,In_1339);
or U1815 (N_1815,In_889,In_2651);
or U1816 (N_1816,In_1048,In_2054);
and U1817 (N_1817,In_39,In_1149);
nor U1818 (N_1818,In_1695,In_1564);
and U1819 (N_1819,In_2893,In_2722);
nor U1820 (N_1820,In_310,In_317);
xor U1821 (N_1821,In_512,In_472);
nor U1822 (N_1822,In_2149,In_1520);
and U1823 (N_1823,In_1167,In_2951);
or U1824 (N_1824,In_1688,In_1594);
nor U1825 (N_1825,In_1143,In_18);
and U1826 (N_1826,In_2317,In_1592);
nand U1827 (N_1827,In_2526,In_10);
or U1828 (N_1828,In_125,In_1785);
or U1829 (N_1829,In_1882,In_358);
or U1830 (N_1830,In_1123,In_2303);
nand U1831 (N_1831,In_1201,In_1011);
xnor U1832 (N_1832,In_598,In_1935);
or U1833 (N_1833,In_1158,In_1540);
xor U1834 (N_1834,In_2337,In_2684);
nand U1835 (N_1835,In_1806,In_2225);
xor U1836 (N_1836,In_1510,In_872);
or U1837 (N_1837,In_2278,In_1476);
xnor U1838 (N_1838,In_2826,In_1572);
or U1839 (N_1839,In_1872,In_924);
nand U1840 (N_1840,In_324,In_1686);
or U1841 (N_1841,In_83,In_1930);
nand U1842 (N_1842,In_389,In_1289);
nand U1843 (N_1843,In_1712,In_477);
xor U1844 (N_1844,In_2156,In_1640);
or U1845 (N_1845,In_2932,In_824);
and U1846 (N_1846,In_419,In_2500);
nand U1847 (N_1847,In_2379,In_1592);
nor U1848 (N_1848,In_366,In_637);
and U1849 (N_1849,In_2128,In_1938);
nor U1850 (N_1850,In_611,In_1464);
xor U1851 (N_1851,In_2921,In_989);
nor U1852 (N_1852,In_832,In_873);
or U1853 (N_1853,In_1930,In_2892);
or U1854 (N_1854,In_320,In_67);
xnor U1855 (N_1855,In_1648,In_2134);
nand U1856 (N_1856,In_1929,In_1202);
and U1857 (N_1857,In_258,In_302);
and U1858 (N_1858,In_1050,In_853);
nor U1859 (N_1859,In_942,In_1202);
nor U1860 (N_1860,In_2268,In_2869);
nor U1861 (N_1861,In_127,In_860);
nand U1862 (N_1862,In_457,In_1606);
and U1863 (N_1863,In_1716,In_2793);
or U1864 (N_1864,In_1009,In_2288);
xnor U1865 (N_1865,In_2613,In_945);
nand U1866 (N_1866,In_1453,In_1661);
or U1867 (N_1867,In_2764,In_1108);
or U1868 (N_1868,In_892,In_2220);
xor U1869 (N_1869,In_2496,In_1597);
nor U1870 (N_1870,In_1155,In_1442);
nor U1871 (N_1871,In_2839,In_1100);
and U1872 (N_1872,In_1693,In_1069);
or U1873 (N_1873,In_2241,In_681);
nand U1874 (N_1874,In_2736,In_1229);
xnor U1875 (N_1875,In_1080,In_1743);
xnor U1876 (N_1876,In_2056,In_836);
nand U1877 (N_1877,In_1301,In_1018);
or U1878 (N_1878,In_2096,In_1770);
nor U1879 (N_1879,In_578,In_69);
xnor U1880 (N_1880,In_2392,In_2826);
and U1881 (N_1881,In_871,In_302);
xnor U1882 (N_1882,In_2934,In_1973);
nand U1883 (N_1883,In_349,In_449);
xor U1884 (N_1884,In_1755,In_1894);
xor U1885 (N_1885,In_2584,In_909);
nor U1886 (N_1886,In_2662,In_1114);
and U1887 (N_1887,In_2459,In_2263);
or U1888 (N_1888,In_192,In_1298);
nor U1889 (N_1889,In_1810,In_1516);
nand U1890 (N_1890,In_1426,In_2293);
or U1891 (N_1891,In_894,In_632);
nand U1892 (N_1892,In_1479,In_2890);
xnor U1893 (N_1893,In_1148,In_2658);
or U1894 (N_1894,In_2384,In_1675);
or U1895 (N_1895,In_1726,In_79);
nor U1896 (N_1896,In_79,In_1437);
nor U1897 (N_1897,In_2227,In_2437);
nand U1898 (N_1898,In_2318,In_2661);
nand U1899 (N_1899,In_2986,In_1842);
nor U1900 (N_1900,In_1230,In_1642);
xnor U1901 (N_1901,In_150,In_1786);
or U1902 (N_1902,In_2644,In_119);
nor U1903 (N_1903,In_2637,In_537);
nand U1904 (N_1904,In_2925,In_2552);
xnor U1905 (N_1905,In_2340,In_575);
and U1906 (N_1906,In_1699,In_489);
or U1907 (N_1907,In_1297,In_27);
xnor U1908 (N_1908,In_1894,In_2628);
nor U1909 (N_1909,In_844,In_626);
xor U1910 (N_1910,In_1323,In_2771);
nand U1911 (N_1911,In_40,In_564);
or U1912 (N_1912,In_2469,In_2175);
nor U1913 (N_1913,In_1318,In_2938);
and U1914 (N_1914,In_223,In_2205);
and U1915 (N_1915,In_2345,In_1476);
xnor U1916 (N_1916,In_447,In_1803);
nor U1917 (N_1917,In_195,In_75);
and U1918 (N_1918,In_51,In_1603);
nor U1919 (N_1919,In_124,In_2347);
nor U1920 (N_1920,In_1590,In_466);
and U1921 (N_1921,In_1818,In_891);
nor U1922 (N_1922,In_459,In_1234);
nand U1923 (N_1923,In_1308,In_2081);
xnor U1924 (N_1924,In_148,In_189);
nor U1925 (N_1925,In_1781,In_1185);
nor U1926 (N_1926,In_1579,In_2811);
nor U1927 (N_1927,In_2151,In_370);
or U1928 (N_1928,In_2518,In_105);
nand U1929 (N_1929,In_2075,In_197);
xor U1930 (N_1930,In_962,In_289);
nor U1931 (N_1931,In_2414,In_129);
nor U1932 (N_1932,In_1186,In_372);
or U1933 (N_1933,In_1017,In_1242);
nor U1934 (N_1934,In_1280,In_1203);
nand U1935 (N_1935,In_450,In_1569);
nand U1936 (N_1936,In_1807,In_1757);
nor U1937 (N_1937,In_129,In_2250);
xnor U1938 (N_1938,In_1264,In_730);
nor U1939 (N_1939,In_2857,In_13);
nand U1940 (N_1940,In_1638,In_1900);
nand U1941 (N_1941,In_2026,In_2979);
nand U1942 (N_1942,In_344,In_2741);
nor U1943 (N_1943,In_671,In_1912);
xor U1944 (N_1944,In_1205,In_1420);
nor U1945 (N_1945,In_2660,In_1632);
xor U1946 (N_1946,In_936,In_165);
xnor U1947 (N_1947,In_2512,In_1520);
and U1948 (N_1948,In_310,In_2000);
nand U1949 (N_1949,In_1923,In_2656);
or U1950 (N_1950,In_2739,In_1749);
nand U1951 (N_1951,In_2509,In_1485);
nor U1952 (N_1952,In_1754,In_1987);
xnor U1953 (N_1953,In_1980,In_2869);
nor U1954 (N_1954,In_2957,In_2696);
nor U1955 (N_1955,In_2465,In_2423);
nand U1956 (N_1956,In_1493,In_1565);
nand U1957 (N_1957,In_2845,In_882);
or U1958 (N_1958,In_2510,In_2172);
nand U1959 (N_1959,In_501,In_2592);
or U1960 (N_1960,In_1409,In_2891);
nand U1961 (N_1961,In_2904,In_1658);
xor U1962 (N_1962,In_315,In_2688);
xor U1963 (N_1963,In_2226,In_2518);
nor U1964 (N_1964,In_962,In_2567);
nor U1965 (N_1965,In_2973,In_1877);
xnor U1966 (N_1966,In_1758,In_602);
nor U1967 (N_1967,In_2601,In_204);
and U1968 (N_1968,In_241,In_1271);
and U1969 (N_1969,In_1589,In_2760);
xnor U1970 (N_1970,In_532,In_331);
xnor U1971 (N_1971,In_2184,In_1557);
or U1972 (N_1972,In_2293,In_2861);
or U1973 (N_1973,In_1913,In_1396);
nor U1974 (N_1974,In_2158,In_1409);
and U1975 (N_1975,In_27,In_1363);
and U1976 (N_1976,In_2610,In_2322);
nand U1977 (N_1977,In_1976,In_1429);
or U1978 (N_1978,In_1008,In_899);
nor U1979 (N_1979,In_887,In_779);
xor U1980 (N_1980,In_2521,In_2469);
nor U1981 (N_1981,In_1825,In_1789);
xor U1982 (N_1982,In_472,In_1185);
or U1983 (N_1983,In_2575,In_2013);
and U1984 (N_1984,In_2880,In_2770);
or U1985 (N_1985,In_2965,In_524);
nor U1986 (N_1986,In_2424,In_2167);
or U1987 (N_1987,In_1568,In_57);
nand U1988 (N_1988,In_906,In_1555);
xnor U1989 (N_1989,In_992,In_536);
xnor U1990 (N_1990,In_701,In_2319);
xor U1991 (N_1991,In_612,In_709);
or U1992 (N_1992,In_910,In_196);
xor U1993 (N_1993,In_783,In_1044);
nor U1994 (N_1994,In_2542,In_1075);
or U1995 (N_1995,In_116,In_1842);
nand U1996 (N_1996,In_1676,In_1854);
xor U1997 (N_1997,In_712,In_1633);
nand U1998 (N_1998,In_1177,In_2328);
or U1999 (N_1999,In_2510,In_2735);
or U2000 (N_2000,N_1434,N_1543);
nor U2001 (N_2001,N_1343,N_820);
and U2002 (N_2002,N_217,N_1266);
nand U2003 (N_2003,N_1707,N_1998);
or U2004 (N_2004,N_706,N_1411);
or U2005 (N_2005,N_829,N_133);
and U2006 (N_2006,N_1648,N_678);
xnor U2007 (N_2007,N_68,N_1645);
xor U2008 (N_2008,N_1808,N_830);
nand U2009 (N_2009,N_651,N_1689);
nand U2010 (N_2010,N_1461,N_42);
nand U2011 (N_2011,N_1951,N_647);
xnor U2012 (N_2012,N_1812,N_306);
nand U2013 (N_2013,N_350,N_1871);
xor U2014 (N_2014,N_1218,N_1379);
xnor U2015 (N_2015,N_578,N_1238);
nor U2016 (N_2016,N_18,N_744);
nor U2017 (N_2017,N_1100,N_40);
and U2018 (N_2018,N_1356,N_274);
nor U2019 (N_2019,N_463,N_1738);
nand U2020 (N_2020,N_432,N_616);
and U2021 (N_2021,N_1083,N_1595);
nand U2022 (N_2022,N_1625,N_1008);
nand U2023 (N_2023,N_1875,N_1937);
xor U2024 (N_2024,N_1601,N_263);
or U2025 (N_2025,N_1448,N_298);
and U2026 (N_2026,N_1373,N_1332);
nand U2027 (N_2027,N_1465,N_392);
and U2028 (N_2028,N_1604,N_1659);
nand U2029 (N_2029,N_1667,N_60);
xnor U2030 (N_2030,N_703,N_165);
nor U2031 (N_2031,N_1039,N_519);
or U2032 (N_2032,N_1413,N_640);
and U2033 (N_2033,N_560,N_445);
or U2034 (N_2034,N_1598,N_351);
nor U2035 (N_2035,N_1251,N_636);
nand U2036 (N_2036,N_1267,N_811);
nand U2037 (N_2037,N_207,N_176);
nand U2038 (N_2038,N_1541,N_924);
or U2039 (N_2039,N_543,N_135);
xnor U2040 (N_2040,N_880,N_1912);
xor U2041 (N_2041,N_1451,N_368);
nor U2042 (N_2042,N_866,N_443);
or U2043 (N_2043,N_1273,N_849);
nor U2044 (N_2044,N_91,N_813);
or U2045 (N_2045,N_1499,N_708);
xor U2046 (N_2046,N_684,N_249);
xor U2047 (N_2047,N_889,N_1695);
nand U2048 (N_2048,N_279,N_272);
nand U2049 (N_2049,N_1114,N_1048);
and U2050 (N_2050,N_1458,N_1926);
or U2051 (N_2051,N_341,N_1693);
xor U2052 (N_2052,N_904,N_733);
xnor U2053 (N_2053,N_81,N_1962);
and U2054 (N_2054,N_1,N_871);
or U2055 (N_2055,N_629,N_1165);
xor U2056 (N_2056,N_762,N_940);
nand U2057 (N_2057,N_1307,N_761);
nor U2058 (N_2058,N_1271,N_1525);
xnor U2059 (N_2059,N_1704,N_1070);
nor U2060 (N_2060,N_688,N_197);
or U2061 (N_2061,N_1119,N_547);
and U2062 (N_2062,N_1925,N_507);
nand U2063 (N_2063,N_527,N_1566);
nor U2064 (N_2064,N_1638,N_1889);
or U2065 (N_2065,N_1453,N_1956);
xor U2066 (N_2066,N_764,N_1291);
and U2067 (N_2067,N_360,N_1662);
and U2068 (N_2068,N_793,N_602);
nor U2069 (N_2069,N_488,N_704);
and U2070 (N_2070,N_637,N_419);
or U2071 (N_2071,N_1553,N_55);
nand U2072 (N_2072,N_1179,N_654);
and U2073 (N_2073,N_789,N_338);
nor U2074 (N_2074,N_57,N_676);
nor U2075 (N_2075,N_1126,N_174);
nand U2076 (N_2076,N_1931,N_1014);
or U2077 (N_2077,N_1372,N_854);
xor U2078 (N_2078,N_246,N_83);
and U2079 (N_2079,N_1462,N_1519);
or U2080 (N_2080,N_968,N_667);
or U2081 (N_2081,N_378,N_426);
xnor U2082 (N_2082,N_1469,N_1574);
xor U2083 (N_2083,N_582,N_1426);
or U2084 (N_2084,N_540,N_1968);
or U2085 (N_2085,N_1801,N_1242);
or U2086 (N_2086,N_1897,N_410);
nand U2087 (N_2087,N_1520,N_606);
and U2088 (N_2088,N_1177,N_1337);
nand U2089 (N_2089,N_427,N_1848);
xnor U2090 (N_2090,N_1018,N_1534);
nand U2091 (N_2091,N_1555,N_1449);
and U2092 (N_2092,N_1533,N_1718);
xnor U2093 (N_2093,N_180,N_1691);
xnor U2094 (N_2094,N_2,N_101);
nand U2095 (N_2095,N_1817,N_1004);
nand U2096 (N_2096,N_1778,N_1585);
nor U2097 (N_2097,N_1651,N_1058);
or U2098 (N_2098,N_917,N_1416);
xor U2099 (N_2099,N_1809,N_1972);
and U2100 (N_2100,N_906,N_960);
nor U2101 (N_2101,N_623,N_280);
nand U2102 (N_2102,N_1980,N_1569);
nor U2103 (N_2103,N_1388,N_70);
nor U2104 (N_2104,N_406,N_873);
or U2105 (N_2105,N_498,N_435);
and U2106 (N_2106,N_120,N_415);
xnor U2107 (N_2107,N_1745,N_586);
nor U2108 (N_2108,N_1876,N_380);
or U2109 (N_2109,N_1163,N_570);
xnor U2110 (N_2110,N_247,N_93);
nand U2111 (N_2111,N_1101,N_1228);
and U2112 (N_2112,N_1118,N_1531);
nor U2113 (N_2113,N_716,N_624);
nor U2114 (N_2114,N_815,N_1109);
and U2115 (N_2115,N_164,N_935);
or U2116 (N_2116,N_134,N_1578);
nor U2117 (N_2117,N_1237,N_662);
or U2118 (N_2118,N_484,N_1514);
xnor U2119 (N_2119,N_1805,N_1679);
nor U2120 (N_2120,N_1011,N_564);
or U2121 (N_2121,N_1121,N_1996);
and U2122 (N_2122,N_1201,N_1522);
nand U2123 (N_2123,N_324,N_1919);
or U2124 (N_2124,N_691,N_1677);
xnor U2125 (N_2125,N_521,N_95);
or U2126 (N_2126,N_1727,N_1144);
or U2127 (N_2127,N_740,N_1846);
nand U2128 (N_2128,N_1496,N_1843);
nand U2129 (N_2129,N_1136,N_140);
and U2130 (N_2130,N_1466,N_1113);
nor U2131 (N_2131,N_1970,N_331);
and U2132 (N_2132,N_1621,N_1974);
and U2133 (N_2133,N_250,N_468);
and U2134 (N_2134,N_574,N_1222);
nand U2135 (N_2135,N_812,N_1867);
or U2136 (N_2136,N_170,N_1432);
and U2137 (N_2137,N_467,N_1103);
nor U2138 (N_2138,N_672,N_1492);
or U2139 (N_2139,N_1747,N_937);
and U2140 (N_2140,N_779,N_151);
or U2141 (N_2141,N_262,N_1976);
xor U2142 (N_2142,N_971,N_1787);
and U2143 (N_2143,N_1297,N_532);
nand U2144 (N_2144,N_625,N_352);
and U2145 (N_2145,N_353,N_1807);
and U2146 (N_2146,N_697,N_1336);
nor U2147 (N_2147,N_215,N_771);
nor U2148 (N_2148,N_124,N_438);
nand U2149 (N_2149,N_491,N_1360);
and U2150 (N_2150,N_307,N_1281);
nor U2151 (N_2151,N_1683,N_660);
nor U2152 (N_2152,N_1920,N_319);
xnor U2153 (N_2153,N_384,N_41);
nor U2154 (N_2154,N_457,N_320);
or U2155 (N_2155,N_1806,N_188);
nor U2156 (N_2156,N_1837,N_518);
nand U2157 (N_2157,N_1841,N_869);
and U2158 (N_2158,N_986,N_1610);
and U2159 (N_2159,N_1736,N_1783);
xor U2160 (N_2160,N_879,N_275);
and U2161 (N_2161,N_1199,N_494);
nor U2162 (N_2162,N_72,N_459);
and U2163 (N_2163,N_760,N_943);
and U2164 (N_2164,N_322,N_1130);
xor U2165 (N_2165,N_853,N_797);
nor U2166 (N_2166,N_712,N_1994);
or U2167 (N_2167,N_816,N_381);
and U2168 (N_2168,N_1486,N_155);
xor U2169 (N_2169,N_257,N_826);
and U2170 (N_2170,N_1879,N_1654);
and U2171 (N_2171,N_219,N_293);
nor U2172 (N_2172,N_1688,N_599);
xor U2173 (N_2173,N_428,N_767);
nor U2174 (N_2174,N_1763,N_1090);
nor U2175 (N_2175,N_213,N_63);
xnor U2176 (N_2176,N_1811,N_798);
or U2177 (N_2177,N_838,N_96);
and U2178 (N_2178,N_303,N_182);
nand U2179 (N_2179,N_572,N_289);
nor U2180 (N_2180,N_1212,N_1717);
nand U2181 (N_2181,N_1795,N_1435);
and U2182 (N_2182,N_115,N_1775);
xnor U2183 (N_2183,N_675,N_828);
nor U2184 (N_2184,N_1229,N_1409);
or U2185 (N_2185,N_1134,N_1915);
and U2186 (N_2186,N_1263,N_1853);
and U2187 (N_2187,N_782,N_845);
xnor U2188 (N_2188,N_1637,N_639);
xor U2189 (N_2189,N_243,N_901);
nand U2190 (N_2190,N_612,N_1636);
or U2191 (N_2191,N_16,N_1731);
and U2192 (N_2192,N_1401,N_551);
and U2193 (N_2193,N_33,N_786);
or U2194 (N_2194,N_1886,N_534);
xor U2195 (N_2195,N_344,N_1646);
nor U2196 (N_2196,N_588,N_1398);
or U2197 (N_2197,N_365,N_915);
nand U2198 (N_2198,N_287,N_1342);
or U2199 (N_2199,N_973,N_372);
nor U2200 (N_2200,N_1989,N_1756);
nor U2201 (N_2201,N_1684,N_1613);
and U2202 (N_2202,N_1794,N_1463);
nor U2203 (N_2203,N_1437,N_868);
nand U2204 (N_2204,N_1949,N_1023);
xor U2205 (N_2205,N_209,N_1026);
or U2206 (N_2206,N_461,N_1608);
and U2207 (N_2207,N_1369,N_1921);
nor U2208 (N_2208,N_1210,N_239);
nand U2209 (N_2209,N_178,N_1712);
and U2210 (N_2210,N_1211,N_942);
nand U2211 (N_2211,N_1836,N_1104);
nor U2212 (N_2212,N_1551,N_1859);
nand U2213 (N_2213,N_1563,N_806);
and U2214 (N_2214,N_536,N_1913);
xor U2215 (N_2215,N_1316,N_1995);
nand U2216 (N_2216,N_1476,N_724);
and U2217 (N_2217,N_150,N_1365);
nor U2218 (N_2218,N_308,N_214);
nand U2219 (N_2219,N_225,N_1855);
nor U2220 (N_2220,N_1154,N_1374);
and U2221 (N_2221,N_1629,N_1133);
or U2222 (N_2222,N_1003,N_1410);
xor U2223 (N_2223,N_430,N_229);
and U2224 (N_2224,N_1623,N_1256);
nor U2225 (N_2225,N_1149,N_557);
nand U2226 (N_2226,N_218,N_183);
xnor U2227 (N_2227,N_1702,N_1538);
and U2228 (N_2228,N_434,N_802);
and U2229 (N_2229,N_642,N_1063);
xor U2230 (N_2230,N_730,N_1363);
nor U2231 (N_2231,N_1813,N_1055);
xor U2232 (N_2232,N_1049,N_58);
nor U2233 (N_2233,N_1067,N_1748);
nor U2234 (N_2234,N_25,N_891);
or U2235 (N_2235,N_1788,N_1184);
xnor U2236 (N_2236,N_997,N_656);
nand U2237 (N_2237,N_1331,N_895);
and U2238 (N_2238,N_181,N_1706);
nand U2239 (N_2239,N_121,N_718);
xnor U2240 (N_2240,N_374,N_326);
nor U2241 (N_2241,N_1181,N_1441);
and U2242 (N_2242,N_1367,N_1554);
nand U2243 (N_2243,N_1112,N_923);
nor U2244 (N_2244,N_846,N_366);
xnor U2245 (N_2245,N_958,N_999);
and U2246 (N_2246,N_423,N_947);
or U2247 (N_2247,N_1376,N_1036);
and U2248 (N_2248,N_728,N_154);
nor U2249 (N_2249,N_126,N_1535);
or U2250 (N_2250,N_687,N_395);
nand U2251 (N_2251,N_1548,N_1078);
and U2252 (N_2252,N_1399,N_1862);
xor U2253 (N_2253,N_1547,N_1171);
xor U2254 (N_2254,N_737,N_600);
and U2255 (N_2255,N_1091,N_922);
nor U2256 (N_2256,N_817,N_1938);
nand U2257 (N_2257,N_159,N_835);
or U2258 (N_2258,N_455,N_1829);
or U2259 (N_2259,N_1830,N_1733);
xnor U2260 (N_2260,N_502,N_255);
or U2261 (N_2261,N_1059,N_962);
nor U2262 (N_2262,N_334,N_969);
or U2263 (N_2263,N_864,N_1287);
and U2264 (N_2264,N_1849,N_1189);
xnor U2265 (N_2265,N_147,N_389);
and U2266 (N_2266,N_998,N_1657);
xor U2267 (N_2267,N_1137,N_930);
and U2268 (N_2268,N_1270,N_664);
and U2269 (N_2269,N_742,N_1800);
nand U2270 (N_2270,N_773,N_1325);
nor U2271 (N_2271,N_439,N_474);
xor U2272 (N_2272,N_1758,N_1891);
and U2273 (N_2273,N_1445,N_1589);
and U2274 (N_2274,N_1580,N_414);
xnor U2275 (N_2275,N_1289,N_989);
nor U2276 (N_2276,N_1402,N_539);
and U2277 (N_2277,N_985,N_1515);
or U2278 (N_2278,N_1105,N_626);
xor U2279 (N_2279,N_1658,N_1205);
xor U2280 (N_2280,N_1456,N_984);
or U2281 (N_2281,N_825,N_591);
or U2282 (N_2282,N_1279,N_107);
nor U2283 (N_2283,N_1570,N_240);
or U2284 (N_2284,N_1017,N_1286);
xor U2285 (N_2285,N_187,N_291);
and U2286 (N_2286,N_1687,N_189);
or U2287 (N_2287,N_450,N_855);
xor U2288 (N_2288,N_872,N_185);
or U2289 (N_2289,N_1259,N_1042);
nor U2290 (N_2290,N_167,N_799);
nor U2291 (N_2291,N_1768,N_1153);
and U2292 (N_2292,N_822,N_1132);
and U2293 (N_2293,N_71,N_1633);
or U2294 (N_2294,N_1075,N_1564);
xnor U2295 (N_2295,N_1029,N_385);
nor U2296 (N_2296,N_757,N_1529);
nor U2297 (N_2297,N_529,N_517);
nand U2298 (N_2298,N_383,N_210);
xor U2299 (N_2299,N_1999,N_1142);
or U2300 (N_2300,N_333,N_1125);
xnor U2301 (N_2301,N_874,N_1898);
xor U2302 (N_2302,N_24,N_114);
nor U2303 (N_2303,N_1334,N_913);
and U2304 (N_2304,N_28,N_1790);
nand U2305 (N_2305,N_22,N_1810);
nor U2306 (N_2306,N_1725,N_885);
xor U2307 (N_2307,N_184,N_839);
xor U2308 (N_2308,N_1169,N_641);
and U2309 (N_2309,N_583,N_363);
and U2310 (N_2310,N_202,N_1282);
and U2311 (N_2311,N_492,N_512);
nand U2312 (N_2312,N_945,N_248);
nand U2313 (N_2313,N_1164,N_304);
and U2314 (N_2314,N_627,N_1825);
nor U2315 (N_2315,N_108,N_1151);
nor U2316 (N_2316,N_770,N_585);
nor U2317 (N_2317,N_8,N_13);
xnor U2318 (N_2318,N_138,N_886);
and U2319 (N_2319,N_752,N_1539);
xor U2320 (N_2320,N_1793,N_1735);
xor U2321 (N_2321,N_422,N_1935);
xor U2322 (N_2322,N_1387,N_933);
xor U2323 (N_2323,N_501,N_954);
nand U2324 (N_2324,N_1309,N_976);
nand U2325 (N_2325,N_1015,N_38);
nor U2326 (N_2326,N_1508,N_73);
or U2327 (N_2327,N_143,N_1663);
nor U2328 (N_2328,N_315,N_1713);
nand U2329 (N_2329,N_1934,N_1942);
nor U2330 (N_2330,N_859,N_1320);
xor U2331 (N_2331,N_1943,N_1513);
or U2332 (N_2332,N_1089,N_1226);
nor U2333 (N_2333,N_1631,N_1182);
or U2334 (N_2334,N_448,N_309);
xor U2335 (N_2335,N_1174,N_230);
xor U2336 (N_2336,N_1250,N_1827);
or U2337 (N_2337,N_1362,N_1739);
nand U2338 (N_2338,N_1382,N_525);
nand U2339 (N_2339,N_1734,N_1797);
nand U2340 (N_2340,N_1729,N_388);
xnor U2341 (N_2341,N_136,N_446);
nor U2342 (N_2342,N_284,N_888);
nor U2343 (N_2343,N_852,N_122);
or U2344 (N_2344,N_715,N_1714);
and U2345 (N_2345,N_490,N_794);
nor U2346 (N_2346,N_717,N_382);
and U2347 (N_2347,N_1924,N_929);
or U2348 (N_2348,N_1371,N_53);
and U2349 (N_2349,N_566,N_1755);
xor U2350 (N_2350,N_1129,N_302);
or U2351 (N_2351,N_653,N_1436);
nor U2352 (N_2352,N_556,N_1544);
and U2353 (N_2353,N_1819,N_1577);
nand U2354 (N_2354,N_1874,N_301);
or U2355 (N_2355,N_974,N_1583);
xor U2356 (N_2356,N_1959,N_875);
and U2357 (N_2357,N_562,N_192);
and U2358 (N_2358,N_775,N_1244);
and U2359 (N_2359,N_1527,N_701);
xor U2360 (N_2360,N_130,N_580);
or U2361 (N_2361,N_785,N_1301);
nor U2362 (N_2362,N_456,N_371);
and U2363 (N_2363,N_705,N_470);
nor U2364 (N_2364,N_714,N_565);
nand U2365 (N_2365,N_1310,N_818);
or U2366 (N_2366,N_1314,N_781);
xor U2367 (N_2367,N_1878,N_743);
or U2368 (N_2368,N_1258,N_628);
and U2369 (N_2369,N_791,N_833);
and U2370 (N_2370,N_1864,N_1028);
nor U2371 (N_2371,N_1854,N_890);
xor U2372 (N_2372,N_948,N_1045);
and U2373 (N_2373,N_1474,N_1277);
xnor U2374 (N_2374,N_1477,N_768);
and U2375 (N_2375,N_595,N_1283);
and U2376 (N_2376,N_1406,N_801);
and U2377 (N_2377,N_575,N_172);
or U2378 (N_2378,N_1979,N_158);
or U2379 (N_2379,N_1140,N_1170);
nand U2380 (N_2380,N_1760,N_541);
or U2381 (N_2381,N_1319,N_1678);
nor U2382 (N_2382,N_1944,N_1346);
nor U2383 (N_2383,N_824,N_146);
and U2384 (N_2384,N_1599,N_1542);
xor U2385 (N_2385,N_1990,N_1295);
and U2386 (N_2386,N_1575,N_412);
or U2387 (N_2387,N_7,N_991);
or U2388 (N_2388,N_1741,N_222);
and U2389 (N_2389,N_1219,N_269);
and U2390 (N_2390,N_80,N_1716);
or U2391 (N_2391,N_175,N_1611);
nand U2392 (N_2392,N_681,N_1700);
xnor U2393 (N_2393,N_573,N_211);
xor U2394 (N_2394,N_1408,N_283);
nor U2395 (N_2395,N_1641,N_398);
xor U2396 (N_2396,N_1506,N_312);
nand U2397 (N_2397,N_1054,N_466);
nor U2398 (N_2398,N_584,N_1200);
nand U2399 (N_2399,N_1417,N_663);
nand U2400 (N_2400,N_405,N_495);
nand U2401 (N_2401,N_191,N_711);
or U2402 (N_2402,N_516,N_292);
and U2403 (N_2403,N_49,N_1893);
xor U2404 (N_2404,N_1510,N_1987);
and U2405 (N_2405,N_1159,N_836);
nand U2406 (N_2406,N_1487,N_1123);
and U2407 (N_2407,N_112,N_1776);
xor U2408 (N_2408,N_375,N_925);
and U2409 (N_2409,N_1857,N_1888);
nand U2410 (N_2410,N_1072,N_1907);
nand U2411 (N_2411,N_1711,N_515);
and U2412 (N_2412,N_1224,N_478);
and U2413 (N_2413,N_1032,N_561);
and U2414 (N_2414,N_10,N_1779);
and U2415 (N_2415,N_266,N_1586);
or U2416 (N_2416,N_74,N_1967);
xor U2417 (N_2417,N_607,N_399);
or U2418 (N_2418,N_804,N_59);
or U2419 (N_2419,N_858,N_520);
and U2420 (N_2420,N_1973,N_1152);
and U2421 (N_2421,N_1928,N_1318);
nor U2422 (N_2422,N_537,N_1315);
or U2423 (N_2423,N_842,N_1789);
nand U2424 (N_2424,N_970,N_196);
and U2425 (N_2425,N_325,N_169);
nand U2426 (N_2426,N_1644,N_118);
and U2427 (N_2427,N_403,N_1632);
and U2428 (N_2428,N_408,N_1838);
nor U2429 (N_2429,N_669,N_892);
or U2430 (N_2430,N_1188,N_1088);
or U2431 (N_2431,N_729,N_203);
or U2432 (N_2432,N_1145,N_234);
xnor U2433 (N_2433,N_1180,N_509);
nor U2434 (N_2434,N_401,N_361);
xor U2435 (N_2435,N_1491,N_1447);
and U2436 (N_2436,N_1473,N_1961);
nor U2437 (N_2437,N_1518,N_679);
xnor U2438 (N_2438,N_957,N_1781);
xnor U2439 (N_2439,N_1701,N_765);
nor U2440 (N_2440,N_1927,N_1480);
xor U2441 (N_2441,N_1438,N_1617);
nand U2442 (N_2442,N_14,N_772);
nor U2443 (N_2443,N_251,N_297);
or U2444 (N_2444,N_563,N_1918);
and U2445 (N_2445,N_959,N_1459);
nand U2446 (N_2446,N_1526,N_212);
nor U2447 (N_2447,N_803,N_530);
or U2448 (N_2448,N_1626,N_554);
nand U2449 (N_2449,N_850,N_1869);
and U2450 (N_2450,N_1952,N_790);
and U2451 (N_2451,N_1602,N_113);
xnor U2452 (N_2452,N_1954,N_163);
nand U2453 (N_2453,N_1214,N_723);
nor U2454 (N_2454,N_1284,N_603);
nor U2455 (N_2455,N_1840,N_1139);
and U2456 (N_2456,N_1322,N_776);
xnor U2457 (N_2457,N_860,N_503);
or U2458 (N_2458,N_1957,N_533);
xnor U2459 (N_2459,N_483,N_1127);
nor U2460 (N_2460,N_788,N_800);
nor U2461 (N_2461,N_1828,N_30);
and U2462 (N_2462,N_548,N_1593);
and U2463 (N_2463,N_1652,N_898);
nand U2464 (N_2464,N_493,N_1591);
or U2465 (N_2465,N_1705,N_1494);
nor U2466 (N_2466,N_1708,N_104);
xor U2467 (N_2467,N_242,N_171);
nand U2468 (N_2468,N_1528,N_1628);
and U2469 (N_2469,N_916,N_436);
nand U2470 (N_2470,N_1366,N_1020);
nor U2471 (N_2471,N_587,N_1672);
nand U2472 (N_2472,N_1824,N_1080);
and U2473 (N_2473,N_1339,N_102);
nand U2474 (N_2474,N_34,N_926);
nand U2475 (N_2475,N_1969,N_604);
or U2476 (N_2476,N_881,N_1167);
nand U2477 (N_2477,N_1916,N_67);
and U2478 (N_2478,N_1584,N_1349);
xor U2479 (N_2479,N_442,N_1963);
or U2480 (N_2480,N_700,N_82);
xor U2481 (N_2481,N_390,N_1324);
or U2482 (N_2482,N_440,N_1472);
nor U2483 (N_2483,N_77,N_1245);
nand U2484 (N_2484,N_1640,N_1087);
or U2485 (N_2485,N_649,N_832);
nor U2486 (N_2486,N_645,N_1630);
xor U2487 (N_2487,N_1418,N_1723);
nor U2488 (N_2488,N_552,N_847);
nand U2489 (N_2489,N_689,N_12);
or U2490 (N_2490,N_413,N_359);
nor U2491 (N_2491,N_1086,N_615);
or U2492 (N_2492,N_1983,N_245);
and U2493 (N_2493,N_1590,N_499);
nand U2494 (N_2494,N_103,N_226);
nor U2495 (N_2495,N_1537,N_429);
nand U2496 (N_2496,N_1415,N_1930);
xnor U2497 (N_2497,N_1120,N_1818);
or U2498 (N_2498,N_1917,N_1675);
or U2499 (N_2499,N_1350,N_1231);
nand U2500 (N_2500,N_753,N_11);
nand U2501 (N_2501,N_305,N_299);
xnor U2502 (N_2502,N_1006,N_228);
xnor U2503 (N_2503,N_258,N_373);
or U2504 (N_2504,N_1909,N_808);
nor U2505 (N_2505,N_981,N_1155);
nand U2506 (N_2506,N_208,N_1558);
nand U2507 (N_2507,N_1596,N_1051);
and U2508 (N_2508,N_695,N_745);
xor U2509 (N_2509,N_1111,N_1338);
and U2510 (N_2510,N_622,N_914);
or U2511 (N_2511,N_921,N_1383);
and U2512 (N_2512,N_1061,N_23);
and U2513 (N_2513,N_677,N_953);
nor U2514 (N_2514,N_476,N_1428);
nand U2515 (N_2515,N_1467,N_685);
nand U2516 (N_2516,N_1292,N_837);
nor U2517 (N_2517,N_1460,N_992);
or U2518 (N_2518,N_1344,N_505);
nor U2519 (N_2519,N_1880,N_944);
and U2520 (N_2520,N_1908,N_1482);
nor U2521 (N_2521,N_1883,N_290);
nor U2522 (N_2522,N_1784,N_759);
nand U2523 (N_2523,N_894,N_236);
or U2524 (N_2524,N_465,N_1782);
xnor U2525 (N_2525,N_1050,N_611);
and U2526 (N_2526,N_376,N_1353);
or U2527 (N_2527,N_758,N_1618);
and U2528 (N_2528,N_650,N_1481);
nand U2529 (N_2529,N_237,N_931);
xnor U2530 (N_2530,N_553,N_35);
nor U2531 (N_2531,N_694,N_1722);
xor U2532 (N_2532,N_1803,N_1985);
xnor U2533 (N_2533,N_1207,N_558);
or U2534 (N_2534,N_286,N_139);
nand U2535 (N_2535,N_1255,N_1225);
nor U2536 (N_2536,N_6,N_1160);
nor U2537 (N_2537,N_1823,N_1730);
xor U2538 (N_2538,N_152,N_1195);
or U2539 (N_2539,N_1642,N_920);
nand U2540 (N_2540,N_1814,N_982);
nor U2541 (N_2541,N_1699,N_936);
nand U2542 (N_2542,N_1737,N_1031);
nand U2543 (N_2543,N_734,N_1073);
xor U2544 (N_2544,N_1340,N_821);
or U2545 (N_2545,N_129,N_271);
nand U2546 (N_2546,N_1721,N_964);
or U2547 (N_2547,N_421,N_610);
and U2548 (N_2548,N_987,N_156);
and U2549 (N_2549,N_148,N_29);
nor U2550 (N_2550,N_996,N_268);
nand U2551 (N_2551,N_1567,N_1396);
nor U2552 (N_2552,N_932,N_1614);
nand U2553 (N_2553,N_1196,N_949);
xnor U2554 (N_2554,N_177,N_1117);
and U2555 (N_2555,N_1187,N_447);
or U2556 (N_2556,N_1902,N_593);
or U2557 (N_2557,N_1391,N_1161);
xnor U2558 (N_2558,N_655,N_1442);
or U2559 (N_2559,N_1208,N_1414);
nand U2560 (N_2560,N_590,N_1624);
nor U2561 (N_2561,N_335,N_1774);
or U2562 (N_2562,N_1066,N_908);
xnor U2563 (N_2563,N_1786,N_620);
nor U2564 (N_2564,N_231,N_887);
or U2565 (N_2565,N_1220,N_1835);
nand U2566 (N_2566,N_861,N_26);
nor U2567 (N_2567,N_766,N_1268);
nand U2568 (N_2568,N_1490,N_1884);
and U2569 (N_2569,N_1766,N_1903);
nand U2570 (N_2570,N_902,N_1261);
and U2571 (N_2571,N_1065,N_1082);
xnor U2572 (N_2572,N_621,N_967);
nand U2573 (N_2573,N_224,N_1664);
or U2574 (N_2574,N_1052,N_905);
xnor U2575 (N_2575,N_1452,N_0);
nor U2576 (N_2576,N_856,N_1085);
nand U2577 (N_2577,N_1044,N_1749);
xor U2578 (N_2578,N_979,N_179);
nor U2579 (N_2579,N_1172,N_1507);
xnor U2580 (N_2580,N_17,N_1122);
nand U2581 (N_2581,N_1102,N_1582);
nor U2582 (N_2582,N_1572,N_1471);
nand U2583 (N_2583,N_975,N_1639);
nand U2584 (N_2584,N_1666,N_1559);
xor U2585 (N_2585,N_1557,N_1450);
xor U2586 (N_2586,N_195,N_680);
nand U2587 (N_2587,N_1016,N_805);
nand U2588 (N_2588,N_1333,N_1345);
nand U2589 (N_2589,N_990,N_528);
xor U2590 (N_2590,N_1306,N_1190);
xnor U2591 (N_2591,N_480,N_1257);
nand U2592 (N_2592,N_1272,N_267);
or U2593 (N_2593,N_538,N_1455);
nand U2594 (N_2594,N_1260,N_1393);
nand U2595 (N_2595,N_1804,N_1899);
or U2596 (N_2596,N_1265,N_1982);
nand U2597 (N_2597,N_1030,N_748);
nand U2598 (N_2598,N_1115,N_44);
xor U2599 (N_2599,N_424,N_988);
and U2600 (N_2600,N_878,N_1489);
or U2601 (N_2601,N_707,N_1504);
xnor U2602 (N_2602,N_1773,N_370);
nor U2603 (N_2603,N_1881,N_97);
xor U2604 (N_2604,N_61,N_88);
nor U2605 (N_2605,N_1047,N_313);
and U2606 (N_2606,N_1221,N_1204);
or U2607 (N_2607,N_1946,N_1420);
nor U2608 (N_2608,N_1468,N_50);
xor U2609 (N_2609,N_1479,N_1565);
xor U2610 (N_2610,N_1882,N_1965);
or U2611 (N_2611,N_1703,N_1929);
nand U2612 (N_2612,N_285,N_1709);
or U2613 (N_2613,N_1148,N_1213);
nor U2614 (N_2614,N_1351,N_1844);
nand U2615 (N_2615,N_559,N_1743);
nor U2616 (N_2616,N_489,N_281);
or U2617 (N_2617,N_542,N_1524);
or U2618 (N_2618,N_52,N_1690);
xor U2619 (N_2619,N_1873,N_597);
and U2620 (N_2620,N_631,N_409);
and U2621 (N_2621,N_1562,N_98);
and U2622 (N_2622,N_1892,N_342);
and U2623 (N_2623,N_201,N_1512);
nand U2624 (N_2624,N_1355,N_1380);
and U2625 (N_2625,N_1726,N_1950);
nand U2626 (N_2626,N_1833,N_109);
nand U2627 (N_2627,N_749,N_1378);
nand U2628 (N_2628,N_939,N_1327);
nand U2629 (N_2629,N_1839,N_750);
nor U2630 (N_2630,N_241,N_692);
nor U2631 (N_2631,N_1863,N_311);
nand U2632 (N_2632,N_1400,N_327);
or U2633 (N_2633,N_589,N_1311);
and U2634 (N_2634,N_407,N_596);
or U2635 (N_2635,N_755,N_784);
or U2636 (N_2636,N_1936,N_205);
or U2637 (N_2637,N_1488,N_317);
nand U2638 (N_2638,N_1752,N_666);
and U2639 (N_2639,N_1370,N_264);
nand U2640 (N_2640,N_751,N_1057);
nor U2641 (N_2641,N_659,N_1796);
nor U2642 (N_2642,N_1024,N_1203);
and U2643 (N_2643,N_116,N_1754);
and U2644 (N_2644,N_1966,N_496);
and U2645 (N_2645,N_100,N_1649);
xnor U2646 (N_2646,N_123,N_952);
xor U2647 (N_2647,N_1001,N_1719);
nand U2648 (N_2648,N_141,N_1682);
xnor U2649 (N_2649,N_1264,N_1945);
and U2650 (N_2650,N_848,N_1670);
nor U2651 (N_2651,N_1680,N_1619);
or U2652 (N_2652,N_865,N_1381);
nand U2653 (N_2653,N_1278,N_613);
nand U2654 (N_2654,N_1280,N_1603);
and U2655 (N_2655,N_1035,N_1751);
and U2656 (N_2656,N_345,N_1901);
nor U2657 (N_2657,N_956,N_256);
nor U2658 (N_2658,N_1233,N_1183);
xor U2659 (N_2659,N_665,N_508);
nor U2660 (N_2660,N_316,N_1941);
nand U2661 (N_2661,N_1368,N_500);
nand U2662 (N_2662,N_919,N_288);
nand U2663 (N_2663,N_870,N_1832);
nor U2664 (N_2664,N_1275,N_1532);
and U2665 (N_2665,N_356,N_1427);
xnor U2666 (N_2666,N_810,N_809);
or U2667 (N_2667,N_644,N_1254);
or U2668 (N_2668,N_1108,N_683);
and U2669 (N_2669,N_1587,N_1503);
nand U2670 (N_2670,N_244,N_966);
xor U2671 (N_2671,N_1834,N_497);
xnor U2672 (N_2672,N_1252,N_658);
nand U2673 (N_2673,N_1655,N_1012);
or U2674 (N_2674,N_1403,N_76);
or U2675 (N_2675,N_45,N_1106);
and U2676 (N_2676,N_1914,N_978);
xnor U2677 (N_2677,N_1728,N_1227);
or U2678 (N_2678,N_831,N_1313);
or U2679 (N_2679,N_1110,N_1317);
or U2680 (N_2680,N_1724,N_531);
and U2681 (N_2681,N_1240,N_1971);
or U2682 (N_2682,N_963,N_1771);
nand U2683 (N_2683,N_161,N_111);
or U2684 (N_2684,N_282,N_1634);
nand U2685 (N_2685,N_934,N_1269);
and U2686 (N_2686,N_1041,N_1419);
nand U2687 (N_2687,N_568,N_106);
or U2688 (N_2688,N_464,N_1792);
or U2689 (N_2689,N_221,N_1364);
or U2690 (N_2690,N_54,N_1821);
xor U2691 (N_2691,N_1194,N_994);
nor U2692 (N_2692,N_37,N_576);
nor U2693 (N_2693,N_1767,N_1235);
xnor U2694 (N_2694,N_1761,N_1523);
nor U2695 (N_2695,N_1981,N_273);
nand U2696 (N_2696,N_1612,N_1552);
and U2697 (N_2697,N_1753,N_1694);
nor U2698 (N_2698,N_1872,N_1759);
and U2699 (N_2699,N_441,N_605);
nor U2700 (N_2700,N_594,N_571);
nand U2701 (N_2701,N_1686,N_1948);
xor U2702 (N_2702,N_1545,N_844);
nand U2703 (N_2703,N_411,N_577);
and U2704 (N_2704,N_1146,N_513);
nand U2705 (N_2705,N_1561,N_1079);
and U2706 (N_2706,N_431,N_598);
xor U2707 (N_2707,N_896,N_792);
xnor U2708 (N_2708,N_581,N_1138);
or U2709 (N_2709,N_635,N_1290);
xnor U2710 (N_2710,N_36,N_867);
or U2711 (N_2711,N_278,N_39);
or U2712 (N_2712,N_358,N_1988);
or U2713 (N_2713,N_1615,N_857);
and U2714 (N_2714,N_1069,N_1698);
nor U2715 (N_2715,N_1681,N_698);
or U2716 (N_2716,N_1198,N_1423);
or U2717 (N_2717,N_394,N_1019);
or U2718 (N_2718,N_87,N_1581);
xnor U2719 (N_2719,N_1303,N_1158);
nor U2720 (N_2720,N_473,N_1597);
or U2721 (N_2721,N_1093,N_796);
and U2722 (N_2722,N_549,N_261);
nor U2723 (N_2723,N_220,N_1107);
and U2724 (N_2724,N_1958,N_416);
nand U2725 (N_2725,N_3,N_216);
xnor U2726 (N_2726,N_1392,N_638);
nand U2727 (N_2727,N_364,N_1027);
nand U2728 (N_2728,N_1304,N_673);
nor U2729 (N_2729,N_1216,N_506);
and U2730 (N_2730,N_546,N_1517);
nor U2731 (N_2731,N_535,N_819);
nor U2732 (N_2732,N_1890,N_876);
and U2733 (N_2733,N_425,N_94);
nor U2734 (N_2734,N_754,N_1978);
and U2735 (N_2735,N_475,N_1197);
or U2736 (N_2736,N_1984,N_1037);
xnor U2737 (N_2737,N_472,N_1769);
and U2738 (N_2738,N_1594,N_1232);
nand U2739 (N_2739,N_1556,N_1299);
and U2740 (N_2740,N_321,N_1071);
nor U2741 (N_2741,N_1025,N_1906);
nor U2742 (N_2742,N_795,N_47);
xnor U2743 (N_2743,N_223,N_1757);
or U2744 (N_2744,N_1643,N_1822);
xnor U2745 (N_2745,N_1294,N_1870);
xor U2746 (N_2746,N_1247,N_1074);
nor U2747 (N_2747,N_780,N_469);
or U2748 (N_2748,N_485,N_128);
nor U2749 (N_2749,N_168,N_671);
and U2750 (N_2750,N_783,N_1097);
and U2751 (N_2751,N_1298,N_1904);
or U2752 (N_2752,N_652,N_1046);
and U2753 (N_2753,N_1820,N_1673);
and U2754 (N_2754,N_477,N_481);
and U2755 (N_2755,N_1647,N_295);
nand U2756 (N_2756,N_1932,N_1856);
xnor U2757 (N_2757,N_774,N_1484);
nand U2758 (N_2758,N_90,N_340);
nor U2759 (N_2759,N_1521,N_1191);
nand U2760 (N_2760,N_1421,N_618);
and U2761 (N_2761,N_199,N_1799);
nor U2762 (N_2762,N_391,N_1412);
xor U2763 (N_2763,N_763,N_1223);
nand U2764 (N_2764,N_259,N_110);
and U2765 (N_2765,N_670,N_420);
and U2766 (N_2766,N_1860,N_699);
and U2767 (N_2767,N_648,N_1997);
nor U2768 (N_2768,N_1246,N_69);
nor U2769 (N_2769,N_1095,N_1549);
nand U2770 (N_2770,N_1616,N_1852);
nor U2771 (N_2771,N_1770,N_89);
nor U2772 (N_2772,N_479,N_1964);
or U2773 (N_2773,N_1845,N_86);
and U2774 (N_2774,N_1960,N_1395);
or U2775 (N_2775,N_1326,N_1186);
nor U2776 (N_2776,N_592,N_453);
and U2777 (N_2777,N_1992,N_1571);
and U2778 (N_2778,N_523,N_567);
nand U2779 (N_2779,N_1425,N_1676);
and U2780 (N_2780,N_1323,N_713);
xor U2781 (N_2781,N_487,N_482);
nand U2782 (N_2782,N_686,N_137);
and U2783 (N_2783,N_1192,N_1385);
xnor U2784 (N_2784,N_550,N_1464);
or U2785 (N_2785,N_1986,N_1173);
nor U2786 (N_2786,N_1785,N_504);
nand U2787 (N_2787,N_1341,N_1653);
xnor U2788 (N_2788,N_977,N_841);
nor U2789 (N_2789,N_1923,N_1135);
nor U2790 (N_2790,N_32,N_893);
or U2791 (N_2791,N_1605,N_1443);
xor U2792 (N_2792,N_1953,N_48);
or U2793 (N_2793,N_75,N_162);
nand U2794 (N_2794,N_265,N_1084);
nand U2795 (N_2795,N_79,N_238);
or U2796 (N_2796,N_131,N_1147);
and U2797 (N_2797,N_27,N_823);
or U2798 (N_2798,N_1550,N_1896);
xnor U2799 (N_2799,N_166,N_1081);
nand U2800 (N_2800,N_1424,N_1877);
nand U2801 (N_2801,N_186,N_1592);
nand U2802 (N_2802,N_609,N_1540);
and U2803 (N_2803,N_1742,N_1285);
xor U2804 (N_2804,N_1305,N_153);
and U2805 (N_2805,N_343,N_778);
and U2806 (N_2806,N_1389,N_1560);
or U2807 (N_2807,N_1010,N_1092);
nand U2808 (N_2808,N_1485,N_1022);
and U2809 (N_2809,N_1674,N_1894);
nand U2810 (N_2810,N_1444,N_1176);
xor U2811 (N_2811,N_386,N_452);
and U2812 (N_2812,N_397,N_1955);
or U2813 (N_2813,N_19,N_252);
nor U2814 (N_2814,N_1021,N_1791);
xor U2815 (N_2815,N_545,N_884);
and U2816 (N_2816,N_995,N_144);
and U2817 (N_2817,N_193,N_84);
or U2818 (N_2818,N_632,N_840);
nor U2819 (N_2819,N_710,N_1043);
nor U2820 (N_2820,N_349,N_1493);
nand U2821 (N_2821,N_1868,N_1009);
nor U2822 (N_2822,N_1002,N_444);
nand U2823 (N_2823,N_417,N_983);
nor U2824 (N_2824,N_369,N_486);
or U2825 (N_2825,N_1606,N_1397);
nor U2826 (N_2826,N_738,N_260);
nand U2827 (N_2827,N_1034,N_1433);
nor U2828 (N_2828,N_1193,N_1178);
nand U2829 (N_2829,N_1099,N_1060);
xnor U2830 (N_2830,N_1053,N_630);
and U2831 (N_2831,N_736,N_198);
and U2832 (N_2832,N_1939,N_377);
xor U2833 (N_2833,N_827,N_634);
or U2834 (N_2834,N_332,N_1568);
and U2835 (N_2835,N_51,N_1895);
and U2836 (N_2836,N_722,N_310);
or U2837 (N_2837,N_85,N_200);
nand U2838 (N_2838,N_912,N_843);
xor U2839 (N_2839,N_661,N_980);
nor U2840 (N_2840,N_1671,N_1241);
nand U2841 (N_2841,N_927,N_1386);
nor U2842 (N_2842,N_1744,N_1588);
or U2843 (N_2843,N_1861,N_1056);
or U2844 (N_2844,N_270,N_276);
nand U2845 (N_2845,N_1851,N_955);
nor U2846 (N_2846,N_1288,N_646);
and U2847 (N_2847,N_1505,N_1710);
and U2848 (N_2848,N_157,N_1842);
xnor U2849 (N_2849,N_418,N_709);
nor U2850 (N_2850,N_437,N_46);
xnor U2851 (N_2851,N_92,N_643);
xnor U2852 (N_2852,N_1430,N_328);
xor U2853 (N_2853,N_1661,N_253);
or U2854 (N_2854,N_739,N_1013);
xnor U2855 (N_2855,N_911,N_1501);
and U2856 (N_2856,N_1720,N_1390);
nor U2857 (N_2857,N_882,N_909);
nor U2858 (N_2858,N_339,N_693);
nor U2859 (N_2859,N_362,N_1124);
nor U2860 (N_2860,N_1816,N_569);
nor U2861 (N_2861,N_690,N_4);
nor U2862 (N_2862,N_1697,N_132);
and U2863 (N_2863,N_15,N_910);
nand U2864 (N_2864,N_232,N_1217);
or U2865 (N_2865,N_1230,N_721);
xnor U2866 (N_2866,N_938,N_510);
nand U2867 (N_2867,N_787,N_1446);
xnor U2868 (N_2868,N_1202,N_1215);
nor U2869 (N_2869,N_1940,N_1911);
or U2870 (N_2870,N_1422,N_1361);
and U2871 (N_2871,N_777,N_1007);
nor U2872 (N_2872,N_1991,N_1168);
nand U2873 (N_2873,N_608,N_1831);
or U2874 (N_2874,N_142,N_1033);
or U2875 (N_2875,N_993,N_719);
or U2876 (N_2876,N_972,N_1377);
nand U2877 (N_2877,N_318,N_1573);
nand U2878 (N_2878,N_65,N_899);
or U2879 (N_2879,N_127,N_1635);
xor U2880 (N_2880,N_56,N_449);
nor U2881 (N_2881,N_1622,N_1607);
nor U2882 (N_2882,N_1431,N_1576);
nand U2883 (N_2883,N_1887,N_462);
xnor U2884 (N_2884,N_62,N_747);
nand U2885 (N_2885,N_1077,N_1765);
xor U2886 (N_2886,N_1665,N_1405);
and U2887 (N_2887,N_769,N_862);
nand U2888 (N_2888,N_329,N_1308);
and U2889 (N_2889,N_1600,N_1900);
nand U2890 (N_2890,N_1439,N_1669);
and U2891 (N_2891,N_404,N_402);
xor U2892 (N_2892,N_668,N_619);
xnor U2893 (N_2893,N_727,N_1440);
xnor U2894 (N_2894,N_367,N_1096);
and U2895 (N_2895,N_1348,N_1858);
and U2896 (N_2896,N_965,N_544);
xnor U2897 (N_2897,N_254,N_294);
or U2898 (N_2898,N_9,N_735);
and U2899 (N_2899,N_64,N_1750);
nand U2900 (N_2900,N_66,N_357);
xor U2901 (N_2901,N_1502,N_1740);
and U2902 (N_2902,N_1407,N_1329);
nor U2903 (N_2903,N_1530,N_863);
or U2904 (N_2904,N_1076,N_1384);
and U2905 (N_2905,N_1497,N_1300);
xnor U2906 (N_2906,N_160,N_918);
nand U2907 (N_2907,N_1905,N_946);
or U2908 (N_2908,N_883,N_1040);
nand U2909 (N_2909,N_355,N_1933);
nor U2910 (N_2910,N_21,N_897);
nand U2911 (N_2911,N_1162,N_337);
or U2912 (N_2912,N_5,N_1866);
xnor U2913 (N_2913,N_387,N_1116);
nor U2914 (N_2914,N_657,N_1064);
xnor U2915 (N_2915,N_119,N_300);
nor U2916 (N_2916,N_1429,N_903);
xnor U2917 (N_2917,N_1668,N_1495);
nor U2918 (N_2918,N_756,N_941);
and U2919 (N_2919,N_834,N_633);
nand U2920 (N_2920,N_1470,N_99);
xnor U2921 (N_2921,N_1236,N_20);
and U2922 (N_2922,N_1175,N_1094);
and U2923 (N_2923,N_1347,N_732);
xnor U2924 (N_2924,N_682,N_1536);
nor U2925 (N_2925,N_194,N_314);
xnor U2926 (N_2926,N_1475,N_190);
nand U2927 (N_2927,N_393,N_579);
or U2928 (N_2928,N_731,N_1296);
or U2929 (N_2929,N_1131,N_460);
or U2930 (N_2930,N_614,N_1685);
xnor U2931 (N_2931,N_1847,N_1328);
nand U2932 (N_2932,N_1500,N_1865);
or U2933 (N_2933,N_105,N_336);
nand U2934 (N_2934,N_233,N_125);
or U2935 (N_2935,N_1330,N_1764);
or U2936 (N_2936,N_347,N_1498);
nand U2937 (N_2937,N_1815,N_1511);
and U2938 (N_2938,N_1239,N_1922);
nand U2939 (N_2939,N_1038,N_1762);
nand U2940 (N_2940,N_1620,N_1394);
xnor U2941 (N_2941,N_1068,N_1715);
or U2942 (N_2942,N_354,N_1947);
and U2943 (N_2943,N_900,N_400);
or U2944 (N_2944,N_1157,N_526);
nand U2945 (N_2945,N_1656,N_227);
or U2946 (N_2946,N_1354,N_1746);
or U2947 (N_2947,N_1359,N_330);
xnor U2948 (N_2948,N_617,N_555);
or U2949 (N_2949,N_1977,N_1802);
or U2950 (N_2950,N_1609,N_1062);
and U2951 (N_2951,N_1243,N_1274);
nor U2952 (N_2952,N_1248,N_433);
nor U2953 (N_2953,N_1732,N_1234);
nand U2954 (N_2954,N_451,N_1454);
nor U2955 (N_2955,N_741,N_1302);
nand U2956 (N_2956,N_1262,N_348);
nor U2957 (N_2957,N_379,N_907);
xnor U2958 (N_2958,N_1579,N_1798);
nand U2959 (N_2959,N_1166,N_1005);
and U2960 (N_2960,N_43,N_1826);
xnor U2961 (N_2961,N_117,N_1627);
xor U2962 (N_2962,N_746,N_1335);
and U2963 (N_2963,N_277,N_928);
nor U2964 (N_2964,N_1358,N_726);
nor U2965 (N_2965,N_522,N_1150);
and U2966 (N_2966,N_149,N_877);
nand U2967 (N_2967,N_725,N_1276);
xor U2968 (N_2968,N_296,N_702);
xnor U2969 (N_2969,N_454,N_1777);
nor U2970 (N_2970,N_1375,N_206);
nand U2971 (N_2971,N_31,N_1910);
nand U2972 (N_2972,N_1478,N_323);
nor U2973 (N_2973,N_1206,N_1156);
nor U2974 (N_2974,N_1352,N_720);
nor U2975 (N_2975,N_173,N_1650);
or U2976 (N_2976,N_1850,N_1185);
or U2977 (N_2977,N_1098,N_1404);
nor U2978 (N_2978,N_601,N_458);
xnor U2979 (N_2979,N_961,N_1696);
nor U2980 (N_2980,N_1546,N_1457);
nor U2981 (N_2981,N_1692,N_511);
and U2982 (N_2982,N_1772,N_1357);
nand U2983 (N_2983,N_1253,N_514);
nor U2984 (N_2984,N_524,N_1483);
nor U2985 (N_2985,N_235,N_1000);
and U2986 (N_2986,N_1975,N_346);
or U2987 (N_2987,N_1209,N_696);
nand U2988 (N_2988,N_851,N_396);
nor U2989 (N_2989,N_78,N_1660);
or U2990 (N_2990,N_1509,N_674);
and U2991 (N_2991,N_471,N_1885);
nand U2992 (N_2992,N_204,N_814);
or U2993 (N_2993,N_1780,N_145);
nand U2994 (N_2994,N_1141,N_1312);
or U2995 (N_2995,N_1993,N_1128);
or U2996 (N_2996,N_1516,N_807);
nand U2997 (N_2997,N_1143,N_1321);
or U2998 (N_2998,N_1293,N_951);
or U2999 (N_2999,N_950,N_1249);
nand U3000 (N_3000,N_686,N_402);
xnor U3001 (N_3001,N_1530,N_417);
nand U3002 (N_3002,N_450,N_1121);
and U3003 (N_3003,N_188,N_107);
nand U3004 (N_3004,N_1929,N_385);
or U3005 (N_3005,N_1429,N_674);
xnor U3006 (N_3006,N_1589,N_1975);
xnor U3007 (N_3007,N_1806,N_1512);
xor U3008 (N_3008,N_1860,N_852);
xnor U3009 (N_3009,N_27,N_1929);
xnor U3010 (N_3010,N_717,N_1576);
nor U3011 (N_3011,N_622,N_122);
xor U3012 (N_3012,N_1362,N_22);
xor U3013 (N_3013,N_378,N_524);
nand U3014 (N_3014,N_622,N_790);
and U3015 (N_3015,N_1572,N_1418);
and U3016 (N_3016,N_1852,N_746);
xnor U3017 (N_3017,N_1558,N_1875);
nand U3018 (N_3018,N_367,N_769);
and U3019 (N_3019,N_1819,N_659);
and U3020 (N_3020,N_728,N_1999);
xnor U3021 (N_3021,N_1863,N_1213);
or U3022 (N_3022,N_1827,N_432);
nor U3023 (N_3023,N_37,N_1489);
xor U3024 (N_3024,N_393,N_1821);
nand U3025 (N_3025,N_1367,N_889);
nand U3026 (N_3026,N_1369,N_458);
xnor U3027 (N_3027,N_895,N_1469);
nand U3028 (N_3028,N_1747,N_745);
or U3029 (N_3029,N_448,N_1919);
xnor U3030 (N_3030,N_1530,N_1449);
or U3031 (N_3031,N_327,N_496);
and U3032 (N_3032,N_1655,N_1486);
xor U3033 (N_3033,N_1087,N_562);
nor U3034 (N_3034,N_1365,N_267);
nor U3035 (N_3035,N_144,N_1926);
nor U3036 (N_3036,N_636,N_1109);
or U3037 (N_3037,N_217,N_647);
nand U3038 (N_3038,N_461,N_316);
or U3039 (N_3039,N_301,N_1390);
xor U3040 (N_3040,N_1419,N_1154);
and U3041 (N_3041,N_793,N_841);
or U3042 (N_3042,N_1293,N_397);
or U3043 (N_3043,N_470,N_1805);
xnor U3044 (N_3044,N_1571,N_835);
xnor U3045 (N_3045,N_1078,N_591);
nor U3046 (N_3046,N_1465,N_427);
nand U3047 (N_3047,N_81,N_1694);
or U3048 (N_3048,N_1227,N_654);
nor U3049 (N_3049,N_300,N_922);
or U3050 (N_3050,N_873,N_1208);
or U3051 (N_3051,N_854,N_724);
xor U3052 (N_3052,N_1936,N_1745);
or U3053 (N_3053,N_947,N_805);
or U3054 (N_3054,N_1815,N_841);
xor U3055 (N_3055,N_1255,N_1022);
or U3056 (N_3056,N_423,N_1887);
nand U3057 (N_3057,N_945,N_305);
and U3058 (N_3058,N_1082,N_1891);
xnor U3059 (N_3059,N_974,N_1137);
nand U3060 (N_3060,N_1831,N_929);
xnor U3061 (N_3061,N_957,N_554);
or U3062 (N_3062,N_1859,N_1079);
nor U3063 (N_3063,N_1497,N_1841);
nand U3064 (N_3064,N_1515,N_137);
and U3065 (N_3065,N_1724,N_279);
and U3066 (N_3066,N_1381,N_852);
xnor U3067 (N_3067,N_480,N_1868);
nor U3068 (N_3068,N_837,N_104);
or U3069 (N_3069,N_1091,N_1796);
xnor U3070 (N_3070,N_1833,N_1379);
or U3071 (N_3071,N_511,N_1791);
or U3072 (N_3072,N_1907,N_647);
nand U3073 (N_3073,N_977,N_1962);
and U3074 (N_3074,N_1368,N_228);
and U3075 (N_3075,N_750,N_775);
nor U3076 (N_3076,N_280,N_1019);
or U3077 (N_3077,N_219,N_321);
nand U3078 (N_3078,N_946,N_184);
nor U3079 (N_3079,N_1144,N_1232);
xor U3080 (N_3080,N_1796,N_1790);
xor U3081 (N_3081,N_227,N_1032);
xnor U3082 (N_3082,N_25,N_921);
xnor U3083 (N_3083,N_1158,N_476);
and U3084 (N_3084,N_1802,N_1562);
xor U3085 (N_3085,N_1454,N_173);
or U3086 (N_3086,N_292,N_130);
and U3087 (N_3087,N_902,N_867);
nand U3088 (N_3088,N_1466,N_1988);
and U3089 (N_3089,N_1356,N_1294);
nor U3090 (N_3090,N_1968,N_1776);
or U3091 (N_3091,N_86,N_1941);
xor U3092 (N_3092,N_1961,N_869);
xnor U3093 (N_3093,N_272,N_280);
nor U3094 (N_3094,N_1780,N_350);
or U3095 (N_3095,N_535,N_465);
xnor U3096 (N_3096,N_1160,N_870);
and U3097 (N_3097,N_366,N_535);
and U3098 (N_3098,N_1411,N_1620);
nand U3099 (N_3099,N_1612,N_1270);
and U3100 (N_3100,N_364,N_1608);
and U3101 (N_3101,N_1440,N_1374);
nand U3102 (N_3102,N_1835,N_1550);
or U3103 (N_3103,N_962,N_1262);
nand U3104 (N_3104,N_1926,N_1267);
xor U3105 (N_3105,N_1619,N_222);
xnor U3106 (N_3106,N_1545,N_134);
or U3107 (N_3107,N_69,N_1504);
nor U3108 (N_3108,N_746,N_593);
or U3109 (N_3109,N_508,N_140);
nand U3110 (N_3110,N_1150,N_1028);
nor U3111 (N_3111,N_1274,N_853);
xnor U3112 (N_3112,N_1108,N_1819);
and U3113 (N_3113,N_850,N_203);
or U3114 (N_3114,N_1237,N_1672);
or U3115 (N_3115,N_1849,N_501);
and U3116 (N_3116,N_1487,N_313);
or U3117 (N_3117,N_698,N_1835);
nand U3118 (N_3118,N_907,N_861);
nor U3119 (N_3119,N_1062,N_1319);
xor U3120 (N_3120,N_1205,N_1964);
or U3121 (N_3121,N_1709,N_1742);
and U3122 (N_3122,N_91,N_737);
nand U3123 (N_3123,N_666,N_1600);
nand U3124 (N_3124,N_602,N_17);
nor U3125 (N_3125,N_1233,N_494);
and U3126 (N_3126,N_1686,N_1137);
and U3127 (N_3127,N_588,N_989);
or U3128 (N_3128,N_1355,N_1259);
and U3129 (N_3129,N_482,N_391);
nor U3130 (N_3130,N_1656,N_1895);
nand U3131 (N_3131,N_1212,N_58);
xor U3132 (N_3132,N_384,N_1594);
nor U3133 (N_3133,N_1682,N_42);
nor U3134 (N_3134,N_1589,N_1247);
or U3135 (N_3135,N_199,N_1364);
nor U3136 (N_3136,N_548,N_1847);
xnor U3137 (N_3137,N_416,N_1489);
or U3138 (N_3138,N_1796,N_1280);
and U3139 (N_3139,N_702,N_873);
nand U3140 (N_3140,N_275,N_1486);
or U3141 (N_3141,N_1496,N_1435);
nand U3142 (N_3142,N_1948,N_1941);
nand U3143 (N_3143,N_1675,N_1624);
nand U3144 (N_3144,N_377,N_152);
nor U3145 (N_3145,N_312,N_1855);
xor U3146 (N_3146,N_1015,N_617);
nand U3147 (N_3147,N_933,N_1950);
nor U3148 (N_3148,N_1140,N_1989);
or U3149 (N_3149,N_1726,N_169);
nor U3150 (N_3150,N_1971,N_1754);
xnor U3151 (N_3151,N_1061,N_366);
or U3152 (N_3152,N_89,N_232);
nand U3153 (N_3153,N_296,N_904);
nor U3154 (N_3154,N_1370,N_993);
xnor U3155 (N_3155,N_815,N_787);
and U3156 (N_3156,N_254,N_403);
nand U3157 (N_3157,N_380,N_1339);
or U3158 (N_3158,N_1861,N_388);
and U3159 (N_3159,N_284,N_423);
nor U3160 (N_3160,N_89,N_590);
xor U3161 (N_3161,N_1860,N_1649);
xor U3162 (N_3162,N_37,N_1823);
nand U3163 (N_3163,N_1569,N_131);
xor U3164 (N_3164,N_814,N_941);
and U3165 (N_3165,N_836,N_866);
nor U3166 (N_3166,N_44,N_1055);
xnor U3167 (N_3167,N_1022,N_554);
nand U3168 (N_3168,N_742,N_1480);
nor U3169 (N_3169,N_1324,N_951);
nand U3170 (N_3170,N_195,N_1565);
and U3171 (N_3171,N_533,N_717);
nor U3172 (N_3172,N_496,N_160);
xor U3173 (N_3173,N_1214,N_261);
and U3174 (N_3174,N_1186,N_1501);
xnor U3175 (N_3175,N_577,N_1402);
nand U3176 (N_3176,N_174,N_148);
nor U3177 (N_3177,N_1467,N_1809);
or U3178 (N_3178,N_1399,N_1839);
and U3179 (N_3179,N_1703,N_809);
or U3180 (N_3180,N_1729,N_217);
and U3181 (N_3181,N_525,N_1521);
xor U3182 (N_3182,N_572,N_1903);
or U3183 (N_3183,N_1430,N_350);
nor U3184 (N_3184,N_1680,N_522);
nand U3185 (N_3185,N_1612,N_50);
and U3186 (N_3186,N_1164,N_959);
nor U3187 (N_3187,N_1022,N_1437);
and U3188 (N_3188,N_773,N_1439);
or U3189 (N_3189,N_416,N_1679);
nand U3190 (N_3190,N_1400,N_671);
nor U3191 (N_3191,N_1788,N_1904);
xnor U3192 (N_3192,N_647,N_1922);
xor U3193 (N_3193,N_481,N_825);
nor U3194 (N_3194,N_1652,N_1659);
and U3195 (N_3195,N_727,N_1377);
and U3196 (N_3196,N_309,N_1172);
and U3197 (N_3197,N_884,N_1225);
xnor U3198 (N_3198,N_97,N_1451);
and U3199 (N_3199,N_900,N_1633);
and U3200 (N_3200,N_1228,N_117);
nor U3201 (N_3201,N_1103,N_293);
and U3202 (N_3202,N_571,N_1613);
or U3203 (N_3203,N_140,N_1802);
or U3204 (N_3204,N_1447,N_320);
nor U3205 (N_3205,N_478,N_639);
xnor U3206 (N_3206,N_1391,N_310);
xnor U3207 (N_3207,N_760,N_191);
or U3208 (N_3208,N_612,N_1272);
or U3209 (N_3209,N_204,N_293);
or U3210 (N_3210,N_1484,N_501);
nand U3211 (N_3211,N_95,N_1407);
or U3212 (N_3212,N_1698,N_606);
xor U3213 (N_3213,N_880,N_407);
and U3214 (N_3214,N_1470,N_516);
and U3215 (N_3215,N_1966,N_358);
and U3216 (N_3216,N_1911,N_1521);
xor U3217 (N_3217,N_1414,N_242);
nor U3218 (N_3218,N_83,N_584);
nand U3219 (N_3219,N_1232,N_1690);
nor U3220 (N_3220,N_1558,N_1191);
and U3221 (N_3221,N_1206,N_626);
xor U3222 (N_3222,N_792,N_1153);
and U3223 (N_3223,N_255,N_943);
xnor U3224 (N_3224,N_1111,N_315);
and U3225 (N_3225,N_31,N_724);
xnor U3226 (N_3226,N_558,N_976);
and U3227 (N_3227,N_1432,N_1281);
or U3228 (N_3228,N_1976,N_1369);
nor U3229 (N_3229,N_769,N_1610);
nand U3230 (N_3230,N_1660,N_1915);
nand U3231 (N_3231,N_1414,N_1443);
or U3232 (N_3232,N_1925,N_1018);
or U3233 (N_3233,N_564,N_632);
nor U3234 (N_3234,N_1908,N_1794);
and U3235 (N_3235,N_1654,N_1986);
and U3236 (N_3236,N_1219,N_584);
or U3237 (N_3237,N_489,N_1019);
or U3238 (N_3238,N_191,N_641);
xnor U3239 (N_3239,N_1289,N_181);
xor U3240 (N_3240,N_1537,N_1202);
nor U3241 (N_3241,N_1441,N_1195);
nand U3242 (N_3242,N_712,N_926);
or U3243 (N_3243,N_1776,N_86);
xnor U3244 (N_3244,N_1008,N_630);
xnor U3245 (N_3245,N_1225,N_1591);
nand U3246 (N_3246,N_1269,N_1340);
xor U3247 (N_3247,N_1279,N_1473);
xor U3248 (N_3248,N_800,N_1900);
nor U3249 (N_3249,N_953,N_634);
xor U3250 (N_3250,N_1509,N_531);
nor U3251 (N_3251,N_662,N_866);
and U3252 (N_3252,N_1592,N_369);
nor U3253 (N_3253,N_977,N_409);
nor U3254 (N_3254,N_1003,N_1335);
nand U3255 (N_3255,N_1990,N_584);
and U3256 (N_3256,N_1097,N_551);
and U3257 (N_3257,N_850,N_1536);
or U3258 (N_3258,N_1185,N_1438);
and U3259 (N_3259,N_1726,N_4);
and U3260 (N_3260,N_255,N_1005);
xor U3261 (N_3261,N_1389,N_1527);
nor U3262 (N_3262,N_706,N_1166);
and U3263 (N_3263,N_1010,N_1755);
nor U3264 (N_3264,N_1675,N_1609);
nor U3265 (N_3265,N_1003,N_1504);
nor U3266 (N_3266,N_274,N_6);
nor U3267 (N_3267,N_1444,N_553);
or U3268 (N_3268,N_408,N_287);
or U3269 (N_3269,N_1798,N_1158);
nor U3270 (N_3270,N_1625,N_1238);
xnor U3271 (N_3271,N_1086,N_1819);
or U3272 (N_3272,N_1576,N_1910);
and U3273 (N_3273,N_62,N_1936);
xor U3274 (N_3274,N_1944,N_1027);
or U3275 (N_3275,N_167,N_3);
xnor U3276 (N_3276,N_1577,N_1807);
nand U3277 (N_3277,N_786,N_1541);
nand U3278 (N_3278,N_1080,N_559);
nand U3279 (N_3279,N_1768,N_1188);
or U3280 (N_3280,N_1923,N_1109);
xor U3281 (N_3281,N_1102,N_891);
xor U3282 (N_3282,N_210,N_297);
xnor U3283 (N_3283,N_558,N_908);
or U3284 (N_3284,N_1830,N_1653);
and U3285 (N_3285,N_1509,N_10);
nor U3286 (N_3286,N_879,N_271);
and U3287 (N_3287,N_551,N_478);
nor U3288 (N_3288,N_87,N_645);
nor U3289 (N_3289,N_127,N_865);
and U3290 (N_3290,N_892,N_12);
nor U3291 (N_3291,N_1103,N_1468);
xor U3292 (N_3292,N_1484,N_126);
or U3293 (N_3293,N_332,N_532);
or U3294 (N_3294,N_758,N_254);
and U3295 (N_3295,N_481,N_143);
xor U3296 (N_3296,N_688,N_1523);
and U3297 (N_3297,N_1698,N_924);
nor U3298 (N_3298,N_110,N_693);
nand U3299 (N_3299,N_1589,N_721);
nand U3300 (N_3300,N_326,N_725);
and U3301 (N_3301,N_885,N_1630);
and U3302 (N_3302,N_1165,N_1446);
nand U3303 (N_3303,N_991,N_793);
and U3304 (N_3304,N_1609,N_576);
and U3305 (N_3305,N_1984,N_547);
or U3306 (N_3306,N_1473,N_1664);
and U3307 (N_3307,N_988,N_752);
and U3308 (N_3308,N_718,N_1622);
and U3309 (N_3309,N_1254,N_498);
nor U3310 (N_3310,N_381,N_1098);
and U3311 (N_3311,N_473,N_1062);
nand U3312 (N_3312,N_1502,N_819);
and U3313 (N_3313,N_1241,N_447);
and U3314 (N_3314,N_1696,N_1953);
or U3315 (N_3315,N_1255,N_1884);
nand U3316 (N_3316,N_1501,N_1367);
and U3317 (N_3317,N_824,N_848);
and U3318 (N_3318,N_1377,N_784);
nand U3319 (N_3319,N_1129,N_137);
xnor U3320 (N_3320,N_1373,N_1568);
and U3321 (N_3321,N_239,N_1353);
and U3322 (N_3322,N_925,N_1754);
nand U3323 (N_3323,N_1368,N_256);
and U3324 (N_3324,N_1299,N_425);
nor U3325 (N_3325,N_239,N_1185);
nand U3326 (N_3326,N_325,N_1008);
or U3327 (N_3327,N_1684,N_1779);
xnor U3328 (N_3328,N_1992,N_685);
nand U3329 (N_3329,N_1609,N_507);
and U3330 (N_3330,N_157,N_1779);
nand U3331 (N_3331,N_725,N_1142);
or U3332 (N_3332,N_1000,N_288);
xor U3333 (N_3333,N_819,N_1686);
and U3334 (N_3334,N_189,N_694);
nor U3335 (N_3335,N_18,N_358);
nor U3336 (N_3336,N_1395,N_1363);
nand U3337 (N_3337,N_1920,N_1999);
and U3338 (N_3338,N_417,N_358);
or U3339 (N_3339,N_943,N_1422);
xor U3340 (N_3340,N_138,N_282);
and U3341 (N_3341,N_637,N_507);
or U3342 (N_3342,N_979,N_917);
or U3343 (N_3343,N_142,N_1054);
nand U3344 (N_3344,N_413,N_1443);
or U3345 (N_3345,N_380,N_975);
nand U3346 (N_3346,N_1597,N_899);
nand U3347 (N_3347,N_606,N_163);
nand U3348 (N_3348,N_773,N_881);
or U3349 (N_3349,N_1549,N_1885);
nand U3350 (N_3350,N_577,N_1044);
nand U3351 (N_3351,N_238,N_1825);
or U3352 (N_3352,N_734,N_1913);
xnor U3353 (N_3353,N_912,N_202);
xnor U3354 (N_3354,N_532,N_156);
nand U3355 (N_3355,N_617,N_193);
and U3356 (N_3356,N_1678,N_1186);
nor U3357 (N_3357,N_808,N_605);
nand U3358 (N_3358,N_214,N_542);
nor U3359 (N_3359,N_1270,N_106);
nand U3360 (N_3360,N_1964,N_361);
or U3361 (N_3361,N_328,N_1314);
nor U3362 (N_3362,N_1491,N_602);
or U3363 (N_3363,N_148,N_1223);
and U3364 (N_3364,N_1931,N_1399);
nand U3365 (N_3365,N_1019,N_730);
and U3366 (N_3366,N_1342,N_369);
or U3367 (N_3367,N_477,N_149);
or U3368 (N_3368,N_895,N_1493);
or U3369 (N_3369,N_1250,N_1798);
and U3370 (N_3370,N_186,N_791);
nand U3371 (N_3371,N_603,N_1275);
or U3372 (N_3372,N_1919,N_1265);
or U3373 (N_3373,N_1843,N_13);
nand U3374 (N_3374,N_653,N_619);
and U3375 (N_3375,N_1623,N_732);
xor U3376 (N_3376,N_1964,N_383);
xor U3377 (N_3377,N_560,N_358);
and U3378 (N_3378,N_1871,N_1266);
and U3379 (N_3379,N_227,N_1699);
nor U3380 (N_3380,N_328,N_938);
xnor U3381 (N_3381,N_316,N_743);
xnor U3382 (N_3382,N_1043,N_758);
nand U3383 (N_3383,N_1979,N_345);
nand U3384 (N_3384,N_1052,N_1763);
nor U3385 (N_3385,N_196,N_1202);
and U3386 (N_3386,N_145,N_1219);
and U3387 (N_3387,N_58,N_435);
nor U3388 (N_3388,N_1649,N_442);
nand U3389 (N_3389,N_378,N_568);
nor U3390 (N_3390,N_875,N_1884);
or U3391 (N_3391,N_1005,N_482);
nor U3392 (N_3392,N_1702,N_523);
nor U3393 (N_3393,N_542,N_959);
or U3394 (N_3394,N_346,N_619);
xor U3395 (N_3395,N_1193,N_698);
nor U3396 (N_3396,N_1842,N_1489);
nor U3397 (N_3397,N_1567,N_920);
or U3398 (N_3398,N_1807,N_850);
or U3399 (N_3399,N_832,N_1826);
and U3400 (N_3400,N_249,N_1791);
or U3401 (N_3401,N_611,N_596);
or U3402 (N_3402,N_241,N_1618);
xor U3403 (N_3403,N_1847,N_413);
nor U3404 (N_3404,N_842,N_1785);
or U3405 (N_3405,N_1760,N_355);
or U3406 (N_3406,N_1022,N_125);
nor U3407 (N_3407,N_1830,N_1750);
nand U3408 (N_3408,N_15,N_678);
xor U3409 (N_3409,N_101,N_261);
nor U3410 (N_3410,N_356,N_975);
xnor U3411 (N_3411,N_651,N_1453);
nor U3412 (N_3412,N_554,N_1156);
nand U3413 (N_3413,N_472,N_397);
xor U3414 (N_3414,N_1527,N_914);
and U3415 (N_3415,N_437,N_1902);
or U3416 (N_3416,N_357,N_742);
and U3417 (N_3417,N_1480,N_1203);
nand U3418 (N_3418,N_1887,N_411);
and U3419 (N_3419,N_281,N_1766);
xor U3420 (N_3420,N_929,N_376);
xnor U3421 (N_3421,N_1868,N_225);
xor U3422 (N_3422,N_487,N_8);
and U3423 (N_3423,N_1069,N_1055);
nor U3424 (N_3424,N_685,N_1051);
or U3425 (N_3425,N_1109,N_1616);
and U3426 (N_3426,N_6,N_1109);
or U3427 (N_3427,N_1625,N_348);
and U3428 (N_3428,N_675,N_1031);
and U3429 (N_3429,N_1911,N_1491);
xnor U3430 (N_3430,N_1292,N_1396);
xor U3431 (N_3431,N_1017,N_56);
xor U3432 (N_3432,N_98,N_335);
nand U3433 (N_3433,N_1565,N_1646);
and U3434 (N_3434,N_1853,N_1327);
or U3435 (N_3435,N_882,N_881);
and U3436 (N_3436,N_301,N_1793);
nand U3437 (N_3437,N_1566,N_354);
nor U3438 (N_3438,N_731,N_1568);
and U3439 (N_3439,N_685,N_1060);
or U3440 (N_3440,N_217,N_1853);
xor U3441 (N_3441,N_317,N_681);
and U3442 (N_3442,N_405,N_1712);
and U3443 (N_3443,N_277,N_292);
nor U3444 (N_3444,N_1959,N_1702);
or U3445 (N_3445,N_184,N_1223);
or U3446 (N_3446,N_90,N_1387);
or U3447 (N_3447,N_853,N_1019);
nor U3448 (N_3448,N_1416,N_238);
xnor U3449 (N_3449,N_1901,N_1952);
and U3450 (N_3450,N_1190,N_1255);
xnor U3451 (N_3451,N_1439,N_1262);
and U3452 (N_3452,N_1682,N_224);
nor U3453 (N_3453,N_1801,N_1396);
or U3454 (N_3454,N_594,N_1319);
nand U3455 (N_3455,N_1305,N_1027);
and U3456 (N_3456,N_1017,N_1447);
and U3457 (N_3457,N_856,N_381);
xnor U3458 (N_3458,N_1920,N_962);
or U3459 (N_3459,N_702,N_1355);
xnor U3460 (N_3460,N_1325,N_541);
xor U3461 (N_3461,N_378,N_1740);
xor U3462 (N_3462,N_776,N_1104);
nand U3463 (N_3463,N_647,N_630);
xnor U3464 (N_3464,N_399,N_189);
xor U3465 (N_3465,N_38,N_1648);
xnor U3466 (N_3466,N_1115,N_1114);
xor U3467 (N_3467,N_1384,N_980);
and U3468 (N_3468,N_351,N_1130);
or U3469 (N_3469,N_1600,N_1624);
xor U3470 (N_3470,N_1220,N_1344);
nor U3471 (N_3471,N_340,N_495);
and U3472 (N_3472,N_484,N_1745);
and U3473 (N_3473,N_1085,N_1218);
nand U3474 (N_3474,N_797,N_1707);
or U3475 (N_3475,N_656,N_1204);
or U3476 (N_3476,N_453,N_1511);
xnor U3477 (N_3477,N_176,N_140);
or U3478 (N_3478,N_388,N_578);
and U3479 (N_3479,N_775,N_776);
and U3480 (N_3480,N_1533,N_342);
nand U3481 (N_3481,N_393,N_572);
or U3482 (N_3482,N_1069,N_621);
and U3483 (N_3483,N_1553,N_1991);
nand U3484 (N_3484,N_1008,N_623);
and U3485 (N_3485,N_540,N_1742);
nor U3486 (N_3486,N_1451,N_1746);
xnor U3487 (N_3487,N_86,N_108);
nand U3488 (N_3488,N_1219,N_725);
nor U3489 (N_3489,N_1374,N_1641);
nor U3490 (N_3490,N_633,N_1225);
xor U3491 (N_3491,N_106,N_622);
and U3492 (N_3492,N_1071,N_328);
xor U3493 (N_3493,N_295,N_1465);
xor U3494 (N_3494,N_865,N_969);
or U3495 (N_3495,N_108,N_1443);
or U3496 (N_3496,N_1544,N_1274);
xor U3497 (N_3497,N_761,N_1978);
nor U3498 (N_3498,N_119,N_782);
nand U3499 (N_3499,N_1929,N_171);
nand U3500 (N_3500,N_1503,N_1398);
xnor U3501 (N_3501,N_576,N_786);
nor U3502 (N_3502,N_1167,N_861);
nor U3503 (N_3503,N_1121,N_273);
nand U3504 (N_3504,N_1214,N_851);
and U3505 (N_3505,N_813,N_1813);
nand U3506 (N_3506,N_711,N_288);
and U3507 (N_3507,N_627,N_1535);
xor U3508 (N_3508,N_1793,N_1048);
and U3509 (N_3509,N_1582,N_1745);
nor U3510 (N_3510,N_1504,N_927);
or U3511 (N_3511,N_1482,N_1540);
or U3512 (N_3512,N_95,N_1754);
and U3513 (N_3513,N_750,N_440);
nor U3514 (N_3514,N_1231,N_1644);
nor U3515 (N_3515,N_1283,N_417);
and U3516 (N_3516,N_1309,N_293);
nand U3517 (N_3517,N_1102,N_1734);
and U3518 (N_3518,N_238,N_471);
nand U3519 (N_3519,N_258,N_869);
nor U3520 (N_3520,N_72,N_40);
or U3521 (N_3521,N_176,N_1882);
nor U3522 (N_3522,N_560,N_234);
or U3523 (N_3523,N_925,N_1419);
nor U3524 (N_3524,N_155,N_535);
xor U3525 (N_3525,N_1196,N_1624);
xnor U3526 (N_3526,N_1850,N_289);
or U3527 (N_3527,N_1571,N_889);
and U3528 (N_3528,N_1543,N_1702);
or U3529 (N_3529,N_391,N_133);
and U3530 (N_3530,N_806,N_173);
nor U3531 (N_3531,N_1263,N_1044);
xnor U3532 (N_3532,N_1817,N_1154);
and U3533 (N_3533,N_1693,N_1162);
and U3534 (N_3534,N_144,N_855);
or U3535 (N_3535,N_1333,N_1503);
nor U3536 (N_3536,N_65,N_71);
xor U3537 (N_3537,N_1673,N_762);
and U3538 (N_3538,N_580,N_1119);
nand U3539 (N_3539,N_1969,N_1682);
nor U3540 (N_3540,N_1429,N_1914);
nor U3541 (N_3541,N_1134,N_1004);
xnor U3542 (N_3542,N_927,N_1852);
nor U3543 (N_3543,N_1253,N_1869);
or U3544 (N_3544,N_462,N_63);
and U3545 (N_3545,N_567,N_1079);
nand U3546 (N_3546,N_1721,N_1141);
and U3547 (N_3547,N_848,N_770);
nand U3548 (N_3548,N_85,N_131);
xnor U3549 (N_3549,N_1810,N_1483);
nor U3550 (N_3550,N_697,N_1299);
xor U3551 (N_3551,N_1350,N_1522);
xor U3552 (N_3552,N_1977,N_1032);
and U3553 (N_3553,N_1090,N_778);
or U3554 (N_3554,N_1381,N_195);
nand U3555 (N_3555,N_1386,N_990);
or U3556 (N_3556,N_1884,N_295);
nor U3557 (N_3557,N_1083,N_1298);
nand U3558 (N_3558,N_885,N_234);
and U3559 (N_3559,N_474,N_32);
and U3560 (N_3560,N_1255,N_1297);
xnor U3561 (N_3561,N_476,N_1628);
or U3562 (N_3562,N_525,N_1570);
nor U3563 (N_3563,N_507,N_1378);
nor U3564 (N_3564,N_288,N_590);
nand U3565 (N_3565,N_1098,N_613);
and U3566 (N_3566,N_1780,N_422);
nor U3567 (N_3567,N_54,N_1343);
xor U3568 (N_3568,N_1532,N_244);
xnor U3569 (N_3569,N_1894,N_1045);
or U3570 (N_3570,N_156,N_30);
nor U3571 (N_3571,N_1316,N_198);
and U3572 (N_3572,N_1615,N_663);
or U3573 (N_3573,N_815,N_597);
and U3574 (N_3574,N_74,N_695);
or U3575 (N_3575,N_1574,N_1444);
xnor U3576 (N_3576,N_1986,N_1056);
nor U3577 (N_3577,N_1454,N_1643);
or U3578 (N_3578,N_157,N_1000);
xnor U3579 (N_3579,N_639,N_737);
nand U3580 (N_3580,N_1806,N_558);
nand U3581 (N_3581,N_1463,N_1588);
nand U3582 (N_3582,N_559,N_689);
and U3583 (N_3583,N_850,N_1079);
or U3584 (N_3584,N_1728,N_1951);
nand U3585 (N_3585,N_608,N_125);
or U3586 (N_3586,N_468,N_152);
nor U3587 (N_3587,N_780,N_308);
nor U3588 (N_3588,N_1557,N_724);
nor U3589 (N_3589,N_408,N_52);
and U3590 (N_3590,N_1927,N_379);
or U3591 (N_3591,N_1986,N_963);
or U3592 (N_3592,N_253,N_1922);
nand U3593 (N_3593,N_1049,N_634);
nand U3594 (N_3594,N_918,N_1762);
and U3595 (N_3595,N_1679,N_1757);
and U3596 (N_3596,N_1528,N_1221);
and U3597 (N_3597,N_40,N_1310);
xnor U3598 (N_3598,N_1871,N_1077);
or U3599 (N_3599,N_1161,N_966);
nor U3600 (N_3600,N_731,N_62);
nand U3601 (N_3601,N_617,N_75);
or U3602 (N_3602,N_1034,N_325);
and U3603 (N_3603,N_1990,N_1326);
or U3604 (N_3604,N_1265,N_879);
nor U3605 (N_3605,N_1696,N_1353);
nand U3606 (N_3606,N_1128,N_1622);
or U3607 (N_3607,N_259,N_196);
and U3608 (N_3608,N_185,N_1249);
or U3609 (N_3609,N_1537,N_1874);
nand U3610 (N_3610,N_1364,N_739);
nor U3611 (N_3611,N_1731,N_280);
nor U3612 (N_3612,N_935,N_1754);
nor U3613 (N_3613,N_1952,N_1896);
xor U3614 (N_3614,N_9,N_1102);
nor U3615 (N_3615,N_689,N_1537);
and U3616 (N_3616,N_28,N_411);
xnor U3617 (N_3617,N_1651,N_940);
nand U3618 (N_3618,N_72,N_1957);
xnor U3619 (N_3619,N_914,N_437);
or U3620 (N_3620,N_462,N_852);
nand U3621 (N_3621,N_488,N_740);
or U3622 (N_3622,N_1631,N_914);
and U3623 (N_3623,N_1119,N_1658);
and U3624 (N_3624,N_1553,N_491);
or U3625 (N_3625,N_1042,N_449);
nand U3626 (N_3626,N_1036,N_1776);
or U3627 (N_3627,N_1338,N_566);
nor U3628 (N_3628,N_82,N_1522);
and U3629 (N_3629,N_987,N_183);
or U3630 (N_3630,N_1181,N_1752);
and U3631 (N_3631,N_196,N_515);
or U3632 (N_3632,N_1457,N_987);
and U3633 (N_3633,N_471,N_1811);
nand U3634 (N_3634,N_1520,N_880);
and U3635 (N_3635,N_1904,N_714);
xor U3636 (N_3636,N_1793,N_847);
nor U3637 (N_3637,N_1724,N_66);
nor U3638 (N_3638,N_1032,N_1434);
nand U3639 (N_3639,N_764,N_1009);
xor U3640 (N_3640,N_1667,N_1623);
nor U3641 (N_3641,N_1223,N_527);
nand U3642 (N_3642,N_1877,N_1347);
and U3643 (N_3643,N_1847,N_730);
nor U3644 (N_3644,N_829,N_1212);
nand U3645 (N_3645,N_545,N_1731);
or U3646 (N_3646,N_270,N_1059);
or U3647 (N_3647,N_1533,N_284);
or U3648 (N_3648,N_167,N_1910);
or U3649 (N_3649,N_1908,N_619);
xnor U3650 (N_3650,N_735,N_1021);
and U3651 (N_3651,N_1119,N_1129);
and U3652 (N_3652,N_1710,N_793);
and U3653 (N_3653,N_1820,N_1533);
and U3654 (N_3654,N_1432,N_626);
xnor U3655 (N_3655,N_230,N_1543);
xnor U3656 (N_3656,N_468,N_672);
and U3657 (N_3657,N_144,N_62);
xnor U3658 (N_3658,N_1201,N_548);
nand U3659 (N_3659,N_430,N_1386);
xnor U3660 (N_3660,N_855,N_393);
nor U3661 (N_3661,N_199,N_1997);
xor U3662 (N_3662,N_1367,N_1242);
or U3663 (N_3663,N_392,N_1689);
nand U3664 (N_3664,N_1156,N_50);
or U3665 (N_3665,N_1000,N_1056);
nand U3666 (N_3666,N_1002,N_467);
nand U3667 (N_3667,N_1664,N_1489);
xnor U3668 (N_3668,N_270,N_1455);
and U3669 (N_3669,N_1915,N_50);
nand U3670 (N_3670,N_362,N_253);
and U3671 (N_3671,N_1628,N_221);
nor U3672 (N_3672,N_171,N_46);
nor U3673 (N_3673,N_192,N_155);
nand U3674 (N_3674,N_1615,N_1899);
and U3675 (N_3675,N_693,N_550);
nand U3676 (N_3676,N_1985,N_509);
xor U3677 (N_3677,N_377,N_1175);
and U3678 (N_3678,N_1040,N_666);
nand U3679 (N_3679,N_1689,N_60);
nor U3680 (N_3680,N_1814,N_1974);
xnor U3681 (N_3681,N_1686,N_1133);
and U3682 (N_3682,N_1543,N_514);
or U3683 (N_3683,N_1925,N_182);
nor U3684 (N_3684,N_1160,N_1021);
xnor U3685 (N_3685,N_735,N_933);
nor U3686 (N_3686,N_912,N_1888);
and U3687 (N_3687,N_250,N_1452);
and U3688 (N_3688,N_1154,N_62);
nand U3689 (N_3689,N_136,N_325);
xor U3690 (N_3690,N_779,N_818);
nand U3691 (N_3691,N_196,N_1500);
nor U3692 (N_3692,N_1562,N_940);
or U3693 (N_3693,N_1702,N_273);
or U3694 (N_3694,N_1323,N_1692);
or U3695 (N_3695,N_1607,N_1744);
or U3696 (N_3696,N_1150,N_1164);
and U3697 (N_3697,N_984,N_1361);
nor U3698 (N_3698,N_1841,N_653);
and U3699 (N_3699,N_238,N_338);
and U3700 (N_3700,N_99,N_1206);
nor U3701 (N_3701,N_765,N_942);
nand U3702 (N_3702,N_1809,N_1531);
xor U3703 (N_3703,N_425,N_1550);
and U3704 (N_3704,N_1151,N_479);
and U3705 (N_3705,N_472,N_1980);
or U3706 (N_3706,N_259,N_1002);
nor U3707 (N_3707,N_1611,N_471);
nor U3708 (N_3708,N_1451,N_1720);
nand U3709 (N_3709,N_547,N_1657);
nor U3710 (N_3710,N_542,N_905);
or U3711 (N_3711,N_54,N_708);
xor U3712 (N_3712,N_1360,N_27);
nand U3713 (N_3713,N_464,N_770);
or U3714 (N_3714,N_1464,N_1842);
nand U3715 (N_3715,N_1422,N_1500);
and U3716 (N_3716,N_1179,N_1845);
xor U3717 (N_3717,N_834,N_1358);
nand U3718 (N_3718,N_1098,N_1185);
or U3719 (N_3719,N_291,N_132);
nand U3720 (N_3720,N_1503,N_40);
and U3721 (N_3721,N_1918,N_66);
nand U3722 (N_3722,N_183,N_40);
xor U3723 (N_3723,N_705,N_1683);
and U3724 (N_3724,N_1068,N_1720);
xor U3725 (N_3725,N_324,N_524);
nor U3726 (N_3726,N_521,N_1666);
and U3727 (N_3727,N_1796,N_1402);
and U3728 (N_3728,N_1886,N_562);
or U3729 (N_3729,N_1582,N_1796);
or U3730 (N_3730,N_1465,N_1621);
or U3731 (N_3731,N_1738,N_1216);
and U3732 (N_3732,N_1489,N_1336);
xnor U3733 (N_3733,N_331,N_851);
nor U3734 (N_3734,N_1079,N_939);
nand U3735 (N_3735,N_1801,N_1694);
nand U3736 (N_3736,N_1871,N_1176);
and U3737 (N_3737,N_883,N_1036);
nand U3738 (N_3738,N_765,N_749);
xor U3739 (N_3739,N_705,N_1122);
or U3740 (N_3740,N_400,N_592);
and U3741 (N_3741,N_1394,N_1074);
or U3742 (N_3742,N_1365,N_1183);
nor U3743 (N_3743,N_1884,N_13);
or U3744 (N_3744,N_1026,N_1882);
nor U3745 (N_3745,N_889,N_1779);
xor U3746 (N_3746,N_708,N_1518);
or U3747 (N_3747,N_249,N_889);
and U3748 (N_3748,N_452,N_756);
or U3749 (N_3749,N_1273,N_815);
and U3750 (N_3750,N_1763,N_1037);
and U3751 (N_3751,N_756,N_284);
and U3752 (N_3752,N_630,N_961);
and U3753 (N_3753,N_1375,N_767);
and U3754 (N_3754,N_1108,N_77);
xnor U3755 (N_3755,N_1999,N_345);
nor U3756 (N_3756,N_1666,N_1733);
or U3757 (N_3757,N_1185,N_1670);
xnor U3758 (N_3758,N_956,N_1763);
nand U3759 (N_3759,N_1120,N_1088);
nand U3760 (N_3760,N_693,N_1597);
xnor U3761 (N_3761,N_439,N_30);
or U3762 (N_3762,N_862,N_1675);
and U3763 (N_3763,N_1502,N_239);
and U3764 (N_3764,N_1154,N_1570);
and U3765 (N_3765,N_1055,N_417);
nor U3766 (N_3766,N_1169,N_319);
nor U3767 (N_3767,N_1260,N_1545);
or U3768 (N_3768,N_1846,N_1614);
nor U3769 (N_3769,N_1341,N_748);
and U3770 (N_3770,N_1157,N_1001);
nor U3771 (N_3771,N_796,N_1684);
or U3772 (N_3772,N_1367,N_445);
nor U3773 (N_3773,N_6,N_1309);
nor U3774 (N_3774,N_1495,N_1753);
nor U3775 (N_3775,N_1305,N_423);
or U3776 (N_3776,N_141,N_1087);
and U3777 (N_3777,N_1770,N_904);
nor U3778 (N_3778,N_641,N_1748);
nand U3779 (N_3779,N_156,N_1948);
nor U3780 (N_3780,N_1745,N_297);
nand U3781 (N_3781,N_1390,N_1515);
xor U3782 (N_3782,N_805,N_212);
nor U3783 (N_3783,N_1128,N_891);
xor U3784 (N_3784,N_1615,N_1928);
or U3785 (N_3785,N_1040,N_1896);
and U3786 (N_3786,N_406,N_834);
nand U3787 (N_3787,N_688,N_1422);
xor U3788 (N_3788,N_1758,N_1301);
xnor U3789 (N_3789,N_1463,N_1524);
nand U3790 (N_3790,N_390,N_1979);
nand U3791 (N_3791,N_1404,N_1698);
nor U3792 (N_3792,N_708,N_83);
xnor U3793 (N_3793,N_82,N_1099);
and U3794 (N_3794,N_1318,N_575);
and U3795 (N_3795,N_352,N_1048);
nor U3796 (N_3796,N_1181,N_101);
xor U3797 (N_3797,N_369,N_871);
nor U3798 (N_3798,N_416,N_1464);
nand U3799 (N_3799,N_948,N_1133);
and U3800 (N_3800,N_1648,N_180);
or U3801 (N_3801,N_281,N_483);
xor U3802 (N_3802,N_1361,N_1880);
and U3803 (N_3803,N_777,N_687);
nand U3804 (N_3804,N_1383,N_137);
nand U3805 (N_3805,N_362,N_1179);
nand U3806 (N_3806,N_305,N_1892);
and U3807 (N_3807,N_166,N_1102);
nand U3808 (N_3808,N_42,N_1542);
nor U3809 (N_3809,N_1912,N_48);
nand U3810 (N_3810,N_5,N_1084);
nand U3811 (N_3811,N_428,N_36);
xor U3812 (N_3812,N_610,N_256);
nand U3813 (N_3813,N_772,N_1530);
or U3814 (N_3814,N_805,N_418);
xor U3815 (N_3815,N_1237,N_1964);
xor U3816 (N_3816,N_853,N_87);
xnor U3817 (N_3817,N_1710,N_1844);
xor U3818 (N_3818,N_1316,N_896);
or U3819 (N_3819,N_1607,N_1806);
xor U3820 (N_3820,N_1632,N_584);
and U3821 (N_3821,N_4,N_709);
xor U3822 (N_3822,N_1779,N_689);
nand U3823 (N_3823,N_1183,N_24);
xor U3824 (N_3824,N_1719,N_582);
nand U3825 (N_3825,N_1548,N_486);
or U3826 (N_3826,N_372,N_227);
xnor U3827 (N_3827,N_1737,N_579);
nor U3828 (N_3828,N_65,N_532);
nand U3829 (N_3829,N_1308,N_1225);
xor U3830 (N_3830,N_172,N_606);
xor U3831 (N_3831,N_1772,N_687);
nand U3832 (N_3832,N_1946,N_1781);
xnor U3833 (N_3833,N_868,N_488);
and U3834 (N_3834,N_1156,N_1605);
and U3835 (N_3835,N_1301,N_1490);
xor U3836 (N_3836,N_114,N_253);
or U3837 (N_3837,N_1925,N_209);
nor U3838 (N_3838,N_36,N_1965);
or U3839 (N_3839,N_1164,N_1274);
nor U3840 (N_3840,N_615,N_837);
xor U3841 (N_3841,N_221,N_1957);
nand U3842 (N_3842,N_1682,N_763);
or U3843 (N_3843,N_1672,N_1494);
nor U3844 (N_3844,N_378,N_667);
xor U3845 (N_3845,N_1292,N_724);
nor U3846 (N_3846,N_723,N_1734);
and U3847 (N_3847,N_1183,N_1547);
xor U3848 (N_3848,N_1265,N_1025);
xnor U3849 (N_3849,N_354,N_1695);
and U3850 (N_3850,N_1461,N_1537);
or U3851 (N_3851,N_1824,N_1270);
nand U3852 (N_3852,N_1089,N_1597);
xnor U3853 (N_3853,N_160,N_339);
nand U3854 (N_3854,N_14,N_691);
or U3855 (N_3855,N_1011,N_1836);
xnor U3856 (N_3856,N_282,N_1542);
xnor U3857 (N_3857,N_1515,N_1805);
or U3858 (N_3858,N_1413,N_1410);
xnor U3859 (N_3859,N_872,N_438);
xor U3860 (N_3860,N_622,N_872);
nand U3861 (N_3861,N_733,N_774);
xor U3862 (N_3862,N_98,N_1535);
and U3863 (N_3863,N_1890,N_1439);
and U3864 (N_3864,N_1802,N_401);
nor U3865 (N_3865,N_1196,N_1929);
and U3866 (N_3866,N_1096,N_1670);
nand U3867 (N_3867,N_475,N_1185);
nor U3868 (N_3868,N_1777,N_992);
xor U3869 (N_3869,N_1355,N_115);
nor U3870 (N_3870,N_1948,N_1349);
xnor U3871 (N_3871,N_1837,N_951);
xnor U3872 (N_3872,N_798,N_1115);
and U3873 (N_3873,N_1852,N_706);
nand U3874 (N_3874,N_1842,N_43);
nand U3875 (N_3875,N_877,N_846);
and U3876 (N_3876,N_614,N_801);
and U3877 (N_3877,N_1021,N_1192);
xnor U3878 (N_3878,N_190,N_294);
or U3879 (N_3879,N_1890,N_863);
and U3880 (N_3880,N_1878,N_1311);
and U3881 (N_3881,N_570,N_822);
or U3882 (N_3882,N_1887,N_1084);
nand U3883 (N_3883,N_1933,N_842);
and U3884 (N_3884,N_1439,N_1968);
and U3885 (N_3885,N_1618,N_1711);
xnor U3886 (N_3886,N_103,N_559);
and U3887 (N_3887,N_98,N_940);
and U3888 (N_3888,N_1319,N_244);
xnor U3889 (N_3889,N_1666,N_1363);
nand U3890 (N_3890,N_612,N_1815);
nor U3891 (N_3891,N_779,N_1728);
and U3892 (N_3892,N_1869,N_1630);
or U3893 (N_3893,N_518,N_924);
and U3894 (N_3894,N_1720,N_157);
nor U3895 (N_3895,N_525,N_1124);
nor U3896 (N_3896,N_1951,N_1564);
nand U3897 (N_3897,N_488,N_865);
and U3898 (N_3898,N_425,N_146);
or U3899 (N_3899,N_1537,N_1335);
or U3900 (N_3900,N_1645,N_110);
or U3901 (N_3901,N_1994,N_240);
xor U3902 (N_3902,N_587,N_242);
or U3903 (N_3903,N_8,N_681);
or U3904 (N_3904,N_1502,N_203);
nor U3905 (N_3905,N_363,N_404);
or U3906 (N_3906,N_25,N_361);
or U3907 (N_3907,N_1516,N_39);
nand U3908 (N_3908,N_1553,N_1998);
nor U3909 (N_3909,N_1300,N_585);
nor U3910 (N_3910,N_462,N_1722);
nand U3911 (N_3911,N_1776,N_45);
nor U3912 (N_3912,N_1020,N_1601);
nand U3913 (N_3913,N_1579,N_70);
and U3914 (N_3914,N_1115,N_1630);
nand U3915 (N_3915,N_1994,N_650);
nand U3916 (N_3916,N_795,N_129);
and U3917 (N_3917,N_300,N_984);
xnor U3918 (N_3918,N_1310,N_779);
xor U3919 (N_3919,N_294,N_33);
xnor U3920 (N_3920,N_1735,N_1928);
or U3921 (N_3921,N_225,N_1908);
nand U3922 (N_3922,N_1094,N_317);
nor U3923 (N_3923,N_38,N_1319);
and U3924 (N_3924,N_493,N_272);
or U3925 (N_3925,N_383,N_1662);
and U3926 (N_3926,N_39,N_865);
nand U3927 (N_3927,N_1234,N_1827);
xnor U3928 (N_3928,N_1656,N_536);
and U3929 (N_3929,N_1353,N_1475);
and U3930 (N_3930,N_1881,N_1925);
nor U3931 (N_3931,N_1213,N_1084);
nor U3932 (N_3932,N_408,N_1752);
nand U3933 (N_3933,N_668,N_275);
or U3934 (N_3934,N_1287,N_160);
nand U3935 (N_3935,N_1514,N_1200);
xor U3936 (N_3936,N_758,N_688);
and U3937 (N_3937,N_264,N_931);
and U3938 (N_3938,N_745,N_1904);
nor U3939 (N_3939,N_1149,N_1868);
or U3940 (N_3940,N_1058,N_1502);
or U3941 (N_3941,N_846,N_408);
nor U3942 (N_3942,N_65,N_1423);
and U3943 (N_3943,N_1127,N_1837);
nand U3944 (N_3944,N_488,N_145);
nor U3945 (N_3945,N_831,N_1303);
xnor U3946 (N_3946,N_265,N_1863);
xor U3947 (N_3947,N_487,N_110);
xnor U3948 (N_3948,N_1266,N_1573);
nor U3949 (N_3949,N_1427,N_1929);
and U3950 (N_3950,N_135,N_1432);
and U3951 (N_3951,N_1847,N_897);
or U3952 (N_3952,N_204,N_374);
and U3953 (N_3953,N_1480,N_71);
xor U3954 (N_3954,N_524,N_1427);
xor U3955 (N_3955,N_1905,N_1283);
nor U3956 (N_3956,N_251,N_16);
nor U3957 (N_3957,N_1208,N_1030);
and U3958 (N_3958,N_992,N_908);
nor U3959 (N_3959,N_1120,N_401);
xor U3960 (N_3960,N_10,N_1773);
nand U3961 (N_3961,N_778,N_1360);
nand U3962 (N_3962,N_1014,N_1776);
and U3963 (N_3963,N_1061,N_1226);
xor U3964 (N_3964,N_1551,N_1176);
nor U3965 (N_3965,N_1304,N_1859);
and U3966 (N_3966,N_137,N_1201);
nand U3967 (N_3967,N_198,N_293);
xnor U3968 (N_3968,N_652,N_508);
xnor U3969 (N_3969,N_1603,N_1822);
nand U3970 (N_3970,N_1491,N_1385);
xor U3971 (N_3971,N_611,N_1553);
or U3972 (N_3972,N_599,N_269);
or U3973 (N_3973,N_1988,N_1770);
or U3974 (N_3974,N_1408,N_246);
nor U3975 (N_3975,N_1769,N_1309);
and U3976 (N_3976,N_1916,N_220);
or U3977 (N_3977,N_487,N_1896);
or U3978 (N_3978,N_63,N_156);
nor U3979 (N_3979,N_1707,N_1754);
nor U3980 (N_3980,N_750,N_189);
xnor U3981 (N_3981,N_88,N_1460);
and U3982 (N_3982,N_1170,N_1860);
xor U3983 (N_3983,N_223,N_1033);
nand U3984 (N_3984,N_311,N_1138);
and U3985 (N_3985,N_243,N_394);
or U3986 (N_3986,N_576,N_549);
nor U3987 (N_3987,N_1460,N_319);
nand U3988 (N_3988,N_339,N_174);
xor U3989 (N_3989,N_1188,N_865);
or U3990 (N_3990,N_1209,N_71);
nor U3991 (N_3991,N_902,N_1871);
nor U3992 (N_3992,N_1898,N_1284);
or U3993 (N_3993,N_1496,N_170);
xnor U3994 (N_3994,N_124,N_467);
and U3995 (N_3995,N_1631,N_1562);
and U3996 (N_3996,N_708,N_1460);
nor U3997 (N_3997,N_991,N_1162);
nor U3998 (N_3998,N_1400,N_907);
and U3999 (N_3999,N_1905,N_335);
nand U4000 (N_4000,N_3593,N_2426);
and U4001 (N_4001,N_2531,N_3078);
xor U4002 (N_4002,N_3004,N_3308);
xnor U4003 (N_4003,N_2510,N_2691);
nor U4004 (N_4004,N_2568,N_3226);
xnor U4005 (N_4005,N_2590,N_3755);
or U4006 (N_4006,N_3095,N_2847);
nor U4007 (N_4007,N_3685,N_3702);
and U4008 (N_4008,N_3426,N_3703);
or U4009 (N_4009,N_3201,N_3911);
and U4010 (N_4010,N_2836,N_3990);
nor U4011 (N_4011,N_2898,N_2697);
xnor U4012 (N_4012,N_3175,N_3814);
xnor U4013 (N_4013,N_3794,N_2630);
and U4014 (N_4014,N_3622,N_2550);
nand U4015 (N_4015,N_3745,N_3013);
nand U4016 (N_4016,N_2149,N_3379);
and U4017 (N_4017,N_2798,N_2631);
or U4018 (N_4018,N_3744,N_3443);
nand U4019 (N_4019,N_3097,N_2946);
nand U4020 (N_4020,N_3938,N_2218);
and U4021 (N_4021,N_3139,N_3200);
nor U4022 (N_4022,N_3536,N_3061);
or U4023 (N_4023,N_3040,N_3287);
or U4024 (N_4024,N_2230,N_3583);
or U4025 (N_4025,N_3157,N_2919);
nor U4026 (N_4026,N_2984,N_2301);
nand U4027 (N_4027,N_2615,N_3594);
and U4028 (N_4028,N_3706,N_2057);
and U4029 (N_4029,N_2471,N_2541);
or U4030 (N_4030,N_3230,N_3587);
or U4031 (N_4031,N_3043,N_2011);
xor U4032 (N_4032,N_2704,N_2022);
xor U4033 (N_4033,N_2746,N_2809);
or U4034 (N_4034,N_3380,N_2566);
or U4035 (N_4035,N_3510,N_2019);
xnor U4036 (N_4036,N_2887,N_2014);
xor U4037 (N_4037,N_3974,N_3055);
nor U4038 (N_4038,N_2720,N_2868);
or U4039 (N_4039,N_3016,N_2570);
nand U4040 (N_4040,N_2270,N_2466);
or U4041 (N_4041,N_2760,N_2128);
nor U4042 (N_4042,N_2757,N_2613);
xnor U4043 (N_4043,N_2796,N_3083);
nand U4044 (N_4044,N_3590,N_2652);
or U4045 (N_4045,N_2601,N_2488);
nand U4046 (N_4046,N_2237,N_2944);
xor U4047 (N_4047,N_2647,N_2724);
or U4048 (N_4048,N_2422,N_2533);
and U4049 (N_4049,N_2393,N_2512);
or U4050 (N_4050,N_3614,N_3207);
xor U4051 (N_4051,N_2045,N_2207);
nand U4052 (N_4052,N_2988,N_2794);
nand U4053 (N_4053,N_3035,N_2286);
or U4054 (N_4054,N_3119,N_3565);
or U4055 (N_4055,N_2320,N_3262);
nor U4056 (N_4056,N_3798,N_2227);
nor U4057 (N_4057,N_2986,N_2171);
and U4058 (N_4058,N_3680,N_2279);
nand U4059 (N_4059,N_3978,N_2950);
nor U4060 (N_4060,N_3983,N_2034);
or U4061 (N_4061,N_3563,N_2161);
xor U4062 (N_4062,N_3627,N_2349);
xor U4063 (N_4063,N_3714,N_2818);
nor U4064 (N_4064,N_3481,N_3842);
nand U4065 (N_4065,N_3967,N_2596);
and U4066 (N_4066,N_3792,N_2053);
nand U4067 (N_4067,N_3874,N_3867);
xnor U4068 (N_4068,N_3750,N_2068);
and U4069 (N_4069,N_3721,N_3224);
xnor U4070 (N_4070,N_2852,N_2973);
and U4071 (N_4071,N_3900,N_3446);
nor U4072 (N_4072,N_2626,N_3447);
nor U4073 (N_4073,N_3917,N_3309);
nand U4074 (N_4074,N_2772,N_2485);
or U4075 (N_4075,N_3353,N_3726);
nand U4076 (N_4076,N_3385,N_3599);
nand U4077 (N_4077,N_3766,N_2363);
xnor U4078 (N_4078,N_2591,N_3021);
and U4079 (N_4079,N_2247,N_3144);
or U4080 (N_4080,N_2957,N_3321);
nor U4081 (N_4081,N_3828,N_3610);
nand U4082 (N_4082,N_3646,N_2658);
or U4083 (N_4083,N_3668,N_2403);
nand U4084 (N_4084,N_3752,N_3600);
xnor U4085 (N_4085,N_3860,N_2650);
and U4086 (N_4086,N_2383,N_2390);
nand U4087 (N_4087,N_3241,N_2565);
nand U4088 (N_4088,N_2273,N_3341);
xnor U4089 (N_4089,N_3955,N_3242);
xnor U4090 (N_4090,N_2535,N_2681);
nor U4091 (N_4091,N_3550,N_3468);
xor U4092 (N_4092,N_2049,N_2028);
and U4093 (N_4093,N_3534,N_3538);
and U4094 (N_4094,N_3048,N_2718);
xor U4095 (N_4095,N_2035,N_3044);
and U4096 (N_4096,N_3577,N_3081);
nand U4097 (N_4097,N_2188,N_3107);
nand U4098 (N_4098,N_2085,N_3249);
or U4099 (N_4099,N_2197,N_2127);
xor U4100 (N_4100,N_2972,N_2961);
and U4101 (N_4101,N_3425,N_2835);
nand U4102 (N_4102,N_2705,N_2318);
xnor U4103 (N_4103,N_2117,N_3179);
nand U4104 (N_4104,N_3694,N_3085);
or U4105 (N_4105,N_2220,N_3756);
or U4106 (N_4106,N_3265,N_3025);
nand U4107 (N_4107,N_2747,N_2929);
or U4108 (N_4108,N_3018,N_3225);
xnor U4109 (N_4109,N_3027,N_3497);
or U4110 (N_4110,N_3776,N_3960);
xor U4111 (N_4111,N_2826,N_2181);
and U4112 (N_4112,N_2966,N_3498);
and U4113 (N_4113,N_3011,N_3188);
xnor U4114 (N_4114,N_3979,N_2699);
xor U4115 (N_4115,N_2905,N_2648);
and U4116 (N_4116,N_2058,N_2820);
nand U4117 (N_4117,N_2076,N_2250);
and U4118 (N_4118,N_3396,N_3592);
xor U4119 (N_4119,N_3686,N_3164);
or U4120 (N_4120,N_3029,N_3476);
or U4121 (N_4121,N_3381,N_3108);
nand U4122 (N_4122,N_3524,N_3864);
and U4123 (N_4123,N_3930,N_2176);
xor U4124 (N_4124,N_3958,N_2569);
xnor U4125 (N_4125,N_3961,N_3933);
and U4126 (N_4126,N_2465,N_3305);
nor U4127 (N_4127,N_2433,N_2925);
or U4128 (N_4128,N_3749,N_2748);
and U4129 (N_4129,N_2000,N_2890);
xnor U4130 (N_4130,N_2519,N_3104);
nand U4131 (N_4131,N_3395,N_2116);
nor U4132 (N_4132,N_2345,N_2906);
nand U4133 (N_4133,N_2862,N_3725);
nor U4134 (N_4134,N_3724,N_2195);
and U4135 (N_4135,N_3219,N_2567);
nand U4136 (N_4136,N_2791,N_2480);
nand U4137 (N_4137,N_3068,N_3542);
nor U4138 (N_4138,N_3333,N_2878);
xnor U4139 (N_4139,N_2805,N_2981);
or U4140 (N_4140,N_2606,N_2725);
nand U4141 (N_4141,N_2959,N_2146);
or U4142 (N_4142,N_3269,N_2937);
nand U4143 (N_4143,N_3937,N_3332);
and U4144 (N_4144,N_2416,N_2498);
and U4145 (N_4145,N_3009,N_2499);
nor U4146 (N_4146,N_3282,N_2871);
nor U4147 (N_4147,N_3457,N_2003);
nand U4148 (N_4148,N_3898,N_2579);
nand U4149 (N_4149,N_3343,N_3875);
nor U4150 (N_4150,N_2192,N_2268);
and U4151 (N_4151,N_3169,N_2120);
nand U4152 (N_4152,N_2990,N_2577);
or U4153 (N_4153,N_2995,N_3189);
and U4154 (N_4154,N_2013,N_3963);
xnor U4155 (N_4155,N_2478,N_2209);
nand U4156 (N_4156,N_3066,N_2417);
or U4157 (N_4157,N_2254,N_3045);
nand U4158 (N_4158,N_2656,N_2398);
xor U4159 (N_4159,N_3031,N_2894);
nand U4160 (N_4160,N_2696,N_2684);
nor U4161 (N_4161,N_3196,N_3290);
nor U4162 (N_4162,N_3185,N_3336);
or U4163 (N_4163,N_2501,N_2353);
nand U4164 (N_4164,N_3549,N_3383);
or U4165 (N_4165,N_2583,N_3277);
xnor U4166 (N_4166,N_3485,N_2113);
or U4167 (N_4167,N_2924,N_3530);
xnor U4168 (N_4168,N_3223,N_3783);
or U4169 (N_4169,N_3998,N_2184);
and U4170 (N_4170,N_3178,N_2534);
and U4171 (N_4171,N_3802,N_3500);
or U4172 (N_4172,N_2712,N_2439);
or U4173 (N_4173,N_2634,N_3063);
nor U4174 (N_4174,N_3453,N_2226);
nor U4175 (N_4175,N_2991,N_2710);
nand U4176 (N_4176,N_2344,N_3484);
or U4177 (N_4177,N_2071,N_2105);
and U4178 (N_4178,N_2559,N_3301);
or U4179 (N_4179,N_2319,N_3032);
nor U4180 (N_4180,N_3964,N_2284);
nor U4181 (N_4181,N_3171,N_3826);
or U4182 (N_4182,N_3886,N_2706);
or U4183 (N_4183,N_3366,N_3382);
nor U4184 (N_4184,N_3950,N_3663);
or U4185 (N_4185,N_2743,N_3758);
nand U4186 (N_4186,N_3653,N_3094);
nor U4187 (N_4187,N_2043,N_2915);
and U4188 (N_4188,N_3909,N_3193);
and U4189 (N_4189,N_2661,N_3098);
nor U4190 (N_4190,N_3719,N_3077);
or U4191 (N_4191,N_3138,N_3401);
and U4192 (N_4192,N_3252,N_3625);
nand U4193 (N_4193,N_3556,N_3390);
xor U4194 (N_4194,N_3279,N_3050);
nor U4195 (N_4195,N_2702,N_2208);
xnor U4196 (N_4196,N_2412,N_2593);
nand U4197 (N_4197,N_3299,N_3255);
nand U4198 (N_4198,N_3871,N_3306);
and U4199 (N_4199,N_3822,N_3890);
or U4200 (N_4200,N_2321,N_2303);
or U4201 (N_4201,N_2703,N_2424);
nor U4202 (N_4202,N_2164,N_2777);
or U4203 (N_4203,N_3866,N_3709);
nand U4204 (N_4204,N_3464,N_3629);
or U4205 (N_4205,N_2151,N_2910);
and U4206 (N_4206,N_2482,N_3391);
and U4207 (N_4207,N_3141,N_2467);
nor U4208 (N_4208,N_2719,N_3084);
nand U4209 (N_4209,N_2111,N_3129);
xor U4210 (N_4210,N_3926,N_2930);
nand U4211 (N_4211,N_2296,N_2384);
nor U4212 (N_4212,N_3403,N_3272);
xor U4213 (N_4213,N_2453,N_2726);
nand U4214 (N_4214,N_2030,N_2443);
or U4215 (N_4215,N_3324,N_2430);
and U4216 (N_4216,N_2982,N_2394);
nand U4217 (N_4217,N_2558,N_2886);
and U4218 (N_4218,N_3372,N_2867);
and U4219 (N_4219,N_3980,N_2256);
xor U4220 (N_4220,N_3761,N_2774);
and U4221 (N_4221,N_2845,N_2342);
and U4222 (N_4222,N_3764,N_3222);
nand U4223 (N_4223,N_2936,N_3214);
xor U4224 (N_4224,N_3941,N_3893);
nor U4225 (N_4225,N_3087,N_2114);
xor U4226 (N_4226,N_3595,N_3182);
and U4227 (N_4227,N_2707,N_3820);
or U4228 (N_4228,N_2638,N_2193);
nor U4229 (N_4229,N_2701,N_3942);
xnor U4230 (N_4230,N_3566,N_2367);
nor U4231 (N_4231,N_3099,N_3058);
or U4232 (N_4232,N_2737,N_3804);
or U4233 (N_4233,N_3012,N_2036);
or U4234 (N_4234,N_2215,N_2142);
or U4235 (N_4235,N_2103,N_2643);
nor U4236 (N_4236,N_3397,N_2607);
nor U4237 (N_4237,N_3519,N_2186);
and U4238 (N_4238,N_2716,N_2880);
nand U4239 (N_4239,N_2386,N_2575);
xnor U4240 (N_4240,N_3681,N_3782);
nand U4241 (N_4241,N_2464,N_3121);
nand U4242 (N_4242,N_3975,N_3947);
or U4243 (N_4243,N_3335,N_2627);
or U4244 (N_4244,N_2481,N_3474);
nand U4245 (N_4245,N_3581,N_2330);
nor U4246 (N_4246,N_3502,N_2069);
or U4247 (N_4247,N_3452,N_3995);
and U4248 (N_4248,N_3079,N_2814);
xnor U4249 (N_4249,N_2162,N_3813);
nor U4250 (N_4250,N_2339,N_2776);
and U4251 (N_4251,N_3891,N_3560);
nand U4252 (N_4252,N_3490,N_2900);
nand U4253 (N_4253,N_2877,N_3421);
xnor U4254 (N_4254,N_3451,N_3717);
nor U4255 (N_4255,N_2768,N_2598);
xnor U4256 (N_4256,N_3951,N_3243);
nor U4257 (N_4257,N_3410,N_2262);
and U4258 (N_4258,N_2338,N_2055);
or U4259 (N_4259,N_3959,N_2129);
xor U4260 (N_4260,N_2801,N_3525);
nor U4261 (N_4261,N_2462,N_3000);
nor U4262 (N_4262,N_3812,N_2199);
xor U4263 (N_4263,N_2395,N_2121);
and U4264 (N_4264,N_2597,N_3808);
nand U4265 (N_4265,N_3470,N_3693);
or U4266 (N_4266,N_2897,N_2200);
nand U4267 (N_4267,N_2564,N_3837);
nand U4268 (N_4268,N_2841,N_2362);
xnor U4269 (N_4269,N_3831,N_2198);
nor U4270 (N_4270,N_2913,N_3501);
nand U4271 (N_4271,N_2434,N_3239);
or U4272 (N_4272,N_2765,N_2992);
nor U4273 (N_4273,N_2411,N_3615);
xnor U4274 (N_4274,N_3966,N_3348);
or U4275 (N_4275,N_3675,N_3580);
nand U4276 (N_4276,N_3639,N_3263);
and U4277 (N_4277,N_3117,N_3635);
nand U4278 (N_4278,N_3256,N_3914);
nor U4279 (N_4279,N_3010,N_3628);
or U4280 (N_4280,N_3245,N_2461);
or U4281 (N_4281,N_3020,N_3883);
xnor U4282 (N_4282,N_2334,N_3855);
and U4283 (N_4283,N_3123,N_2548);
xnor U4284 (N_4284,N_3418,N_3863);
nand U4285 (N_4285,N_2054,N_3957);
xnor U4286 (N_4286,N_3739,N_2511);
nor U4287 (N_4287,N_3537,N_2854);
nand U4288 (N_4288,N_2447,N_2675);
nand U4289 (N_4289,N_2266,N_2655);
and U4290 (N_4290,N_2115,N_3969);
nand U4291 (N_4291,N_2849,N_3710);
nand U4292 (N_4292,N_2278,N_3539);
nor U4293 (N_4293,N_3658,N_2624);
and U4294 (N_4294,N_3340,N_2314);
nand U4295 (N_4295,N_3849,N_3146);
xor U4296 (N_4296,N_3924,N_2828);
xnor U4297 (N_4297,N_3575,N_3167);
or U4298 (N_4298,N_3494,N_3641);
and U4299 (N_4299,N_3375,N_2970);
xor U4300 (N_4300,N_3902,N_2274);
and U4301 (N_4301,N_3161,N_2246);
and U4302 (N_4302,N_2689,N_2327);
xor U4303 (N_4303,N_2152,N_3130);
or U4304 (N_4304,N_3358,N_3271);
xor U4305 (N_4305,N_2491,N_3832);
xnor U4306 (N_4306,N_2557,N_2140);
nor U4307 (N_4307,N_2884,N_3848);
nand U4308 (N_4308,N_2029,N_2917);
or U4309 (N_4309,N_3100,N_2104);
and U4310 (N_4310,N_2123,N_2110);
nand U4311 (N_4311,N_3439,N_3112);
and U4312 (N_4312,N_3696,N_2432);
and U4313 (N_4313,N_2442,N_2914);
xor U4314 (N_4314,N_2031,N_2388);
and U4315 (N_4315,N_3729,N_2585);
nand U4316 (N_4316,N_2484,N_2934);
and U4317 (N_4317,N_3503,N_2025);
nor U4318 (N_4318,N_3830,N_3799);
nor U4319 (N_4319,N_3073,N_3511);
nor U4320 (N_4320,N_3151,N_2322);
nand U4321 (N_4321,N_2964,N_3643);
or U4322 (N_4322,N_3617,N_3904);
xnor U4323 (N_4323,N_2124,N_2295);
or U4324 (N_4324,N_2389,N_3977);
nand U4325 (N_4325,N_3888,N_2665);
nand U4326 (N_4326,N_2538,N_2026);
and U4327 (N_4327,N_3131,N_3499);
or U4328 (N_4328,N_3062,N_2232);
nand U4329 (N_4329,N_2660,N_2470);
nand U4330 (N_4330,N_2359,N_3313);
nand U4331 (N_4331,N_3649,N_2891);
nor U4332 (N_4332,N_3777,N_2281);
nor U4333 (N_4333,N_3338,N_3730);
xor U4334 (N_4334,N_3846,N_3785);
nand U4335 (N_4335,N_2431,N_2893);
and U4336 (N_4336,N_3953,N_2778);
and U4337 (N_4337,N_3405,N_3296);
nor U4338 (N_4338,N_3994,N_2739);
or U4339 (N_4339,N_2083,N_2135);
nor U4340 (N_4340,N_2185,N_3697);
or U4341 (N_4341,N_3734,N_3912);
xnor U4342 (N_4342,N_3127,N_3765);
nand U4343 (N_4343,N_3543,N_2945);
xnor U4344 (N_4344,N_3297,N_3492);
nor U4345 (N_4345,N_2632,N_3330);
nor U4346 (N_4346,N_3442,N_3971);
nand U4347 (N_4347,N_3988,N_3093);
xnor U4348 (N_4348,N_3150,N_2493);
and U4349 (N_4349,N_3847,N_3682);
nand U4350 (N_4350,N_3602,N_3419);
nor U4351 (N_4351,N_2487,N_3790);
or U4352 (N_4352,N_3195,N_2549);
nor U4353 (N_4353,N_3266,N_3248);
nand U4354 (N_4354,N_3985,N_2381);
or U4355 (N_4355,N_2799,N_3041);
xor U4356 (N_4356,N_3124,N_3125);
nand U4357 (N_4357,N_3486,N_3905);
xnor U4358 (N_4358,N_2793,N_2452);
or U4359 (N_4359,N_3722,N_3645);
or U4360 (N_4360,N_3364,N_3868);
nand U4361 (N_4361,N_3173,N_2380);
xor U4362 (N_4362,N_3152,N_2908);
and U4363 (N_4363,N_2806,N_2122);
nor U4364 (N_4364,N_3763,N_2245);
or U4365 (N_4365,N_3787,N_3295);
or U4366 (N_4366,N_2370,N_2317);
nor U4367 (N_4367,N_2088,N_3895);
nand U4368 (N_4368,N_2502,N_2879);
nand U4369 (N_4369,N_3954,N_2108);
or U4370 (N_4370,N_2821,N_2474);
nor U4371 (N_4371,N_2637,N_3992);
nor U4372 (N_4372,N_2271,N_3322);
nand U4373 (N_4373,N_2436,N_3319);
nand U4374 (N_4374,N_3708,N_2969);
or U4375 (N_4375,N_2267,N_2587);
or U4376 (N_4376,N_3976,N_3835);
nand U4377 (N_4377,N_2335,N_3292);
or U4378 (N_4378,N_2721,N_2476);
nand U4379 (N_4379,N_3387,N_2225);
or U4380 (N_4380,N_2407,N_3238);
nand U4381 (N_4381,N_2328,N_3889);
xnor U4382 (N_4382,N_2832,N_2039);
and U4383 (N_4383,N_3943,N_3005);
nor U4384 (N_4384,N_2130,N_2479);
and U4385 (N_4385,N_2304,N_3732);
xor U4386 (N_4386,N_3267,N_3505);
or U4387 (N_4387,N_3612,N_2574);
or U4388 (N_4388,N_3217,N_2931);
nand U4389 (N_4389,N_3775,N_3430);
nand U4390 (N_4390,N_2001,N_2933);
xor U4391 (N_4391,N_2428,N_2280);
nor U4392 (N_4392,N_3345,N_2833);
or U4393 (N_4393,N_2400,N_3283);
nor U4394 (N_4394,N_3619,N_3836);
xnor U4395 (N_4395,N_3467,N_3149);
or U4396 (N_4396,N_3356,N_2843);
and U4397 (N_4397,N_2610,N_2755);
xor U4398 (N_4398,N_2297,N_2525);
and U4399 (N_4399,N_3573,N_3731);
or U4400 (N_4400,N_2939,N_2157);
xor U4401 (N_4401,N_3240,N_3054);
and U4402 (N_4402,N_3270,N_2817);
nor U4403 (N_4403,N_2903,N_3588);
xnor U4404 (N_4404,N_2236,N_3377);
and U4405 (N_4405,N_2883,N_2770);
and U4406 (N_4406,N_3047,N_3861);
and U4407 (N_4407,N_2438,N_2662);
xnor U4408 (N_4408,N_3071,N_3554);
and U4409 (N_4409,N_2955,N_2680);
or U4410 (N_4410,N_3906,N_3650);
and U4411 (N_4411,N_2050,N_2997);
xnor U4412 (N_4412,N_3584,N_2714);
and U4413 (N_4413,N_3570,N_3212);
nor U4414 (N_4414,N_3192,N_3591);
xnor U4415 (N_4415,N_3370,N_2985);
nor U4416 (N_4416,N_2508,N_2239);
nand U4417 (N_4417,N_2537,N_2563);
or U4418 (N_4418,N_2248,N_3609);
nor U4419 (N_4419,N_2763,N_3317);
nand U4420 (N_4420,N_3571,N_3999);
xor U4421 (N_4421,N_2842,N_2473);
and U4422 (N_4422,N_2611,N_3360);
or U4423 (N_4423,N_3298,N_2787);
nor U4424 (N_4424,N_3608,N_3065);
and U4425 (N_4425,N_2823,N_2639);
nor U4426 (N_4426,N_2562,N_2918);
nor U4427 (N_4427,N_2736,N_2580);
nor U4428 (N_4428,N_2644,N_2299);
nor U4429 (N_4429,N_3626,N_2175);
and U4430 (N_4430,N_2010,N_2090);
nand U4431 (N_4431,N_3671,N_2855);
xor U4432 (N_4432,N_2668,N_2628);
xor U4433 (N_4433,N_2773,N_3378);
xnor U4434 (N_4434,N_2514,N_3823);
or U4435 (N_4435,N_3285,N_2635);
and U4436 (N_4436,N_3274,N_3228);
or U4437 (N_4437,N_2163,N_2457);
or U4438 (N_4438,N_2722,N_3872);
xnor U4439 (N_4439,N_2376,N_2751);
and U4440 (N_4440,N_2958,N_3651);
nand U4441 (N_4441,N_3878,N_2839);
and U4442 (N_4442,N_2560,N_2860);
or U4443 (N_4443,N_3815,N_3284);
nand U4444 (N_4444,N_3092,N_3705);
xnor U4445 (N_4445,N_2998,N_2695);
or U4446 (N_4446,N_3251,N_3038);
or U4447 (N_4447,N_3657,N_3408);
and U4448 (N_4448,N_2965,N_3740);
xnor U4449 (N_4449,N_2977,N_2015);
and U4450 (N_4450,N_3655,N_3487);
nand U4451 (N_4451,N_2708,N_3916);
xnor U4452 (N_4452,N_2735,N_2265);
nand U4453 (N_4453,N_3116,N_2455);
nand U4454 (N_4454,N_2576,N_2895);
nand U4455 (N_4455,N_2094,N_3140);
nand U4456 (N_4456,N_2131,N_2364);
and U4457 (N_4457,N_3033,N_3552);
and U4458 (N_4458,N_2160,N_3762);
or U4459 (N_4459,N_3115,N_3496);
nand U4460 (N_4460,N_3393,N_2834);
or U4461 (N_4461,N_3704,N_2269);
or U4462 (N_4462,N_2405,N_2179);
and U4463 (N_4463,N_2779,N_3771);
xnor U4464 (N_4464,N_2172,N_2745);
nand U4465 (N_4465,N_3523,N_2858);
or U4466 (N_4466,N_3384,N_3850);
nor U4467 (N_4467,N_3120,N_2781);
or U4468 (N_4468,N_2496,N_3795);
and U4469 (N_4469,N_3275,N_2948);
or U4470 (N_4470,N_3234,N_2404);
and U4471 (N_4471,N_3278,N_2622);
or U4472 (N_4472,N_2653,N_2926);
and U4473 (N_4473,N_2264,N_3126);
xor U4474 (N_4474,N_3293,N_2048);
or U4475 (N_4475,N_3064,N_2229);
and U4476 (N_4476,N_3133,N_2979);
and U4477 (N_4477,N_3773,N_3699);
xnor U4478 (N_4478,N_2410,N_2904);
or U4479 (N_4479,N_3965,N_2646);
xnor U4480 (N_4480,N_3407,N_2521);
nor U4481 (N_4481,N_2844,N_3323);
nor U4482 (N_4482,N_3199,N_3076);
nor U4483 (N_4483,N_2348,N_2976);
nand U4484 (N_4484,N_3767,N_2804);
nor U4485 (N_4485,N_3136,N_3513);
or U4486 (N_4486,N_2940,N_3354);
and U4487 (N_4487,N_2202,N_3876);
xor U4488 (N_4488,N_2594,N_2522);
nor U4489 (N_4489,N_3737,N_2978);
or U4490 (N_4490,N_2633,N_2686);
nor U4491 (N_4491,N_3286,N_2378);
and U4492 (N_4492,N_3844,N_3259);
nand U4493 (N_4493,N_3897,N_2951);
xnor U4494 (N_4494,N_3198,N_3618);
nand U4495 (N_4495,N_3637,N_2608);
xor U4496 (N_4496,N_3070,N_3023);
xor U4497 (N_4497,N_2837,N_3647);
nor U4498 (N_4498,N_3945,N_3253);
nor U4499 (N_4499,N_3392,N_3105);
or U4500 (N_4500,N_2024,N_3520);
nand U4501 (N_4501,N_3544,N_2542);
xor U4502 (N_4502,N_3851,N_3736);
xnor U4503 (N_4503,N_2063,N_2365);
nor U4504 (N_4504,N_2874,N_3197);
xor U4505 (N_4505,N_3733,N_2073);
xor U4506 (N_4506,N_3039,N_3956);
nor U4507 (N_4507,N_3359,N_3887);
nand U4508 (N_4508,N_2372,N_2807);
nor U4509 (N_4509,N_2974,N_3521);
and U4510 (N_4510,N_2141,N_2037);
nand U4511 (N_4511,N_3462,N_2641);
or U4512 (N_4512,N_3052,N_2619);
xor U4513 (N_4513,N_2089,N_3746);
nor U4514 (N_4514,N_2881,N_2305);
xor U4515 (N_4515,N_3803,N_3949);
nor U4516 (N_4516,N_2223,N_2308);
or U4517 (N_4517,N_2093,N_2840);
nor U4518 (N_4518,N_2674,N_2810);
and U4519 (N_4519,N_3002,N_2125);
or U4520 (N_4520,N_2406,N_2667);
or U4521 (N_4521,N_3925,N_3624);
nor U4522 (N_4522,N_3232,N_3143);
xor U4523 (N_4523,N_3174,N_2856);
xnor U4524 (N_4524,N_3770,N_3669);
nor U4525 (N_4525,N_2351,N_3611);
or U4526 (N_4526,N_2853,N_2340);
or U4527 (N_4527,N_2573,N_2518);
xnor U4528 (N_4528,N_3110,N_3469);
nor U4529 (N_4529,N_3082,N_2033);
and U4530 (N_4530,N_2358,N_3482);
xnor U4531 (N_4531,N_2784,N_3991);
and U4532 (N_4532,N_3919,N_2960);
xnor U4533 (N_4533,N_2692,N_3090);
xnor U4534 (N_4534,N_3970,N_2901);
or U4535 (N_4535,N_2070,N_3202);
and U4536 (N_4536,N_2261,N_2170);
nor U4537 (N_4537,N_2288,N_3362);
nand U4538 (N_4538,N_3689,N_2545);
and U4539 (N_4539,N_3922,N_3670);
nor U4540 (N_4540,N_2194,N_2588);
nor U4541 (N_4541,N_2741,N_3852);
nor U4542 (N_4542,N_2838,N_2206);
or U4543 (N_4543,N_3491,N_3546);
xor U4544 (N_4544,N_2079,N_2540);
xor U4545 (N_4545,N_3024,N_2107);
nor U4546 (N_4546,N_2556,N_2932);
nand U4547 (N_4547,N_2375,N_2444);
nor U4548 (N_4548,N_3788,N_3948);
or U4549 (N_4549,N_2651,N_3006);
or U4550 (N_4550,N_3008,N_2258);
and U4551 (N_4551,N_2252,N_3122);
nor U4552 (N_4552,N_3042,N_3142);
and U4553 (N_4553,N_3528,N_2769);
nor U4554 (N_4554,N_3723,N_3982);
nor U4555 (N_4555,N_2682,N_3996);
and U4556 (N_4556,N_3210,N_3526);
nor U4557 (N_4557,N_2771,N_2397);
and U4558 (N_4558,N_3454,N_2516);
xnor U4559 (N_4559,N_3597,N_2762);
nand U4560 (N_4560,N_2870,N_3662);
and U4561 (N_4561,N_3825,N_3398);
or U4562 (N_4562,N_2399,N_3921);
xor U4563 (N_4563,N_3165,N_2645);
or U4564 (N_4564,N_2477,N_3780);
and U4565 (N_4565,N_2401,N_3310);
nor U4566 (N_4566,N_3944,N_2214);
and U4567 (N_4567,N_3057,N_2715);
and U4568 (N_4568,N_3910,N_2782);
xor U4569 (N_4569,N_2500,N_3508);
nor U4570 (N_4570,N_2341,N_3727);
xnor U4571 (N_4571,N_3877,N_3483);
nand U4572 (N_4572,N_2582,N_3579);
xnor U4573 (N_4573,N_3137,N_2310);
or U4574 (N_4574,N_2761,N_2963);
nand U4575 (N_4575,N_3091,N_2909);
or U4576 (N_4576,N_3318,N_3128);
nor U4577 (N_4577,N_2329,N_2600);
and U4578 (N_4578,N_3854,N_3972);
nor U4579 (N_4579,N_2307,N_2572);
nand U4580 (N_4580,N_2561,N_2989);
xor U4581 (N_4581,N_2490,N_3168);
nor U4582 (N_4582,N_2872,N_3388);
nand U4583 (N_4583,N_2993,N_2683);
nand U4584 (N_4584,N_2242,N_2293);
nand U4585 (N_4585,N_3477,N_3772);
xor U4586 (N_4586,N_3415,N_2051);
and U4587 (N_4587,N_3400,N_3701);
xnor U4588 (N_4588,N_2623,N_3118);
and U4589 (N_4589,N_2419,N_3720);
nand U4590 (N_4590,N_3585,N_2996);
nor U4591 (N_4591,N_3735,N_3751);
and U4592 (N_4592,N_2873,N_2052);
nor U4593 (N_4593,N_3300,N_3331);
and U4594 (N_4594,N_2727,N_2469);
nor U4595 (N_4595,N_3489,N_3172);
xor U4596 (N_4596,N_3406,N_2584);
nand U4597 (N_4597,N_2065,N_2007);
xor U4598 (N_4598,N_2306,N_3315);
xor U4599 (N_4599,N_3316,N_3069);
nand U4600 (N_4600,N_3827,N_3307);
nor U4601 (N_4601,N_3993,N_2888);
or U4602 (N_4602,N_3962,N_3644);
nand U4603 (N_4603,N_3461,N_2238);
nor U4604 (N_4604,N_3676,N_2938);
nor U4605 (N_4605,N_2109,N_3433);
or U4606 (N_4606,N_3824,N_2078);
nand U4607 (N_4607,N_2091,N_2953);
xnor U4608 (N_4608,N_3281,N_2544);
or U4609 (N_4609,N_3342,N_2792);
nor U4610 (N_4610,N_2234,N_3328);
xor U4611 (N_4611,N_2350,N_2942);
and U4612 (N_4612,N_3572,N_3604);
and U4613 (N_4613,N_2396,N_3404);
xnor U4614 (N_4614,N_2723,N_2213);
and U4615 (N_4615,N_2592,N_2257);
nor U4616 (N_4616,N_2009,N_2402);
xor U4617 (N_4617,N_2167,N_2313);
nor U4618 (N_4618,N_2337,N_3899);
nand U4619 (N_4619,N_3495,N_2098);
and U4620 (N_4620,N_3664,N_2201);
xnor U4621 (N_4621,N_3934,N_3488);
xnor U4622 (N_4622,N_3504,N_3923);
and U4623 (N_4623,N_3294,N_2694);
and U4624 (N_4624,N_2092,N_3191);
nand U4625 (N_4625,N_3134,N_3314);
or U4626 (N_4626,N_3894,N_3640);
nor U4627 (N_4627,N_2625,N_2520);
and U4628 (N_4628,N_2427,N_3557);
and U4629 (N_4629,N_3367,N_2687);
or U4630 (N_4630,N_3420,N_2077);
nand U4631 (N_4631,N_3673,N_2864);
or U4632 (N_4632,N_2138,N_2355);
or U4633 (N_4633,N_2636,N_3231);
or U4634 (N_4634,N_2042,N_2315);
xnor U4635 (N_4635,N_3621,N_2289);
nand U4636 (N_4636,N_2732,N_3261);
and U4637 (N_4637,N_3450,N_3793);
and U4638 (N_4638,N_2666,N_2456);
nand U4639 (N_4639,N_3247,N_3989);
xor U4640 (N_4640,N_2212,N_3371);
or U4641 (N_4641,N_2106,N_3203);
or U4642 (N_4642,N_3636,N_2016);
or U4643 (N_4643,N_2118,N_2620);
nor U4644 (N_4644,N_2374,N_3334);
nand U4645 (N_4645,N_3677,N_2190);
or U4646 (N_4646,N_2552,N_2415);
nand U4647 (N_4647,N_3715,N_2693);
or U4648 (N_4648,N_2159,N_3857);
nor U4649 (N_4649,N_2409,N_3683);
nand U4650 (N_4650,N_2272,N_2137);
nor U4651 (N_4651,N_2713,N_3394);
or U4652 (N_4652,N_3797,N_2731);
or U4653 (N_4653,N_3034,N_3598);
nor U4654 (N_4654,N_2038,N_3414);
or U4655 (N_4655,N_2495,N_3236);
nor U4656 (N_4656,N_2578,N_3417);
nor U4657 (N_4657,N_3623,N_2080);
nand U4658 (N_4658,N_2676,N_3691);
nand U4659 (N_4659,N_2790,N_3412);
xor U4660 (N_4660,N_2032,N_2061);
or U4661 (N_4661,N_2454,N_2505);
or U4662 (N_4662,N_2312,N_3471);
and U4663 (N_4663,N_3929,N_2609);
nand U4664 (N_4664,N_3344,N_2581);
and U4665 (N_4665,N_2017,N_2882);
or U4666 (N_4666,N_3880,N_3885);
or U4667 (N_4667,N_2154,N_3791);
or U4668 (N_4668,N_2309,N_2815);
nand U4669 (N_4669,N_3870,N_2589);
nand U4670 (N_4670,N_3936,N_3060);
xnor U4671 (N_4671,N_2441,N_3166);
nor U4672 (N_4672,N_2440,N_3633);
nand U4673 (N_4673,N_3456,N_3089);
nand U4674 (N_4674,N_3227,N_3760);
nor U4675 (N_4675,N_2967,N_2528);
nand U4676 (N_4676,N_2361,N_3748);
nand U4677 (N_4677,N_2046,N_3700);
and U4678 (N_4678,N_2827,N_3350);
nor U4679 (N_4679,N_2529,N_2387);
nand U4680 (N_4680,N_2354,N_2515);
nand U4681 (N_4681,N_2458,N_2673);
and U4682 (N_4682,N_2685,N_2775);
nand U4683 (N_4683,N_3984,N_3472);
nor U4684 (N_4684,N_3564,N_2216);
or U4685 (N_4685,N_2571,N_3357);
or U4686 (N_4686,N_3789,N_2018);
xnor U4687 (N_4687,N_3059,N_3548);
and U4688 (N_4688,N_3908,N_3246);
and U4689 (N_4689,N_2277,N_3007);
xnor U4690 (N_4690,N_3754,N_2911);
nand U4691 (N_4691,N_2971,N_3774);
and U4692 (N_4692,N_2962,N_2059);
or U4693 (N_4693,N_2012,N_2283);
and U4694 (N_4694,N_2983,N_3506);
and U4695 (N_4695,N_3235,N_2764);
or U4696 (N_4696,N_2155,N_2324);
and U4697 (N_4697,N_3840,N_2899);
nand U4698 (N_4698,N_2885,N_3997);
nor U4699 (N_4699,N_2664,N_2795);
and U4700 (N_4700,N_3541,N_2829);
and U4701 (N_4701,N_2087,N_2825);
xor U4702 (N_4702,N_3514,N_2177);
and U4703 (N_4703,N_2102,N_2928);
or U4704 (N_4704,N_2850,N_2331);
xor U4705 (N_4705,N_3547,N_2086);
nor U4706 (N_4706,N_2486,N_3545);
nand U4707 (N_4707,N_2021,N_3352);
or U4708 (N_4708,N_3692,N_2371);
and U4709 (N_4709,N_2654,N_2408);
and U4710 (N_4710,N_2980,N_3209);
xor U4711 (N_4711,N_2733,N_3509);
nand U4712 (N_4712,N_3183,N_2789);
or U4713 (N_4713,N_2097,N_3440);
or U4714 (N_4714,N_2912,N_2147);
and U4715 (N_4715,N_2547,N_3913);
nand U4716 (N_4716,N_3103,N_2203);
xnor U4717 (N_4717,N_3268,N_2366);
xnor U4718 (N_4718,N_3402,N_2492);
xnor U4719 (N_4719,N_2112,N_2333);
and U4720 (N_4720,N_3431,N_2224);
or U4721 (N_4721,N_3821,N_2169);
and U4722 (N_4722,N_3102,N_3858);
or U4723 (N_4723,N_2002,N_3156);
xor U4724 (N_4724,N_2205,N_3555);
and U4725 (N_4725,N_2526,N_2767);
nand U4726 (N_4726,N_2717,N_2425);
nand U4727 (N_4727,N_2811,N_3516);
and U4728 (N_4728,N_3022,N_2249);
nand U4729 (N_4729,N_3688,N_2943);
nand U4730 (N_4730,N_3153,N_2730);
and U4731 (N_4731,N_2744,N_3512);
or U4732 (N_4732,N_2008,N_2586);
nand U4733 (N_4733,N_2604,N_3427);
and U4734 (N_4734,N_3028,N_3409);
nor U4735 (N_4735,N_3667,N_3533);
xor U4736 (N_4736,N_2217,N_3698);
nor U4737 (N_4737,N_2463,N_2251);
nor U4738 (N_4738,N_2326,N_2196);
nor U4739 (N_4739,N_2642,N_3441);
nor U4740 (N_4740,N_2657,N_2148);
nand U4741 (N_4741,N_3229,N_3687);
and U4742 (N_4742,N_3892,N_3154);
and U4743 (N_4743,N_2902,N_2347);
xor U4744 (N_4744,N_3805,N_2921);
or U4745 (N_4745,N_3845,N_2614);
and U4746 (N_4746,N_3053,N_3373);
or U4747 (N_4747,N_2134,N_3086);
nor U4748 (N_4748,N_2144,N_2437);
and U4749 (N_4749,N_2368,N_2047);
nor U4750 (N_4750,N_3416,N_2126);
nor U4751 (N_4751,N_3932,N_2802);
nor U4752 (N_4752,N_2231,N_3304);
nand U4753 (N_4753,N_3001,N_3928);
and U4754 (N_4754,N_2527,N_2649);
nand U4755 (N_4755,N_3347,N_3535);
and U4756 (N_4756,N_2153,N_2056);
nand U4757 (N_4757,N_3728,N_3642);
nand U4758 (N_4758,N_2166,N_3205);
xor U4759 (N_4759,N_3288,N_3672);
and U4760 (N_4760,N_3465,N_2968);
or U4761 (N_4761,N_3903,N_3741);
nand U4762 (N_4762,N_2812,N_3424);
and U4763 (N_4763,N_2907,N_2859);
nand U4764 (N_4764,N_3147,N_3291);
nor U4765 (N_4765,N_3656,N_3839);
nand U4766 (N_4766,N_3036,N_2532);
xor U4767 (N_4767,N_3015,N_3429);
or U4768 (N_4768,N_2178,N_2875);
xnor U4769 (N_4769,N_2494,N_2819);
and U4770 (N_4770,N_2243,N_3080);
nand U4771 (N_4771,N_3796,N_3631);
nor U4772 (N_4772,N_2483,N_2783);
xnor U4773 (N_4773,N_2460,N_3473);
and U4774 (N_4774,N_3273,N_3480);
nor U4775 (N_4775,N_3460,N_2445);
and U4776 (N_4776,N_3280,N_2233);
and U4777 (N_4777,N_3711,N_3220);
xor U4778 (N_4778,N_2189,N_3918);
or U4779 (N_4779,N_2543,N_2133);
nor U4780 (N_4780,N_2027,N_3769);
nand U4781 (N_4781,N_2603,N_3551);
and U4782 (N_4782,N_3630,N_2332);
and U4783 (N_4783,N_3049,N_3652);
and U4784 (N_4784,N_2391,N_2861);
or U4785 (N_4785,N_3529,N_2290);
nand U4786 (N_4786,N_2174,N_2539);
nand U4787 (N_4787,N_3896,N_3257);
or U4788 (N_4788,N_3135,N_2678);
xnor U4789 (N_4789,N_3026,N_3037);
and U4790 (N_4790,N_3216,N_3101);
and U4791 (N_4791,N_3927,N_2259);
xor U4792 (N_4792,N_2803,N_3386);
and U4793 (N_4793,N_3303,N_3106);
and U4794 (N_4794,N_3507,N_3448);
nand U4795 (N_4795,N_2659,N_2863);
nand U4796 (N_4796,N_2263,N_2679);
and U4797 (N_4797,N_3531,N_2005);
nor U4798 (N_4798,N_2987,N_3111);
or U4799 (N_4799,N_2785,N_2489);
nor U4800 (N_4800,N_3190,N_3302);
and U4801 (N_4801,N_3389,N_3569);
and U4802 (N_4802,N_3363,N_2824);
xor U4803 (N_4803,N_2294,N_2728);
nor U4804 (N_4804,N_3437,N_2800);
or U4805 (N_4805,N_2448,N_3648);
and U4806 (N_4806,N_2451,N_2067);
and U4807 (N_4807,N_3184,N_3753);
nand U4808 (N_4808,N_3784,N_2738);
or U4809 (N_4809,N_3289,N_2612);
xnor U4810 (N_4810,N_2740,N_2346);
xnor U4811 (N_4811,N_3155,N_3873);
nor U4812 (N_4812,N_2756,N_2323);
and U4813 (N_4813,N_3939,N_3311);
nor U4814 (N_4814,N_3865,N_2421);
xnor U4815 (N_4815,N_3809,N_3369);
and U4816 (N_4816,N_3423,N_3145);
xor U4817 (N_4817,N_3616,N_2435);
or U4818 (N_4818,N_3684,N_2749);
nor U4819 (N_4819,N_2605,N_2429);
nand U4820 (N_4820,N_3638,N_3337);
nand U4821 (N_4821,N_3072,N_3665);
nor U4822 (N_4822,N_2831,N_2506);
nor U4823 (N_4823,N_2449,N_2357);
xnor U4824 (N_4824,N_3713,N_3607);
nor U4825 (N_4825,N_2621,N_3162);
xor U4826 (N_4826,N_3562,N_2507);
nor U4827 (N_4827,N_3660,N_3659);
or U4828 (N_4828,N_2413,N_3329);
nand U4829 (N_4829,N_3208,N_2896);
nor U4830 (N_4830,N_3674,N_2287);
or U4831 (N_4831,N_3869,N_2139);
and U4832 (N_4832,N_3712,N_3132);
nor U4833 (N_4833,N_3019,N_3180);
nand U4834 (N_4834,N_2064,N_3856);
xor U4835 (N_4835,N_3163,N_2095);
nand U4836 (N_4836,N_2292,N_3634);
nand U4837 (N_4837,N_2360,N_2754);
and U4838 (N_4838,N_3879,N_2857);
nor U4839 (N_4839,N_3920,N_3351);
nand U4840 (N_4840,N_3260,N_2758);
or U4841 (N_4841,N_2211,N_3833);
nor U4842 (N_4842,N_3987,N_2060);
or U4843 (N_4843,N_2865,N_2074);
or U4844 (N_4844,N_3935,N_3466);
xor U4845 (N_4845,N_2044,N_2446);
nand U4846 (N_4846,N_3759,N_3312);
and U4847 (N_4847,N_2553,N_3187);
xor U4848 (N_4848,N_3718,N_2040);
nor U4849 (N_4849,N_3170,N_2173);
nor U4850 (N_4850,N_2099,N_2311);
xor U4851 (N_4851,N_2356,N_2285);
nor U4852 (N_4852,N_3067,N_2182);
xnor U4853 (N_4853,N_2497,N_3096);
or U4854 (N_4854,N_3522,N_3109);
nand U4855 (N_4855,N_2062,N_2551);
nand U4856 (N_4856,N_2150,N_2669);
nor U4857 (N_4857,N_2734,N_3915);
xnor U4858 (N_4858,N_3603,N_2920);
nor U4859 (N_4859,N_3361,N_3074);
or U4860 (N_4860,N_2780,N_3349);
and U4861 (N_4861,N_2235,N_2629);
xor U4862 (N_4862,N_2892,N_2183);
or U4863 (N_4863,N_3113,N_2640);
nor U4864 (N_4864,N_2808,N_2373);
nor U4865 (N_4865,N_2927,N_2677);
or U4866 (N_4866,N_3413,N_2101);
xor U4867 (N_4867,N_2082,N_2023);
or U4868 (N_4868,N_2670,N_3432);
and U4869 (N_4869,N_3518,N_3743);
or U4870 (N_4870,N_3159,N_3819);
nand U4871 (N_4871,N_3632,N_3365);
nand U4872 (N_4872,N_3952,N_2698);
or U4873 (N_4873,N_2132,N_2711);
and U4874 (N_4874,N_2952,N_2846);
or U4875 (N_4875,N_2253,N_3003);
or U4876 (N_4876,N_3986,N_2688);
nor U4877 (N_4877,N_2750,N_2187);
and U4878 (N_4878,N_2369,N_3213);
nor U4879 (N_4879,N_2282,N_3558);
or U4880 (N_4880,N_3559,N_2536);
xor U4881 (N_4881,N_2291,N_2096);
nand U4882 (N_4882,N_3853,N_2851);
nand U4883 (N_4883,N_3436,N_3586);
nor U4884 (N_4884,N_3030,N_2316);
nand U4885 (N_4885,N_3578,N_3186);
or U4886 (N_4886,N_3411,N_2240);
nand U4887 (N_4887,N_3786,N_3218);
nand U4888 (N_4888,N_2923,N_3695);
nand U4889 (N_4889,N_2753,N_2418);
nor U4890 (N_4890,N_3075,N_2941);
nand U4891 (N_4891,N_3325,N_3455);
nand U4892 (N_4892,N_3747,N_3757);
and U4893 (N_4893,N_2509,N_2119);
nand U4894 (N_4894,N_2221,N_3778);
nor U4895 (N_4895,N_2423,N_3596);
nand U4896 (N_4896,N_3768,N_3742);
or U4897 (N_4897,N_3046,N_2916);
nand U4898 (N_4898,N_2617,N_3244);
xor U4899 (N_4899,N_3605,N_3678);
nor U4900 (N_4900,N_2081,N_2788);
and U4901 (N_4901,N_2994,N_2513);
nor U4902 (N_4902,N_3661,N_3264);
xor U4903 (N_4903,N_2672,N_3206);
nand U4904 (N_4904,N_2595,N_2700);
or U4905 (N_4905,N_3884,N_3463);
nor U4906 (N_4906,N_3973,N_2947);
and U4907 (N_4907,N_2690,N_2219);
or U4908 (N_4908,N_2145,N_2759);
xor U4909 (N_4909,N_2379,N_3233);
nand U4910 (N_4910,N_2414,N_2523);
nand U4911 (N_4911,N_2165,N_3017);
nand U4912 (N_4912,N_3428,N_3606);
or U4913 (N_4913,N_3882,N_3114);
nand U4914 (N_4914,N_3177,N_3679);
or U4915 (N_4915,N_3981,N_2876);
xnor U4916 (N_4916,N_2956,N_2382);
and U4917 (N_4917,N_2813,N_3707);
and U4918 (N_4918,N_3829,N_3237);
nand U4919 (N_4919,N_3326,N_2336);
nand U4920 (N_4920,N_3194,N_3807);
nand U4921 (N_4921,N_3479,N_2599);
or U4922 (N_4922,N_2922,N_3176);
nor U4923 (N_4923,N_2503,N_2546);
and U4924 (N_4924,N_3435,N_3567);
and U4925 (N_4925,N_2204,N_3738);
xor U4926 (N_4926,N_3160,N_3445);
nand U4927 (N_4927,N_2041,N_3666);
and U4928 (N_4928,N_2816,N_3834);
or U4929 (N_4929,N_2663,N_2084);
and U4930 (N_4930,N_3250,N_2671);
nor U4931 (N_4931,N_3810,N_3368);
or U4932 (N_4932,N_2530,N_3327);
nor U4933 (N_4933,N_2616,N_2158);
nor U4934 (N_4934,N_2260,N_2385);
xnor U4935 (N_4935,N_2020,N_3493);
or U4936 (N_4936,N_2935,N_2392);
and U4937 (N_4937,N_2298,N_2300);
and U4938 (N_4938,N_2276,N_3781);
and U4939 (N_4939,N_2241,N_2954);
and U4940 (N_4940,N_2468,N_2156);
xnor U4941 (N_4941,N_3374,N_3818);
xor U4942 (N_4942,N_2504,N_3613);
nor U4943 (N_4943,N_3148,N_3254);
and U4944 (N_4944,N_3527,N_3801);
and U4945 (N_4945,N_2006,N_2602);
nor U4946 (N_4946,N_3014,N_3204);
and U4947 (N_4947,N_2343,N_2302);
xor U4948 (N_4948,N_3158,N_3459);
xor U4949 (N_4949,N_2066,N_2228);
xor U4950 (N_4950,N_3601,N_3276);
and U4951 (N_4951,N_2136,N_2786);
or U4952 (N_4952,N_3940,N_3574);
and U4953 (N_4953,N_3806,N_3540);
nand U4954 (N_4954,N_3478,N_2255);
and U4955 (N_4955,N_3620,N_3215);
xor U4956 (N_4956,N_3346,N_2729);
or U4957 (N_4957,N_2949,N_2420);
nor U4958 (N_4958,N_3589,N_2075);
nor U4959 (N_4959,N_2999,N_3654);
nor U4960 (N_4960,N_3056,N_3088);
nor U4961 (N_4961,N_2869,N_2244);
or U4962 (N_4962,N_3399,N_2450);
xnor U4963 (N_4963,N_2222,N_3475);
nor U4964 (N_4964,N_3901,N_3838);
nor U4965 (N_4965,N_3422,N_3320);
xnor U4966 (N_4966,N_2352,N_2618);
xnor U4967 (N_4967,N_2848,N_3355);
or U4968 (N_4968,N_3434,N_2475);
and U4969 (N_4969,N_2866,N_2766);
nand U4970 (N_4970,N_2517,N_3716);
nand U4971 (N_4971,N_3449,N_3800);
xor U4972 (N_4972,N_2275,N_3946);
xor U4973 (N_4973,N_3051,N_3968);
nand U4974 (N_4974,N_2168,N_3553);
or U4975 (N_4975,N_3859,N_3862);
and U4976 (N_4976,N_2377,N_3444);
nand U4977 (N_4977,N_3817,N_2830);
or U4978 (N_4978,N_3690,N_3532);
nor U4979 (N_4979,N_3515,N_2742);
nor U4980 (N_4980,N_2325,N_3582);
or U4981 (N_4981,N_3181,N_2004);
nand U4982 (N_4982,N_2889,N_3211);
and U4983 (N_4983,N_2709,N_3816);
xor U4984 (N_4984,N_3258,N_2191);
nor U4985 (N_4985,N_3907,N_3779);
nor U4986 (N_4986,N_3931,N_2555);
and U4987 (N_4987,N_3881,N_3517);
nor U4988 (N_4988,N_2975,N_3843);
or U4989 (N_4989,N_2210,N_3568);
and U4990 (N_4990,N_3376,N_2100);
xor U4991 (N_4991,N_2180,N_2143);
nor U4992 (N_4992,N_2472,N_3841);
xor U4993 (N_4993,N_2072,N_3561);
or U4994 (N_4994,N_3438,N_3458);
xor U4995 (N_4995,N_3811,N_3576);
xor U4996 (N_4996,N_2752,N_2524);
and U4997 (N_4997,N_2459,N_2797);
and U4998 (N_4998,N_3339,N_2554);
and U4999 (N_4999,N_3221,N_2822);
nor U5000 (N_5000,N_3580,N_3770);
and U5001 (N_5001,N_2188,N_3436);
nand U5002 (N_5002,N_3688,N_2273);
or U5003 (N_5003,N_2608,N_2135);
or U5004 (N_5004,N_3811,N_3451);
nor U5005 (N_5005,N_2529,N_2593);
or U5006 (N_5006,N_2905,N_2939);
nand U5007 (N_5007,N_2473,N_3939);
nor U5008 (N_5008,N_3032,N_2133);
or U5009 (N_5009,N_3761,N_3795);
nand U5010 (N_5010,N_2961,N_3667);
nor U5011 (N_5011,N_2686,N_2304);
nor U5012 (N_5012,N_2468,N_3993);
and U5013 (N_5013,N_2372,N_2241);
or U5014 (N_5014,N_2974,N_3289);
and U5015 (N_5015,N_2052,N_3687);
xor U5016 (N_5016,N_2425,N_2641);
or U5017 (N_5017,N_3899,N_2296);
nand U5018 (N_5018,N_2123,N_3528);
or U5019 (N_5019,N_3004,N_2513);
nand U5020 (N_5020,N_3347,N_3833);
nor U5021 (N_5021,N_2733,N_3668);
nand U5022 (N_5022,N_2486,N_2845);
nor U5023 (N_5023,N_3392,N_3561);
nand U5024 (N_5024,N_2853,N_2286);
and U5025 (N_5025,N_2783,N_2327);
or U5026 (N_5026,N_3909,N_2219);
and U5027 (N_5027,N_3243,N_2229);
or U5028 (N_5028,N_3466,N_2462);
nand U5029 (N_5029,N_2005,N_2782);
nor U5030 (N_5030,N_3055,N_3808);
or U5031 (N_5031,N_3580,N_2774);
and U5032 (N_5032,N_3713,N_3248);
nand U5033 (N_5033,N_3048,N_3971);
and U5034 (N_5034,N_3551,N_2617);
or U5035 (N_5035,N_2299,N_3954);
xor U5036 (N_5036,N_3697,N_3652);
nor U5037 (N_5037,N_2363,N_2616);
xor U5038 (N_5038,N_2899,N_2441);
nand U5039 (N_5039,N_3599,N_2454);
or U5040 (N_5040,N_2479,N_2400);
and U5041 (N_5041,N_2973,N_3794);
nand U5042 (N_5042,N_3944,N_3956);
xor U5043 (N_5043,N_2988,N_3362);
nand U5044 (N_5044,N_3570,N_2157);
nor U5045 (N_5045,N_3440,N_2692);
and U5046 (N_5046,N_3079,N_3731);
xnor U5047 (N_5047,N_2093,N_3164);
nor U5048 (N_5048,N_3575,N_2124);
xnor U5049 (N_5049,N_2890,N_2402);
or U5050 (N_5050,N_3086,N_2646);
and U5051 (N_5051,N_3806,N_3613);
nand U5052 (N_5052,N_2744,N_2932);
nand U5053 (N_5053,N_3229,N_2064);
or U5054 (N_5054,N_2161,N_2909);
or U5055 (N_5055,N_3230,N_2703);
and U5056 (N_5056,N_3711,N_3196);
nor U5057 (N_5057,N_2898,N_3257);
or U5058 (N_5058,N_2310,N_2402);
nor U5059 (N_5059,N_3049,N_2532);
xor U5060 (N_5060,N_2805,N_3906);
nand U5061 (N_5061,N_3795,N_3468);
nor U5062 (N_5062,N_2531,N_3205);
or U5063 (N_5063,N_2660,N_2413);
xnor U5064 (N_5064,N_3610,N_3961);
nor U5065 (N_5065,N_3277,N_2727);
nor U5066 (N_5066,N_3017,N_2831);
nand U5067 (N_5067,N_2126,N_2392);
or U5068 (N_5068,N_2254,N_2645);
or U5069 (N_5069,N_2536,N_2555);
nor U5070 (N_5070,N_3335,N_3818);
nor U5071 (N_5071,N_3290,N_2012);
xnor U5072 (N_5072,N_3181,N_2587);
nand U5073 (N_5073,N_2973,N_3171);
nand U5074 (N_5074,N_3994,N_2849);
or U5075 (N_5075,N_2234,N_3202);
or U5076 (N_5076,N_2406,N_2751);
nand U5077 (N_5077,N_2595,N_2040);
or U5078 (N_5078,N_2440,N_3794);
nand U5079 (N_5079,N_3303,N_3455);
and U5080 (N_5080,N_2348,N_3685);
or U5081 (N_5081,N_2313,N_2414);
nand U5082 (N_5082,N_3058,N_3333);
or U5083 (N_5083,N_3705,N_2057);
nor U5084 (N_5084,N_3226,N_3781);
xor U5085 (N_5085,N_3338,N_2995);
nor U5086 (N_5086,N_3537,N_3930);
nand U5087 (N_5087,N_2951,N_3513);
or U5088 (N_5088,N_2604,N_2603);
xor U5089 (N_5089,N_2985,N_3095);
or U5090 (N_5090,N_2959,N_3861);
xor U5091 (N_5091,N_3873,N_3830);
nor U5092 (N_5092,N_2944,N_3425);
nand U5093 (N_5093,N_2012,N_2385);
nor U5094 (N_5094,N_3236,N_2373);
or U5095 (N_5095,N_3622,N_2662);
nand U5096 (N_5096,N_2348,N_3055);
xor U5097 (N_5097,N_2973,N_2266);
xnor U5098 (N_5098,N_2761,N_2227);
and U5099 (N_5099,N_3832,N_2264);
xor U5100 (N_5100,N_3532,N_3667);
and U5101 (N_5101,N_2223,N_2438);
nor U5102 (N_5102,N_2118,N_2586);
nand U5103 (N_5103,N_3912,N_2318);
nor U5104 (N_5104,N_3572,N_3494);
and U5105 (N_5105,N_2805,N_3637);
xnor U5106 (N_5106,N_3374,N_3267);
xor U5107 (N_5107,N_3612,N_3089);
xor U5108 (N_5108,N_2146,N_3468);
nor U5109 (N_5109,N_2836,N_3001);
nand U5110 (N_5110,N_3908,N_3440);
and U5111 (N_5111,N_2824,N_3514);
or U5112 (N_5112,N_3897,N_2251);
xor U5113 (N_5113,N_2200,N_2731);
and U5114 (N_5114,N_3676,N_2193);
nor U5115 (N_5115,N_2575,N_3665);
xor U5116 (N_5116,N_2628,N_2262);
or U5117 (N_5117,N_2345,N_3920);
nor U5118 (N_5118,N_2400,N_3155);
and U5119 (N_5119,N_2302,N_3018);
xnor U5120 (N_5120,N_3573,N_3322);
or U5121 (N_5121,N_3590,N_3091);
nand U5122 (N_5122,N_2577,N_3938);
nor U5123 (N_5123,N_2086,N_2119);
nor U5124 (N_5124,N_2332,N_3434);
or U5125 (N_5125,N_3079,N_3213);
nand U5126 (N_5126,N_2730,N_2182);
nand U5127 (N_5127,N_2685,N_3667);
xnor U5128 (N_5128,N_2580,N_2937);
nor U5129 (N_5129,N_2650,N_2588);
nor U5130 (N_5130,N_2868,N_3169);
nand U5131 (N_5131,N_3146,N_3479);
and U5132 (N_5132,N_3120,N_2524);
nor U5133 (N_5133,N_2458,N_2692);
nor U5134 (N_5134,N_2129,N_2015);
xnor U5135 (N_5135,N_2754,N_2370);
xor U5136 (N_5136,N_3567,N_3189);
xnor U5137 (N_5137,N_3954,N_3167);
and U5138 (N_5138,N_3358,N_2408);
nor U5139 (N_5139,N_2953,N_3088);
and U5140 (N_5140,N_3859,N_3754);
nand U5141 (N_5141,N_2335,N_3052);
nand U5142 (N_5142,N_3936,N_3409);
and U5143 (N_5143,N_3303,N_2888);
nand U5144 (N_5144,N_2345,N_3767);
and U5145 (N_5145,N_3308,N_2308);
nand U5146 (N_5146,N_3057,N_3395);
or U5147 (N_5147,N_2294,N_3087);
and U5148 (N_5148,N_2581,N_2400);
nor U5149 (N_5149,N_2991,N_2658);
or U5150 (N_5150,N_2503,N_3023);
xor U5151 (N_5151,N_2601,N_2703);
xor U5152 (N_5152,N_3597,N_2951);
nand U5153 (N_5153,N_3735,N_2678);
nand U5154 (N_5154,N_2087,N_3951);
or U5155 (N_5155,N_2961,N_3638);
nand U5156 (N_5156,N_2474,N_2459);
and U5157 (N_5157,N_3479,N_2446);
xor U5158 (N_5158,N_2822,N_2118);
xor U5159 (N_5159,N_2557,N_2780);
xnor U5160 (N_5160,N_3443,N_3258);
or U5161 (N_5161,N_3089,N_3447);
nor U5162 (N_5162,N_2736,N_2429);
nor U5163 (N_5163,N_2401,N_2425);
nand U5164 (N_5164,N_2062,N_3310);
or U5165 (N_5165,N_3110,N_2235);
and U5166 (N_5166,N_2941,N_2835);
or U5167 (N_5167,N_2156,N_3722);
nor U5168 (N_5168,N_2790,N_3986);
nor U5169 (N_5169,N_2089,N_2047);
or U5170 (N_5170,N_3021,N_2535);
or U5171 (N_5171,N_3085,N_3022);
or U5172 (N_5172,N_2043,N_3271);
and U5173 (N_5173,N_3938,N_2643);
xor U5174 (N_5174,N_3273,N_2728);
nor U5175 (N_5175,N_3779,N_3730);
or U5176 (N_5176,N_3726,N_2639);
or U5177 (N_5177,N_3439,N_3630);
or U5178 (N_5178,N_3287,N_3403);
or U5179 (N_5179,N_2063,N_2986);
or U5180 (N_5180,N_3058,N_3509);
and U5181 (N_5181,N_2544,N_2498);
nor U5182 (N_5182,N_2962,N_2977);
xor U5183 (N_5183,N_2189,N_2429);
and U5184 (N_5184,N_2546,N_2001);
xor U5185 (N_5185,N_3235,N_2967);
xor U5186 (N_5186,N_3776,N_2820);
nor U5187 (N_5187,N_2319,N_2347);
or U5188 (N_5188,N_3725,N_3304);
nand U5189 (N_5189,N_2770,N_3239);
or U5190 (N_5190,N_2720,N_2895);
and U5191 (N_5191,N_3939,N_2941);
nand U5192 (N_5192,N_2988,N_2400);
or U5193 (N_5193,N_3882,N_3131);
nor U5194 (N_5194,N_2996,N_3679);
xnor U5195 (N_5195,N_2698,N_3501);
nor U5196 (N_5196,N_2184,N_2375);
or U5197 (N_5197,N_3875,N_3842);
or U5198 (N_5198,N_3259,N_2554);
and U5199 (N_5199,N_2211,N_2031);
nand U5200 (N_5200,N_2177,N_3359);
and U5201 (N_5201,N_2581,N_3176);
xor U5202 (N_5202,N_2104,N_2179);
and U5203 (N_5203,N_2971,N_3938);
nor U5204 (N_5204,N_3399,N_2395);
xnor U5205 (N_5205,N_3766,N_3638);
and U5206 (N_5206,N_3762,N_2121);
and U5207 (N_5207,N_2511,N_3749);
nor U5208 (N_5208,N_3353,N_3499);
xnor U5209 (N_5209,N_2497,N_2495);
or U5210 (N_5210,N_2507,N_2043);
nand U5211 (N_5211,N_3048,N_2095);
and U5212 (N_5212,N_2038,N_2876);
nand U5213 (N_5213,N_2229,N_3987);
and U5214 (N_5214,N_2167,N_3680);
nor U5215 (N_5215,N_3082,N_3081);
nand U5216 (N_5216,N_2070,N_3880);
or U5217 (N_5217,N_2579,N_3529);
or U5218 (N_5218,N_3067,N_2308);
or U5219 (N_5219,N_2008,N_3164);
and U5220 (N_5220,N_3736,N_3358);
xor U5221 (N_5221,N_2251,N_3420);
or U5222 (N_5222,N_2743,N_3339);
xor U5223 (N_5223,N_3981,N_3097);
nand U5224 (N_5224,N_3900,N_3453);
nand U5225 (N_5225,N_3537,N_2419);
xnor U5226 (N_5226,N_3012,N_3435);
xor U5227 (N_5227,N_2506,N_3628);
or U5228 (N_5228,N_3418,N_2521);
nand U5229 (N_5229,N_3086,N_2698);
nor U5230 (N_5230,N_3508,N_3463);
xor U5231 (N_5231,N_2954,N_3259);
nand U5232 (N_5232,N_2813,N_3299);
nand U5233 (N_5233,N_2209,N_3595);
or U5234 (N_5234,N_3659,N_2443);
nand U5235 (N_5235,N_2128,N_2763);
and U5236 (N_5236,N_3592,N_2310);
nand U5237 (N_5237,N_2147,N_3899);
or U5238 (N_5238,N_3751,N_3937);
nor U5239 (N_5239,N_2489,N_2693);
nor U5240 (N_5240,N_3058,N_2931);
nor U5241 (N_5241,N_3412,N_3606);
xnor U5242 (N_5242,N_2580,N_2950);
xnor U5243 (N_5243,N_3536,N_2209);
xnor U5244 (N_5244,N_2697,N_2446);
or U5245 (N_5245,N_3264,N_2158);
xnor U5246 (N_5246,N_3714,N_2670);
and U5247 (N_5247,N_3221,N_3821);
nor U5248 (N_5248,N_2410,N_3341);
nor U5249 (N_5249,N_3364,N_2149);
and U5250 (N_5250,N_3881,N_2840);
nor U5251 (N_5251,N_2976,N_2439);
nand U5252 (N_5252,N_3180,N_2489);
nor U5253 (N_5253,N_3643,N_3578);
nand U5254 (N_5254,N_2893,N_3881);
nor U5255 (N_5255,N_2232,N_2904);
nand U5256 (N_5256,N_2888,N_2763);
nand U5257 (N_5257,N_2535,N_2000);
nand U5258 (N_5258,N_3181,N_3872);
or U5259 (N_5259,N_3240,N_3405);
and U5260 (N_5260,N_2311,N_2407);
and U5261 (N_5261,N_2740,N_3128);
xor U5262 (N_5262,N_3730,N_2172);
nand U5263 (N_5263,N_2806,N_2860);
or U5264 (N_5264,N_2989,N_3974);
xnor U5265 (N_5265,N_3035,N_2735);
nor U5266 (N_5266,N_3904,N_3959);
xnor U5267 (N_5267,N_2192,N_3130);
or U5268 (N_5268,N_3636,N_3131);
or U5269 (N_5269,N_2296,N_3907);
xor U5270 (N_5270,N_2162,N_3132);
nand U5271 (N_5271,N_3782,N_2791);
nor U5272 (N_5272,N_3451,N_3886);
or U5273 (N_5273,N_3339,N_2411);
or U5274 (N_5274,N_3296,N_2873);
nor U5275 (N_5275,N_3113,N_3134);
xnor U5276 (N_5276,N_2278,N_2657);
nor U5277 (N_5277,N_2590,N_2077);
xnor U5278 (N_5278,N_2867,N_2172);
nand U5279 (N_5279,N_3625,N_2698);
xnor U5280 (N_5280,N_3522,N_2646);
nand U5281 (N_5281,N_3497,N_3573);
or U5282 (N_5282,N_2303,N_2142);
or U5283 (N_5283,N_2496,N_3331);
or U5284 (N_5284,N_3434,N_2045);
or U5285 (N_5285,N_3561,N_2025);
xor U5286 (N_5286,N_2245,N_2962);
and U5287 (N_5287,N_3768,N_2364);
xnor U5288 (N_5288,N_3031,N_3194);
nor U5289 (N_5289,N_3820,N_2090);
xnor U5290 (N_5290,N_3680,N_3370);
nand U5291 (N_5291,N_3421,N_3112);
or U5292 (N_5292,N_3928,N_3926);
or U5293 (N_5293,N_2501,N_2207);
and U5294 (N_5294,N_3658,N_3412);
xnor U5295 (N_5295,N_3337,N_2623);
nand U5296 (N_5296,N_3869,N_3626);
nor U5297 (N_5297,N_3136,N_2500);
xor U5298 (N_5298,N_3822,N_2012);
nor U5299 (N_5299,N_3386,N_3785);
xor U5300 (N_5300,N_3986,N_3914);
xnor U5301 (N_5301,N_2546,N_3428);
and U5302 (N_5302,N_2164,N_2373);
nor U5303 (N_5303,N_2572,N_2915);
nor U5304 (N_5304,N_3555,N_2070);
and U5305 (N_5305,N_2035,N_2405);
xor U5306 (N_5306,N_2480,N_3891);
nand U5307 (N_5307,N_3934,N_2122);
and U5308 (N_5308,N_2795,N_3722);
xor U5309 (N_5309,N_3505,N_3553);
nand U5310 (N_5310,N_2934,N_2981);
xnor U5311 (N_5311,N_2934,N_2168);
xnor U5312 (N_5312,N_3115,N_3064);
nand U5313 (N_5313,N_3343,N_2883);
and U5314 (N_5314,N_2538,N_2242);
nand U5315 (N_5315,N_2095,N_2782);
and U5316 (N_5316,N_2993,N_2236);
and U5317 (N_5317,N_2808,N_2419);
nor U5318 (N_5318,N_2243,N_3991);
or U5319 (N_5319,N_2667,N_2719);
or U5320 (N_5320,N_3875,N_3822);
or U5321 (N_5321,N_2254,N_2238);
or U5322 (N_5322,N_3724,N_3773);
xor U5323 (N_5323,N_3971,N_3999);
nand U5324 (N_5324,N_3757,N_3217);
and U5325 (N_5325,N_3744,N_2280);
xor U5326 (N_5326,N_2956,N_2710);
or U5327 (N_5327,N_2745,N_2553);
and U5328 (N_5328,N_3793,N_2846);
or U5329 (N_5329,N_2791,N_3464);
nor U5330 (N_5330,N_2163,N_2600);
nand U5331 (N_5331,N_3167,N_3407);
xnor U5332 (N_5332,N_3224,N_2050);
or U5333 (N_5333,N_3304,N_3583);
or U5334 (N_5334,N_3571,N_3113);
nand U5335 (N_5335,N_3335,N_2036);
xnor U5336 (N_5336,N_2891,N_2631);
xnor U5337 (N_5337,N_3470,N_2436);
nand U5338 (N_5338,N_3961,N_3584);
nor U5339 (N_5339,N_3124,N_2587);
or U5340 (N_5340,N_2230,N_3157);
or U5341 (N_5341,N_3315,N_3100);
nand U5342 (N_5342,N_2585,N_2055);
or U5343 (N_5343,N_2194,N_2642);
xnor U5344 (N_5344,N_3357,N_2017);
xor U5345 (N_5345,N_3494,N_3613);
and U5346 (N_5346,N_2429,N_3525);
xor U5347 (N_5347,N_2121,N_3443);
nand U5348 (N_5348,N_3493,N_3546);
nor U5349 (N_5349,N_3387,N_2635);
xnor U5350 (N_5350,N_3477,N_3853);
nand U5351 (N_5351,N_2559,N_2252);
xnor U5352 (N_5352,N_2351,N_2102);
nand U5353 (N_5353,N_2847,N_3775);
xor U5354 (N_5354,N_2229,N_2998);
or U5355 (N_5355,N_3214,N_3135);
and U5356 (N_5356,N_2933,N_3367);
or U5357 (N_5357,N_3598,N_3676);
nand U5358 (N_5358,N_2931,N_2813);
nand U5359 (N_5359,N_3263,N_2788);
nor U5360 (N_5360,N_3831,N_3897);
nand U5361 (N_5361,N_3861,N_2806);
and U5362 (N_5362,N_3600,N_3387);
or U5363 (N_5363,N_3539,N_3548);
nor U5364 (N_5364,N_3691,N_3549);
nand U5365 (N_5365,N_3104,N_2854);
xor U5366 (N_5366,N_2829,N_2798);
nand U5367 (N_5367,N_3291,N_3753);
nor U5368 (N_5368,N_2463,N_3372);
xor U5369 (N_5369,N_2661,N_2823);
or U5370 (N_5370,N_2566,N_2239);
nor U5371 (N_5371,N_2663,N_2743);
and U5372 (N_5372,N_3954,N_3890);
nand U5373 (N_5373,N_2856,N_2253);
nor U5374 (N_5374,N_3676,N_3617);
nand U5375 (N_5375,N_3806,N_2907);
nand U5376 (N_5376,N_2636,N_3770);
or U5377 (N_5377,N_3175,N_3100);
and U5378 (N_5378,N_3879,N_2962);
xnor U5379 (N_5379,N_2934,N_2290);
and U5380 (N_5380,N_3788,N_3125);
xnor U5381 (N_5381,N_2751,N_3365);
nand U5382 (N_5382,N_3715,N_3643);
nor U5383 (N_5383,N_2527,N_3670);
nand U5384 (N_5384,N_3664,N_2381);
xor U5385 (N_5385,N_2925,N_3107);
nand U5386 (N_5386,N_3737,N_2465);
or U5387 (N_5387,N_2562,N_2556);
nand U5388 (N_5388,N_2962,N_2128);
nand U5389 (N_5389,N_2774,N_2903);
or U5390 (N_5390,N_3247,N_2783);
nor U5391 (N_5391,N_3454,N_2247);
nand U5392 (N_5392,N_2601,N_3976);
nor U5393 (N_5393,N_2928,N_3208);
xor U5394 (N_5394,N_2067,N_3672);
nor U5395 (N_5395,N_3741,N_3152);
and U5396 (N_5396,N_2653,N_2508);
or U5397 (N_5397,N_3372,N_2132);
nand U5398 (N_5398,N_2122,N_3444);
xor U5399 (N_5399,N_3754,N_2120);
nor U5400 (N_5400,N_2387,N_3740);
and U5401 (N_5401,N_3194,N_2227);
nor U5402 (N_5402,N_2510,N_2480);
or U5403 (N_5403,N_3957,N_3552);
xor U5404 (N_5404,N_3376,N_3290);
xnor U5405 (N_5405,N_3774,N_3643);
nand U5406 (N_5406,N_2939,N_2799);
xor U5407 (N_5407,N_3727,N_2434);
xnor U5408 (N_5408,N_3811,N_2189);
xnor U5409 (N_5409,N_3500,N_3789);
nand U5410 (N_5410,N_2417,N_2737);
and U5411 (N_5411,N_2784,N_3185);
xnor U5412 (N_5412,N_2210,N_2503);
nand U5413 (N_5413,N_2802,N_3802);
and U5414 (N_5414,N_2192,N_2613);
xor U5415 (N_5415,N_3941,N_3917);
and U5416 (N_5416,N_2926,N_3477);
nand U5417 (N_5417,N_2331,N_2497);
xnor U5418 (N_5418,N_3457,N_2936);
nand U5419 (N_5419,N_2593,N_2311);
nor U5420 (N_5420,N_3970,N_3067);
and U5421 (N_5421,N_3786,N_3100);
or U5422 (N_5422,N_2685,N_2363);
nor U5423 (N_5423,N_3629,N_2510);
nand U5424 (N_5424,N_2795,N_2439);
nor U5425 (N_5425,N_2862,N_3210);
or U5426 (N_5426,N_2766,N_2486);
xor U5427 (N_5427,N_3209,N_3142);
xor U5428 (N_5428,N_3841,N_2501);
nand U5429 (N_5429,N_3746,N_3145);
nor U5430 (N_5430,N_2491,N_2313);
and U5431 (N_5431,N_2209,N_3594);
and U5432 (N_5432,N_2687,N_2738);
nand U5433 (N_5433,N_2753,N_2416);
or U5434 (N_5434,N_2804,N_2507);
or U5435 (N_5435,N_3112,N_2088);
or U5436 (N_5436,N_3129,N_2478);
or U5437 (N_5437,N_3016,N_2186);
nand U5438 (N_5438,N_3373,N_2715);
nor U5439 (N_5439,N_3290,N_2797);
nor U5440 (N_5440,N_2488,N_2519);
or U5441 (N_5441,N_2601,N_2330);
or U5442 (N_5442,N_3272,N_3487);
nor U5443 (N_5443,N_2545,N_3462);
xnor U5444 (N_5444,N_3187,N_2730);
or U5445 (N_5445,N_3147,N_3924);
nor U5446 (N_5446,N_3956,N_2797);
nor U5447 (N_5447,N_3188,N_2252);
or U5448 (N_5448,N_2656,N_2785);
or U5449 (N_5449,N_3241,N_2177);
nand U5450 (N_5450,N_3067,N_2716);
nand U5451 (N_5451,N_3806,N_2195);
or U5452 (N_5452,N_3615,N_3013);
and U5453 (N_5453,N_3716,N_2542);
and U5454 (N_5454,N_3183,N_3095);
nand U5455 (N_5455,N_3488,N_3263);
nand U5456 (N_5456,N_2917,N_2470);
nor U5457 (N_5457,N_2240,N_2644);
and U5458 (N_5458,N_2823,N_3039);
nor U5459 (N_5459,N_2555,N_3442);
nor U5460 (N_5460,N_3078,N_3277);
nor U5461 (N_5461,N_3751,N_2578);
and U5462 (N_5462,N_2264,N_2262);
nor U5463 (N_5463,N_2848,N_3137);
nor U5464 (N_5464,N_3549,N_3351);
xor U5465 (N_5465,N_3477,N_3601);
and U5466 (N_5466,N_2602,N_3926);
and U5467 (N_5467,N_3221,N_2353);
xor U5468 (N_5468,N_2258,N_3900);
and U5469 (N_5469,N_3319,N_3581);
nor U5470 (N_5470,N_2947,N_3087);
nor U5471 (N_5471,N_2123,N_3542);
or U5472 (N_5472,N_3263,N_2621);
xnor U5473 (N_5473,N_3620,N_2231);
and U5474 (N_5474,N_2884,N_3007);
or U5475 (N_5475,N_2099,N_3741);
and U5476 (N_5476,N_3937,N_3852);
xor U5477 (N_5477,N_2457,N_3872);
xnor U5478 (N_5478,N_2538,N_3647);
and U5479 (N_5479,N_2541,N_3505);
xnor U5480 (N_5480,N_2393,N_2396);
nor U5481 (N_5481,N_2265,N_3310);
or U5482 (N_5482,N_2719,N_2852);
nand U5483 (N_5483,N_3619,N_3758);
nor U5484 (N_5484,N_3760,N_2135);
nor U5485 (N_5485,N_3925,N_2880);
nand U5486 (N_5486,N_3676,N_2180);
nand U5487 (N_5487,N_2991,N_3871);
xnor U5488 (N_5488,N_3422,N_2516);
or U5489 (N_5489,N_3449,N_2864);
xnor U5490 (N_5490,N_2698,N_3995);
nand U5491 (N_5491,N_2447,N_2804);
or U5492 (N_5492,N_2053,N_3320);
xor U5493 (N_5493,N_2938,N_3268);
nor U5494 (N_5494,N_3033,N_3326);
and U5495 (N_5495,N_3751,N_2315);
nand U5496 (N_5496,N_2958,N_2154);
nand U5497 (N_5497,N_2415,N_3723);
and U5498 (N_5498,N_3377,N_3597);
nand U5499 (N_5499,N_3172,N_3380);
xor U5500 (N_5500,N_2370,N_3414);
nor U5501 (N_5501,N_2797,N_3016);
and U5502 (N_5502,N_3970,N_2435);
nand U5503 (N_5503,N_2707,N_2215);
nor U5504 (N_5504,N_2033,N_2868);
and U5505 (N_5505,N_2509,N_3250);
and U5506 (N_5506,N_3943,N_3298);
nor U5507 (N_5507,N_3904,N_3375);
xnor U5508 (N_5508,N_2082,N_2906);
or U5509 (N_5509,N_2342,N_3394);
nor U5510 (N_5510,N_3254,N_3845);
xnor U5511 (N_5511,N_3444,N_2222);
or U5512 (N_5512,N_2970,N_3171);
nor U5513 (N_5513,N_2897,N_3645);
and U5514 (N_5514,N_2856,N_2729);
and U5515 (N_5515,N_2171,N_2608);
nor U5516 (N_5516,N_2650,N_2570);
and U5517 (N_5517,N_2441,N_3639);
and U5518 (N_5518,N_2893,N_2044);
nor U5519 (N_5519,N_2877,N_3865);
xor U5520 (N_5520,N_2137,N_2140);
and U5521 (N_5521,N_2742,N_3193);
or U5522 (N_5522,N_3412,N_2245);
and U5523 (N_5523,N_3946,N_3045);
xor U5524 (N_5524,N_2572,N_3044);
xnor U5525 (N_5525,N_2641,N_3120);
and U5526 (N_5526,N_3171,N_2027);
nand U5527 (N_5527,N_3038,N_2392);
and U5528 (N_5528,N_2752,N_2367);
or U5529 (N_5529,N_2301,N_3827);
nor U5530 (N_5530,N_3719,N_3456);
nand U5531 (N_5531,N_3338,N_3556);
and U5532 (N_5532,N_3957,N_2991);
xor U5533 (N_5533,N_2611,N_2301);
or U5534 (N_5534,N_3301,N_2134);
nand U5535 (N_5535,N_3671,N_2758);
nor U5536 (N_5536,N_3300,N_2425);
and U5537 (N_5537,N_3675,N_2627);
nor U5538 (N_5538,N_2610,N_3413);
or U5539 (N_5539,N_3390,N_2103);
and U5540 (N_5540,N_2122,N_2916);
nand U5541 (N_5541,N_2712,N_3720);
nor U5542 (N_5542,N_2762,N_3407);
nor U5543 (N_5543,N_3651,N_2705);
nand U5544 (N_5544,N_3172,N_3946);
nor U5545 (N_5545,N_3550,N_2245);
xnor U5546 (N_5546,N_2954,N_2874);
nor U5547 (N_5547,N_2136,N_2747);
or U5548 (N_5548,N_2553,N_2297);
nor U5549 (N_5549,N_3085,N_2521);
nor U5550 (N_5550,N_2134,N_2627);
xnor U5551 (N_5551,N_2562,N_2233);
nand U5552 (N_5552,N_3217,N_2869);
nand U5553 (N_5553,N_3208,N_2608);
nand U5554 (N_5554,N_2622,N_3131);
or U5555 (N_5555,N_2225,N_3302);
and U5556 (N_5556,N_3018,N_3026);
xor U5557 (N_5557,N_3043,N_3625);
and U5558 (N_5558,N_2277,N_2883);
or U5559 (N_5559,N_3415,N_2158);
and U5560 (N_5560,N_2790,N_2916);
nor U5561 (N_5561,N_2888,N_2399);
or U5562 (N_5562,N_3708,N_2133);
and U5563 (N_5563,N_3519,N_2489);
or U5564 (N_5564,N_3761,N_3387);
xor U5565 (N_5565,N_3257,N_3351);
and U5566 (N_5566,N_3901,N_2928);
nor U5567 (N_5567,N_2197,N_2775);
nand U5568 (N_5568,N_2284,N_3315);
and U5569 (N_5569,N_2288,N_2947);
or U5570 (N_5570,N_3609,N_3039);
nand U5571 (N_5571,N_3626,N_2385);
xor U5572 (N_5572,N_3280,N_3054);
xor U5573 (N_5573,N_2824,N_2373);
nand U5574 (N_5574,N_3532,N_2264);
and U5575 (N_5575,N_2034,N_3564);
xnor U5576 (N_5576,N_2385,N_2519);
and U5577 (N_5577,N_2037,N_2174);
or U5578 (N_5578,N_3629,N_2841);
and U5579 (N_5579,N_2536,N_2291);
nor U5580 (N_5580,N_2706,N_3837);
xor U5581 (N_5581,N_3816,N_2402);
nor U5582 (N_5582,N_2463,N_3611);
or U5583 (N_5583,N_3363,N_3620);
nor U5584 (N_5584,N_3631,N_3729);
nor U5585 (N_5585,N_3801,N_3093);
and U5586 (N_5586,N_2012,N_2072);
and U5587 (N_5587,N_3825,N_3529);
or U5588 (N_5588,N_2695,N_2356);
nor U5589 (N_5589,N_2675,N_3043);
nor U5590 (N_5590,N_3627,N_2615);
or U5591 (N_5591,N_3922,N_3691);
nor U5592 (N_5592,N_3457,N_2237);
and U5593 (N_5593,N_2851,N_2539);
or U5594 (N_5594,N_3480,N_2686);
xor U5595 (N_5595,N_3485,N_2722);
and U5596 (N_5596,N_2691,N_2851);
nor U5597 (N_5597,N_2406,N_2388);
nor U5598 (N_5598,N_2111,N_2598);
xor U5599 (N_5599,N_3906,N_2191);
nand U5600 (N_5600,N_2633,N_3072);
nand U5601 (N_5601,N_2248,N_3769);
or U5602 (N_5602,N_2869,N_3158);
xnor U5603 (N_5603,N_3434,N_2308);
xnor U5604 (N_5604,N_3349,N_2335);
xor U5605 (N_5605,N_3193,N_3508);
xnor U5606 (N_5606,N_3212,N_3404);
nor U5607 (N_5607,N_3664,N_3079);
xor U5608 (N_5608,N_3619,N_3158);
and U5609 (N_5609,N_3459,N_2605);
nor U5610 (N_5610,N_3768,N_2165);
or U5611 (N_5611,N_3339,N_2479);
or U5612 (N_5612,N_2709,N_3395);
nand U5613 (N_5613,N_2359,N_3494);
or U5614 (N_5614,N_2582,N_2646);
nand U5615 (N_5615,N_2334,N_2074);
xnor U5616 (N_5616,N_2840,N_2536);
xor U5617 (N_5617,N_3927,N_2413);
nor U5618 (N_5618,N_2184,N_3200);
xor U5619 (N_5619,N_2120,N_3365);
xor U5620 (N_5620,N_3173,N_3278);
nor U5621 (N_5621,N_3128,N_3666);
and U5622 (N_5622,N_3480,N_2537);
xor U5623 (N_5623,N_3384,N_2339);
xor U5624 (N_5624,N_3084,N_3785);
nand U5625 (N_5625,N_3101,N_3296);
or U5626 (N_5626,N_2364,N_2170);
nand U5627 (N_5627,N_2636,N_3813);
or U5628 (N_5628,N_3606,N_3478);
and U5629 (N_5629,N_2765,N_2317);
and U5630 (N_5630,N_2700,N_2187);
xnor U5631 (N_5631,N_2267,N_3988);
nand U5632 (N_5632,N_2257,N_2169);
nand U5633 (N_5633,N_3113,N_3204);
xnor U5634 (N_5634,N_3555,N_3355);
nand U5635 (N_5635,N_3141,N_2152);
xnor U5636 (N_5636,N_3496,N_3751);
and U5637 (N_5637,N_2189,N_2843);
and U5638 (N_5638,N_3778,N_3360);
or U5639 (N_5639,N_3829,N_3313);
nand U5640 (N_5640,N_2357,N_2429);
and U5641 (N_5641,N_2614,N_2731);
and U5642 (N_5642,N_2945,N_3236);
nand U5643 (N_5643,N_2283,N_2057);
or U5644 (N_5644,N_2736,N_2086);
nor U5645 (N_5645,N_3276,N_2922);
nand U5646 (N_5646,N_3814,N_3959);
xor U5647 (N_5647,N_2893,N_2757);
and U5648 (N_5648,N_2407,N_3044);
and U5649 (N_5649,N_2933,N_2658);
nor U5650 (N_5650,N_2454,N_3047);
or U5651 (N_5651,N_2503,N_2742);
xnor U5652 (N_5652,N_3282,N_2857);
nand U5653 (N_5653,N_2352,N_3055);
nor U5654 (N_5654,N_2830,N_2586);
nand U5655 (N_5655,N_3146,N_2058);
or U5656 (N_5656,N_2257,N_3879);
or U5657 (N_5657,N_3531,N_2680);
and U5658 (N_5658,N_3495,N_3365);
and U5659 (N_5659,N_2894,N_2718);
nor U5660 (N_5660,N_3711,N_2403);
and U5661 (N_5661,N_2978,N_2957);
xor U5662 (N_5662,N_3004,N_2226);
nand U5663 (N_5663,N_2937,N_3888);
xor U5664 (N_5664,N_2588,N_3071);
nor U5665 (N_5665,N_2946,N_2309);
and U5666 (N_5666,N_3011,N_2373);
nand U5667 (N_5667,N_3599,N_3791);
or U5668 (N_5668,N_3728,N_2916);
nand U5669 (N_5669,N_3549,N_2551);
xnor U5670 (N_5670,N_2744,N_2549);
nor U5671 (N_5671,N_2627,N_3309);
or U5672 (N_5672,N_2627,N_3203);
and U5673 (N_5673,N_3037,N_2501);
nand U5674 (N_5674,N_2240,N_2514);
nand U5675 (N_5675,N_2213,N_2606);
or U5676 (N_5676,N_3245,N_2483);
nand U5677 (N_5677,N_2578,N_2327);
nand U5678 (N_5678,N_3931,N_2329);
xor U5679 (N_5679,N_3384,N_3131);
xnor U5680 (N_5680,N_3380,N_3154);
and U5681 (N_5681,N_2557,N_2179);
or U5682 (N_5682,N_3461,N_2068);
xor U5683 (N_5683,N_2145,N_3800);
and U5684 (N_5684,N_2700,N_3979);
or U5685 (N_5685,N_3818,N_3832);
xnor U5686 (N_5686,N_3937,N_3991);
and U5687 (N_5687,N_2163,N_3296);
nand U5688 (N_5688,N_3991,N_2336);
and U5689 (N_5689,N_3469,N_3247);
nand U5690 (N_5690,N_3399,N_3409);
xor U5691 (N_5691,N_3683,N_2114);
or U5692 (N_5692,N_3050,N_2328);
and U5693 (N_5693,N_2497,N_2511);
and U5694 (N_5694,N_2049,N_3598);
xnor U5695 (N_5695,N_3372,N_2722);
and U5696 (N_5696,N_2064,N_2962);
xor U5697 (N_5697,N_2866,N_2893);
or U5698 (N_5698,N_2716,N_2811);
or U5699 (N_5699,N_2521,N_2365);
nand U5700 (N_5700,N_3616,N_3259);
nand U5701 (N_5701,N_2442,N_2540);
and U5702 (N_5702,N_2843,N_3121);
xor U5703 (N_5703,N_2066,N_3935);
nor U5704 (N_5704,N_2497,N_3616);
nand U5705 (N_5705,N_2219,N_2114);
and U5706 (N_5706,N_3202,N_3704);
nand U5707 (N_5707,N_3940,N_2312);
and U5708 (N_5708,N_3122,N_3537);
and U5709 (N_5709,N_2517,N_3033);
and U5710 (N_5710,N_3225,N_2448);
and U5711 (N_5711,N_3544,N_3960);
and U5712 (N_5712,N_2060,N_3686);
nor U5713 (N_5713,N_3877,N_2020);
xor U5714 (N_5714,N_3251,N_2160);
xnor U5715 (N_5715,N_3797,N_2796);
and U5716 (N_5716,N_3610,N_2044);
and U5717 (N_5717,N_2557,N_2696);
and U5718 (N_5718,N_2925,N_3707);
nand U5719 (N_5719,N_3249,N_3518);
and U5720 (N_5720,N_3397,N_3382);
or U5721 (N_5721,N_3210,N_2320);
and U5722 (N_5722,N_3891,N_3376);
nor U5723 (N_5723,N_3293,N_3042);
nor U5724 (N_5724,N_3472,N_3444);
or U5725 (N_5725,N_2853,N_3263);
or U5726 (N_5726,N_2123,N_3608);
nand U5727 (N_5727,N_2594,N_3695);
xnor U5728 (N_5728,N_3454,N_2388);
nor U5729 (N_5729,N_3929,N_3902);
nand U5730 (N_5730,N_2585,N_2803);
nand U5731 (N_5731,N_3473,N_3728);
xnor U5732 (N_5732,N_2473,N_2874);
xnor U5733 (N_5733,N_2801,N_3429);
and U5734 (N_5734,N_2955,N_3429);
or U5735 (N_5735,N_3250,N_2018);
xor U5736 (N_5736,N_3022,N_2238);
and U5737 (N_5737,N_3264,N_2704);
nor U5738 (N_5738,N_3178,N_2642);
nand U5739 (N_5739,N_3431,N_3516);
and U5740 (N_5740,N_2209,N_2002);
nand U5741 (N_5741,N_3951,N_2880);
nor U5742 (N_5742,N_3806,N_2935);
or U5743 (N_5743,N_3191,N_2142);
and U5744 (N_5744,N_3404,N_2702);
nand U5745 (N_5745,N_2622,N_2960);
and U5746 (N_5746,N_2641,N_3099);
and U5747 (N_5747,N_3394,N_2316);
xnor U5748 (N_5748,N_2304,N_2782);
or U5749 (N_5749,N_2723,N_3656);
or U5750 (N_5750,N_2222,N_2013);
and U5751 (N_5751,N_2560,N_3697);
nand U5752 (N_5752,N_3296,N_3235);
nor U5753 (N_5753,N_3368,N_2319);
xnor U5754 (N_5754,N_2737,N_2935);
xor U5755 (N_5755,N_3166,N_3476);
nor U5756 (N_5756,N_2625,N_2178);
and U5757 (N_5757,N_3277,N_3002);
and U5758 (N_5758,N_3649,N_3054);
nor U5759 (N_5759,N_3737,N_2173);
nor U5760 (N_5760,N_2611,N_2199);
and U5761 (N_5761,N_2138,N_2123);
xor U5762 (N_5762,N_2851,N_3214);
nor U5763 (N_5763,N_2863,N_2426);
or U5764 (N_5764,N_3794,N_2131);
nand U5765 (N_5765,N_2307,N_3729);
and U5766 (N_5766,N_2420,N_3401);
and U5767 (N_5767,N_2740,N_2963);
nand U5768 (N_5768,N_3055,N_3990);
nand U5769 (N_5769,N_2707,N_3655);
nand U5770 (N_5770,N_3260,N_3810);
xor U5771 (N_5771,N_2433,N_3940);
nor U5772 (N_5772,N_2525,N_3232);
and U5773 (N_5773,N_2874,N_3881);
nor U5774 (N_5774,N_2615,N_2876);
xor U5775 (N_5775,N_3500,N_3262);
nor U5776 (N_5776,N_2694,N_3510);
and U5777 (N_5777,N_2772,N_3261);
and U5778 (N_5778,N_2012,N_3976);
nor U5779 (N_5779,N_2175,N_2769);
nor U5780 (N_5780,N_2053,N_3849);
xor U5781 (N_5781,N_3695,N_2376);
or U5782 (N_5782,N_2417,N_3634);
nor U5783 (N_5783,N_2322,N_2864);
nor U5784 (N_5784,N_3845,N_3283);
nand U5785 (N_5785,N_3389,N_2207);
nand U5786 (N_5786,N_2916,N_3109);
and U5787 (N_5787,N_3396,N_2972);
and U5788 (N_5788,N_2207,N_2181);
nand U5789 (N_5789,N_3127,N_2764);
or U5790 (N_5790,N_2805,N_2619);
or U5791 (N_5791,N_3657,N_3854);
nor U5792 (N_5792,N_3819,N_3244);
xor U5793 (N_5793,N_2739,N_3908);
nand U5794 (N_5794,N_2564,N_2326);
nor U5795 (N_5795,N_2453,N_2317);
or U5796 (N_5796,N_3717,N_2586);
nand U5797 (N_5797,N_3118,N_3147);
nor U5798 (N_5798,N_2121,N_2097);
or U5799 (N_5799,N_2297,N_2626);
nand U5800 (N_5800,N_3578,N_2820);
nand U5801 (N_5801,N_3814,N_3385);
or U5802 (N_5802,N_3424,N_2074);
xor U5803 (N_5803,N_2869,N_3002);
xnor U5804 (N_5804,N_2021,N_3968);
xnor U5805 (N_5805,N_3580,N_3225);
and U5806 (N_5806,N_3829,N_3638);
xnor U5807 (N_5807,N_2948,N_3792);
or U5808 (N_5808,N_3755,N_3174);
or U5809 (N_5809,N_2144,N_2059);
and U5810 (N_5810,N_2347,N_2535);
nand U5811 (N_5811,N_2441,N_3575);
or U5812 (N_5812,N_3968,N_3971);
or U5813 (N_5813,N_2621,N_2976);
and U5814 (N_5814,N_3156,N_3855);
and U5815 (N_5815,N_3881,N_3417);
nand U5816 (N_5816,N_3929,N_3380);
and U5817 (N_5817,N_2520,N_2326);
and U5818 (N_5818,N_3733,N_3597);
and U5819 (N_5819,N_3860,N_3601);
nor U5820 (N_5820,N_2439,N_3989);
and U5821 (N_5821,N_3368,N_2340);
nand U5822 (N_5822,N_2615,N_3992);
xnor U5823 (N_5823,N_2396,N_2763);
and U5824 (N_5824,N_3305,N_3245);
nor U5825 (N_5825,N_2355,N_3163);
nand U5826 (N_5826,N_3578,N_2153);
nand U5827 (N_5827,N_2531,N_3483);
and U5828 (N_5828,N_3966,N_2084);
xor U5829 (N_5829,N_2112,N_3224);
or U5830 (N_5830,N_3962,N_2171);
or U5831 (N_5831,N_3885,N_2916);
nor U5832 (N_5832,N_3818,N_3296);
and U5833 (N_5833,N_3979,N_3726);
and U5834 (N_5834,N_3945,N_2817);
or U5835 (N_5835,N_2815,N_3964);
nand U5836 (N_5836,N_2902,N_3408);
or U5837 (N_5837,N_3109,N_2721);
xnor U5838 (N_5838,N_3492,N_3595);
and U5839 (N_5839,N_2226,N_2434);
xnor U5840 (N_5840,N_2689,N_2267);
or U5841 (N_5841,N_2920,N_2084);
nand U5842 (N_5842,N_2374,N_3150);
xor U5843 (N_5843,N_2367,N_2654);
nand U5844 (N_5844,N_3222,N_3997);
nor U5845 (N_5845,N_2222,N_3214);
and U5846 (N_5846,N_2486,N_3219);
or U5847 (N_5847,N_3712,N_2694);
xnor U5848 (N_5848,N_2246,N_3660);
xor U5849 (N_5849,N_2785,N_2372);
and U5850 (N_5850,N_2722,N_2768);
and U5851 (N_5851,N_3032,N_3561);
nand U5852 (N_5852,N_2211,N_2318);
or U5853 (N_5853,N_2585,N_2744);
and U5854 (N_5854,N_3084,N_2325);
xor U5855 (N_5855,N_3609,N_3164);
nor U5856 (N_5856,N_2991,N_3091);
xor U5857 (N_5857,N_3071,N_3068);
xor U5858 (N_5858,N_2999,N_2902);
xnor U5859 (N_5859,N_2310,N_3547);
and U5860 (N_5860,N_3372,N_3991);
or U5861 (N_5861,N_3159,N_3920);
xnor U5862 (N_5862,N_3977,N_2016);
xnor U5863 (N_5863,N_3472,N_3609);
nand U5864 (N_5864,N_3093,N_2865);
or U5865 (N_5865,N_3773,N_2082);
and U5866 (N_5866,N_2883,N_3508);
and U5867 (N_5867,N_2036,N_2297);
and U5868 (N_5868,N_2841,N_2206);
nand U5869 (N_5869,N_3761,N_3894);
xnor U5870 (N_5870,N_3962,N_2857);
and U5871 (N_5871,N_2236,N_2788);
nand U5872 (N_5872,N_3659,N_2928);
nand U5873 (N_5873,N_2600,N_3612);
and U5874 (N_5874,N_2876,N_2879);
xor U5875 (N_5875,N_2073,N_2956);
xnor U5876 (N_5876,N_2702,N_3658);
and U5877 (N_5877,N_2826,N_2120);
or U5878 (N_5878,N_3329,N_2391);
nand U5879 (N_5879,N_3481,N_2622);
xor U5880 (N_5880,N_2763,N_3796);
nand U5881 (N_5881,N_2966,N_3579);
xor U5882 (N_5882,N_2139,N_2701);
and U5883 (N_5883,N_2189,N_2490);
nand U5884 (N_5884,N_2199,N_3217);
nand U5885 (N_5885,N_2456,N_3035);
or U5886 (N_5886,N_2911,N_2559);
or U5887 (N_5887,N_2343,N_3896);
and U5888 (N_5888,N_3529,N_3149);
or U5889 (N_5889,N_2499,N_3846);
or U5890 (N_5890,N_2563,N_3147);
nand U5891 (N_5891,N_2862,N_2672);
and U5892 (N_5892,N_3674,N_3974);
xor U5893 (N_5893,N_2195,N_2960);
nor U5894 (N_5894,N_3758,N_2940);
nor U5895 (N_5895,N_2511,N_2526);
nor U5896 (N_5896,N_2086,N_3596);
xor U5897 (N_5897,N_2757,N_2744);
nor U5898 (N_5898,N_2291,N_3704);
and U5899 (N_5899,N_3008,N_2133);
xor U5900 (N_5900,N_3243,N_2576);
and U5901 (N_5901,N_3170,N_2617);
and U5902 (N_5902,N_2866,N_2056);
nand U5903 (N_5903,N_3126,N_3475);
nand U5904 (N_5904,N_2274,N_3899);
nor U5905 (N_5905,N_2858,N_3145);
nand U5906 (N_5906,N_3837,N_3189);
xor U5907 (N_5907,N_3344,N_3517);
and U5908 (N_5908,N_2574,N_3057);
or U5909 (N_5909,N_2911,N_3171);
and U5910 (N_5910,N_2075,N_2399);
xnor U5911 (N_5911,N_3824,N_2775);
nor U5912 (N_5912,N_2485,N_3807);
or U5913 (N_5913,N_3062,N_3944);
and U5914 (N_5914,N_2557,N_2184);
nand U5915 (N_5915,N_3988,N_2212);
and U5916 (N_5916,N_2053,N_3196);
nand U5917 (N_5917,N_3028,N_3727);
nor U5918 (N_5918,N_3788,N_3219);
and U5919 (N_5919,N_3793,N_3558);
and U5920 (N_5920,N_3045,N_2197);
xnor U5921 (N_5921,N_2210,N_3514);
or U5922 (N_5922,N_3540,N_3686);
nor U5923 (N_5923,N_2738,N_3363);
nor U5924 (N_5924,N_2507,N_3460);
or U5925 (N_5925,N_2430,N_2547);
nand U5926 (N_5926,N_2239,N_3304);
xnor U5927 (N_5927,N_3778,N_2304);
nor U5928 (N_5928,N_2162,N_3894);
nand U5929 (N_5929,N_3988,N_3285);
nand U5930 (N_5930,N_3496,N_3649);
and U5931 (N_5931,N_3710,N_2753);
or U5932 (N_5932,N_3238,N_2748);
xor U5933 (N_5933,N_3885,N_3419);
and U5934 (N_5934,N_2010,N_2468);
or U5935 (N_5935,N_3682,N_2101);
nor U5936 (N_5936,N_3022,N_3114);
and U5937 (N_5937,N_3734,N_2753);
nand U5938 (N_5938,N_3468,N_3357);
nand U5939 (N_5939,N_2360,N_3547);
or U5940 (N_5940,N_2680,N_2938);
nand U5941 (N_5941,N_3615,N_3149);
or U5942 (N_5942,N_2242,N_2967);
nand U5943 (N_5943,N_3504,N_3819);
and U5944 (N_5944,N_3527,N_3149);
xnor U5945 (N_5945,N_2039,N_2685);
xnor U5946 (N_5946,N_2599,N_3575);
xnor U5947 (N_5947,N_3451,N_2782);
nand U5948 (N_5948,N_2454,N_3797);
or U5949 (N_5949,N_2799,N_2844);
xor U5950 (N_5950,N_3176,N_2388);
and U5951 (N_5951,N_2489,N_2510);
and U5952 (N_5952,N_2506,N_2786);
nor U5953 (N_5953,N_3955,N_2418);
and U5954 (N_5954,N_2626,N_2269);
or U5955 (N_5955,N_2619,N_2806);
xnor U5956 (N_5956,N_3749,N_2731);
xor U5957 (N_5957,N_2614,N_2344);
or U5958 (N_5958,N_3910,N_3874);
and U5959 (N_5959,N_2410,N_2040);
nand U5960 (N_5960,N_2492,N_2518);
xor U5961 (N_5961,N_2015,N_2835);
xor U5962 (N_5962,N_2585,N_2648);
nand U5963 (N_5963,N_2349,N_3740);
or U5964 (N_5964,N_3959,N_3184);
and U5965 (N_5965,N_2243,N_3665);
and U5966 (N_5966,N_2162,N_2627);
or U5967 (N_5967,N_2406,N_3616);
nor U5968 (N_5968,N_2426,N_2015);
xnor U5969 (N_5969,N_3873,N_2326);
and U5970 (N_5970,N_3825,N_3863);
nor U5971 (N_5971,N_3156,N_3716);
nor U5972 (N_5972,N_2279,N_3451);
or U5973 (N_5973,N_2414,N_2732);
nor U5974 (N_5974,N_3414,N_2677);
nand U5975 (N_5975,N_2982,N_2829);
xnor U5976 (N_5976,N_3817,N_2844);
nand U5977 (N_5977,N_3252,N_3388);
xnor U5978 (N_5978,N_3465,N_2093);
nand U5979 (N_5979,N_3584,N_3272);
and U5980 (N_5980,N_2118,N_3269);
nor U5981 (N_5981,N_3951,N_2282);
xnor U5982 (N_5982,N_3920,N_2054);
xnor U5983 (N_5983,N_2655,N_2319);
xnor U5984 (N_5984,N_3095,N_3759);
and U5985 (N_5985,N_2828,N_3879);
and U5986 (N_5986,N_3662,N_3174);
xor U5987 (N_5987,N_2472,N_2944);
nor U5988 (N_5988,N_3781,N_3684);
nor U5989 (N_5989,N_2373,N_2189);
nor U5990 (N_5990,N_2294,N_2997);
or U5991 (N_5991,N_2582,N_3350);
or U5992 (N_5992,N_3256,N_3766);
xnor U5993 (N_5993,N_3863,N_2374);
nand U5994 (N_5994,N_2895,N_2800);
or U5995 (N_5995,N_2308,N_3044);
nor U5996 (N_5996,N_2554,N_2340);
nand U5997 (N_5997,N_3192,N_3516);
xor U5998 (N_5998,N_2282,N_2908);
xor U5999 (N_5999,N_3824,N_2766);
nand U6000 (N_6000,N_4662,N_4634);
or U6001 (N_6001,N_4270,N_4961);
and U6002 (N_6002,N_4033,N_5497);
nand U6003 (N_6003,N_4404,N_5081);
nand U6004 (N_6004,N_5971,N_4975);
or U6005 (N_6005,N_4292,N_5920);
xor U6006 (N_6006,N_4916,N_5605);
nor U6007 (N_6007,N_4632,N_4527);
xnor U6008 (N_6008,N_4150,N_4598);
nor U6009 (N_6009,N_4650,N_5615);
xnor U6010 (N_6010,N_4848,N_5431);
nor U6011 (N_6011,N_4436,N_4992);
and U6012 (N_6012,N_5612,N_5536);
and U6013 (N_6013,N_4308,N_4883);
nor U6014 (N_6014,N_5298,N_5618);
nand U6015 (N_6015,N_4291,N_5991);
nand U6016 (N_6016,N_5566,N_5983);
and U6017 (N_6017,N_5011,N_5411);
and U6018 (N_6018,N_4329,N_4686);
and U6019 (N_6019,N_5044,N_4091);
xor U6020 (N_6020,N_4532,N_5811);
and U6021 (N_6021,N_4027,N_4197);
nor U6022 (N_6022,N_5316,N_4928);
xnor U6023 (N_6023,N_4281,N_4149);
nand U6024 (N_6024,N_4242,N_5053);
or U6025 (N_6025,N_4415,N_4639);
and U6026 (N_6026,N_5821,N_5279);
nor U6027 (N_6027,N_4118,N_5548);
nand U6028 (N_6028,N_5870,N_5491);
or U6029 (N_6029,N_4919,N_5947);
nand U6030 (N_6030,N_5052,N_5659);
and U6031 (N_6031,N_5132,N_4352);
or U6032 (N_6032,N_4971,N_4227);
xnor U6033 (N_6033,N_4955,N_5614);
and U6034 (N_6034,N_4534,N_5623);
and U6035 (N_6035,N_4178,N_5399);
and U6036 (N_6036,N_5265,N_5394);
xor U6037 (N_6037,N_4438,N_4705);
or U6038 (N_6038,N_4768,N_4183);
and U6039 (N_6039,N_5606,N_4185);
or U6040 (N_6040,N_4714,N_4805);
xor U6041 (N_6041,N_5848,N_5508);
xnor U6042 (N_6042,N_5185,N_5350);
and U6043 (N_6043,N_4278,N_5672);
nand U6044 (N_6044,N_5123,N_5900);
xnor U6045 (N_6045,N_5713,N_4342);
nand U6046 (N_6046,N_4029,N_4924);
and U6047 (N_6047,N_5752,N_5965);
nand U6048 (N_6048,N_4968,N_4383);
xnor U6049 (N_6049,N_4010,N_5238);
xnor U6050 (N_6050,N_5217,N_4229);
and U6051 (N_6051,N_4012,N_4897);
and U6052 (N_6052,N_4794,N_4796);
and U6053 (N_6053,N_4721,N_5529);
nor U6054 (N_6054,N_5578,N_4170);
nand U6055 (N_6055,N_5302,N_5162);
xor U6056 (N_6056,N_4320,N_4996);
xor U6057 (N_6057,N_4943,N_5251);
xnor U6058 (N_6058,N_4604,N_4315);
xnor U6059 (N_6059,N_5173,N_5013);
or U6060 (N_6060,N_5658,N_4513);
or U6061 (N_6061,N_4195,N_5640);
and U6062 (N_6062,N_4437,N_5914);
nor U6063 (N_6063,N_5239,N_4387);
or U6064 (N_6064,N_4323,N_4059);
or U6065 (N_6065,N_4665,N_4833);
nor U6066 (N_6066,N_4316,N_5791);
or U6067 (N_6067,N_5740,N_5595);
or U6068 (N_6068,N_5480,N_4479);
nor U6069 (N_6069,N_4396,N_5747);
nor U6070 (N_6070,N_4093,N_4138);
and U6071 (N_6071,N_4300,N_4073);
or U6072 (N_6072,N_5264,N_4452);
nand U6073 (N_6073,N_5363,N_4930);
nand U6074 (N_6074,N_4487,N_5976);
and U6075 (N_6075,N_4976,N_5987);
xnor U6076 (N_6076,N_5113,N_5768);
nor U6077 (N_6077,N_4477,N_5581);
or U6078 (N_6078,N_4755,N_5027);
or U6079 (N_6079,N_5864,N_4542);
nor U6080 (N_6080,N_5634,N_5693);
and U6081 (N_6081,N_5242,N_4793);
nor U6082 (N_6082,N_5125,N_4243);
or U6083 (N_6083,N_4496,N_5170);
and U6084 (N_6084,N_5405,N_4787);
xor U6085 (N_6085,N_5921,N_5200);
nand U6086 (N_6086,N_5923,N_4162);
and U6087 (N_6087,N_4753,N_5649);
xnor U6088 (N_6088,N_4819,N_4483);
xor U6089 (N_6089,N_5136,N_5002);
and U6090 (N_6090,N_4004,N_5168);
nor U6091 (N_6091,N_4917,N_4552);
or U6092 (N_6092,N_5797,N_5447);
or U6093 (N_6093,N_4600,N_4792);
xor U6094 (N_6094,N_4578,N_5674);
and U6095 (N_6095,N_4458,N_4279);
nor U6096 (N_6096,N_5771,N_5131);
xnor U6097 (N_6097,N_5365,N_4869);
nand U6098 (N_6098,N_4934,N_5155);
nand U6099 (N_6099,N_4133,N_5677);
nor U6100 (N_6100,N_4922,N_4077);
and U6101 (N_6101,N_5189,N_5515);
and U6102 (N_6102,N_4453,N_5819);
nand U6103 (N_6103,N_5330,N_4645);
nor U6104 (N_6104,N_4669,N_4354);
and U6105 (N_6105,N_5435,N_5580);
or U6106 (N_6106,N_5641,N_4122);
nand U6107 (N_6107,N_5776,N_4704);
nor U6108 (N_6108,N_4121,N_4672);
nor U6109 (N_6109,N_5942,N_4759);
nor U6110 (N_6110,N_4506,N_5390);
xor U6111 (N_6111,N_4574,N_5021);
xnor U6112 (N_6112,N_5552,N_5868);
or U6113 (N_6113,N_4584,N_4555);
nand U6114 (N_6114,N_4030,N_4865);
and U6115 (N_6115,N_5831,N_4245);
nor U6116 (N_6116,N_4336,N_5652);
or U6117 (N_6117,N_4023,N_4790);
xor U6118 (N_6118,N_4457,N_5761);
or U6119 (N_6119,N_5010,N_4969);
nor U6120 (N_6120,N_4215,N_4096);
or U6121 (N_6121,N_5250,N_4006);
or U6122 (N_6122,N_5312,N_4493);
or U6123 (N_6123,N_4207,N_5470);
nand U6124 (N_6124,N_4439,N_4823);
or U6125 (N_6125,N_4680,N_4046);
nor U6126 (N_6126,N_5826,N_5386);
or U6127 (N_6127,N_5009,N_5025);
nor U6128 (N_6128,N_4657,N_4938);
and U6129 (N_6129,N_5725,N_4827);
nand U6130 (N_6130,N_4560,N_4406);
and U6131 (N_6131,N_4289,N_4852);
or U6132 (N_6132,N_4663,N_5378);
xor U6133 (N_6133,N_5423,N_4495);
nor U6134 (N_6134,N_4689,N_4511);
nand U6135 (N_6135,N_4967,N_4053);
xor U6136 (N_6136,N_4719,N_4576);
and U6137 (N_6137,N_4143,N_5486);
or U6138 (N_6138,N_5099,N_5899);
xnor U6139 (N_6139,N_4656,N_5089);
nor U6140 (N_6140,N_5161,N_5715);
or U6141 (N_6141,N_4379,N_5562);
nand U6142 (N_6142,N_5880,N_4690);
and U6143 (N_6143,N_4168,N_5610);
nor U6144 (N_6144,N_4959,N_5318);
nor U6145 (N_6145,N_5661,N_4522);
nand U6146 (N_6146,N_5818,N_4175);
xor U6147 (N_6147,N_4814,N_5893);
nand U6148 (N_6148,N_5925,N_5400);
xnor U6149 (N_6149,N_5982,N_4764);
or U6150 (N_6150,N_5753,N_5549);
or U6151 (N_6151,N_5072,N_5257);
xor U6152 (N_6152,N_5256,N_4572);
xnor U6153 (N_6153,N_4824,N_4675);
and U6154 (N_6154,N_5457,N_4985);
nand U6155 (N_6155,N_5222,N_5449);
and U6156 (N_6156,N_4622,N_4365);
nor U6157 (N_6157,N_4879,N_4200);
nor U6158 (N_6158,N_4582,N_4945);
or U6159 (N_6159,N_5700,N_5563);
and U6160 (N_6160,N_5575,N_4082);
or U6161 (N_6161,N_4203,N_4119);
nor U6162 (N_6162,N_4911,N_4025);
nor U6163 (N_6163,N_4523,N_4981);
xnor U6164 (N_6164,N_5703,N_5973);
and U6165 (N_6165,N_4909,N_5273);
nand U6166 (N_6166,N_5858,N_5387);
and U6167 (N_6167,N_5499,N_4345);
and U6168 (N_6168,N_5970,N_4948);
xor U6169 (N_6169,N_4616,N_5084);
nor U6170 (N_6170,N_5984,N_4593);
xor U6171 (N_6171,N_4462,N_5056);
and U6172 (N_6172,N_5346,N_5382);
and U6173 (N_6173,N_5739,N_4654);
or U6174 (N_6174,N_5936,N_4927);
nor U6175 (N_6175,N_5259,N_4258);
xnor U6176 (N_6176,N_4842,N_4234);
xnor U6177 (N_6177,N_5816,N_4051);
and U6178 (N_6178,N_4060,N_5897);
nor U6179 (N_6179,N_5024,N_5154);
or U6180 (N_6180,N_4519,N_4867);
nand U6181 (N_6181,N_4209,N_5721);
nor U6182 (N_6182,N_5019,N_5175);
xor U6183 (N_6183,N_4633,N_5326);
nor U6184 (N_6184,N_5050,N_4433);
nor U6185 (N_6185,N_4647,N_5832);
nand U6186 (N_6186,N_4319,N_4710);
xnor U6187 (N_6187,N_5957,N_5074);
or U6188 (N_6188,N_5188,N_4001);
or U6189 (N_6189,N_5780,N_5590);
xnor U6190 (N_6190,N_4125,N_5028);
xor U6191 (N_6191,N_4249,N_4525);
nand U6192 (N_6192,N_4065,N_4039);
nand U6193 (N_6193,N_5235,N_5774);
xnor U6194 (N_6194,N_4233,N_4649);
xor U6195 (N_6195,N_4638,N_4161);
and U6196 (N_6196,N_4546,N_4817);
and U6197 (N_6197,N_4703,N_4765);
or U6198 (N_6198,N_4044,N_4318);
nor U6199 (N_6199,N_4864,N_4957);
xor U6200 (N_6200,N_5967,N_5037);
and U6201 (N_6201,N_4346,N_4761);
or U6202 (N_6202,N_5637,N_4936);
nand U6203 (N_6203,N_4488,N_5938);
nand U6204 (N_6204,N_4344,N_4129);
or U6205 (N_6205,N_5202,N_5960);
or U6206 (N_6206,N_5146,N_4235);
xor U6207 (N_6207,N_5334,N_5626);
and U6208 (N_6208,N_4196,N_4490);
and U6209 (N_6209,N_4984,N_4664);
or U6210 (N_6210,N_4325,N_5018);
xnor U6211 (N_6211,N_4543,N_5432);
nor U6212 (N_6212,N_4414,N_5461);
nand U6213 (N_6213,N_5783,N_4536);
and U6214 (N_6214,N_4956,N_5696);
nand U6215 (N_6215,N_5230,N_5600);
nor U6216 (N_6216,N_5246,N_5471);
or U6217 (N_6217,N_5134,N_4559);
and U6218 (N_6218,N_5793,N_5398);
nor U6219 (N_6219,N_5803,N_4421);
nand U6220 (N_6220,N_4013,N_4641);
nor U6221 (N_6221,N_4268,N_5221);
nand U6222 (N_6222,N_4244,N_5116);
nor U6223 (N_6223,N_4591,N_4731);
nand U6224 (N_6224,N_5359,N_4226);
xnor U6225 (N_6225,N_5118,N_4861);
nor U6226 (N_6226,N_5453,N_4217);
xor U6227 (N_6227,N_4707,N_4095);
nor U6228 (N_6228,N_5687,N_5100);
or U6229 (N_6229,N_5697,N_5139);
or U6230 (N_6230,N_5214,N_5758);
nand U6231 (N_6231,N_5607,N_4213);
xor U6232 (N_6232,N_5502,N_5931);
nor U6233 (N_6233,N_4169,N_4070);
nand U6234 (N_6234,N_5723,N_4424);
nor U6235 (N_6235,N_5477,N_4020);
xnor U6236 (N_6236,N_4628,N_4862);
or U6237 (N_6237,N_4331,N_5441);
and U6238 (N_6238,N_5518,N_5244);
nor U6239 (N_6239,N_4114,N_4771);
xnor U6240 (N_6240,N_5822,N_5717);
or U6241 (N_6241,N_4391,N_4940);
and U6242 (N_6242,N_5726,N_5974);
xor U6243 (N_6243,N_4442,N_4154);
nand U6244 (N_6244,N_5682,N_4274);
nor U6245 (N_6245,N_4648,N_5665);
nor U6246 (N_6246,N_4614,N_5488);
nor U6247 (N_6247,N_5422,N_4964);
nand U6248 (N_6248,N_4000,N_4470);
or U6249 (N_6249,N_4850,N_5571);
or U6250 (N_6250,N_5408,N_4124);
nor U6251 (N_6251,N_5532,N_4533);
nor U6252 (N_6252,N_4958,N_5836);
xnor U6253 (N_6253,N_4729,N_5380);
and U6254 (N_6254,N_5340,N_5760);
nor U6255 (N_6255,N_5732,N_5085);
and U6256 (N_6256,N_4577,N_4142);
xnor U6257 (N_6257,N_4742,N_4653);
nand U6258 (N_6258,N_4158,N_5782);
nor U6259 (N_6259,N_4811,N_4290);
and U6260 (N_6260,N_4637,N_5775);
and U6261 (N_6261,N_4579,N_4722);
nand U6262 (N_6262,N_4518,N_5097);
nand U6263 (N_6263,N_5598,N_5333);
and U6264 (N_6264,N_5918,N_4531);
nor U6265 (N_6265,N_5218,N_5465);
or U6266 (N_6266,N_4825,N_4165);
nand U6267 (N_6267,N_4809,N_4120);
and U6268 (N_6268,N_4199,N_4427);
or U6269 (N_6269,N_5859,N_4899);
xnor U6270 (N_6270,N_4715,N_5625);
nor U6271 (N_6271,N_5962,N_5287);
and U6272 (N_6272,N_5809,N_4224);
and U6273 (N_6273,N_5337,N_5988);
or U6274 (N_6274,N_4454,N_4803);
and U6275 (N_6275,N_4146,N_4997);
and U6276 (N_6276,N_4949,N_4720);
or U6277 (N_6277,N_5820,N_5841);
or U6278 (N_6278,N_4284,N_5927);
xnor U6279 (N_6279,N_5736,N_5035);
nor U6280 (N_6280,N_4569,N_4031);
nand U6281 (N_6281,N_4418,N_5345);
nand U6282 (N_6282,N_4747,N_5787);
or U6283 (N_6283,N_4241,N_4965);
nor U6284 (N_6284,N_5255,N_4152);
nor U6285 (N_6285,N_5487,N_4484);
nand U6286 (N_6286,N_4630,N_4448);
and U6287 (N_6287,N_4791,N_4882);
nand U6288 (N_6288,N_5286,N_5303);
nor U6289 (N_6289,N_4918,N_4566);
or U6290 (N_6290,N_4334,N_5850);
and U6291 (N_6291,N_5180,N_5468);
and U6292 (N_6292,N_4401,N_4181);
and U6293 (N_6293,N_5907,N_5424);
or U6294 (N_6294,N_4907,N_4423);
xnor U6295 (N_6295,N_4520,N_5117);
nand U6296 (N_6296,N_5898,N_5299);
and U6297 (N_6297,N_5702,N_4371);
or U6298 (N_6298,N_4335,N_4507);
xnor U6299 (N_6299,N_4079,N_5000);
nor U6300 (N_6300,N_5915,N_4563);
and U6301 (N_6301,N_5057,N_5140);
nand U6302 (N_6302,N_4605,N_5065);
or U6303 (N_6303,N_5639,N_5585);
xor U6304 (N_6304,N_5628,N_5838);
nand U6305 (N_6305,N_5356,N_5428);
or U6306 (N_6306,N_4854,N_4540);
and U6307 (N_6307,N_5216,N_4109);
nand U6308 (N_6308,N_4989,N_4789);
nor U6309 (N_6309,N_5828,N_4966);
or U6310 (N_6310,N_4545,N_5190);
or U6311 (N_6311,N_5855,N_5643);
or U6312 (N_6312,N_4257,N_4333);
or U6313 (N_6313,N_4986,N_5601);
nand U6314 (N_6314,N_4581,N_5521);
xor U6315 (N_6315,N_5716,N_5889);
nor U6316 (N_6316,N_5023,N_4795);
and U6317 (N_6317,N_4878,N_5924);
nand U6318 (N_6318,N_5778,N_5773);
nor U6319 (N_6319,N_5544,N_4313);
and U6320 (N_6320,N_4309,N_4906);
nor U6321 (N_6321,N_5410,N_4667);
xnor U6322 (N_6322,N_4627,N_5135);
or U6323 (N_6323,N_4845,N_4238);
or U6324 (N_6324,N_4028,N_5501);
and U6325 (N_6325,N_4009,N_4855);
or U6326 (N_6326,N_5274,N_5223);
and U6327 (N_6327,N_5569,N_4763);
and U6328 (N_6328,N_4330,N_4987);
and U6329 (N_6329,N_4974,N_5762);
or U6330 (N_6330,N_5622,N_5485);
and U6331 (N_6331,N_5698,N_5062);
and U6332 (N_6332,N_4367,N_5254);
and U6333 (N_6333,N_5517,N_4944);
xnor U6334 (N_6334,N_5041,N_5944);
nor U6335 (N_6335,N_5434,N_5121);
or U6336 (N_6336,N_5750,N_4314);
and U6337 (N_6337,N_5737,N_4145);
nand U6338 (N_6338,N_4735,N_5751);
or U6339 (N_6339,N_4888,N_4980);
or U6340 (N_6340,N_5300,N_4038);
nor U6341 (N_6341,N_5808,N_5690);
nor U6342 (N_6342,N_5695,N_4252);
nand U6343 (N_6343,N_5741,N_4456);
xor U6344 (N_6344,N_5888,N_5051);
or U6345 (N_6345,N_5391,N_5955);
or U6346 (N_6346,N_4822,N_4561);
and U6347 (N_6347,N_4048,N_5533);
nor U6348 (N_6348,N_4251,N_4127);
and U6349 (N_6349,N_5219,N_5781);
xor U6350 (N_6350,N_5474,N_5416);
xnor U6351 (N_6351,N_4429,N_4230);
or U6352 (N_6352,N_4692,N_5141);
and U6353 (N_6353,N_4126,N_4036);
nand U6354 (N_6354,N_5296,N_5080);
nor U6355 (N_6355,N_5063,N_5712);
or U6356 (N_6356,N_5379,N_5842);
or U6357 (N_6357,N_5020,N_4613);
or U6358 (N_6358,N_5413,N_4491);
nand U6359 (N_6359,N_4434,N_5472);
and U6360 (N_6360,N_4360,N_4405);
or U6361 (N_6361,N_5964,N_4256);
nor U6362 (N_6362,N_4500,N_4410);
nor U6363 (N_6363,N_5669,N_5489);
nor U6364 (N_6364,N_4564,N_4166);
nand U6365 (N_6365,N_5156,N_4392);
or U6366 (N_6366,N_4858,N_5397);
or U6367 (N_6367,N_4709,N_4570);
and U6368 (N_6368,N_5556,N_5396);
and U6369 (N_6369,N_5655,N_5182);
and U6370 (N_6370,N_4688,N_5290);
xor U6371 (N_6371,N_4592,N_4187);
or U6372 (N_6372,N_4282,N_5660);
nand U6373 (N_6373,N_5930,N_4332);
and U6374 (N_6374,N_4035,N_4248);
xnor U6375 (N_6375,N_4698,N_5232);
xor U6376 (N_6376,N_4537,N_4380);
and U6377 (N_6377,N_5371,N_4762);
xnor U6378 (N_6378,N_5040,N_5194);
and U6379 (N_6379,N_4697,N_5986);
xor U6380 (N_6380,N_4273,N_4349);
or U6381 (N_6381,N_4337,N_5070);
nand U6382 (N_6382,N_4902,N_5483);
nor U6383 (N_6383,N_5817,N_4901);
or U6384 (N_6384,N_5181,N_5565);
or U6385 (N_6385,N_5090,N_4440);
nand U6386 (N_6386,N_4485,N_5956);
and U6387 (N_6387,N_5127,N_4461);
nor U6388 (N_6388,N_4615,N_4358);
or U6389 (N_6389,N_4781,N_4123);
nand U6390 (N_6390,N_4419,N_5343);
or U6391 (N_6391,N_4014,N_5314);
nand U6392 (N_6392,N_4877,N_5573);
nand U6393 (N_6393,N_4366,N_4375);
and U6394 (N_6394,N_5513,N_5381);
and U6395 (N_6395,N_5805,N_4113);
or U6396 (N_6396,N_5507,N_4341);
and U6397 (N_6397,N_5912,N_5861);
or U6398 (N_6398,N_5177,N_5228);
xor U6399 (N_6399,N_5935,N_5852);
and U6400 (N_6400,N_5635,N_4857);
xnor U6401 (N_6401,N_5479,N_4111);
and U6402 (N_6402,N_5790,N_5550);
xor U6403 (N_6403,N_4348,N_4198);
xor U6404 (N_6404,N_4478,N_5594);
xor U6405 (N_6405,N_5476,N_5484);
nand U6406 (N_6406,N_4946,N_4602);
xor U6407 (N_6407,N_4651,N_4843);
nand U6408 (N_6408,N_4002,N_4844);
nand U6409 (N_6409,N_5149,N_4914);
xnor U6410 (N_6410,N_4164,N_5886);
nand U6411 (N_6411,N_4887,N_4212);
xnor U6412 (N_6412,N_5420,N_4317);
xnor U6413 (N_6413,N_5017,N_5577);
xnor U6414 (N_6414,N_4034,N_5464);
nand U6415 (N_6415,N_4388,N_4473);
and U6416 (N_6416,N_5005,N_4110);
nor U6417 (N_6417,N_4767,N_4874);
and U6418 (N_6418,N_5516,N_4502);
and U6419 (N_6419,N_5240,N_5361);
nor U6420 (N_6420,N_5106,N_4047);
nand U6421 (N_6421,N_5767,N_5749);
nor U6422 (N_6422,N_4192,N_4116);
xor U6423 (N_6423,N_4254,N_5153);
nand U6424 (N_6424,N_5327,N_5895);
nor U6425 (N_6425,N_4135,N_5685);
xnor U6426 (N_6426,N_5032,N_5977);
xnor U6427 (N_6427,N_4469,N_4193);
xnor U6428 (N_6428,N_5348,N_5830);
or U6429 (N_6429,N_4713,N_4237);
or U6430 (N_6430,N_5404,N_5347);
nand U6431 (N_6431,N_5328,N_5367);
or U6432 (N_6432,N_5187,N_5266);
nand U6433 (N_6433,N_4117,N_5949);
and U6434 (N_6434,N_5042,N_4580);
nor U6435 (N_6435,N_4952,N_4625);
or U6436 (N_6436,N_4770,N_4571);
nand U6437 (N_6437,N_4104,N_4216);
and U6438 (N_6438,N_5718,N_5812);
nor U6439 (N_6439,N_4214,N_5212);
xnor U6440 (N_6440,N_4210,N_5588);
or U6441 (N_6441,N_4050,N_4061);
or U6442 (N_6442,N_4272,N_4400);
xor U6443 (N_6443,N_5112,N_5530);
nand U6444 (N_6444,N_5657,N_5102);
nand U6445 (N_6445,N_4003,N_5126);
or U6446 (N_6446,N_5527,N_4514);
nand U6447 (N_6447,N_5492,N_4652);
nor U6448 (N_6448,N_5285,N_4859);
xor U6449 (N_6449,N_5883,N_5746);
or U6450 (N_6450,N_5849,N_5710);
nand U6451 (N_6451,N_4139,N_4100);
and U6452 (N_6452,N_4293,N_5128);
or U6453 (N_6453,N_5528,N_5520);
nand U6454 (N_6454,N_4750,N_5352);
or U6455 (N_6455,N_4838,N_4026);
or U6456 (N_6456,N_5183,N_5210);
nand U6457 (N_6457,N_4994,N_5060);
or U6458 (N_6458,N_4695,N_4626);
nor U6459 (N_6459,N_5884,N_4459);
nand U6460 (N_6460,N_4884,N_5777);
nand U6461 (N_6461,N_4903,N_5846);
and U6462 (N_6462,N_4766,N_5932);
xor U6463 (N_6463,N_4983,N_5389);
nand U6464 (N_6464,N_4264,N_4058);
xor U6465 (N_6465,N_5872,N_5107);
and U6466 (N_6466,N_5211,N_5731);
xor U6467 (N_6467,N_4737,N_4206);
and U6468 (N_6468,N_5624,N_5950);
nand U6469 (N_6469,N_4913,N_4057);
or U6470 (N_6470,N_4147,N_4933);
nor U6471 (N_6471,N_4191,N_5373);
or U6472 (N_6472,N_4711,N_5509);
or U6473 (N_6473,N_5727,N_5460);
nor U6474 (N_6474,N_5459,N_5798);
nand U6475 (N_6475,N_4476,N_4910);
xnor U6476 (N_6476,N_5415,N_5851);
nand U6477 (N_6477,N_5757,N_5887);
nor U6478 (N_6478,N_4299,N_5262);
and U6479 (N_6479,N_5892,N_4225);
and U6480 (N_6480,N_5061,N_5744);
nor U6481 (N_6481,N_4587,N_4505);
and U6482 (N_6482,N_5443,N_4081);
and U6483 (N_6483,N_4807,N_5277);
and U6484 (N_6484,N_5814,N_4468);
and U6485 (N_6485,N_5946,N_4995);
nor U6486 (N_6486,N_4420,N_4373);
or U6487 (N_6487,N_4190,N_4895);
or U6488 (N_6488,N_4849,N_5675);
nor U6489 (N_6489,N_5586,N_4723);
and U6490 (N_6490,N_5445,N_5806);
or U6491 (N_6491,N_4370,N_5505);
and U6492 (N_6492,N_4835,N_4159);
or U6493 (N_6493,N_4055,N_4236);
nand U6494 (N_6494,N_4670,N_4881);
and U6495 (N_6495,N_5874,N_5802);
or U6496 (N_6496,N_5272,N_4512);
and U6497 (N_6497,N_4797,N_5978);
and U6498 (N_6498,N_5092,N_4603);
and U6499 (N_6499,N_4089,N_5455);
nor U6500 (N_6500,N_4947,N_5030);
and U6501 (N_6501,N_5364,N_4482);
nand U6502 (N_6502,N_4094,N_4451);
and U6503 (N_6503,N_5705,N_4084);
or U6504 (N_6504,N_4595,N_5336);
and U6505 (N_6505,N_4880,N_5231);
xnor U6506 (N_6506,N_5093,N_5825);
and U6507 (N_6507,N_5335,N_4635);
or U6508 (N_6508,N_5007,N_5226);
nand U6509 (N_6509,N_5357,N_4778);
nand U6510 (N_6510,N_5463,N_4810);
nand U6511 (N_6511,N_4751,N_5593);
and U6512 (N_6512,N_4860,N_4799);
xnor U6513 (N_6513,N_4492,N_4338);
and U6514 (N_6514,N_5358,N_5281);
nor U6515 (N_6515,N_5096,N_5064);
xnor U6516 (N_6516,N_5688,N_5342);
and U6517 (N_6517,N_5192,N_4384);
xor U6518 (N_6518,N_5524,N_4005);
and U6519 (N_6519,N_4450,N_4042);
nor U6520 (N_6520,N_5512,N_5111);
nand U6521 (N_6521,N_5759,N_5704);
and U6522 (N_6522,N_5220,N_5807);
and U6523 (N_6523,N_4385,N_4745);
or U6524 (N_6524,N_5213,N_4350);
nor U6525 (N_6525,N_5894,N_5616);
or U6526 (N_6526,N_5179,N_5253);
nand U6527 (N_6527,N_4585,N_4586);
xnor U6528 (N_6528,N_4472,N_5109);
nand U6529 (N_6529,N_5772,N_4151);
or U6530 (N_6530,N_5903,N_4460);
and U6531 (N_6531,N_4374,N_5143);
nand U6532 (N_6532,N_4951,N_5878);
xnor U6533 (N_6533,N_4549,N_5144);
xnor U6534 (N_6534,N_4941,N_5539);
and U6535 (N_6535,N_4774,N_5174);
and U6536 (N_6536,N_5503,N_4678);
nand U6537 (N_6537,N_5278,N_4873);
and U6538 (N_6538,N_5869,N_5191);
nand U6539 (N_6539,N_5769,N_4757);
nor U6540 (N_6540,N_5667,N_4661);
nand U6541 (N_6541,N_5701,N_5055);
and U6542 (N_6542,N_5436,N_4301);
xnor U6543 (N_6543,N_5523,N_4993);
and U6544 (N_6544,N_4724,N_4693);
or U6545 (N_6545,N_4021,N_4890);
xnor U6546 (N_6546,N_5966,N_5227);
nor U6547 (N_6547,N_5733,N_5788);
xnor U6548 (N_6548,N_4538,N_4306);
xnor U6549 (N_6549,N_5766,N_4428);
nor U6550 (N_6550,N_4136,N_4445);
or U6551 (N_6551,N_5748,N_4802);
and U6552 (N_6552,N_4772,N_4263);
nand U6553 (N_6553,N_4754,N_5843);
and U6554 (N_6554,N_4359,N_5969);
xor U6555 (N_6555,N_4736,N_4925);
or U6556 (N_6556,N_5172,N_4395);
and U6557 (N_6557,N_5165,N_5860);
or U6558 (N_6558,N_4606,N_4889);
xor U6559 (N_6559,N_5321,N_5167);
or U6560 (N_6560,N_4979,N_5066);
nor U6561 (N_6561,N_5708,N_5215);
nor U6562 (N_6562,N_5075,N_5467);
nand U6563 (N_6563,N_5995,N_5647);
nor U6564 (N_6564,N_5103,N_4818);
or U6565 (N_6565,N_5115,N_5114);
or U6566 (N_6566,N_4265,N_5305);
or U6567 (N_6567,N_4872,N_4155);
and U6568 (N_6568,N_5147,N_5724);
or U6569 (N_6569,N_5638,N_5570);
and U6570 (N_6570,N_4471,N_5130);
and U6571 (N_6571,N_5673,N_5994);
xor U6572 (N_6572,N_5917,N_5840);
nor U6573 (N_6573,N_4101,N_5417);
xor U6574 (N_6574,N_4307,N_5260);
and U6575 (N_6575,N_5928,N_5730);
nor U6576 (N_6576,N_4846,N_4937);
xor U6577 (N_6577,N_4748,N_5271);
or U6578 (N_6578,N_4172,N_4624);
and U6579 (N_6579,N_4871,N_4153);
or U6580 (N_6580,N_4261,N_5785);
nand U6581 (N_6581,N_5046,N_5763);
and U6582 (N_6582,N_4340,N_5429);
or U6583 (N_6583,N_5105,N_4182);
nand U6584 (N_6584,N_4932,N_5008);
and U6585 (N_6585,N_4287,N_4892);
or U6586 (N_6586,N_5369,N_4728);
or U6587 (N_6587,N_5451,N_4904);
nor U6588 (N_6588,N_5514,N_5313);
xor U6589 (N_6589,N_5526,N_4556);
or U6590 (N_6590,N_5603,N_4298);
xor U6591 (N_6591,N_5953,N_4054);
and U6592 (N_6592,N_5591,N_5043);
and U6593 (N_6593,N_4551,N_4016);
or U6594 (N_6594,N_4435,N_5998);
or U6595 (N_6595,N_5067,N_4660);
nor U6596 (N_6596,N_5629,N_5686);
and U6597 (N_6597,N_5794,N_4176);
nand U6598 (N_6598,N_4510,N_4908);
nand U6599 (N_6599,N_5026,N_5707);
and U6600 (N_6600,N_5755,N_4390);
xor U6601 (N_6601,N_5684,N_4529);
xnor U6602 (N_6602,N_4277,N_5073);
and U6603 (N_6603,N_4607,N_5729);
nor U6604 (N_6604,N_5368,N_4726);
or U6605 (N_6605,N_4978,N_4779);
nand U6606 (N_6606,N_4621,N_4088);
nor U6607 (N_6607,N_4072,N_5972);
or U6608 (N_6608,N_4250,N_4950);
nand U6609 (N_6609,N_5482,N_4851);
or U6610 (N_6610,N_4022,N_4939);
xnor U6611 (N_6611,N_5679,N_5504);
nor U6612 (N_6612,N_4931,N_4891);
nand U6613 (N_6613,N_5004,N_4267);
xnor U6614 (N_6614,N_5442,N_5996);
nor U6615 (N_6615,N_4475,N_5554);
xor U6616 (N_6616,N_5203,N_4378);
or U6617 (N_6617,N_4610,N_4321);
nand U6618 (N_6618,N_5534,N_4481);
nand U6619 (N_6619,N_4411,N_4463);
xnor U6620 (N_6620,N_4826,N_4364);
or U6621 (N_6621,N_4524,N_5908);
nand U6622 (N_6622,N_5108,N_5885);
or U6623 (N_6623,N_4163,N_4960);
xor U6624 (N_6624,N_4239,N_5958);
and U6625 (N_6625,N_4548,N_5754);
xnor U6626 (N_6626,N_5940,N_4443);
and U6627 (N_6627,N_4064,N_5403);
xor U6628 (N_6628,N_5653,N_4550);
xnor U6629 (N_6629,N_5670,N_5939);
nand U6630 (N_6630,N_5295,N_4696);
or U6631 (N_6631,N_4631,N_4876);
or U6632 (N_6632,N_5280,N_4999);
xnor U6633 (N_6633,N_4056,N_4489);
nand U6634 (N_6634,N_4773,N_5481);
nand U6635 (N_6635,N_4963,N_5426);
or U6636 (N_6636,N_5662,N_5943);
nand U6637 (N_6637,N_4134,N_4156);
nand U6638 (N_6638,N_5650,N_5016);
nand U6639 (N_6639,N_5620,N_5234);
nor U6640 (N_6640,N_4885,N_4804);
nor U6641 (N_6641,N_5558,N_4106);
nor U6642 (N_6642,N_4174,N_5425);
or U6643 (N_6643,N_4953,N_4353);
or U6644 (N_6644,N_4798,N_4738);
and U6645 (N_6645,N_4032,N_4682);
or U6646 (N_6646,N_5195,N_5283);
nor U6647 (N_6647,N_5439,N_5245);
nand U6648 (N_6648,N_5913,N_5493);
nor U6649 (N_6649,N_5087,N_4386);
or U6650 (N_6650,N_5546,N_4866);
or U6651 (N_6651,N_4255,N_5289);
nor U6652 (N_6652,N_5385,N_4194);
or U6653 (N_6653,N_5613,N_5576);
or U6654 (N_6654,N_4467,N_5159);
and U6655 (N_6655,N_5275,N_4777);
nand U6656 (N_6656,N_4188,N_5633);
nor U6657 (N_6657,N_4184,N_4567);
or U6658 (N_6658,N_5496,N_5354);
and U6659 (N_6659,N_4393,N_4644);
xnor U6660 (N_6660,N_4868,N_4780);
nor U6661 (N_6661,N_4821,N_5490);
xnor U6662 (N_6662,N_5088,N_5466);
xor U6663 (N_6663,N_5596,N_5862);
or U6664 (N_6664,N_4744,N_5568);
nand U6665 (N_6665,N_4691,N_4497);
xor U6666 (N_6666,N_5383,N_5545);
nor U6667 (N_6667,N_5433,N_5664);
xnor U6668 (N_6668,N_5418,N_5876);
nor U6669 (N_6669,N_4205,N_4839);
nor U6670 (N_6670,N_5993,N_5877);
xnor U6671 (N_6671,N_4528,N_4102);
nor U6672 (N_6672,N_5572,N_5241);
or U6673 (N_6673,N_5511,N_4052);
xnor U6674 (N_6674,N_5979,N_5743);
nand U6675 (N_6675,N_5209,N_5975);
and U6676 (N_6676,N_4087,N_5666);
or U6677 (N_6677,N_4128,N_5564);
nor U6678 (N_6678,N_4935,N_5770);
xor U6679 (N_6679,N_5631,N_4565);
or U6680 (N_6680,N_5609,N_4220);
nor U6681 (N_6681,N_5048,N_5919);
xor U6682 (N_6682,N_5765,N_4407);
and U6683 (N_6683,N_5689,N_5452);
nand U6684 (N_6684,N_4743,N_5879);
or U6685 (N_6685,N_4363,N_5284);
nor U6686 (N_6686,N_4776,N_5039);
or U6687 (N_6687,N_5054,N_5229);
nor U6688 (N_6688,N_4403,N_4099);
or U6689 (N_6689,N_5325,N_4733);
xor U6690 (N_6690,N_4732,N_5098);
nand U6691 (N_6691,N_4008,N_5003);
nand U6692 (N_6692,N_4137,N_4526);
or U6693 (N_6693,N_5448,N_4700);
xnor U6694 (N_6694,N_5654,N_5082);
or U6695 (N_6695,N_4464,N_5437);
and U6696 (N_6696,N_5792,N_5407);
xor U6697 (N_6697,N_5269,N_4828);
and U6698 (N_6698,N_5095,N_5856);
nor U6699 (N_6699,N_4413,N_4179);
nor U6700 (N_6700,N_4756,N_4501);
nor U6701 (N_6701,N_5735,N_5789);
xor U6702 (N_6702,N_4727,N_5992);
or U6703 (N_6703,N_5344,N_4847);
nand U6704 (N_6704,N_5906,N_5169);
xor U6705 (N_6705,N_4486,N_4816);
or U6706 (N_6706,N_5555,N_5989);
and U6707 (N_6707,N_4590,N_4112);
xor U6708 (N_6708,N_4372,N_5863);
and U6709 (N_6709,N_4024,N_5362);
xnor U6710 (N_6710,N_5444,N_5207);
xor U6711 (N_6711,N_4801,N_5745);
and U6712 (N_6712,N_5071,N_4148);
nand U6713 (N_6713,N_5589,N_5500);
nand U6714 (N_6714,N_5525,N_4544);
xor U6715 (N_6715,N_5542,N_5308);
nand U6716 (N_6716,N_5261,N_5120);
or U6717 (N_6717,N_5671,N_4201);
and U6718 (N_6718,N_5276,N_4417);
or U6719 (N_6719,N_4831,N_5164);
or U6720 (N_6720,N_4741,N_5237);
xor U6721 (N_6721,N_4702,N_4718);
xnor U6722 (N_6722,N_4019,N_5980);
nor U6723 (N_6723,N_5377,N_4841);
nor U6724 (N_6724,N_5045,N_5249);
xnor U6725 (N_6725,N_4232,N_4076);
and U6726 (N_6726,N_4066,N_4712);
and U6727 (N_6727,N_5678,N_4222);
or U6728 (N_6728,N_4328,N_4962);
or U6729 (N_6729,N_4045,N_4666);
and U6730 (N_6730,N_5642,N_5122);
and U6731 (N_6731,N_5409,N_5929);
or U6732 (N_6732,N_5012,N_5845);
and U6733 (N_6733,N_5148,N_5178);
and U6734 (N_6734,N_4347,N_4998);
nand U6735 (N_6735,N_5881,N_4204);
nor U6736 (N_6736,N_5311,N_4562);
nor U6737 (N_6737,N_5355,N_4305);
nor U6738 (N_6738,N_5157,N_4708);
nand U6739 (N_6739,N_4398,N_4017);
nor U6740 (N_6740,N_5873,N_4361);
or U6741 (N_6741,N_4382,N_5796);
and U6742 (N_6742,N_5630,N_5225);
nand U6743 (N_6743,N_4588,N_4597);
or U6744 (N_6744,N_4357,N_4408);
nand U6745 (N_6745,N_4508,N_5049);
nand U6746 (N_6746,N_4080,N_4219);
nor U6747 (N_6747,N_4609,N_4749);
nor U6748 (N_6748,N_4785,N_4769);
nand U6749 (N_6749,N_5694,N_4706);
nor U6750 (N_6750,N_5719,N_4180);
and U6751 (N_6751,N_5388,N_4465);
or U6752 (N_6752,N_5427,N_5981);
xnor U6753 (N_6753,N_5632,N_4140);
or U6754 (N_6754,N_4642,N_4425);
and U6755 (N_6755,N_5651,N_5199);
or U6756 (N_6756,N_4800,N_5531);
xnor U6757 (N_6757,N_5854,N_5036);
xnor U6758 (N_6758,N_5810,N_5985);
nand U6759 (N_6759,N_5309,N_5857);
xor U6760 (N_6760,N_4870,N_4432);
nand U6761 (N_6761,N_4611,N_5412);
and U6762 (N_6762,N_4351,N_4262);
or U6763 (N_6763,N_4304,N_5933);
xnor U6764 (N_6764,N_5317,N_5583);
and U6765 (N_6765,N_5456,N_5668);
xnor U6766 (N_6766,N_5376,N_4679);
and U6767 (N_6767,N_5094,N_5421);
nor U6768 (N_6768,N_5068,N_5833);
or U6769 (N_6769,N_5091,N_4905);
or U6770 (N_6770,N_5401,N_5617);
nand U6771 (N_6771,N_5680,N_4815);
nor U6772 (N_6772,N_5475,N_5910);
nor U6773 (N_6773,N_5522,N_5291);
or U6774 (N_6774,N_4269,N_4573);
and U6775 (N_6775,N_4640,N_4658);
nand U6776 (N_6776,N_4362,N_4015);
nand U6777 (N_6777,N_5551,N_5997);
and U6778 (N_6778,N_5393,N_4808);
xnor U6779 (N_6779,N_5248,N_4832);
and U6780 (N_6780,N_4601,N_5233);
or U6781 (N_6781,N_5882,N_5469);
or U6782 (N_6782,N_5152,N_5948);
and U6783 (N_6783,N_5959,N_5478);
or U6784 (N_6784,N_4090,N_5208);
or U6785 (N_6785,N_5205,N_4494);
nand U6786 (N_6786,N_4422,N_4900);
xor U6787 (N_6787,N_5069,N_4310);
xor U6788 (N_6788,N_4097,N_4107);
and U6789 (N_6789,N_4977,N_5078);
xor U6790 (N_6790,N_5547,N_4541);
xnor U6791 (N_6791,N_4674,N_4671);
or U6792 (N_6792,N_5402,N_4617);
xnor U6793 (N_6793,N_4171,N_4498);
nor U6794 (N_6794,N_5331,N_5813);
or U6795 (N_6795,N_5137,N_5375);
or U6796 (N_6796,N_5599,N_4683);
nand U6797 (N_6797,N_5619,N_5395);
nor U6798 (N_6798,N_4141,N_4535);
and U6799 (N_6799,N_5204,N_5963);
or U6800 (N_6800,N_4397,N_4177);
or U6801 (N_6801,N_5406,N_4075);
nor U6802 (N_6802,N_4915,N_5077);
nand U6803 (N_6803,N_5734,N_5709);
xor U6804 (N_6804,N_4758,N_4247);
nand U6805 (N_6805,N_5867,N_5644);
nand U6806 (N_6806,N_4474,N_5663);
xor U6807 (N_6807,N_4740,N_4988);
nor U6808 (N_6808,N_4040,N_4894);
nand U6809 (N_6809,N_5292,N_4098);
and U6810 (N_6810,N_4211,N_5224);
nand U6811 (N_6811,N_4921,N_5133);
xor U6812 (N_6812,N_4253,N_4694);
and U6813 (N_6813,N_5926,N_5837);
or U6814 (N_6814,N_5866,N_5142);
xor U6815 (N_6815,N_4160,N_4295);
nand U6816 (N_6816,N_5597,N_4186);
xor U6817 (N_6817,N_4699,N_5645);
nor U6818 (N_6818,N_5014,N_4739);
xor U6819 (N_6819,N_5904,N_4018);
or U6820 (N_6820,N_4836,N_5158);
xor U6821 (N_6821,N_4929,N_4455);
or U6822 (N_6822,N_4416,N_4240);
nor U6823 (N_6823,N_5151,N_4381);
or U6824 (N_6824,N_5374,N_4912);
nand U6825 (N_6825,N_4982,N_5288);
nand U6826 (N_6826,N_5890,N_4589);
nor U6827 (N_6827,N_5372,N_5891);
nand U6828 (N_6828,N_5186,N_4409);
nor U6829 (N_6829,N_5922,N_4530);
nor U6830 (N_6830,N_4837,N_4283);
or U6831 (N_6831,N_5150,N_4517);
xor U6832 (N_6832,N_5961,N_5648);
nor U6833 (N_6833,N_5519,N_5258);
nand U6834 (N_6834,N_4266,N_4132);
or U6835 (N_6835,N_4246,N_5446);
nor U6836 (N_6836,N_4619,N_4568);
nand U6837 (N_6837,N_4942,N_5310);
or U6838 (N_6838,N_4775,N_5553);
or U6839 (N_6839,N_5243,N_5307);
or U6840 (N_6840,N_5901,N_4355);
or U6841 (N_6841,N_5627,N_4260);
nand U6842 (N_6842,N_5083,N_4734);
xnor U6843 (N_6843,N_5823,N_5329);
xnor U6844 (N_6844,N_5252,N_5498);
nand U6845 (N_6845,N_4539,N_4806);
nand U6846 (N_6846,N_4063,N_5304);
xnor U6847 (N_6847,N_4840,N_5268);
nand U6848 (N_6848,N_5535,N_4157);
xnor U6849 (N_6849,N_4643,N_4043);
xor U6850 (N_6850,N_5332,N_5270);
xnor U6851 (N_6851,N_4228,N_4599);
or U6852 (N_6852,N_5579,N_5557);
and U6853 (N_6853,N_4218,N_5902);
or U6854 (N_6854,N_5495,N_4288);
and U6855 (N_6855,N_4829,N_5592);
or U6856 (N_6856,N_4259,N_4973);
nor U6857 (N_6857,N_4368,N_5764);
or U6858 (N_6858,N_4322,N_5543);
and U6859 (N_6859,N_5015,N_5323);
or U6860 (N_6860,N_5267,N_4612);
or U6861 (N_6861,N_5263,N_5059);
xnor U6862 (N_6862,N_4521,N_4115);
nand U6863 (N_6863,N_4923,N_4746);
nor U6864 (N_6864,N_5184,N_4886);
or U6865 (N_6865,N_5033,N_5315);
and U6866 (N_6866,N_5720,N_4813);
and U6867 (N_6867,N_4596,N_5206);
and U6868 (N_6868,N_5297,N_5795);
or U6869 (N_6869,N_5722,N_5699);
or U6870 (N_6870,N_5951,N_5440);
nor U6871 (N_6871,N_5353,N_4725);
and U6872 (N_6872,N_5079,N_5236);
and U6873 (N_6873,N_5201,N_5800);
and U6874 (N_6874,N_4717,N_4788);
nor U6875 (N_6875,N_5756,N_5909);
and U6876 (N_6876,N_4853,N_5414);
or U6877 (N_6877,N_4701,N_4685);
nand U6878 (N_6878,N_4594,N_4990);
nor U6879 (N_6879,N_4954,N_5990);
nand U6880 (N_6880,N_4499,N_5324);
xor U6881 (N_6881,N_5871,N_4583);
nor U6882 (N_6882,N_4515,N_5506);
xor U6883 (N_6883,N_4629,N_4067);
nand U6884 (N_6884,N_4830,N_5022);
nand U6885 (N_6885,N_5738,N_4668);
nand U6886 (N_6886,N_4898,N_5166);
nand U6887 (N_6887,N_4553,N_5784);
and U6888 (N_6888,N_5865,N_4007);
or U6889 (N_6889,N_4311,N_5104);
xor U6890 (N_6890,N_5034,N_5282);
nand U6891 (N_6891,N_5567,N_5322);
nand U6892 (N_6892,N_5611,N_4896);
nand U6893 (N_6893,N_4503,N_5293);
nand U6894 (N_6894,N_4516,N_5129);
or U6895 (N_6895,N_4730,N_5124);
xnor U6896 (N_6896,N_4608,N_4108);
xnor U6897 (N_6897,N_4326,N_4389);
nor U6898 (N_6898,N_4271,N_4302);
xnor U6899 (N_6899,N_5338,N_4131);
nand U6900 (N_6900,N_5031,N_5621);
nand U6901 (N_6901,N_4716,N_5656);
nand U6902 (N_6902,N_4285,N_4575);
or U6903 (N_6903,N_4441,N_5538);
xnor U6904 (N_6904,N_4426,N_5916);
nand U6905 (N_6905,N_4920,N_4677);
nor U6906 (N_6906,N_4655,N_4376);
or U6907 (N_6907,N_4074,N_5834);
or U6908 (N_6908,N_5839,N_4303);
and U6909 (N_6909,N_5001,N_5646);
nand U6910 (N_6910,N_4444,N_5676);
nand U6911 (N_6911,N_5934,N_4636);
or U6912 (N_6912,N_5047,N_4068);
xnor U6913 (N_6913,N_4144,N_5602);
nand U6914 (N_6914,N_4684,N_5711);
xnor U6915 (N_6915,N_4504,N_5827);
and U6916 (N_6916,N_4676,N_4480);
nand U6917 (N_6917,N_5604,N_4085);
nand U6918 (N_6918,N_5306,N_5728);
nand U6919 (N_6919,N_4041,N_5835);
xnor U6920 (N_6920,N_4339,N_4069);
xor U6921 (N_6921,N_5911,N_5319);
xnor U6922 (N_6922,N_5587,N_5968);
or U6923 (N_6923,N_4130,N_5683);
or U6924 (N_6924,N_5006,N_5829);
nor U6925 (N_6925,N_5608,N_5341);
nor U6926 (N_6926,N_5145,N_5110);
nand U6927 (N_6927,N_4062,N_4875);
nand U6928 (N_6928,N_5636,N_4231);
or U6929 (N_6929,N_5086,N_4466);
nand U6930 (N_6930,N_5454,N_4343);
or U6931 (N_6931,N_5294,N_4071);
xor U6932 (N_6932,N_5952,N_5038);
nand U6933 (N_6933,N_5714,N_5076);
xor U6934 (N_6934,N_4083,N_5494);
nand U6935 (N_6935,N_5198,N_5320);
nor U6936 (N_6936,N_5875,N_5574);
and U6937 (N_6937,N_4972,N_4783);
nand U6938 (N_6938,N_5349,N_4167);
and U6939 (N_6939,N_4296,N_4618);
or U6940 (N_6940,N_4280,N_5681);
and U6941 (N_6941,N_5691,N_4369);
nand U6942 (N_6942,N_5160,N_5561);
nand U6943 (N_6943,N_4646,N_4173);
and U6944 (N_6944,N_4687,N_4202);
nand U6945 (N_6945,N_4431,N_4275);
or U6946 (N_6946,N_4208,N_5559);
nand U6947 (N_6947,N_5196,N_5247);
xor U6948 (N_6948,N_5301,N_5742);
and U6949 (N_6949,N_4558,N_5101);
and U6950 (N_6950,N_4659,N_4991);
xnor U6951 (N_6951,N_4078,N_5799);
nor U6952 (N_6952,N_5540,N_5999);
and U6953 (N_6953,N_5896,N_4399);
nand U6954 (N_6954,N_5905,N_5171);
xor U6955 (N_6955,N_5029,N_5458);
xnor U6956 (N_6956,N_4623,N_4297);
xnor U6957 (N_6957,N_4105,N_4221);
xnor U6958 (N_6958,N_4092,N_5392);
or U6959 (N_6959,N_5541,N_4402);
and U6960 (N_6960,N_5847,N_5853);
and U6961 (N_6961,N_4812,N_4446);
xnor U6962 (N_6962,N_5954,N_5197);
and U6963 (N_6963,N_4760,N_4893);
nor U6964 (N_6964,N_5119,N_4294);
and U6965 (N_6965,N_5384,N_4103);
nand U6966 (N_6966,N_4509,N_4673);
and U6967 (N_6967,N_5370,N_4324);
nor U6968 (N_6968,N_4286,N_5193);
or U6969 (N_6969,N_5339,N_4276);
nor U6970 (N_6970,N_5584,N_5804);
xor U6971 (N_6971,N_4786,N_4412);
nand U6972 (N_6972,N_4782,N_4547);
nor U6973 (N_6973,N_4970,N_5438);
or U6974 (N_6974,N_5351,N_5786);
and U6975 (N_6975,N_4086,N_4784);
and U6976 (N_6976,N_4926,N_5537);
nor U6977 (N_6977,N_4449,N_4834);
nand U6978 (N_6978,N_5360,N_4356);
xnor U6979 (N_6979,N_4620,N_5366);
and U6980 (N_6980,N_4394,N_4681);
nand U6981 (N_6981,N_5937,N_4430);
or U6982 (N_6982,N_5941,N_5462);
nor U6983 (N_6983,N_5138,N_5824);
and U6984 (N_6984,N_5510,N_4037);
nor U6985 (N_6985,N_5692,N_5450);
and U6986 (N_6986,N_5473,N_5430);
nor U6987 (N_6987,N_5582,N_4863);
xnor U6988 (N_6988,N_4223,N_4189);
nand U6989 (N_6989,N_5815,N_5801);
or U6990 (N_6990,N_5706,N_5163);
nand U6991 (N_6991,N_4752,N_5176);
nor U6992 (N_6992,N_5945,N_4327);
xor U6993 (N_6993,N_4011,N_4557);
or U6994 (N_6994,N_5844,N_5560);
and U6995 (N_6995,N_4049,N_4377);
or U6996 (N_6996,N_4447,N_4312);
and U6997 (N_6997,N_4856,N_4554);
nor U6998 (N_6998,N_5419,N_5779);
xor U6999 (N_6999,N_5058,N_4820);
or U7000 (N_7000,N_4455,N_5275);
and U7001 (N_7001,N_5424,N_4514);
and U7002 (N_7002,N_5973,N_5320);
or U7003 (N_7003,N_5407,N_4067);
xnor U7004 (N_7004,N_5126,N_4751);
nand U7005 (N_7005,N_4394,N_4125);
or U7006 (N_7006,N_5341,N_5291);
xor U7007 (N_7007,N_4157,N_5684);
xnor U7008 (N_7008,N_4698,N_5601);
and U7009 (N_7009,N_5654,N_4618);
and U7010 (N_7010,N_5280,N_5622);
or U7011 (N_7011,N_5951,N_5509);
xnor U7012 (N_7012,N_5528,N_4891);
and U7013 (N_7013,N_5654,N_4422);
and U7014 (N_7014,N_5298,N_4960);
nand U7015 (N_7015,N_5737,N_4760);
or U7016 (N_7016,N_4384,N_5050);
xor U7017 (N_7017,N_5886,N_4846);
nor U7018 (N_7018,N_5466,N_5438);
nor U7019 (N_7019,N_5319,N_5459);
or U7020 (N_7020,N_5389,N_4023);
xor U7021 (N_7021,N_4460,N_4838);
xnor U7022 (N_7022,N_5017,N_5024);
nand U7023 (N_7023,N_4817,N_5073);
and U7024 (N_7024,N_4874,N_5253);
or U7025 (N_7025,N_5250,N_5998);
and U7026 (N_7026,N_5901,N_4952);
xnor U7027 (N_7027,N_5409,N_4526);
xor U7028 (N_7028,N_4092,N_5810);
and U7029 (N_7029,N_5209,N_5650);
nand U7030 (N_7030,N_4128,N_5901);
xor U7031 (N_7031,N_5727,N_5556);
nor U7032 (N_7032,N_4279,N_5284);
nand U7033 (N_7033,N_5194,N_5457);
nand U7034 (N_7034,N_4596,N_4344);
and U7035 (N_7035,N_4519,N_5313);
nor U7036 (N_7036,N_5030,N_5764);
nor U7037 (N_7037,N_5072,N_5687);
nand U7038 (N_7038,N_5416,N_5829);
or U7039 (N_7039,N_5835,N_4349);
xnor U7040 (N_7040,N_4054,N_5055);
and U7041 (N_7041,N_4034,N_4795);
or U7042 (N_7042,N_4128,N_5612);
or U7043 (N_7043,N_4661,N_4356);
xnor U7044 (N_7044,N_5715,N_5924);
xnor U7045 (N_7045,N_5396,N_5438);
nor U7046 (N_7046,N_4058,N_5339);
nor U7047 (N_7047,N_5216,N_5194);
nor U7048 (N_7048,N_5704,N_4329);
or U7049 (N_7049,N_5871,N_5177);
or U7050 (N_7050,N_5394,N_4500);
nor U7051 (N_7051,N_4114,N_4700);
nand U7052 (N_7052,N_5433,N_5311);
and U7053 (N_7053,N_4561,N_5577);
xor U7054 (N_7054,N_4860,N_4467);
or U7055 (N_7055,N_5165,N_5413);
nor U7056 (N_7056,N_4270,N_4211);
and U7057 (N_7057,N_4007,N_4032);
or U7058 (N_7058,N_5470,N_5075);
nand U7059 (N_7059,N_4701,N_5561);
and U7060 (N_7060,N_5989,N_4670);
and U7061 (N_7061,N_5462,N_5743);
nor U7062 (N_7062,N_5859,N_4910);
xor U7063 (N_7063,N_4858,N_4464);
nand U7064 (N_7064,N_5607,N_5890);
nand U7065 (N_7065,N_4278,N_4631);
and U7066 (N_7066,N_4795,N_4842);
and U7067 (N_7067,N_5469,N_4643);
nand U7068 (N_7068,N_4155,N_5170);
nor U7069 (N_7069,N_5474,N_5012);
and U7070 (N_7070,N_4294,N_4843);
xnor U7071 (N_7071,N_4644,N_4531);
and U7072 (N_7072,N_5214,N_5578);
nand U7073 (N_7073,N_4850,N_5139);
and U7074 (N_7074,N_5717,N_4402);
and U7075 (N_7075,N_4830,N_4106);
xor U7076 (N_7076,N_5925,N_4609);
or U7077 (N_7077,N_5473,N_5429);
and U7078 (N_7078,N_4737,N_5774);
nor U7079 (N_7079,N_5143,N_4581);
xnor U7080 (N_7080,N_5941,N_4041);
or U7081 (N_7081,N_5692,N_4401);
or U7082 (N_7082,N_4173,N_4697);
and U7083 (N_7083,N_5028,N_5057);
xor U7084 (N_7084,N_4279,N_4092);
nand U7085 (N_7085,N_4094,N_5227);
xnor U7086 (N_7086,N_4494,N_5490);
nor U7087 (N_7087,N_5047,N_4940);
and U7088 (N_7088,N_4778,N_5086);
xor U7089 (N_7089,N_4005,N_5684);
xor U7090 (N_7090,N_5265,N_5342);
or U7091 (N_7091,N_5026,N_4486);
or U7092 (N_7092,N_4146,N_4483);
nor U7093 (N_7093,N_4969,N_5987);
nor U7094 (N_7094,N_5706,N_4480);
and U7095 (N_7095,N_4661,N_4081);
nand U7096 (N_7096,N_5333,N_4754);
xnor U7097 (N_7097,N_4488,N_4794);
xor U7098 (N_7098,N_4392,N_4518);
or U7099 (N_7099,N_5682,N_4262);
and U7100 (N_7100,N_5551,N_4641);
or U7101 (N_7101,N_4678,N_4323);
xnor U7102 (N_7102,N_4116,N_4311);
xnor U7103 (N_7103,N_4758,N_5047);
nor U7104 (N_7104,N_5909,N_5916);
or U7105 (N_7105,N_4209,N_5719);
nor U7106 (N_7106,N_4038,N_4729);
and U7107 (N_7107,N_5966,N_5443);
and U7108 (N_7108,N_4736,N_5276);
xor U7109 (N_7109,N_4905,N_5484);
nand U7110 (N_7110,N_4748,N_4062);
nor U7111 (N_7111,N_4422,N_4736);
nor U7112 (N_7112,N_5099,N_4935);
nand U7113 (N_7113,N_4912,N_4661);
nor U7114 (N_7114,N_5405,N_4192);
nor U7115 (N_7115,N_5319,N_5155);
and U7116 (N_7116,N_4732,N_4068);
nor U7117 (N_7117,N_5531,N_4099);
nand U7118 (N_7118,N_5468,N_5714);
and U7119 (N_7119,N_5159,N_4528);
nor U7120 (N_7120,N_5218,N_4373);
nand U7121 (N_7121,N_4339,N_5424);
or U7122 (N_7122,N_5629,N_4120);
and U7123 (N_7123,N_5357,N_5941);
and U7124 (N_7124,N_4889,N_5562);
xnor U7125 (N_7125,N_4863,N_5539);
or U7126 (N_7126,N_5379,N_4001);
nor U7127 (N_7127,N_4613,N_4740);
xnor U7128 (N_7128,N_5174,N_4252);
xnor U7129 (N_7129,N_4876,N_5083);
xor U7130 (N_7130,N_4219,N_4624);
xnor U7131 (N_7131,N_4774,N_4139);
nor U7132 (N_7132,N_5670,N_5571);
or U7133 (N_7133,N_5838,N_4151);
or U7134 (N_7134,N_5397,N_5729);
and U7135 (N_7135,N_4807,N_5596);
xor U7136 (N_7136,N_4529,N_5223);
and U7137 (N_7137,N_5561,N_4252);
or U7138 (N_7138,N_5121,N_5207);
xor U7139 (N_7139,N_4467,N_5339);
xnor U7140 (N_7140,N_4013,N_4847);
nor U7141 (N_7141,N_4758,N_4974);
or U7142 (N_7142,N_5168,N_4934);
xnor U7143 (N_7143,N_4844,N_4103);
xor U7144 (N_7144,N_5063,N_4926);
nor U7145 (N_7145,N_4116,N_4603);
nand U7146 (N_7146,N_4893,N_5897);
or U7147 (N_7147,N_4754,N_4047);
or U7148 (N_7148,N_4373,N_5940);
nand U7149 (N_7149,N_5875,N_4401);
xor U7150 (N_7150,N_5975,N_4053);
and U7151 (N_7151,N_4083,N_5054);
xnor U7152 (N_7152,N_5572,N_5915);
or U7153 (N_7153,N_5762,N_5295);
nor U7154 (N_7154,N_4541,N_4284);
or U7155 (N_7155,N_4786,N_5743);
or U7156 (N_7156,N_4128,N_5894);
and U7157 (N_7157,N_5815,N_4530);
or U7158 (N_7158,N_5895,N_4957);
or U7159 (N_7159,N_5092,N_5519);
nand U7160 (N_7160,N_4622,N_4856);
nor U7161 (N_7161,N_5713,N_5920);
xor U7162 (N_7162,N_5933,N_5806);
xnor U7163 (N_7163,N_4659,N_5983);
and U7164 (N_7164,N_5639,N_4930);
nand U7165 (N_7165,N_5579,N_5674);
xor U7166 (N_7166,N_5456,N_4809);
or U7167 (N_7167,N_5639,N_5951);
nor U7168 (N_7168,N_4714,N_4210);
nand U7169 (N_7169,N_4158,N_4207);
xnor U7170 (N_7170,N_5522,N_5274);
nand U7171 (N_7171,N_5949,N_4695);
xor U7172 (N_7172,N_4624,N_5797);
nand U7173 (N_7173,N_4418,N_5699);
xnor U7174 (N_7174,N_5814,N_5223);
or U7175 (N_7175,N_5979,N_4910);
or U7176 (N_7176,N_5799,N_5374);
or U7177 (N_7177,N_4655,N_4183);
nand U7178 (N_7178,N_5919,N_4283);
xor U7179 (N_7179,N_5346,N_4002);
and U7180 (N_7180,N_5499,N_5123);
and U7181 (N_7181,N_4067,N_4180);
nor U7182 (N_7182,N_5412,N_4083);
xnor U7183 (N_7183,N_5257,N_5532);
nand U7184 (N_7184,N_5368,N_5860);
xor U7185 (N_7185,N_5846,N_5949);
nor U7186 (N_7186,N_5941,N_5602);
or U7187 (N_7187,N_5429,N_5065);
and U7188 (N_7188,N_4475,N_5947);
and U7189 (N_7189,N_4479,N_5805);
nor U7190 (N_7190,N_5660,N_5852);
nor U7191 (N_7191,N_4950,N_4831);
and U7192 (N_7192,N_4144,N_5684);
and U7193 (N_7193,N_4440,N_5355);
or U7194 (N_7194,N_4569,N_4344);
nand U7195 (N_7195,N_4872,N_4741);
and U7196 (N_7196,N_4929,N_4520);
or U7197 (N_7197,N_4591,N_4043);
nand U7198 (N_7198,N_5650,N_4188);
xor U7199 (N_7199,N_5456,N_4127);
or U7200 (N_7200,N_4559,N_5423);
nor U7201 (N_7201,N_4072,N_5486);
xnor U7202 (N_7202,N_4642,N_5308);
or U7203 (N_7203,N_5227,N_5716);
xor U7204 (N_7204,N_5986,N_5779);
nand U7205 (N_7205,N_4983,N_5879);
nor U7206 (N_7206,N_5135,N_5336);
or U7207 (N_7207,N_5760,N_4610);
xnor U7208 (N_7208,N_4948,N_5700);
or U7209 (N_7209,N_4587,N_5154);
and U7210 (N_7210,N_5135,N_4830);
nand U7211 (N_7211,N_4207,N_4672);
and U7212 (N_7212,N_5387,N_4584);
xnor U7213 (N_7213,N_5498,N_4932);
and U7214 (N_7214,N_5033,N_4456);
and U7215 (N_7215,N_4357,N_5377);
or U7216 (N_7216,N_5261,N_5143);
xnor U7217 (N_7217,N_5377,N_5138);
nand U7218 (N_7218,N_5043,N_4157);
or U7219 (N_7219,N_4093,N_4876);
xnor U7220 (N_7220,N_5699,N_4121);
and U7221 (N_7221,N_4841,N_4891);
xor U7222 (N_7222,N_4057,N_4888);
nand U7223 (N_7223,N_4602,N_5530);
or U7224 (N_7224,N_4907,N_4277);
and U7225 (N_7225,N_4209,N_5016);
and U7226 (N_7226,N_4418,N_4372);
or U7227 (N_7227,N_5507,N_5794);
nand U7228 (N_7228,N_4903,N_5068);
and U7229 (N_7229,N_5727,N_5892);
or U7230 (N_7230,N_4435,N_5330);
and U7231 (N_7231,N_5915,N_5565);
or U7232 (N_7232,N_5867,N_4264);
nor U7233 (N_7233,N_4328,N_5069);
or U7234 (N_7234,N_4412,N_4187);
or U7235 (N_7235,N_5582,N_5946);
nand U7236 (N_7236,N_5818,N_5008);
and U7237 (N_7237,N_4545,N_5777);
or U7238 (N_7238,N_5907,N_5037);
xnor U7239 (N_7239,N_4801,N_5540);
and U7240 (N_7240,N_5452,N_4604);
nor U7241 (N_7241,N_5581,N_5598);
xnor U7242 (N_7242,N_5290,N_4573);
xnor U7243 (N_7243,N_4659,N_4617);
nand U7244 (N_7244,N_5018,N_4691);
nand U7245 (N_7245,N_5073,N_5112);
nand U7246 (N_7246,N_4738,N_5264);
or U7247 (N_7247,N_5967,N_5050);
nand U7248 (N_7248,N_4468,N_4620);
nor U7249 (N_7249,N_4306,N_5298);
xor U7250 (N_7250,N_5565,N_4269);
nor U7251 (N_7251,N_4847,N_5448);
and U7252 (N_7252,N_5163,N_4589);
or U7253 (N_7253,N_4990,N_4472);
nand U7254 (N_7254,N_4539,N_4555);
nand U7255 (N_7255,N_4889,N_5688);
nand U7256 (N_7256,N_4339,N_5987);
and U7257 (N_7257,N_4774,N_4301);
and U7258 (N_7258,N_5972,N_5942);
and U7259 (N_7259,N_4974,N_4270);
nor U7260 (N_7260,N_5506,N_5482);
xor U7261 (N_7261,N_4121,N_4774);
or U7262 (N_7262,N_5163,N_5255);
nand U7263 (N_7263,N_4614,N_5156);
or U7264 (N_7264,N_5426,N_5199);
or U7265 (N_7265,N_4922,N_5844);
xor U7266 (N_7266,N_4102,N_4364);
xor U7267 (N_7267,N_5128,N_5477);
nor U7268 (N_7268,N_4931,N_4309);
or U7269 (N_7269,N_5408,N_4144);
and U7270 (N_7270,N_5860,N_4748);
nand U7271 (N_7271,N_4070,N_4174);
and U7272 (N_7272,N_4503,N_5632);
xor U7273 (N_7273,N_4660,N_5652);
nor U7274 (N_7274,N_4045,N_5592);
or U7275 (N_7275,N_4700,N_4018);
or U7276 (N_7276,N_4670,N_4809);
and U7277 (N_7277,N_5797,N_4152);
xnor U7278 (N_7278,N_4309,N_4639);
nor U7279 (N_7279,N_5970,N_5832);
and U7280 (N_7280,N_5079,N_4216);
and U7281 (N_7281,N_5349,N_5788);
and U7282 (N_7282,N_4867,N_5042);
nand U7283 (N_7283,N_4596,N_4107);
or U7284 (N_7284,N_4105,N_4553);
or U7285 (N_7285,N_5544,N_5886);
and U7286 (N_7286,N_5748,N_4170);
xor U7287 (N_7287,N_4554,N_5118);
and U7288 (N_7288,N_5881,N_4514);
and U7289 (N_7289,N_4026,N_5228);
nor U7290 (N_7290,N_5668,N_5685);
and U7291 (N_7291,N_5503,N_4063);
or U7292 (N_7292,N_5921,N_4720);
nand U7293 (N_7293,N_5230,N_5559);
nand U7294 (N_7294,N_5186,N_5117);
nand U7295 (N_7295,N_5724,N_5571);
nor U7296 (N_7296,N_4018,N_4332);
and U7297 (N_7297,N_5477,N_4550);
nand U7298 (N_7298,N_4186,N_5097);
xnor U7299 (N_7299,N_5554,N_4241);
or U7300 (N_7300,N_4548,N_4545);
nor U7301 (N_7301,N_5016,N_5468);
nor U7302 (N_7302,N_5627,N_5718);
nor U7303 (N_7303,N_4169,N_5681);
xor U7304 (N_7304,N_5901,N_4522);
and U7305 (N_7305,N_4572,N_5447);
xnor U7306 (N_7306,N_4123,N_4266);
xnor U7307 (N_7307,N_5408,N_4005);
nor U7308 (N_7308,N_4346,N_4582);
and U7309 (N_7309,N_5105,N_5465);
nand U7310 (N_7310,N_4523,N_4730);
or U7311 (N_7311,N_5660,N_5099);
or U7312 (N_7312,N_5936,N_5614);
nor U7313 (N_7313,N_5210,N_5096);
xnor U7314 (N_7314,N_5477,N_4644);
xnor U7315 (N_7315,N_4027,N_5042);
nand U7316 (N_7316,N_4782,N_4938);
nor U7317 (N_7317,N_5585,N_4298);
nor U7318 (N_7318,N_5341,N_4091);
nand U7319 (N_7319,N_4248,N_4128);
nor U7320 (N_7320,N_4736,N_4375);
nor U7321 (N_7321,N_4803,N_5939);
nand U7322 (N_7322,N_4158,N_5470);
nor U7323 (N_7323,N_4119,N_5828);
and U7324 (N_7324,N_5574,N_4607);
nand U7325 (N_7325,N_5867,N_5689);
or U7326 (N_7326,N_5985,N_5157);
and U7327 (N_7327,N_4622,N_4246);
and U7328 (N_7328,N_4525,N_4256);
nor U7329 (N_7329,N_5999,N_4158);
or U7330 (N_7330,N_5370,N_5409);
nor U7331 (N_7331,N_5904,N_5777);
nand U7332 (N_7332,N_4337,N_5743);
and U7333 (N_7333,N_5768,N_4440);
or U7334 (N_7334,N_4318,N_5089);
xnor U7335 (N_7335,N_4349,N_5887);
and U7336 (N_7336,N_5691,N_4687);
or U7337 (N_7337,N_4701,N_4013);
and U7338 (N_7338,N_4819,N_4328);
and U7339 (N_7339,N_5553,N_5957);
nand U7340 (N_7340,N_5943,N_5476);
nand U7341 (N_7341,N_5537,N_4334);
or U7342 (N_7342,N_4754,N_4509);
and U7343 (N_7343,N_4357,N_4494);
xnor U7344 (N_7344,N_4019,N_4064);
xnor U7345 (N_7345,N_4256,N_5786);
xnor U7346 (N_7346,N_4585,N_4375);
xor U7347 (N_7347,N_5262,N_5509);
or U7348 (N_7348,N_4074,N_5912);
xnor U7349 (N_7349,N_5620,N_4979);
nand U7350 (N_7350,N_4177,N_5547);
nand U7351 (N_7351,N_5260,N_4570);
nand U7352 (N_7352,N_5833,N_5112);
or U7353 (N_7353,N_4918,N_5550);
xor U7354 (N_7354,N_4852,N_4394);
nand U7355 (N_7355,N_4719,N_4682);
xor U7356 (N_7356,N_5701,N_4557);
and U7357 (N_7357,N_5510,N_5621);
and U7358 (N_7358,N_4043,N_4992);
and U7359 (N_7359,N_5047,N_4770);
nor U7360 (N_7360,N_4797,N_5658);
nor U7361 (N_7361,N_5265,N_5228);
and U7362 (N_7362,N_5582,N_4901);
xor U7363 (N_7363,N_5857,N_5037);
and U7364 (N_7364,N_4056,N_4850);
nor U7365 (N_7365,N_4746,N_4026);
and U7366 (N_7366,N_4760,N_5363);
or U7367 (N_7367,N_5963,N_4723);
nand U7368 (N_7368,N_4130,N_4565);
nor U7369 (N_7369,N_4899,N_4755);
nand U7370 (N_7370,N_4514,N_5962);
and U7371 (N_7371,N_4795,N_4232);
xnor U7372 (N_7372,N_5750,N_5363);
nor U7373 (N_7373,N_5813,N_4101);
xnor U7374 (N_7374,N_5449,N_4843);
or U7375 (N_7375,N_5572,N_5234);
or U7376 (N_7376,N_5462,N_4526);
xnor U7377 (N_7377,N_5493,N_4426);
or U7378 (N_7378,N_5680,N_4722);
nand U7379 (N_7379,N_5690,N_4434);
and U7380 (N_7380,N_5524,N_4049);
nand U7381 (N_7381,N_5582,N_5992);
nand U7382 (N_7382,N_5819,N_4226);
xnor U7383 (N_7383,N_4321,N_5119);
xnor U7384 (N_7384,N_5631,N_5794);
and U7385 (N_7385,N_4885,N_5838);
and U7386 (N_7386,N_4630,N_5716);
nand U7387 (N_7387,N_5135,N_5933);
nand U7388 (N_7388,N_4489,N_4233);
and U7389 (N_7389,N_5144,N_4880);
and U7390 (N_7390,N_4301,N_4345);
and U7391 (N_7391,N_5619,N_5419);
xor U7392 (N_7392,N_4579,N_5948);
xnor U7393 (N_7393,N_4408,N_4148);
nand U7394 (N_7394,N_5982,N_4234);
or U7395 (N_7395,N_5129,N_4080);
xor U7396 (N_7396,N_4549,N_4780);
xnor U7397 (N_7397,N_5971,N_4662);
nand U7398 (N_7398,N_4357,N_5746);
xnor U7399 (N_7399,N_5234,N_5344);
nor U7400 (N_7400,N_5585,N_4792);
nor U7401 (N_7401,N_4989,N_4889);
or U7402 (N_7402,N_4722,N_5544);
or U7403 (N_7403,N_4851,N_5123);
xor U7404 (N_7404,N_4149,N_5428);
xor U7405 (N_7405,N_5165,N_4953);
and U7406 (N_7406,N_4046,N_4515);
or U7407 (N_7407,N_4697,N_4133);
nor U7408 (N_7408,N_4505,N_5609);
and U7409 (N_7409,N_5501,N_5334);
nand U7410 (N_7410,N_4308,N_5030);
xor U7411 (N_7411,N_5045,N_4894);
nand U7412 (N_7412,N_5220,N_5982);
nor U7413 (N_7413,N_5538,N_5032);
xor U7414 (N_7414,N_4039,N_5949);
and U7415 (N_7415,N_5588,N_5855);
xnor U7416 (N_7416,N_5102,N_4821);
or U7417 (N_7417,N_4833,N_4221);
nand U7418 (N_7418,N_4644,N_4045);
and U7419 (N_7419,N_5343,N_5455);
nor U7420 (N_7420,N_5085,N_4412);
and U7421 (N_7421,N_5619,N_4998);
or U7422 (N_7422,N_5754,N_5923);
or U7423 (N_7423,N_4403,N_5339);
nor U7424 (N_7424,N_4529,N_5025);
and U7425 (N_7425,N_4942,N_5035);
or U7426 (N_7426,N_5159,N_4896);
nand U7427 (N_7427,N_5239,N_5168);
and U7428 (N_7428,N_4541,N_5275);
xnor U7429 (N_7429,N_5690,N_4708);
and U7430 (N_7430,N_4895,N_5221);
and U7431 (N_7431,N_5538,N_4281);
nor U7432 (N_7432,N_5511,N_4067);
and U7433 (N_7433,N_5813,N_4637);
or U7434 (N_7434,N_5378,N_5938);
nor U7435 (N_7435,N_4818,N_4971);
or U7436 (N_7436,N_5468,N_5640);
and U7437 (N_7437,N_4943,N_4283);
nand U7438 (N_7438,N_5834,N_5892);
and U7439 (N_7439,N_4529,N_4557);
or U7440 (N_7440,N_4287,N_4911);
nand U7441 (N_7441,N_4376,N_4496);
and U7442 (N_7442,N_5661,N_4187);
and U7443 (N_7443,N_5174,N_5618);
xor U7444 (N_7444,N_4121,N_4905);
nand U7445 (N_7445,N_5082,N_5975);
or U7446 (N_7446,N_5832,N_5804);
nor U7447 (N_7447,N_5716,N_4167);
xnor U7448 (N_7448,N_5437,N_5584);
nor U7449 (N_7449,N_5384,N_4864);
or U7450 (N_7450,N_4034,N_4337);
or U7451 (N_7451,N_4306,N_4335);
and U7452 (N_7452,N_4195,N_5304);
or U7453 (N_7453,N_5753,N_5601);
nand U7454 (N_7454,N_4656,N_5605);
or U7455 (N_7455,N_4218,N_4909);
nand U7456 (N_7456,N_5538,N_4022);
and U7457 (N_7457,N_4788,N_4520);
nor U7458 (N_7458,N_4833,N_5028);
xor U7459 (N_7459,N_5446,N_4844);
and U7460 (N_7460,N_4340,N_5802);
or U7461 (N_7461,N_4523,N_4907);
nor U7462 (N_7462,N_5248,N_5838);
nand U7463 (N_7463,N_4218,N_5517);
or U7464 (N_7464,N_5294,N_5288);
nor U7465 (N_7465,N_4605,N_4097);
xor U7466 (N_7466,N_4594,N_5480);
xor U7467 (N_7467,N_5749,N_4505);
or U7468 (N_7468,N_4913,N_5288);
xor U7469 (N_7469,N_4115,N_5567);
nor U7470 (N_7470,N_4283,N_5290);
or U7471 (N_7471,N_5751,N_5289);
and U7472 (N_7472,N_5033,N_5307);
nor U7473 (N_7473,N_4809,N_4494);
nor U7474 (N_7474,N_4782,N_5339);
nor U7475 (N_7475,N_4914,N_5729);
or U7476 (N_7476,N_4876,N_4688);
xnor U7477 (N_7477,N_5549,N_4840);
and U7478 (N_7478,N_5112,N_5991);
or U7479 (N_7479,N_5606,N_5510);
or U7480 (N_7480,N_4739,N_4091);
and U7481 (N_7481,N_5445,N_4292);
or U7482 (N_7482,N_5822,N_5317);
xor U7483 (N_7483,N_4274,N_4340);
xor U7484 (N_7484,N_5792,N_5145);
xnor U7485 (N_7485,N_4820,N_5812);
and U7486 (N_7486,N_5998,N_4409);
xor U7487 (N_7487,N_5069,N_5725);
nand U7488 (N_7488,N_5948,N_5308);
and U7489 (N_7489,N_4020,N_5184);
xor U7490 (N_7490,N_5786,N_5863);
or U7491 (N_7491,N_4059,N_5304);
and U7492 (N_7492,N_5805,N_4406);
nand U7493 (N_7493,N_4820,N_5241);
or U7494 (N_7494,N_5189,N_4856);
xor U7495 (N_7495,N_5550,N_5807);
xor U7496 (N_7496,N_5540,N_4212);
xnor U7497 (N_7497,N_4573,N_4523);
and U7498 (N_7498,N_5842,N_4494);
and U7499 (N_7499,N_5259,N_4324);
xor U7500 (N_7500,N_5431,N_5447);
nor U7501 (N_7501,N_4609,N_5669);
nor U7502 (N_7502,N_4519,N_4173);
or U7503 (N_7503,N_4735,N_5699);
and U7504 (N_7504,N_4317,N_5599);
nor U7505 (N_7505,N_5293,N_5140);
xor U7506 (N_7506,N_5760,N_5775);
or U7507 (N_7507,N_5907,N_5302);
or U7508 (N_7508,N_4868,N_4640);
or U7509 (N_7509,N_4587,N_4712);
or U7510 (N_7510,N_4241,N_5943);
nand U7511 (N_7511,N_5079,N_4154);
xnor U7512 (N_7512,N_5133,N_5449);
and U7513 (N_7513,N_5246,N_5123);
and U7514 (N_7514,N_4234,N_5732);
nand U7515 (N_7515,N_4886,N_4997);
nor U7516 (N_7516,N_4910,N_5655);
nor U7517 (N_7517,N_5722,N_5853);
and U7518 (N_7518,N_4315,N_5655);
nand U7519 (N_7519,N_5370,N_5949);
xnor U7520 (N_7520,N_4733,N_4573);
xnor U7521 (N_7521,N_4843,N_5398);
or U7522 (N_7522,N_4095,N_4428);
and U7523 (N_7523,N_5372,N_4316);
and U7524 (N_7524,N_5181,N_5064);
nand U7525 (N_7525,N_4222,N_4409);
xor U7526 (N_7526,N_5156,N_5110);
nor U7527 (N_7527,N_5079,N_5274);
xnor U7528 (N_7528,N_5435,N_4470);
nand U7529 (N_7529,N_4607,N_4474);
nand U7530 (N_7530,N_4493,N_4018);
nor U7531 (N_7531,N_4674,N_5190);
nand U7532 (N_7532,N_5148,N_5929);
nand U7533 (N_7533,N_5692,N_5010);
nor U7534 (N_7534,N_5580,N_4518);
nand U7535 (N_7535,N_5374,N_4438);
and U7536 (N_7536,N_5777,N_4441);
xor U7537 (N_7537,N_4816,N_4452);
nor U7538 (N_7538,N_5178,N_5521);
and U7539 (N_7539,N_4423,N_5176);
and U7540 (N_7540,N_4375,N_5451);
nand U7541 (N_7541,N_5789,N_5122);
or U7542 (N_7542,N_4788,N_4457);
or U7543 (N_7543,N_4416,N_5111);
and U7544 (N_7544,N_5968,N_4663);
nor U7545 (N_7545,N_5747,N_4609);
and U7546 (N_7546,N_5516,N_4892);
xnor U7547 (N_7547,N_5883,N_5016);
and U7548 (N_7548,N_5816,N_4863);
nor U7549 (N_7549,N_4499,N_4393);
xor U7550 (N_7550,N_4585,N_5662);
or U7551 (N_7551,N_5239,N_5849);
xor U7552 (N_7552,N_4994,N_4300);
nand U7553 (N_7553,N_5961,N_4139);
nand U7554 (N_7554,N_4565,N_5913);
or U7555 (N_7555,N_5445,N_4990);
xnor U7556 (N_7556,N_4658,N_4024);
xor U7557 (N_7557,N_5343,N_4003);
and U7558 (N_7558,N_5058,N_4482);
and U7559 (N_7559,N_4017,N_5929);
nand U7560 (N_7560,N_4036,N_5242);
nand U7561 (N_7561,N_5213,N_5057);
or U7562 (N_7562,N_4862,N_5258);
xnor U7563 (N_7563,N_5119,N_5370);
or U7564 (N_7564,N_4388,N_4083);
and U7565 (N_7565,N_5138,N_4122);
xor U7566 (N_7566,N_4023,N_5222);
and U7567 (N_7567,N_4200,N_5822);
xnor U7568 (N_7568,N_4539,N_5991);
nand U7569 (N_7569,N_5487,N_4867);
nand U7570 (N_7570,N_4685,N_5815);
xor U7571 (N_7571,N_4009,N_5583);
or U7572 (N_7572,N_5986,N_5675);
nand U7573 (N_7573,N_4729,N_4548);
nand U7574 (N_7574,N_4544,N_5917);
xor U7575 (N_7575,N_4250,N_4913);
nor U7576 (N_7576,N_5031,N_4293);
and U7577 (N_7577,N_4386,N_5191);
nor U7578 (N_7578,N_4809,N_4297);
nor U7579 (N_7579,N_4940,N_5055);
xor U7580 (N_7580,N_5726,N_5020);
xor U7581 (N_7581,N_5920,N_4352);
or U7582 (N_7582,N_5155,N_5390);
nand U7583 (N_7583,N_5844,N_4115);
nor U7584 (N_7584,N_4553,N_4869);
and U7585 (N_7585,N_5214,N_5154);
or U7586 (N_7586,N_5113,N_4160);
nor U7587 (N_7587,N_4715,N_4362);
or U7588 (N_7588,N_4879,N_4805);
nor U7589 (N_7589,N_5419,N_5052);
xnor U7590 (N_7590,N_5821,N_5370);
or U7591 (N_7591,N_5078,N_4525);
and U7592 (N_7592,N_4924,N_5546);
xor U7593 (N_7593,N_4631,N_5105);
and U7594 (N_7594,N_5547,N_5191);
nand U7595 (N_7595,N_4704,N_4525);
nor U7596 (N_7596,N_4306,N_5903);
nand U7597 (N_7597,N_5179,N_5217);
and U7598 (N_7598,N_4466,N_4328);
or U7599 (N_7599,N_5897,N_4742);
nor U7600 (N_7600,N_5991,N_5807);
and U7601 (N_7601,N_5673,N_5151);
or U7602 (N_7602,N_5525,N_4396);
and U7603 (N_7603,N_4266,N_5677);
and U7604 (N_7604,N_5161,N_4336);
xor U7605 (N_7605,N_4618,N_5221);
xor U7606 (N_7606,N_4432,N_5572);
or U7607 (N_7607,N_5209,N_4083);
and U7608 (N_7608,N_5886,N_5319);
xnor U7609 (N_7609,N_5638,N_5602);
or U7610 (N_7610,N_5043,N_4040);
or U7611 (N_7611,N_4178,N_5652);
nand U7612 (N_7612,N_5668,N_5502);
or U7613 (N_7613,N_5916,N_4907);
nand U7614 (N_7614,N_5606,N_5347);
xnor U7615 (N_7615,N_4835,N_4171);
nand U7616 (N_7616,N_4371,N_5837);
and U7617 (N_7617,N_4064,N_5932);
nand U7618 (N_7618,N_5647,N_5257);
or U7619 (N_7619,N_5854,N_4848);
and U7620 (N_7620,N_5853,N_4854);
and U7621 (N_7621,N_4173,N_4712);
xor U7622 (N_7622,N_5325,N_5904);
xnor U7623 (N_7623,N_5478,N_4862);
xor U7624 (N_7624,N_5686,N_4169);
and U7625 (N_7625,N_4809,N_5172);
xor U7626 (N_7626,N_4074,N_5328);
nor U7627 (N_7627,N_4859,N_5500);
and U7628 (N_7628,N_5565,N_5019);
or U7629 (N_7629,N_5855,N_4969);
nor U7630 (N_7630,N_4034,N_5236);
xnor U7631 (N_7631,N_5542,N_4481);
nor U7632 (N_7632,N_5431,N_4727);
or U7633 (N_7633,N_5932,N_5661);
and U7634 (N_7634,N_4765,N_5767);
nor U7635 (N_7635,N_4110,N_4376);
xor U7636 (N_7636,N_5850,N_4964);
or U7637 (N_7637,N_4977,N_5159);
or U7638 (N_7638,N_4676,N_4150);
xnor U7639 (N_7639,N_4154,N_5196);
xnor U7640 (N_7640,N_4934,N_4173);
nor U7641 (N_7641,N_4865,N_5621);
xor U7642 (N_7642,N_4224,N_4761);
and U7643 (N_7643,N_4436,N_4774);
nor U7644 (N_7644,N_5783,N_4417);
nand U7645 (N_7645,N_4725,N_4215);
or U7646 (N_7646,N_5046,N_5547);
nand U7647 (N_7647,N_5962,N_5508);
or U7648 (N_7648,N_5983,N_4256);
and U7649 (N_7649,N_4146,N_4696);
nand U7650 (N_7650,N_5583,N_5214);
nand U7651 (N_7651,N_4504,N_5468);
xnor U7652 (N_7652,N_5258,N_5339);
nand U7653 (N_7653,N_4130,N_4690);
or U7654 (N_7654,N_4172,N_4255);
nand U7655 (N_7655,N_5243,N_5207);
nand U7656 (N_7656,N_5369,N_4866);
and U7657 (N_7657,N_5678,N_5713);
or U7658 (N_7658,N_5331,N_4585);
nor U7659 (N_7659,N_4689,N_5439);
nor U7660 (N_7660,N_4978,N_5530);
nand U7661 (N_7661,N_5176,N_4081);
or U7662 (N_7662,N_5963,N_4038);
or U7663 (N_7663,N_4532,N_5445);
xnor U7664 (N_7664,N_4413,N_5240);
nand U7665 (N_7665,N_5076,N_5013);
nand U7666 (N_7666,N_4400,N_5747);
nand U7667 (N_7667,N_5869,N_4417);
nor U7668 (N_7668,N_4432,N_5558);
or U7669 (N_7669,N_4965,N_4022);
nand U7670 (N_7670,N_4518,N_4763);
and U7671 (N_7671,N_5595,N_5824);
nor U7672 (N_7672,N_4846,N_5242);
and U7673 (N_7673,N_5528,N_5873);
and U7674 (N_7674,N_5371,N_5992);
xnor U7675 (N_7675,N_5468,N_5769);
xor U7676 (N_7676,N_4983,N_5882);
or U7677 (N_7677,N_4400,N_5827);
and U7678 (N_7678,N_5093,N_4517);
or U7679 (N_7679,N_4623,N_5272);
or U7680 (N_7680,N_5392,N_4224);
nand U7681 (N_7681,N_5742,N_4531);
nor U7682 (N_7682,N_4156,N_5017);
nor U7683 (N_7683,N_4362,N_5612);
or U7684 (N_7684,N_5204,N_5601);
and U7685 (N_7685,N_5623,N_4519);
xnor U7686 (N_7686,N_4096,N_5908);
or U7687 (N_7687,N_4150,N_5471);
nor U7688 (N_7688,N_5380,N_4187);
nor U7689 (N_7689,N_4009,N_5195);
and U7690 (N_7690,N_4787,N_4414);
or U7691 (N_7691,N_4342,N_5020);
nand U7692 (N_7692,N_5749,N_5091);
nor U7693 (N_7693,N_5904,N_5330);
or U7694 (N_7694,N_4110,N_4112);
nor U7695 (N_7695,N_4892,N_4665);
nor U7696 (N_7696,N_5984,N_4932);
or U7697 (N_7697,N_4954,N_5895);
xnor U7698 (N_7698,N_4649,N_4240);
and U7699 (N_7699,N_4434,N_4668);
xor U7700 (N_7700,N_4088,N_4995);
or U7701 (N_7701,N_5699,N_4075);
and U7702 (N_7702,N_4101,N_4699);
and U7703 (N_7703,N_4604,N_5937);
nor U7704 (N_7704,N_4092,N_4700);
nor U7705 (N_7705,N_5434,N_4754);
xnor U7706 (N_7706,N_5866,N_4356);
or U7707 (N_7707,N_4184,N_4050);
and U7708 (N_7708,N_5137,N_4941);
nor U7709 (N_7709,N_4330,N_4094);
nor U7710 (N_7710,N_4136,N_5904);
nor U7711 (N_7711,N_5048,N_5453);
and U7712 (N_7712,N_5643,N_5585);
or U7713 (N_7713,N_5203,N_5095);
and U7714 (N_7714,N_4453,N_5122);
nor U7715 (N_7715,N_5758,N_5189);
nand U7716 (N_7716,N_5719,N_4109);
nor U7717 (N_7717,N_5031,N_5258);
and U7718 (N_7718,N_5711,N_4138);
nand U7719 (N_7719,N_5575,N_4099);
nand U7720 (N_7720,N_4626,N_5945);
or U7721 (N_7721,N_5656,N_5671);
nor U7722 (N_7722,N_5286,N_4714);
nor U7723 (N_7723,N_5175,N_5598);
and U7724 (N_7724,N_5169,N_4180);
xor U7725 (N_7725,N_5802,N_4380);
nor U7726 (N_7726,N_5339,N_5164);
nand U7727 (N_7727,N_4151,N_4495);
nor U7728 (N_7728,N_4284,N_4495);
xor U7729 (N_7729,N_5770,N_4365);
xor U7730 (N_7730,N_4477,N_4123);
nand U7731 (N_7731,N_4444,N_5362);
and U7732 (N_7732,N_4914,N_5103);
xor U7733 (N_7733,N_5614,N_5550);
nor U7734 (N_7734,N_4772,N_4774);
nand U7735 (N_7735,N_4141,N_4285);
xnor U7736 (N_7736,N_4583,N_5369);
nand U7737 (N_7737,N_4403,N_4165);
nor U7738 (N_7738,N_5329,N_5306);
nor U7739 (N_7739,N_5641,N_4631);
nor U7740 (N_7740,N_4931,N_5989);
nand U7741 (N_7741,N_5235,N_4620);
nand U7742 (N_7742,N_4221,N_4583);
and U7743 (N_7743,N_4637,N_5849);
xor U7744 (N_7744,N_5230,N_4841);
nand U7745 (N_7745,N_5147,N_5547);
nor U7746 (N_7746,N_5431,N_4457);
or U7747 (N_7747,N_4329,N_4451);
and U7748 (N_7748,N_4737,N_5629);
xor U7749 (N_7749,N_5255,N_4362);
and U7750 (N_7750,N_4667,N_5852);
and U7751 (N_7751,N_4805,N_5954);
nand U7752 (N_7752,N_5894,N_4469);
nand U7753 (N_7753,N_5725,N_5762);
nor U7754 (N_7754,N_5372,N_5041);
nand U7755 (N_7755,N_4105,N_4791);
or U7756 (N_7756,N_5358,N_4729);
or U7757 (N_7757,N_5306,N_4700);
and U7758 (N_7758,N_5104,N_5878);
xor U7759 (N_7759,N_5958,N_5055);
nand U7760 (N_7760,N_4645,N_5072);
and U7761 (N_7761,N_4075,N_5726);
nand U7762 (N_7762,N_5778,N_5289);
xor U7763 (N_7763,N_5986,N_4784);
nand U7764 (N_7764,N_5607,N_5457);
nand U7765 (N_7765,N_4858,N_4910);
nand U7766 (N_7766,N_5563,N_4987);
nand U7767 (N_7767,N_4251,N_4497);
or U7768 (N_7768,N_4664,N_4044);
nand U7769 (N_7769,N_5676,N_5387);
or U7770 (N_7770,N_4078,N_4695);
or U7771 (N_7771,N_5949,N_5274);
nand U7772 (N_7772,N_5188,N_5028);
nand U7773 (N_7773,N_5799,N_5693);
or U7774 (N_7774,N_4528,N_4168);
nand U7775 (N_7775,N_4279,N_5695);
or U7776 (N_7776,N_4437,N_5371);
nand U7777 (N_7777,N_5014,N_4937);
xor U7778 (N_7778,N_5635,N_4029);
nand U7779 (N_7779,N_5759,N_5743);
nand U7780 (N_7780,N_4395,N_4963);
or U7781 (N_7781,N_4468,N_5352);
nand U7782 (N_7782,N_5826,N_4285);
nor U7783 (N_7783,N_4525,N_5646);
xor U7784 (N_7784,N_5378,N_4263);
xor U7785 (N_7785,N_5978,N_4914);
xnor U7786 (N_7786,N_5412,N_4870);
and U7787 (N_7787,N_4202,N_4218);
and U7788 (N_7788,N_5375,N_4217);
nor U7789 (N_7789,N_5461,N_4269);
nor U7790 (N_7790,N_4147,N_5494);
nor U7791 (N_7791,N_5680,N_4156);
and U7792 (N_7792,N_4142,N_4241);
xnor U7793 (N_7793,N_5586,N_4942);
nand U7794 (N_7794,N_5361,N_5164);
nor U7795 (N_7795,N_4436,N_4296);
xor U7796 (N_7796,N_4981,N_4904);
xnor U7797 (N_7797,N_5942,N_5394);
or U7798 (N_7798,N_4431,N_5518);
xnor U7799 (N_7799,N_4730,N_4336);
nand U7800 (N_7800,N_5443,N_5592);
or U7801 (N_7801,N_5871,N_5628);
nand U7802 (N_7802,N_5581,N_5134);
xor U7803 (N_7803,N_5673,N_4378);
or U7804 (N_7804,N_4482,N_5299);
nor U7805 (N_7805,N_5552,N_4731);
xnor U7806 (N_7806,N_4973,N_4777);
xnor U7807 (N_7807,N_5774,N_5900);
nor U7808 (N_7808,N_5676,N_5903);
and U7809 (N_7809,N_5519,N_4508);
or U7810 (N_7810,N_4437,N_5606);
or U7811 (N_7811,N_5080,N_5652);
nand U7812 (N_7812,N_5124,N_5401);
or U7813 (N_7813,N_5896,N_4173);
nand U7814 (N_7814,N_5255,N_5518);
or U7815 (N_7815,N_5472,N_4440);
and U7816 (N_7816,N_5417,N_5520);
xnor U7817 (N_7817,N_4993,N_5231);
xnor U7818 (N_7818,N_5256,N_5529);
or U7819 (N_7819,N_5755,N_5856);
xnor U7820 (N_7820,N_5613,N_4331);
xnor U7821 (N_7821,N_4720,N_5909);
nand U7822 (N_7822,N_4846,N_5769);
nand U7823 (N_7823,N_4841,N_4881);
and U7824 (N_7824,N_4578,N_5244);
nor U7825 (N_7825,N_5813,N_5577);
or U7826 (N_7826,N_5299,N_4319);
and U7827 (N_7827,N_4893,N_4252);
xor U7828 (N_7828,N_5192,N_4041);
xnor U7829 (N_7829,N_5117,N_5520);
or U7830 (N_7830,N_5945,N_4217);
nand U7831 (N_7831,N_4028,N_4942);
xnor U7832 (N_7832,N_4149,N_4852);
and U7833 (N_7833,N_5832,N_5739);
xnor U7834 (N_7834,N_4114,N_5892);
and U7835 (N_7835,N_4873,N_5159);
nand U7836 (N_7836,N_4586,N_4232);
xnor U7837 (N_7837,N_5553,N_4282);
nand U7838 (N_7838,N_5443,N_4405);
or U7839 (N_7839,N_5462,N_5087);
xnor U7840 (N_7840,N_4541,N_4374);
nor U7841 (N_7841,N_5265,N_4201);
xnor U7842 (N_7842,N_4421,N_5354);
and U7843 (N_7843,N_5566,N_4132);
xor U7844 (N_7844,N_4685,N_4499);
xor U7845 (N_7845,N_5965,N_4582);
nor U7846 (N_7846,N_4664,N_4769);
xor U7847 (N_7847,N_4394,N_5526);
xnor U7848 (N_7848,N_5993,N_4576);
nand U7849 (N_7849,N_4996,N_5785);
nor U7850 (N_7850,N_5749,N_5976);
nand U7851 (N_7851,N_4940,N_4190);
nand U7852 (N_7852,N_5399,N_4618);
and U7853 (N_7853,N_5378,N_5874);
nor U7854 (N_7854,N_4918,N_4436);
nor U7855 (N_7855,N_5625,N_4431);
nor U7856 (N_7856,N_5991,N_4070);
xnor U7857 (N_7857,N_4399,N_5877);
or U7858 (N_7858,N_5093,N_4207);
xnor U7859 (N_7859,N_4604,N_5944);
nand U7860 (N_7860,N_5542,N_4739);
and U7861 (N_7861,N_4683,N_4361);
nor U7862 (N_7862,N_4780,N_5008);
nor U7863 (N_7863,N_5818,N_4383);
nand U7864 (N_7864,N_5141,N_4845);
or U7865 (N_7865,N_4030,N_4409);
nor U7866 (N_7866,N_5199,N_4516);
or U7867 (N_7867,N_5306,N_4976);
nor U7868 (N_7868,N_4116,N_5669);
or U7869 (N_7869,N_4153,N_4438);
or U7870 (N_7870,N_5181,N_5242);
nand U7871 (N_7871,N_5280,N_4527);
and U7872 (N_7872,N_4618,N_5317);
or U7873 (N_7873,N_5406,N_4454);
or U7874 (N_7874,N_5225,N_5022);
xor U7875 (N_7875,N_5070,N_5983);
or U7876 (N_7876,N_4003,N_4214);
and U7877 (N_7877,N_4179,N_4825);
nor U7878 (N_7878,N_5255,N_4419);
and U7879 (N_7879,N_5979,N_4176);
xor U7880 (N_7880,N_5929,N_5685);
nand U7881 (N_7881,N_4623,N_5851);
xnor U7882 (N_7882,N_5768,N_5003);
or U7883 (N_7883,N_4873,N_5633);
nor U7884 (N_7884,N_5563,N_4977);
nand U7885 (N_7885,N_5238,N_4885);
or U7886 (N_7886,N_5083,N_5886);
xor U7887 (N_7887,N_5013,N_4578);
and U7888 (N_7888,N_5447,N_5278);
xor U7889 (N_7889,N_4264,N_5068);
xnor U7890 (N_7890,N_4257,N_5171);
or U7891 (N_7891,N_4727,N_4491);
and U7892 (N_7892,N_4020,N_4225);
xor U7893 (N_7893,N_4053,N_5630);
nor U7894 (N_7894,N_5030,N_4420);
xnor U7895 (N_7895,N_4148,N_4381);
nor U7896 (N_7896,N_5141,N_4880);
nor U7897 (N_7897,N_4547,N_5174);
nor U7898 (N_7898,N_5727,N_4346);
and U7899 (N_7899,N_5137,N_5643);
and U7900 (N_7900,N_4225,N_4319);
nor U7901 (N_7901,N_5534,N_4497);
or U7902 (N_7902,N_4254,N_5046);
or U7903 (N_7903,N_4621,N_5222);
and U7904 (N_7904,N_4673,N_5182);
or U7905 (N_7905,N_5748,N_5329);
nand U7906 (N_7906,N_5498,N_4955);
nor U7907 (N_7907,N_4182,N_4665);
xnor U7908 (N_7908,N_4566,N_5613);
xor U7909 (N_7909,N_5423,N_4094);
and U7910 (N_7910,N_5062,N_4564);
nor U7911 (N_7911,N_4039,N_4818);
nand U7912 (N_7912,N_5945,N_4645);
nor U7913 (N_7913,N_4114,N_4088);
xor U7914 (N_7914,N_4617,N_4990);
nand U7915 (N_7915,N_4501,N_4688);
nand U7916 (N_7916,N_4404,N_5782);
nand U7917 (N_7917,N_4988,N_4306);
nor U7918 (N_7918,N_4228,N_5355);
or U7919 (N_7919,N_4782,N_5062);
nand U7920 (N_7920,N_4077,N_5130);
xnor U7921 (N_7921,N_5759,N_4853);
or U7922 (N_7922,N_5260,N_5823);
nor U7923 (N_7923,N_4601,N_4250);
nor U7924 (N_7924,N_5609,N_4780);
or U7925 (N_7925,N_5669,N_5224);
or U7926 (N_7926,N_4397,N_4392);
and U7927 (N_7927,N_4147,N_5064);
and U7928 (N_7928,N_4373,N_4033);
xor U7929 (N_7929,N_5848,N_5359);
xor U7930 (N_7930,N_5834,N_5273);
xor U7931 (N_7931,N_4231,N_5892);
nand U7932 (N_7932,N_4814,N_5124);
or U7933 (N_7933,N_4776,N_4174);
nor U7934 (N_7934,N_5018,N_4618);
or U7935 (N_7935,N_4021,N_5163);
xor U7936 (N_7936,N_5696,N_4985);
or U7937 (N_7937,N_5671,N_5378);
xnor U7938 (N_7938,N_5891,N_5046);
nor U7939 (N_7939,N_4186,N_5302);
nor U7940 (N_7940,N_4278,N_5827);
or U7941 (N_7941,N_5065,N_5524);
or U7942 (N_7942,N_5072,N_4130);
nand U7943 (N_7943,N_4676,N_4008);
nor U7944 (N_7944,N_4705,N_5689);
xnor U7945 (N_7945,N_4734,N_4499);
xnor U7946 (N_7946,N_5631,N_5232);
xor U7947 (N_7947,N_4446,N_4110);
or U7948 (N_7948,N_5112,N_4390);
nor U7949 (N_7949,N_4055,N_4812);
xor U7950 (N_7950,N_4901,N_5366);
nor U7951 (N_7951,N_5827,N_5118);
nor U7952 (N_7952,N_4704,N_5063);
and U7953 (N_7953,N_4873,N_4632);
and U7954 (N_7954,N_4649,N_5534);
nor U7955 (N_7955,N_5159,N_5303);
and U7956 (N_7956,N_4226,N_5416);
nor U7957 (N_7957,N_5338,N_4173);
and U7958 (N_7958,N_5632,N_5175);
and U7959 (N_7959,N_4556,N_5235);
and U7960 (N_7960,N_4399,N_4233);
nand U7961 (N_7961,N_4208,N_5905);
or U7962 (N_7962,N_5262,N_5755);
nand U7963 (N_7963,N_4451,N_5963);
nor U7964 (N_7964,N_5360,N_4747);
or U7965 (N_7965,N_4683,N_4307);
nand U7966 (N_7966,N_5676,N_5747);
xor U7967 (N_7967,N_4244,N_5535);
and U7968 (N_7968,N_5093,N_5061);
nor U7969 (N_7969,N_5885,N_5406);
or U7970 (N_7970,N_4486,N_4139);
xor U7971 (N_7971,N_4214,N_5385);
nand U7972 (N_7972,N_4938,N_4715);
nor U7973 (N_7973,N_5290,N_5226);
nand U7974 (N_7974,N_5239,N_4579);
nand U7975 (N_7975,N_5509,N_5891);
and U7976 (N_7976,N_4366,N_4111);
nand U7977 (N_7977,N_4207,N_4323);
and U7978 (N_7978,N_4388,N_4505);
or U7979 (N_7979,N_4945,N_5357);
or U7980 (N_7980,N_5198,N_4906);
nand U7981 (N_7981,N_5902,N_5261);
or U7982 (N_7982,N_4353,N_4410);
and U7983 (N_7983,N_4948,N_5909);
nand U7984 (N_7984,N_4192,N_5958);
nor U7985 (N_7985,N_5599,N_5833);
nor U7986 (N_7986,N_5158,N_5689);
or U7987 (N_7987,N_5628,N_5457);
or U7988 (N_7988,N_5168,N_4806);
xnor U7989 (N_7989,N_5402,N_4358);
nor U7990 (N_7990,N_5393,N_5902);
xnor U7991 (N_7991,N_4719,N_5276);
nand U7992 (N_7992,N_4990,N_5085);
nor U7993 (N_7993,N_4418,N_5165);
xnor U7994 (N_7994,N_5387,N_4028);
or U7995 (N_7995,N_5107,N_4797);
xnor U7996 (N_7996,N_4061,N_5368);
and U7997 (N_7997,N_4697,N_5723);
xor U7998 (N_7998,N_5697,N_5921);
nor U7999 (N_7999,N_4538,N_4016);
nor U8000 (N_8000,N_6711,N_7850);
xnor U8001 (N_8001,N_7014,N_6139);
nand U8002 (N_8002,N_7409,N_7773);
nand U8003 (N_8003,N_7351,N_7815);
nor U8004 (N_8004,N_7548,N_6461);
nand U8005 (N_8005,N_7027,N_6322);
nor U8006 (N_8006,N_6213,N_7478);
and U8007 (N_8007,N_6613,N_6190);
nor U8008 (N_8008,N_7368,N_7326);
nand U8009 (N_8009,N_6527,N_6567);
or U8010 (N_8010,N_6379,N_7606);
or U8011 (N_8011,N_6976,N_7986);
or U8012 (N_8012,N_6353,N_6437);
nor U8013 (N_8013,N_6151,N_6229);
xnor U8014 (N_8014,N_7953,N_6834);
nand U8015 (N_8015,N_7428,N_6180);
nor U8016 (N_8016,N_7455,N_6061);
and U8017 (N_8017,N_7041,N_7821);
and U8018 (N_8018,N_7392,N_6842);
and U8019 (N_8019,N_6645,N_6354);
nor U8020 (N_8020,N_7774,N_6175);
and U8021 (N_8021,N_7020,N_6516);
or U8022 (N_8022,N_6221,N_6673);
xor U8023 (N_8023,N_7658,N_7803);
nand U8024 (N_8024,N_6226,N_7964);
and U8025 (N_8025,N_6975,N_6666);
or U8026 (N_8026,N_7141,N_7012);
xnor U8027 (N_8027,N_7627,N_6133);
and U8028 (N_8028,N_7717,N_7491);
nor U8029 (N_8029,N_6668,N_7034);
nand U8030 (N_8030,N_7445,N_7853);
or U8031 (N_8031,N_6212,N_6074);
and U8032 (N_8032,N_7019,N_7301);
and U8033 (N_8033,N_7458,N_6559);
and U8034 (N_8034,N_6857,N_7680);
xor U8035 (N_8035,N_7831,N_6441);
and U8036 (N_8036,N_6535,N_6433);
nand U8037 (N_8037,N_7299,N_7010);
or U8038 (N_8038,N_6858,N_6701);
nor U8039 (N_8039,N_7473,N_6272);
nor U8040 (N_8040,N_6562,N_6906);
xor U8041 (N_8041,N_6145,N_7394);
nor U8042 (N_8042,N_6128,N_7250);
xnor U8043 (N_8043,N_6800,N_7227);
nand U8044 (N_8044,N_7684,N_6949);
and U8045 (N_8045,N_7566,N_6455);
xor U8046 (N_8046,N_7869,N_7882);
xnor U8047 (N_8047,N_6291,N_7788);
xor U8048 (N_8048,N_6044,N_7765);
nor U8049 (N_8049,N_7556,N_6189);
nand U8050 (N_8050,N_6958,N_6629);
or U8051 (N_8051,N_6094,N_6801);
or U8052 (N_8052,N_7811,N_6714);
or U8053 (N_8053,N_7183,N_7649);
or U8054 (N_8054,N_7160,N_7600);
xor U8055 (N_8055,N_6928,N_7192);
xnor U8056 (N_8056,N_6796,N_7139);
and U8057 (N_8057,N_7482,N_6258);
nand U8058 (N_8058,N_7834,N_6684);
xnor U8059 (N_8059,N_6112,N_6118);
xnor U8060 (N_8060,N_6298,N_7745);
nand U8061 (N_8061,N_7185,N_7565);
and U8062 (N_8062,N_7492,N_7642);
nor U8063 (N_8063,N_7497,N_7057);
nor U8064 (N_8064,N_6797,N_7637);
and U8065 (N_8065,N_7676,N_6955);
nand U8066 (N_8066,N_7363,N_7349);
nor U8067 (N_8067,N_7925,N_7142);
and U8068 (N_8068,N_6582,N_7345);
and U8069 (N_8069,N_7645,N_7901);
xnor U8070 (N_8070,N_6308,N_6307);
or U8071 (N_8071,N_7650,N_6265);
and U8072 (N_8072,N_6075,N_6847);
xnor U8073 (N_8073,N_7422,N_7644);
nand U8074 (N_8074,N_7885,N_6588);
nand U8075 (N_8075,N_7878,N_6736);
nor U8076 (N_8076,N_6692,N_6373);
and U8077 (N_8077,N_7673,N_6498);
xor U8078 (N_8078,N_7224,N_7144);
nor U8079 (N_8079,N_6843,N_7304);
or U8080 (N_8080,N_7951,N_6695);
or U8081 (N_8081,N_7451,N_7841);
xor U8082 (N_8082,N_6867,N_6915);
or U8083 (N_8083,N_7119,N_7354);
nor U8084 (N_8084,N_7073,N_6886);
or U8085 (N_8085,N_7985,N_6382);
or U8086 (N_8086,N_7694,N_7564);
nor U8087 (N_8087,N_7804,N_7824);
xnor U8088 (N_8088,N_7038,N_6972);
nand U8089 (N_8089,N_6443,N_6740);
and U8090 (N_8090,N_6885,N_7753);
xnor U8091 (N_8091,N_7614,N_7103);
xnor U8092 (N_8092,N_6077,N_7883);
xor U8093 (N_8093,N_7604,N_7947);
nor U8094 (N_8094,N_7782,N_7801);
xor U8095 (N_8095,N_6934,N_6698);
nor U8096 (N_8096,N_6616,N_7714);
or U8097 (N_8097,N_6520,N_6859);
and U8098 (N_8098,N_6158,N_7932);
or U8099 (N_8099,N_6297,N_7449);
or U8100 (N_8100,N_7259,N_7919);
nor U8101 (N_8101,N_6046,N_7091);
or U8102 (N_8102,N_7122,N_6578);
nor U8103 (N_8103,N_7770,N_7105);
nand U8104 (N_8104,N_6770,N_7866);
and U8105 (N_8105,N_7366,N_7311);
and U8106 (N_8106,N_6254,N_6971);
nand U8107 (N_8107,N_7934,N_7738);
nand U8108 (N_8108,N_7570,N_7044);
or U8109 (N_8109,N_7899,N_7598);
and U8110 (N_8110,N_7191,N_6950);
nor U8111 (N_8111,N_6248,N_7529);
nor U8112 (N_8112,N_7987,N_7728);
or U8113 (N_8113,N_7494,N_7337);
or U8114 (N_8114,N_6721,N_7835);
xor U8115 (N_8115,N_7381,N_6123);
xnor U8116 (N_8116,N_6444,N_6561);
and U8117 (N_8117,N_7195,N_6415);
xor U8118 (N_8118,N_6171,N_7528);
nand U8119 (N_8119,N_6596,N_6276);
nor U8120 (N_8120,N_6193,N_6486);
xnor U8121 (N_8121,N_6737,N_6547);
nand U8122 (N_8122,N_6918,N_6533);
nand U8123 (N_8123,N_7416,N_6388);
and U8124 (N_8124,N_7228,N_6176);
nor U8125 (N_8125,N_7164,N_7240);
nor U8126 (N_8126,N_6453,N_7184);
xnor U8127 (N_8127,N_6474,N_6957);
nand U8128 (N_8128,N_6473,N_6984);
xnor U8129 (N_8129,N_7218,N_6321);
and U8130 (N_8130,N_6244,N_7075);
or U8131 (N_8131,N_6704,N_7253);
xor U8132 (N_8132,N_6085,N_7891);
or U8133 (N_8133,N_6787,N_7131);
nor U8134 (N_8134,N_6155,N_6706);
or U8135 (N_8135,N_6497,N_6919);
or U8136 (N_8136,N_6960,N_6925);
nand U8137 (N_8137,N_7467,N_6850);
nand U8138 (N_8138,N_7291,N_7813);
or U8139 (N_8139,N_7173,N_7104);
or U8140 (N_8140,N_6799,N_7531);
nand U8141 (N_8141,N_6700,N_7968);
nor U8142 (N_8142,N_6674,N_7223);
xor U8143 (N_8143,N_6196,N_7602);
xnor U8144 (N_8144,N_6182,N_6439);
or U8145 (N_8145,N_6008,N_6476);
nand U8146 (N_8146,N_7156,N_6006);
nand U8147 (N_8147,N_6719,N_6568);
nor U8148 (N_8148,N_7226,N_6767);
nand U8149 (N_8149,N_7759,N_6048);
nand U8150 (N_8150,N_7630,N_6177);
nor U8151 (N_8151,N_7561,N_7942);
nand U8152 (N_8152,N_6862,N_6848);
nor U8153 (N_8153,N_6785,N_6153);
nor U8154 (N_8154,N_6451,N_6705);
xor U8155 (N_8155,N_6246,N_7403);
or U8156 (N_8156,N_6037,N_7407);
or U8157 (N_8157,N_7360,N_7113);
nand U8158 (N_8158,N_7419,N_7661);
nand U8159 (N_8159,N_6689,N_6198);
nand U8160 (N_8160,N_6845,N_7702);
and U8161 (N_8161,N_6661,N_7065);
nand U8162 (N_8162,N_7413,N_6428);
and U8163 (N_8163,N_7961,N_6286);
nor U8164 (N_8164,N_7646,N_6168);
or U8165 (N_8165,N_6768,N_6129);
nand U8166 (N_8166,N_7359,N_7050);
xnor U8167 (N_8167,N_7999,N_6585);
nand U8168 (N_8168,N_6948,N_7198);
or U8169 (N_8169,N_7798,N_6249);
nor U8170 (N_8170,N_7997,N_6600);
or U8171 (N_8171,N_7086,N_6968);
nor U8172 (N_8172,N_7254,N_7635);
nor U8173 (N_8173,N_7486,N_7468);
nor U8174 (N_8174,N_7314,N_6266);
nor U8175 (N_8175,N_7082,N_6977);
xor U8176 (N_8176,N_6894,N_6622);
or U8177 (N_8177,N_7682,N_7390);
nand U8178 (N_8178,N_7816,N_7843);
or U8179 (N_8179,N_6664,N_6269);
nor U8180 (N_8180,N_7926,N_6369);
or U8181 (N_8181,N_7527,N_6728);
xnor U8182 (N_8182,N_6983,N_7282);
and U8183 (N_8183,N_6341,N_6466);
nand U8184 (N_8184,N_7576,N_7537);
or U8185 (N_8185,N_7387,N_6835);
nor U8186 (N_8186,N_6335,N_6795);
and U8187 (N_8187,N_7775,N_7053);
and U8188 (N_8188,N_6323,N_7323);
xor U8189 (N_8189,N_7006,N_6457);
nand U8190 (N_8190,N_7352,N_6993);
nor U8191 (N_8191,N_7618,N_7232);
nor U8192 (N_8192,N_7205,N_6065);
and U8193 (N_8193,N_7480,N_7905);
and U8194 (N_8194,N_7890,N_6069);
or U8195 (N_8195,N_6927,N_7622);
nor U8196 (N_8196,N_6230,N_7398);
xor U8197 (N_8197,N_6693,N_6606);
or U8198 (N_8198,N_6271,N_7851);
nand U8199 (N_8199,N_6345,N_7791);
nand U8200 (N_8200,N_6691,N_6480);
xor U8201 (N_8201,N_6518,N_6277);
and U8202 (N_8202,N_6270,N_7581);
nor U8203 (N_8203,N_6091,N_6288);
nor U8204 (N_8204,N_7763,N_6199);
nand U8205 (N_8205,N_7330,N_6316);
xnor U8206 (N_8206,N_6510,N_7509);
nand U8207 (N_8207,N_6367,N_6363);
xor U8208 (N_8208,N_6222,N_6365);
xor U8209 (N_8209,N_7401,N_6115);
nor U8210 (N_8210,N_7532,N_7723);
or U8211 (N_8211,N_6471,N_7585);
xnor U8212 (N_8212,N_6519,N_7133);
nand U8213 (N_8213,N_6338,N_6462);
or U8214 (N_8214,N_6765,N_7977);
or U8215 (N_8215,N_7744,N_7426);
nand U8216 (N_8216,N_6334,N_7109);
or U8217 (N_8217,N_7596,N_6192);
xnor U8218 (N_8218,N_6550,N_6206);
nor U8219 (N_8219,N_7251,N_6079);
nand U8220 (N_8220,N_6884,N_7615);
nand U8221 (N_8221,N_7081,N_6090);
nor U8222 (N_8222,N_6106,N_7067);
nand U8223 (N_8223,N_6963,N_7466);
and U8224 (N_8224,N_7263,N_7462);
nor U8225 (N_8225,N_7573,N_7132);
and U8226 (N_8226,N_7167,N_7002);
xor U8227 (N_8227,N_7981,N_6101);
nor U8228 (N_8228,N_6723,N_6598);
and U8229 (N_8229,N_6617,N_7713);
nor U8230 (N_8230,N_7196,N_7092);
xnor U8231 (N_8231,N_7471,N_6463);
nand U8232 (N_8232,N_6204,N_6947);
and U8233 (N_8233,N_6494,N_6408);
nand U8234 (N_8234,N_6836,N_7580);
xnor U8235 (N_8235,N_7209,N_6374);
xnor U8236 (N_8236,N_6003,N_7889);
nand U8237 (N_8237,N_6011,N_6887);
and U8238 (N_8238,N_7178,N_7583);
nand U8239 (N_8239,N_6743,N_7464);
xnor U8240 (N_8240,N_7652,N_7781);
xnor U8241 (N_8241,N_6620,N_7829);
xor U8242 (N_8242,N_7944,N_7767);
nand U8243 (N_8243,N_7000,N_6724);
nand U8244 (N_8244,N_7447,N_7474);
or U8245 (N_8245,N_7219,N_6357);
nor U8246 (N_8246,N_7562,N_7230);
and U8247 (N_8247,N_7921,N_7172);
or U8248 (N_8248,N_7089,N_7749);
nor U8249 (N_8249,N_7538,N_7785);
xor U8250 (N_8250,N_6150,N_6911);
or U8251 (N_8251,N_7024,N_6121);
nand U8252 (N_8252,N_6589,N_6402);
or U8253 (N_8253,N_7935,N_6360);
and U8254 (N_8254,N_7830,N_6166);
and U8255 (N_8255,N_7040,N_6852);
nand U8256 (N_8256,N_6839,N_6031);
or U8257 (N_8257,N_6019,N_7318);
and U8258 (N_8258,N_6794,N_6289);
or U8259 (N_8259,N_7917,N_7106);
or U8260 (N_8260,N_7212,N_6076);
nand U8261 (N_8261,N_7430,N_7324);
or U8262 (N_8262,N_7971,N_6012);
nor U8263 (N_8263,N_6855,N_6105);
xnor U8264 (N_8264,N_6487,N_7856);
nor U8265 (N_8265,N_7595,N_6667);
nor U8266 (N_8266,N_6776,N_6401);
nor U8267 (N_8267,N_7849,N_6631);
nor U8268 (N_8268,N_7707,N_7085);
or U8269 (N_8269,N_7696,N_7769);
or U8270 (N_8270,N_7820,N_6619);
and U8271 (N_8271,N_7377,N_7292);
and U8272 (N_8272,N_7364,N_6570);
xnor U8273 (N_8273,N_7171,N_7382);
or U8274 (N_8274,N_7275,N_6235);
and U8275 (N_8275,N_7779,N_7632);
or U8276 (N_8276,N_7285,N_6716);
nor U8277 (N_8277,N_7698,N_7424);
and U8278 (N_8278,N_6318,N_7385);
or U8279 (N_8279,N_7055,N_7018);
nand U8280 (N_8280,N_6278,N_6515);
or U8281 (N_8281,N_6086,N_7094);
and U8282 (N_8282,N_6897,N_6029);
and U8283 (N_8283,N_7303,N_7189);
and U8284 (N_8284,N_7780,N_7827);
and U8285 (N_8285,N_7099,N_7454);
and U8286 (N_8286,N_6059,N_7902);
nand U8287 (N_8287,N_6904,N_6362);
xor U8288 (N_8288,N_7530,N_6371);
and U8289 (N_8289,N_6707,N_7796);
nor U8290 (N_8290,N_7578,N_6344);
and U8291 (N_8291,N_6818,N_6813);
nor U8292 (N_8292,N_7975,N_7751);
nor U8293 (N_8293,N_6389,N_7490);
and U8294 (N_8294,N_7470,N_7411);
or U8295 (N_8295,N_6750,N_7236);
xnor U8296 (N_8296,N_7641,N_7438);
nand U8297 (N_8297,N_7166,N_6311);
nor U8298 (N_8298,N_6917,N_6505);
xor U8299 (N_8299,N_7158,N_6423);
nand U8300 (N_8300,N_7743,N_6220);
nor U8301 (N_8301,N_6305,N_7152);
xor U8302 (N_8302,N_6791,N_7408);
nor U8303 (N_8303,N_6045,N_7003);
nand U8304 (N_8304,N_7249,N_7266);
nand U8305 (N_8305,N_7720,N_7435);
nor U8306 (N_8306,N_6370,N_7983);
nand U8307 (N_8307,N_6060,N_6679);
or U8308 (N_8308,N_6986,N_7629);
nand U8309 (N_8309,N_6580,N_6552);
nand U8310 (N_8310,N_7998,N_6162);
nor U8311 (N_8311,N_6681,N_7907);
and U8312 (N_8312,N_6876,N_7147);
and U8313 (N_8313,N_6969,N_6109);
nand U8314 (N_8314,N_6898,N_6581);
nor U8315 (N_8315,N_6541,N_7735);
nand U8316 (N_8316,N_6556,N_7153);
xor U8317 (N_8317,N_7710,N_7208);
and U8318 (N_8318,N_6283,N_6087);
and U8319 (N_8319,N_6202,N_7693);
or U8320 (N_8320,N_6590,N_7872);
xor U8321 (N_8321,N_6997,N_7193);
xnor U8322 (N_8322,N_6440,N_6763);
nor U8323 (N_8323,N_6426,N_7362);
nor U8324 (N_8324,N_6393,N_6024);
and U8325 (N_8325,N_7453,N_6290);
and U8326 (N_8326,N_6981,N_7063);
nand U8327 (N_8327,N_6865,N_6407);
xnor U8328 (N_8328,N_7700,N_6047);
xnor U8329 (N_8329,N_7076,N_6766);
xor U8330 (N_8330,N_6951,N_7916);
nor U8331 (N_8331,N_6781,N_7023);
xor U8332 (N_8332,N_7125,N_7313);
or U8333 (N_8333,N_6712,N_6895);
nand U8334 (N_8334,N_7732,N_6201);
nand U8335 (N_8335,N_7356,N_7107);
nor U8336 (N_8336,N_6495,N_6452);
xnor U8337 (N_8337,N_7847,N_7761);
xor U8338 (N_8338,N_6054,N_7129);
and U8339 (N_8339,N_7182,N_6195);
nor U8340 (N_8340,N_7518,N_7064);
xnor U8341 (N_8341,N_7534,N_6064);
nand U8342 (N_8342,N_7268,N_6049);
and U8343 (N_8343,N_6250,N_6038);
xnor U8344 (N_8344,N_7683,N_6654);
and U8345 (N_8345,N_6348,N_7140);
and U8346 (N_8346,N_7339,N_6186);
xor U8347 (N_8347,N_6964,N_7298);
and U8348 (N_8348,N_7135,N_6417);
and U8349 (N_8349,N_6092,N_6853);
or U8350 (N_8350,N_6146,N_7358);
or U8351 (N_8351,N_7786,N_6741);
xnor U8352 (N_8352,N_7659,N_6544);
nor U8353 (N_8353,N_6209,N_7657);
nand U8354 (N_8354,N_7756,N_7599);
nand U8355 (N_8355,N_7194,N_6722);
nor U8356 (N_8356,N_6241,N_6144);
and U8357 (N_8357,N_6694,N_7648);
nor U8358 (N_8358,N_7687,N_6647);
nor U8359 (N_8359,N_7505,N_7060);
or U8360 (N_8360,N_6041,N_7818);
and U8361 (N_8361,N_6952,N_6342);
nand U8362 (N_8362,N_7283,N_6814);
and U8363 (N_8363,N_6788,N_6583);
nand U8364 (N_8364,N_6989,N_6772);
xnor U8365 (N_8365,N_6746,N_7443);
xor U8366 (N_8366,N_7582,N_6352);
nor U8367 (N_8367,N_6251,N_7608);
nand U8368 (N_8368,N_6413,N_6509);
nor U8369 (N_8369,N_7035,N_7825);
nor U8370 (N_8370,N_6866,N_7248);
and U8371 (N_8371,N_7372,N_7789);
or U8372 (N_8372,N_6935,N_7974);
nand U8373 (N_8373,N_6830,N_7111);
nor U8374 (N_8374,N_6187,N_7016);
xor U8375 (N_8375,N_6071,N_7090);
and U8376 (N_8376,N_6604,N_7202);
or U8377 (N_8377,N_7118,N_6688);
xnor U8378 (N_8378,N_7543,N_7072);
and U8379 (N_8379,N_7281,N_7681);
xnor U8380 (N_8380,N_6184,N_7897);
xnor U8381 (N_8381,N_7258,N_6657);
nand U8382 (N_8382,N_6526,N_7279);
nand U8383 (N_8383,N_7145,N_7854);
nor U8384 (N_8384,N_7535,N_6881);
nand U8385 (N_8385,N_6394,N_7046);
nor U8386 (N_8386,N_7665,N_7873);
xor U8387 (N_8387,N_7724,N_6923);
and U8388 (N_8388,N_7026,N_6420);
xor U8389 (N_8389,N_6485,N_7848);
and U8390 (N_8390,N_6543,N_7952);
and U8391 (N_8391,N_6546,N_7487);
nor U8392 (N_8392,N_7375,N_6760);
nand U8393 (N_8393,N_7540,N_6844);
nand U8394 (N_8394,N_7077,N_6970);
and U8395 (N_8395,N_7887,N_7293);
nor U8396 (N_8396,N_6178,N_7868);
nor U8397 (N_8397,N_7795,N_6194);
or U8398 (N_8398,N_6577,N_7146);
nand U8399 (N_8399,N_6333,N_7437);
nand U8400 (N_8400,N_7725,N_7619);
nor U8401 (N_8401,N_7674,N_7984);
and U8402 (N_8402,N_7071,N_7879);
xnor U8403 (N_8403,N_6135,N_7817);
xnor U8404 (N_8404,N_6988,N_6777);
nand U8405 (N_8405,N_7787,N_7880);
nor U8406 (N_8406,N_7277,N_6243);
nand U8407 (N_8407,N_7061,N_7488);
and U8408 (N_8408,N_7481,N_7931);
nor U8409 (N_8409,N_7078,N_7591);
and U8410 (N_8410,N_6662,N_7716);
or U8411 (N_8411,N_6142,N_6165);
and U8412 (N_8412,N_6409,N_7484);
or U8413 (N_8413,N_7169,N_6941);
xor U8414 (N_8414,N_6754,N_6125);
and U8415 (N_8415,N_7783,N_6504);
nor U8416 (N_8416,N_7877,N_7956);
xor U8417 (N_8417,N_6104,N_6749);
xnor U8418 (N_8418,N_6875,N_6942);
nand U8419 (N_8419,N_6331,N_6554);
nand U8420 (N_8420,N_6715,N_6637);
nand U8421 (N_8421,N_6310,N_7525);
xnor U8422 (N_8422,N_7594,N_6001);
and U8423 (N_8423,N_7669,N_7689);
or U8424 (N_8424,N_7549,N_6686);
nor U8425 (N_8425,N_7327,N_7643);
nand U8426 (N_8426,N_7870,N_6639);
xnor U8427 (N_8427,N_7727,N_7601);
or U8428 (N_8428,N_6097,N_6912);
or U8429 (N_8429,N_6672,N_7489);
xnor U8430 (N_8430,N_7871,N_6682);
and U8431 (N_8431,N_6524,N_6214);
nand U8432 (N_8432,N_6521,N_7894);
nand U8433 (N_8433,N_6810,N_7545);
nand U8434 (N_8434,N_7960,N_6783);
xor U8435 (N_8435,N_6010,N_6663);
or U8436 (N_8436,N_6558,N_6748);
nor U8437 (N_8437,N_6821,N_6878);
and U8438 (N_8438,N_6207,N_6566);
nand U8439 (N_8439,N_7826,N_7404);
or U8440 (N_8440,N_6157,N_6874);
and U8441 (N_8441,N_7513,N_6421);
and U8442 (N_8442,N_7425,N_6675);
nand U8443 (N_8443,N_6890,N_7333);
nand U8444 (N_8444,N_6636,N_7544);
nand U8445 (N_8445,N_7721,N_6326);
nor U8446 (N_8446,N_6169,N_7009);
nor U8447 (N_8447,N_6922,N_7033);
nand U8448 (N_8448,N_6475,N_6312);
nand U8449 (N_8449,N_7990,N_6227);
nand U8450 (N_8450,N_7864,N_7030);
xor U8451 (N_8451,N_7768,N_7331);
xnor U8452 (N_8452,N_6016,N_6380);
nand U8453 (N_8453,N_7739,N_6808);
and U8454 (N_8454,N_6924,N_6826);
nand U8455 (N_8455,N_7367,N_6738);
nand U8456 (N_8456,N_7320,N_7346);
nand U8457 (N_8457,N_6501,N_7348);
and U8458 (N_8458,N_7719,N_7740);
nor U8459 (N_8459,N_6376,N_7469);
or U8460 (N_8460,N_7412,N_6827);
nor U8461 (N_8461,N_6493,N_6152);
xnor U8462 (N_8462,N_6436,N_6320);
and U8463 (N_8463,N_6603,N_7836);
xnor U8464 (N_8464,N_6240,N_6998);
xor U8465 (N_8465,N_7475,N_6319);
and U8466 (N_8466,N_6687,N_7128);
nor U8467 (N_8467,N_6764,N_6962);
and U8468 (N_8468,N_7450,N_7855);
or U8469 (N_8469,N_6478,N_7045);
xnor U8470 (N_8470,N_6774,N_7148);
nor U8471 (N_8471,N_6840,N_6396);
nor U8472 (N_8472,N_6517,N_7628);
xor U8473 (N_8473,N_7199,N_7151);
nor U8474 (N_8474,N_7634,N_7114);
or U8475 (N_8475,N_6729,N_6231);
and U8476 (N_8476,N_6039,N_6930);
nand U8477 (N_8477,N_6287,N_6996);
nand U8478 (N_8478,N_6445,N_7519);
and U8479 (N_8479,N_7691,N_6938);
xnor U8480 (N_8480,N_7308,N_7638);
nor U8481 (N_8481,N_6584,N_7571);
nand U8482 (N_8482,N_6678,N_7459);
xor U8483 (N_8483,N_7668,N_7965);
nor U8484 (N_8484,N_7609,N_6792);
and U8485 (N_8485,N_6696,N_7559);
and U8486 (N_8486,N_7052,N_7216);
nor U8487 (N_8487,N_6921,N_7733);
xnor U8488 (N_8488,N_6782,N_7746);
nand U8489 (N_8489,N_6030,N_6500);
xor U8490 (N_8490,N_7149,N_6490);
nor U8491 (N_8491,N_7752,N_7605);
nand U8492 (N_8492,N_6368,N_6817);
or U8493 (N_8493,N_6837,N_7909);
nand U8494 (N_8494,N_7962,N_7342);
or U8495 (N_8495,N_7371,N_6780);
or U8496 (N_8496,N_6872,N_7340);
xor U8497 (N_8497,N_6978,N_7465);
nand U8498 (N_8498,N_6597,N_6236);
or U8499 (N_8499,N_6913,N_7705);
and U8500 (N_8500,N_7886,N_7123);
and U8501 (N_8501,N_7507,N_6386);
and U8502 (N_8502,N_7592,N_6789);
xnor U8503 (N_8503,N_7819,N_6889);
nor U8504 (N_8504,N_7706,N_6004);
and U8505 (N_8505,N_6138,N_6506);
xor U8506 (N_8506,N_7402,N_6400);
and U8507 (N_8507,N_7515,N_6624);
nor U8508 (N_8508,N_7210,N_6653);
xor U8509 (N_8509,N_6005,N_7059);
or U8510 (N_8510,N_6974,N_6946);
nor U8511 (N_8511,N_6651,N_7993);
or U8512 (N_8512,N_7797,N_7589);
xor U8513 (N_8513,N_6908,N_7247);
or U8514 (N_8514,N_6804,N_7432);
nor U8515 (N_8515,N_7666,N_6325);
nand U8516 (N_8516,N_6395,N_7307);
nand U8517 (N_8517,N_6416,N_7521);
nand U8518 (N_8518,N_7512,N_6083);
xnor U8519 (N_8519,N_6683,N_7558);
xor U8520 (N_8520,N_7058,N_6185);
nand U8521 (N_8521,N_7954,N_6300);
nand U8522 (N_8522,N_7656,N_6815);
and U8523 (N_8523,N_7911,N_6429);
nor U8524 (N_8524,N_6119,N_6136);
and U8525 (N_8525,N_6990,N_6247);
or U8526 (N_8526,N_7100,N_7966);
nor U8527 (N_8527,N_7718,N_6891);
nand U8528 (N_8528,N_7690,N_7287);
xor U8529 (N_8529,N_7844,N_6082);
or U8530 (N_8530,N_7043,N_7150);
xor U8531 (N_8531,N_6784,N_7579);
xor U8532 (N_8532,N_7378,N_6484);
nand U8533 (N_8533,N_7776,N_7280);
nand U8534 (N_8534,N_7211,N_6264);
nor U8535 (N_8535,N_6900,N_7572);
or U8536 (N_8536,N_6831,N_7711);
xnor U8537 (N_8537,N_6205,N_6513);
or U8538 (N_8538,N_6179,N_6279);
xnor U8539 (N_8539,N_6468,N_7472);
or U8540 (N_8540,N_7370,N_7495);
or U8541 (N_8541,N_6390,N_6502);
nand U8542 (N_8542,N_7321,N_6914);
xnor U8543 (N_8543,N_6931,N_6642);
nand U8544 (N_8544,N_7697,N_7625);
and U8545 (N_8545,N_6708,N_7022);
or U8546 (N_8546,N_7021,N_6607);
and U8547 (N_8547,N_7238,N_7037);
xnor U8548 (N_8548,N_6555,N_6572);
xor U8549 (N_8549,N_6477,N_6649);
xnor U8550 (N_8550,N_7336,N_7994);
or U8551 (N_8551,N_7093,N_7215);
nor U8552 (N_8552,N_6591,N_6491);
and U8553 (N_8553,N_6841,N_6055);
nor U8554 (N_8554,N_7137,N_6351);
nand U8555 (N_8555,N_6739,N_6174);
xor U8556 (N_8556,N_7812,N_6419);
and U8557 (N_8557,N_6592,N_7322);
nand U8558 (N_8558,N_6434,N_7203);
xor U8559 (N_8559,N_6628,N_7315);
or U8560 (N_8560,N_6391,N_7516);
and U8561 (N_8561,N_7671,N_6405);
nand U8562 (N_8562,N_7499,N_7241);
nor U8563 (N_8563,N_7460,N_7217);
nor U8564 (N_8564,N_7912,N_7244);
and U8565 (N_8565,N_7406,N_6599);
nor U8566 (N_8566,N_6328,N_6650);
nand U8567 (N_8567,N_6089,N_6259);
nor U8568 (N_8568,N_6255,N_6458);
and U8569 (N_8569,N_7273,N_6245);
or U8570 (N_8570,N_7444,N_6903);
and U8571 (N_8571,N_7302,N_6411);
or U8572 (N_8572,N_6734,N_6459);
and U8573 (N_8573,N_6758,N_7923);
xor U8574 (N_8574,N_6051,N_7084);
xor U8575 (N_8575,N_7893,N_6638);
or U8576 (N_8576,N_7049,N_6350);
nand U8577 (N_8577,N_7025,N_6803);
or U8578 (N_8578,N_6216,N_7784);
nor U8579 (N_8579,N_7373,N_6143);
and U8580 (N_8580,N_7833,N_7457);
nor U8581 (N_8581,N_6612,N_7214);
nand U8582 (N_8582,N_6378,N_7914);
xor U8583 (N_8583,N_6991,N_6757);
nand U8584 (N_8584,N_7688,N_6081);
and U8585 (N_8585,N_7504,N_7440);
xnor U8586 (N_8586,N_7278,N_7485);
or U8587 (N_8587,N_7162,N_6761);
or U8588 (N_8588,N_7039,N_7828);
or U8589 (N_8589,N_7959,N_7712);
and U8590 (N_8590,N_6752,N_7068);
xor U8591 (N_8591,N_7522,N_6210);
nor U8592 (N_8592,N_6838,N_7334);
or U8593 (N_8593,N_7800,N_6542);
xor U8594 (N_8594,N_6685,N_7456);
nor U8595 (N_8595,N_6147,N_6822);
nand U8596 (N_8596,N_7588,N_7701);
nor U8597 (N_8597,N_6117,N_6860);
and U8598 (N_8598,N_6882,N_6658);
nor U8599 (N_8599,N_7631,N_6730);
and U8600 (N_8600,N_6197,N_7881);
nand U8601 (N_8601,N_6026,N_7463);
xnor U8602 (N_8602,N_7264,N_7500);
and U8603 (N_8603,N_7611,N_7910);
nand U8604 (N_8604,N_7127,N_7865);
or U8605 (N_8605,N_7286,N_7434);
xor U8606 (N_8606,N_6013,N_6242);
nand U8607 (N_8607,N_6633,N_6422);
nor U8608 (N_8608,N_7483,N_6183);
and U8609 (N_8609,N_7350,N_7187);
nor U8610 (N_8610,N_7290,N_6744);
and U8611 (N_8611,N_7695,N_7943);
xor U8612 (N_8612,N_7180,N_6809);
nand U8613 (N_8613,N_7653,N_6188);
nor U8614 (N_8614,N_7032,N_7070);
xnor U8615 (N_8615,N_6481,N_7257);
nor U8616 (N_8616,N_7161,N_6438);
or U8617 (N_8617,N_6387,N_7388);
xor U8618 (N_8618,N_7120,N_7992);
or U8619 (N_8619,N_7708,N_6273);
and U8620 (N_8620,N_7730,N_6551);
nand U8621 (N_8621,N_7159,N_7341);
or U8622 (N_8622,N_6745,N_6805);
nor U8623 (N_8623,N_6790,N_6238);
nor U8624 (N_8624,N_7317,N_6358);
or U8625 (N_8625,N_7329,N_7414);
and U8626 (N_8626,N_6656,N_6586);
nor U8627 (N_8627,N_6534,N_6798);
or U8628 (N_8628,N_7042,N_7860);
xor U8629 (N_8629,N_7731,N_7884);
and U8630 (N_8630,N_7929,N_6870);
nand U8631 (N_8631,N_7802,N_6713);
or U8632 (N_8632,N_7017,N_6992);
and U8633 (N_8633,N_7452,N_7206);
nand U8634 (N_8634,N_7996,N_6025);
xnor U8635 (N_8635,N_7062,N_6863);
and U8636 (N_8636,N_7269,N_7647);
nor U8637 (N_8637,N_6779,N_7651);
xnor U8638 (N_8638,N_6292,N_6040);
nor U8639 (N_8639,N_7757,N_7237);
or U8640 (N_8640,N_6910,N_7726);
or U8641 (N_8641,N_7108,N_7577);
or U8642 (N_8642,N_7102,N_7305);
and U8643 (N_8643,N_7771,N_6871);
and U8644 (N_8644,N_7640,N_6557);
nand U8645 (N_8645,N_6710,N_6052);
and U8646 (N_8646,N_7121,N_7704);
nand U8647 (N_8647,N_6072,N_6228);
nand U8648 (N_8648,N_7748,N_7918);
xnor U8649 (N_8649,N_6671,N_7777);
xor U8650 (N_8650,N_7270,N_7574);
nor U8651 (N_8651,N_7036,N_6160);
xor U8652 (N_8652,N_7709,N_7005);
or U8653 (N_8653,N_7520,N_6553);
nand U8654 (N_8654,N_7309,N_6448);
xor U8655 (N_8655,N_7429,N_7995);
xnor U8656 (N_8656,N_6096,N_6940);
and U8657 (N_8657,N_6641,N_7703);
nand U8658 (N_8658,N_6816,N_7664);
and U8659 (N_8659,N_6080,N_7514);
or U8660 (N_8660,N_6861,N_6833);
and U8661 (N_8661,N_6676,N_6595);
and U8662 (N_8662,N_6717,N_6593);
nand U8663 (N_8663,N_6141,N_6067);
nor U8664 (N_8664,N_7755,N_6635);
nor U8665 (N_8665,N_6233,N_7343);
nand U8666 (N_8666,N_7945,N_7832);
xnor U8667 (N_8667,N_7928,N_7239);
xnor U8668 (N_8668,N_7799,N_6953);
or U8669 (N_8669,N_7207,N_7288);
or U8670 (N_8670,N_7502,N_7165);
nand U8671 (N_8671,N_6601,N_7575);
nand U8672 (N_8672,N_7715,N_7410);
nor U8673 (N_8673,N_6253,N_7415);
nand U8674 (N_8674,N_6099,N_7616);
nand U8675 (N_8675,N_7134,N_6454);
or U8676 (N_8676,N_7526,N_6965);
and U8677 (N_8677,N_6503,N_7660);
nand U8678 (N_8678,N_7477,N_6538);
nand U8679 (N_8679,N_7620,N_6893);
and U8680 (N_8680,N_6340,N_6644);
xnor U8681 (N_8681,N_7110,N_7937);
xor U8682 (N_8682,N_7946,N_7235);
xnor U8683 (N_8683,N_6430,N_7421);
or U8684 (N_8684,N_7355,N_6512);
xnor U8685 (N_8685,N_7117,N_7436);
xnor U8686 (N_8686,N_7175,N_6027);
nand U8687 (N_8687,N_6769,N_7976);
nand U8688 (N_8688,N_7949,N_6873);
or U8689 (N_8689,N_6937,N_7242);
and U8690 (N_8690,N_7736,N_7418);
nor U8691 (N_8691,N_7555,N_6224);
nor U8692 (N_8692,N_6869,N_7400);
and U8693 (N_8693,N_6435,N_6614);
and U8694 (N_8694,N_6304,N_6431);
xor U8695 (N_8695,N_7221,N_7220);
and U8696 (N_8696,N_6314,N_7626);
or U8697 (N_8697,N_7295,N_7888);
xnor U8698 (N_8698,N_6066,N_7262);
or U8699 (N_8699,N_6018,N_7261);
xor U8700 (N_8700,N_7510,N_7007);
nand U8701 (N_8701,N_6134,N_7136);
xnor U8702 (N_8702,N_6618,N_7383);
or U8703 (N_8703,N_6356,N_6961);
xor U8704 (N_8704,N_6539,N_6530);
xor U8705 (N_8705,N_6508,N_6313);
or U8706 (N_8706,N_7846,N_6424);
and U8707 (N_8707,N_7431,N_6973);
nand U8708 (N_8708,N_7096,N_6677);
nand U8709 (N_8709,N_7679,N_7245);
or U8710 (N_8710,N_6404,N_7551);
xnor U8711 (N_8711,N_7379,N_6470);
nor U8712 (N_8712,N_6315,N_6625);
and U8713 (N_8713,N_7524,N_6130);
or U8714 (N_8714,N_6828,N_6303);
and U8715 (N_8715,N_7442,N_6995);
and U8716 (N_8716,N_6496,N_6043);
nor U8717 (N_8717,N_7479,N_7174);
xnor U8718 (N_8718,N_7233,N_6324);
nand U8719 (N_8719,N_7380,N_6295);
or U8720 (N_8720,N_7806,N_7920);
nor U8721 (N_8721,N_7675,N_7417);
and U8722 (N_8722,N_6732,N_7567);
xnor U8723 (N_8723,N_7066,N_6933);
nor U8724 (N_8724,N_7623,N_6093);
and U8725 (N_8725,N_6812,N_6102);
nor U8726 (N_8726,N_7176,N_6449);
xnor U8727 (N_8727,N_7384,N_6173);
and U8728 (N_8728,N_6762,N_7810);
nand U8729 (N_8729,N_6406,N_7560);
and U8730 (N_8730,N_6883,N_7098);
xor U8731 (N_8731,N_7607,N_7201);
or U8732 (N_8732,N_7423,N_6223);
and U8733 (N_8733,N_6945,N_7550);
xor U8734 (N_8734,N_6058,N_7517);
nand U8735 (N_8735,N_7852,N_7289);
or U8736 (N_8736,N_6697,N_7967);
nand U8737 (N_8737,N_7328,N_7274);
xor U8738 (N_8738,N_7386,N_6703);
and U8739 (N_8739,N_7876,N_7310);
or U8740 (N_8740,N_7554,N_6699);
xnor U8741 (N_8741,N_7255,N_7734);
nor U8742 (N_8742,N_7814,N_6293);
nor U8743 (N_8743,N_6892,N_7361);
or U8744 (N_8744,N_6164,N_6587);
or U8745 (N_8745,N_6225,N_6576);
xnor U8746 (N_8746,N_6646,N_7405);
or U8747 (N_8747,N_6615,N_7225);
nand U8748 (N_8748,N_7163,N_6100);
nor U8749 (N_8749,N_6999,N_7940);
nand U8750 (N_8750,N_7861,N_7927);
xor U8751 (N_8751,N_6073,N_6514);
or U8752 (N_8752,N_7737,N_7862);
and U8753 (N_8753,N_7741,N_7272);
or U8754 (N_8754,N_7822,N_7446);
nor U8755 (N_8755,N_6632,N_7325);
xnor U8756 (N_8756,N_6200,N_6170);
or U8757 (N_8757,N_6098,N_6215);
nor U8758 (N_8758,N_6339,N_7772);
xnor U8759 (N_8759,N_7988,N_7941);
or U8760 (N_8760,N_7957,N_6442);
xnor U8761 (N_8761,N_7958,N_7420);
or U8762 (N_8762,N_6472,N_6479);
nor U8763 (N_8763,N_6208,N_7476);
or U8764 (N_8764,N_6905,N_6751);
and U8765 (N_8765,N_6849,N_7115);
and U8766 (N_8766,N_7859,N_6456);
nand U8767 (N_8767,N_6523,N_6181);
or U8768 (N_8768,N_6237,N_7533);
and U8769 (N_8769,N_7823,N_6720);
nand U8770 (N_8770,N_7501,N_6680);
nor U8771 (N_8771,N_6621,N_6605);
xnor U8772 (N_8772,N_6285,N_6327);
xnor U8773 (N_8773,N_7011,N_7809);
nor U8774 (N_8774,N_6901,N_6034);
or U8775 (N_8775,N_7654,N_7590);
or U8776 (N_8776,N_7508,N_7074);
xor U8777 (N_8777,N_6020,N_6888);
and U8778 (N_8778,N_7686,N_6163);
xor U8779 (N_8779,N_7297,N_7124);
and U8780 (N_8780,N_6966,N_6114);
xor U8781 (N_8781,N_6127,N_7015);
nand U8782 (N_8782,N_6522,N_7922);
xnor U8783 (N_8783,N_6294,N_6381);
or U8784 (N_8784,N_7613,N_7267);
nand U8785 (N_8785,N_7186,N_7276);
or U8786 (N_8786,N_7858,N_7838);
xor U8787 (N_8787,N_7874,N_6499);
xor U8788 (N_8788,N_6464,N_7722);
nand U8789 (N_8789,N_7316,N_7794);
xor U8790 (N_8790,N_6050,N_6256);
nand U8791 (N_8791,N_7955,N_7048);
or U8792 (N_8792,N_6203,N_6747);
nand U8793 (N_8793,N_7793,N_6122);
xnor U8794 (N_8794,N_7088,N_6610);
and U8795 (N_8795,N_6375,N_6009);
or U8796 (N_8796,N_7991,N_7969);
nor U8797 (N_8797,N_7204,N_7593);
xor U8798 (N_8798,N_6820,N_7938);
nor U8799 (N_8799,N_6926,N_7805);
and U8800 (N_8800,N_6469,N_7008);
and U8801 (N_8801,N_6346,N_6343);
nand U8802 (N_8802,N_6652,N_6802);
xor U8803 (N_8803,N_7296,N_6113);
and U8804 (N_8804,N_7461,N_6648);
xnor U8805 (N_8805,N_7792,N_6528);
or U8806 (N_8806,N_6239,N_6807);
nand U8807 (N_8807,N_7662,N_7655);
nand U8808 (N_8808,N_6731,N_7083);
nand U8809 (N_8809,N_6880,N_7950);
nor U8810 (N_8810,N_6103,N_6856);
nand U8811 (N_8811,N_7930,N_6536);
or U8812 (N_8812,N_7503,N_7839);
xor U8813 (N_8813,N_6002,N_6359);
or U8814 (N_8814,N_6851,N_6511);
xnor U8815 (N_8815,N_7750,N_7633);
nor U8816 (N_8816,N_6260,N_6084);
nand U8817 (N_8817,N_7395,N_6771);
xor U8818 (N_8818,N_6361,N_6309);
and U8819 (N_8819,N_7692,N_7857);
and U8820 (N_8820,N_6131,N_6302);
nand U8821 (N_8821,N_7584,N_7213);
or U8822 (N_8822,N_7536,N_6793);
xnor U8823 (N_8823,N_6140,N_7294);
or U8824 (N_8824,N_6846,N_6028);
xnor U8825 (N_8825,N_7948,N_6349);
and U8826 (N_8826,N_6702,N_6532);
or U8827 (N_8827,N_6733,N_6364);
nor U8828 (N_8828,N_7552,N_6126);
or U8829 (N_8829,N_6718,N_6575);
and U8830 (N_8830,N_7097,N_7903);
xnor U8831 (N_8831,N_7924,N_7353);
or U8832 (N_8832,N_6056,N_7778);
xnor U8833 (N_8833,N_6111,N_7029);
and U8834 (N_8834,N_6057,N_6410);
xnor U8835 (N_8835,N_6626,N_6301);
nand U8836 (N_8836,N_7319,N_7001);
and U8837 (N_8837,N_7079,N_7758);
and U8838 (N_8838,N_7374,N_6868);
nor U8839 (N_8839,N_7112,N_6824);
or U8840 (N_8840,N_6643,N_7177);
nand U8841 (N_8841,N_7243,N_6979);
xnor U8842 (N_8842,N_6725,N_7170);
and U8843 (N_8843,N_7840,N_6611);
xnor U8844 (N_8844,N_7229,N_6877);
nor U8845 (N_8845,N_7980,N_6529);
xor U8846 (N_8846,N_6021,N_7222);
xnor U8847 (N_8847,N_6488,N_7678);
or U8848 (N_8848,N_6336,N_7300);
xor U8849 (N_8849,N_6015,N_6267);
xnor U8850 (N_8850,N_6124,N_7396);
or U8851 (N_8851,N_7979,N_7908);
or U8852 (N_8852,N_6159,N_6756);
nand U8853 (N_8853,N_6489,N_6033);
or U8854 (N_8854,N_7898,N_7939);
nand U8855 (N_8855,N_6573,N_6191);
nor U8856 (N_8856,N_7116,N_6571);
or U8857 (N_8857,N_6372,N_6659);
nor U8858 (N_8858,N_6660,N_7729);
nor U8859 (N_8859,N_6811,N_7200);
nand U8860 (N_8860,N_7612,N_7357);
and U8861 (N_8861,N_7393,N_7338);
and U8862 (N_8862,N_7904,N_6425);
nor U8863 (N_8863,N_6967,N_6602);
and U8864 (N_8864,N_7511,N_7028);
xnor U8865 (N_8865,N_6281,N_7933);
or U8866 (N_8866,N_6956,N_6403);
or U8867 (N_8867,N_7808,N_7179);
or U8868 (N_8868,N_6916,N_7427);
or U8869 (N_8869,N_6332,N_6384);
nor U8870 (N_8870,N_6537,N_7742);
xor U8871 (N_8871,N_6132,N_7439);
xor U8872 (N_8872,N_6108,N_6929);
nor U8873 (N_8873,N_7670,N_7047);
or U8874 (N_8874,N_7875,N_7563);
xor U8875 (N_8875,N_6854,N_7541);
and U8876 (N_8876,N_6022,N_7389);
and U8877 (N_8877,N_7915,N_6907);
nand U8878 (N_8878,N_7188,N_7369);
or U8879 (N_8879,N_7306,N_6954);
and U8880 (N_8880,N_6399,N_6219);
or U8881 (N_8881,N_6330,N_6161);
and U8882 (N_8882,N_7764,N_6726);
nor U8883 (N_8883,N_6565,N_6579);
nand U8884 (N_8884,N_6282,N_7568);
nor U8885 (N_8885,N_7842,N_7252);
xnor U8886 (N_8886,N_6397,N_7344);
nand U8887 (N_8887,N_7667,N_6167);
nor U8888 (N_8888,N_6014,N_6392);
and U8889 (N_8889,N_6943,N_6232);
nand U8890 (N_8890,N_6564,N_6507);
nor U8891 (N_8891,N_7013,N_6594);
and U8892 (N_8892,N_7539,N_6899);
xor U8893 (N_8893,N_7335,N_6864);
or U8894 (N_8894,N_7597,N_7181);
nand U8895 (N_8895,N_7080,N_6920);
and U8896 (N_8896,N_7095,N_7138);
nor U8897 (N_8897,N_6709,N_7448);
and U8898 (N_8898,N_7260,N_7973);
xnor U8899 (N_8899,N_7989,N_6385);
nor U8900 (N_8900,N_7157,N_6280);
and U8901 (N_8901,N_6263,N_7542);
or U8902 (N_8902,N_6299,N_6563);
nor U8903 (N_8903,N_7906,N_7399);
xor U8904 (N_8904,N_6078,N_6068);
or U8905 (N_8905,N_6735,N_7970);
or U8906 (N_8906,N_7256,N_6317);
nor U8907 (N_8907,N_6985,N_6095);
nand U8908 (N_8908,N_6690,N_7569);
xnor U8909 (N_8909,N_7087,N_7126);
or U8910 (N_8910,N_7913,N_7790);
nor U8911 (N_8911,N_6120,N_7863);
nor U8912 (N_8912,N_7101,N_7234);
or U8913 (N_8913,N_6902,N_6982);
nand U8914 (N_8914,N_7754,N_6450);
or U8915 (N_8915,N_6825,N_7586);
nand U8916 (N_8916,N_6042,N_7699);
or U8917 (N_8917,N_7762,N_6896);
or U8918 (N_8918,N_7867,N_7051);
and U8919 (N_8919,N_7433,N_7154);
nand U8920 (N_8920,N_7677,N_7498);
xnor U8921 (N_8921,N_7391,N_6548);
nand U8922 (N_8922,N_7639,N_7031);
nand U8923 (N_8923,N_6261,N_6832);
nor U8924 (N_8924,N_7332,N_6531);
nor U8925 (N_8925,N_7624,N_6366);
and U8926 (N_8926,N_7190,N_6337);
and U8927 (N_8927,N_6987,N_6755);
nand U8928 (N_8928,N_6414,N_7663);
nor U8929 (N_8929,N_6492,N_7231);
or U8930 (N_8930,N_7197,N_7603);
and U8931 (N_8931,N_6465,N_7621);
or U8932 (N_8932,N_7895,N_6432);
nor U8933 (N_8933,N_6634,N_6296);
or U8934 (N_8934,N_6560,N_7807);
nor U8935 (N_8935,N_6823,N_6007);
and U8936 (N_8936,N_6609,N_7547);
and U8937 (N_8937,N_7900,N_7982);
xnor U8938 (N_8938,N_6932,N_7963);
and U8939 (N_8939,N_6549,N_6819);
or U8940 (N_8940,N_7155,N_7557);
and U8941 (N_8941,N_6806,N_6936);
xnor U8942 (N_8942,N_6483,N_7069);
and U8943 (N_8943,N_7936,N_7837);
nand U8944 (N_8944,N_6053,N_6116);
nor U8945 (N_8945,N_6234,N_7246);
nor U8946 (N_8946,N_7143,N_6306);
xor U8947 (N_8947,N_6217,N_6110);
and U8948 (N_8948,N_6154,N_7376);
nand U8949 (N_8949,N_6377,N_7587);
nand U8950 (N_8950,N_6252,N_7493);
nor U8951 (N_8951,N_7617,N_6446);
xnor U8952 (N_8952,N_7365,N_6467);
xor U8953 (N_8953,N_6035,N_7636);
nor U8954 (N_8954,N_6786,N_6329);
or U8955 (N_8955,N_7845,N_6665);
and U8956 (N_8956,N_6980,N_7546);
or U8957 (N_8957,N_6630,N_6655);
xor U8958 (N_8958,N_7506,N_6460);
nor U8959 (N_8959,N_7312,N_7054);
and U8960 (N_8960,N_6383,N_6670);
nand U8961 (N_8961,N_6257,N_6412);
nor U8962 (N_8962,N_6627,N_6727);
nor U8963 (N_8963,N_7397,N_6569);
and U8964 (N_8964,N_7685,N_6218);
nor U8965 (N_8965,N_6211,N_7760);
xnor U8966 (N_8966,N_6284,N_6879);
nor U8967 (N_8967,N_6023,N_6909);
nand U8968 (N_8968,N_7892,N_6107);
nand U8969 (N_8969,N_7972,N_7978);
or U8970 (N_8970,N_7896,N_7553);
nand U8971 (N_8971,N_6149,N_6063);
xnor U8972 (N_8972,N_7747,N_6623);
xnor U8973 (N_8973,N_6775,N_6939);
nor U8974 (N_8974,N_7284,N_7496);
xnor U8975 (N_8975,N_6172,N_6525);
and U8976 (N_8976,N_6944,N_6062);
and U8977 (N_8977,N_6608,N_6959);
and U8978 (N_8978,N_7610,N_6753);
nor U8979 (N_8979,N_7672,N_6742);
and U8980 (N_8980,N_7056,N_6000);
nor U8981 (N_8981,N_7347,N_6482);
xnor U8982 (N_8982,N_7523,N_7168);
xnor U8983 (N_8983,N_6032,N_6994);
or U8984 (N_8984,N_6829,N_6574);
and U8985 (N_8985,N_7441,N_6447);
and U8986 (N_8986,N_6275,N_6418);
xnor U8987 (N_8987,N_6427,N_7265);
nor U8988 (N_8988,N_6540,N_6156);
and U8989 (N_8989,N_6274,N_6036);
and U8990 (N_8990,N_6262,N_6347);
and U8991 (N_8991,N_7271,N_6398);
nand U8992 (N_8992,N_6148,N_6640);
nor U8993 (N_8993,N_6070,N_6759);
or U8994 (N_8994,N_6778,N_6773);
or U8995 (N_8995,N_6088,N_7766);
nand U8996 (N_8996,N_6017,N_7004);
nand U8997 (N_8997,N_6137,N_6268);
and U8998 (N_8998,N_6545,N_6355);
xnor U8999 (N_8999,N_6669,N_7130);
nand U9000 (N_9000,N_7042,N_7111);
and U9001 (N_9001,N_7822,N_6048);
and U9002 (N_9002,N_7152,N_7067);
and U9003 (N_9003,N_7880,N_7703);
or U9004 (N_9004,N_7648,N_7920);
xnor U9005 (N_9005,N_7621,N_6142);
nand U9006 (N_9006,N_7701,N_7555);
and U9007 (N_9007,N_7514,N_7477);
nand U9008 (N_9008,N_7407,N_6247);
nand U9009 (N_9009,N_7101,N_7629);
nand U9010 (N_9010,N_6743,N_6207);
or U9011 (N_9011,N_6082,N_6145);
xnor U9012 (N_9012,N_7781,N_7212);
or U9013 (N_9013,N_6706,N_7291);
nor U9014 (N_9014,N_7264,N_6777);
and U9015 (N_9015,N_7737,N_6917);
nor U9016 (N_9016,N_7432,N_6681);
xnor U9017 (N_9017,N_6398,N_7792);
nor U9018 (N_9018,N_7780,N_7398);
nor U9019 (N_9019,N_6361,N_7139);
xnor U9020 (N_9020,N_7447,N_7833);
nor U9021 (N_9021,N_6040,N_7742);
xnor U9022 (N_9022,N_7830,N_6138);
xnor U9023 (N_9023,N_7812,N_6230);
or U9024 (N_9024,N_7503,N_7389);
or U9025 (N_9025,N_7947,N_7749);
or U9026 (N_9026,N_6510,N_7789);
or U9027 (N_9027,N_7361,N_7813);
or U9028 (N_9028,N_6113,N_7245);
or U9029 (N_9029,N_7987,N_7202);
nand U9030 (N_9030,N_6223,N_7975);
xor U9031 (N_9031,N_6228,N_7018);
nor U9032 (N_9032,N_7221,N_6931);
nor U9033 (N_9033,N_7517,N_6374);
xor U9034 (N_9034,N_6503,N_7359);
or U9035 (N_9035,N_6331,N_7609);
or U9036 (N_9036,N_7038,N_6722);
nor U9037 (N_9037,N_7750,N_6486);
or U9038 (N_9038,N_6717,N_6896);
and U9039 (N_9039,N_7919,N_6791);
nand U9040 (N_9040,N_7656,N_7392);
nand U9041 (N_9041,N_6661,N_7967);
xnor U9042 (N_9042,N_6220,N_6888);
and U9043 (N_9043,N_6224,N_7493);
xor U9044 (N_9044,N_6513,N_6245);
xnor U9045 (N_9045,N_6143,N_6658);
nor U9046 (N_9046,N_6476,N_6709);
and U9047 (N_9047,N_7749,N_7193);
nor U9048 (N_9048,N_7086,N_7558);
and U9049 (N_9049,N_7414,N_7238);
and U9050 (N_9050,N_6707,N_6340);
nand U9051 (N_9051,N_6148,N_6417);
or U9052 (N_9052,N_6585,N_7857);
xnor U9053 (N_9053,N_7588,N_7771);
or U9054 (N_9054,N_7786,N_7056);
and U9055 (N_9055,N_6624,N_6407);
and U9056 (N_9056,N_6646,N_6420);
nand U9057 (N_9057,N_7164,N_6355);
xnor U9058 (N_9058,N_6810,N_6349);
xor U9059 (N_9059,N_6921,N_7947);
xor U9060 (N_9060,N_7060,N_7278);
nor U9061 (N_9061,N_7994,N_7825);
nor U9062 (N_9062,N_6743,N_6062);
and U9063 (N_9063,N_7650,N_7245);
nand U9064 (N_9064,N_7136,N_7995);
nand U9065 (N_9065,N_7099,N_7785);
xor U9066 (N_9066,N_7580,N_6556);
nor U9067 (N_9067,N_7037,N_7772);
nand U9068 (N_9068,N_6469,N_7455);
nor U9069 (N_9069,N_7242,N_7406);
and U9070 (N_9070,N_7032,N_7942);
and U9071 (N_9071,N_6396,N_6665);
nor U9072 (N_9072,N_7428,N_6087);
nand U9073 (N_9073,N_6897,N_7866);
and U9074 (N_9074,N_6588,N_6552);
nor U9075 (N_9075,N_7834,N_7773);
nor U9076 (N_9076,N_6345,N_6428);
nor U9077 (N_9077,N_6199,N_6968);
or U9078 (N_9078,N_6613,N_6383);
xor U9079 (N_9079,N_6661,N_7130);
xor U9080 (N_9080,N_6203,N_6869);
and U9081 (N_9081,N_7053,N_6650);
and U9082 (N_9082,N_7533,N_7333);
nand U9083 (N_9083,N_7092,N_6985);
or U9084 (N_9084,N_6077,N_6167);
and U9085 (N_9085,N_6277,N_7259);
nand U9086 (N_9086,N_7122,N_6344);
nand U9087 (N_9087,N_7396,N_7996);
or U9088 (N_9088,N_7802,N_7403);
nor U9089 (N_9089,N_6253,N_6165);
nor U9090 (N_9090,N_7439,N_7938);
or U9091 (N_9091,N_7630,N_6850);
nand U9092 (N_9092,N_6123,N_7850);
and U9093 (N_9093,N_7493,N_7115);
or U9094 (N_9094,N_7830,N_6699);
nor U9095 (N_9095,N_6587,N_6053);
nor U9096 (N_9096,N_6399,N_7626);
nand U9097 (N_9097,N_7675,N_7370);
xnor U9098 (N_9098,N_6762,N_7473);
xnor U9099 (N_9099,N_7580,N_6897);
and U9100 (N_9100,N_7502,N_7114);
xor U9101 (N_9101,N_6435,N_6622);
and U9102 (N_9102,N_6396,N_6205);
xor U9103 (N_9103,N_6455,N_6700);
and U9104 (N_9104,N_7178,N_7408);
xnor U9105 (N_9105,N_6246,N_6481);
nand U9106 (N_9106,N_6488,N_6883);
nand U9107 (N_9107,N_7013,N_6259);
xnor U9108 (N_9108,N_6415,N_7107);
or U9109 (N_9109,N_6944,N_7297);
or U9110 (N_9110,N_6443,N_7645);
and U9111 (N_9111,N_7469,N_7238);
and U9112 (N_9112,N_7374,N_6092);
nor U9113 (N_9113,N_6871,N_6751);
nor U9114 (N_9114,N_7873,N_7566);
nor U9115 (N_9115,N_7840,N_6570);
nand U9116 (N_9116,N_7840,N_6973);
or U9117 (N_9117,N_7339,N_6051);
or U9118 (N_9118,N_6789,N_6464);
and U9119 (N_9119,N_7016,N_6113);
xnor U9120 (N_9120,N_6686,N_7816);
or U9121 (N_9121,N_7401,N_6183);
or U9122 (N_9122,N_7068,N_7803);
or U9123 (N_9123,N_6059,N_6639);
or U9124 (N_9124,N_6865,N_6168);
xnor U9125 (N_9125,N_6093,N_6583);
xor U9126 (N_9126,N_7191,N_7080);
or U9127 (N_9127,N_6765,N_6954);
nor U9128 (N_9128,N_7565,N_7161);
nor U9129 (N_9129,N_7889,N_6974);
and U9130 (N_9130,N_6933,N_6682);
nor U9131 (N_9131,N_6987,N_6973);
nor U9132 (N_9132,N_7151,N_6185);
or U9133 (N_9133,N_6717,N_6575);
nor U9134 (N_9134,N_7170,N_6047);
xor U9135 (N_9135,N_6249,N_6845);
or U9136 (N_9136,N_7892,N_6125);
and U9137 (N_9137,N_7141,N_6081);
and U9138 (N_9138,N_7027,N_6501);
nor U9139 (N_9139,N_6473,N_6699);
nor U9140 (N_9140,N_6098,N_7273);
nand U9141 (N_9141,N_7317,N_6014);
and U9142 (N_9142,N_7789,N_7617);
xor U9143 (N_9143,N_7822,N_6470);
nor U9144 (N_9144,N_7651,N_6458);
or U9145 (N_9145,N_7094,N_7609);
nor U9146 (N_9146,N_6246,N_6873);
nor U9147 (N_9147,N_7363,N_6143);
xnor U9148 (N_9148,N_7058,N_6768);
or U9149 (N_9149,N_6744,N_6677);
xor U9150 (N_9150,N_7916,N_7710);
nor U9151 (N_9151,N_7755,N_6202);
nand U9152 (N_9152,N_7439,N_6693);
and U9153 (N_9153,N_7851,N_7095);
xnor U9154 (N_9154,N_7667,N_7777);
nor U9155 (N_9155,N_7277,N_7008);
or U9156 (N_9156,N_7574,N_7692);
nand U9157 (N_9157,N_6688,N_6623);
xor U9158 (N_9158,N_6135,N_6685);
or U9159 (N_9159,N_6216,N_6549);
nand U9160 (N_9160,N_7261,N_7890);
nand U9161 (N_9161,N_7615,N_6158);
nand U9162 (N_9162,N_7288,N_7429);
and U9163 (N_9163,N_7585,N_6234);
nor U9164 (N_9164,N_6602,N_7460);
xnor U9165 (N_9165,N_6433,N_6098);
nand U9166 (N_9166,N_7672,N_7819);
nor U9167 (N_9167,N_6401,N_7557);
nor U9168 (N_9168,N_7066,N_6173);
xnor U9169 (N_9169,N_7962,N_6039);
xnor U9170 (N_9170,N_7604,N_6342);
or U9171 (N_9171,N_7862,N_7519);
or U9172 (N_9172,N_6576,N_6398);
nor U9173 (N_9173,N_6325,N_6647);
nand U9174 (N_9174,N_7333,N_6865);
nand U9175 (N_9175,N_7647,N_7922);
and U9176 (N_9176,N_6578,N_7631);
nand U9177 (N_9177,N_7666,N_6349);
nand U9178 (N_9178,N_6409,N_6010);
nor U9179 (N_9179,N_6865,N_6874);
xor U9180 (N_9180,N_6380,N_6461);
and U9181 (N_9181,N_6223,N_6334);
xor U9182 (N_9182,N_6866,N_7479);
and U9183 (N_9183,N_6062,N_7881);
nand U9184 (N_9184,N_7484,N_7608);
nor U9185 (N_9185,N_7445,N_6415);
xnor U9186 (N_9186,N_6849,N_7366);
nand U9187 (N_9187,N_6701,N_6164);
xor U9188 (N_9188,N_7216,N_7915);
nand U9189 (N_9189,N_7938,N_6427);
and U9190 (N_9190,N_6061,N_6513);
nand U9191 (N_9191,N_6627,N_6120);
nand U9192 (N_9192,N_7554,N_7970);
nand U9193 (N_9193,N_6662,N_6709);
nand U9194 (N_9194,N_6583,N_6416);
nand U9195 (N_9195,N_7943,N_7487);
nor U9196 (N_9196,N_7589,N_7366);
nand U9197 (N_9197,N_7007,N_6602);
and U9198 (N_9198,N_6428,N_7690);
xor U9199 (N_9199,N_6265,N_6984);
and U9200 (N_9200,N_7089,N_7668);
nand U9201 (N_9201,N_7031,N_6019);
nand U9202 (N_9202,N_7127,N_6357);
or U9203 (N_9203,N_7370,N_7803);
nor U9204 (N_9204,N_7001,N_7844);
or U9205 (N_9205,N_7842,N_6295);
and U9206 (N_9206,N_6390,N_6839);
or U9207 (N_9207,N_6232,N_6419);
xnor U9208 (N_9208,N_6691,N_7428);
nand U9209 (N_9209,N_6428,N_6494);
and U9210 (N_9210,N_7967,N_6852);
nor U9211 (N_9211,N_7140,N_7696);
or U9212 (N_9212,N_7506,N_6980);
and U9213 (N_9213,N_6803,N_7408);
or U9214 (N_9214,N_6756,N_6713);
nor U9215 (N_9215,N_6623,N_6736);
xor U9216 (N_9216,N_7840,N_6635);
nor U9217 (N_9217,N_6680,N_7911);
or U9218 (N_9218,N_6998,N_7670);
and U9219 (N_9219,N_7984,N_7358);
xor U9220 (N_9220,N_7645,N_6180);
xnor U9221 (N_9221,N_6653,N_7162);
nand U9222 (N_9222,N_7162,N_6380);
nor U9223 (N_9223,N_7695,N_7818);
nor U9224 (N_9224,N_6293,N_7775);
and U9225 (N_9225,N_7654,N_6355);
and U9226 (N_9226,N_6886,N_7252);
nand U9227 (N_9227,N_6220,N_7826);
xnor U9228 (N_9228,N_6475,N_6101);
and U9229 (N_9229,N_6671,N_7497);
nand U9230 (N_9230,N_6527,N_7706);
and U9231 (N_9231,N_7061,N_7759);
nand U9232 (N_9232,N_7007,N_7430);
xor U9233 (N_9233,N_6188,N_6460);
and U9234 (N_9234,N_6866,N_6730);
or U9235 (N_9235,N_7019,N_6024);
nand U9236 (N_9236,N_7819,N_7524);
xnor U9237 (N_9237,N_6104,N_6443);
nor U9238 (N_9238,N_7079,N_6896);
and U9239 (N_9239,N_7140,N_7945);
or U9240 (N_9240,N_7880,N_6911);
nand U9241 (N_9241,N_6365,N_7068);
xor U9242 (N_9242,N_6681,N_6184);
nor U9243 (N_9243,N_7706,N_7640);
or U9244 (N_9244,N_7535,N_7074);
or U9245 (N_9245,N_7659,N_6476);
nand U9246 (N_9246,N_7063,N_7013);
or U9247 (N_9247,N_7633,N_6469);
nor U9248 (N_9248,N_7355,N_6929);
xor U9249 (N_9249,N_7675,N_7730);
xnor U9250 (N_9250,N_6735,N_6397);
xor U9251 (N_9251,N_6903,N_7977);
xnor U9252 (N_9252,N_7643,N_6535);
xor U9253 (N_9253,N_6635,N_7275);
and U9254 (N_9254,N_7747,N_6807);
and U9255 (N_9255,N_7880,N_7800);
or U9256 (N_9256,N_6987,N_7026);
nor U9257 (N_9257,N_7617,N_7033);
nand U9258 (N_9258,N_7170,N_6836);
xor U9259 (N_9259,N_7199,N_6870);
or U9260 (N_9260,N_7321,N_6074);
nand U9261 (N_9261,N_6444,N_6498);
nor U9262 (N_9262,N_7738,N_7830);
nand U9263 (N_9263,N_7115,N_7574);
and U9264 (N_9264,N_6308,N_7973);
or U9265 (N_9265,N_6942,N_6476);
or U9266 (N_9266,N_7719,N_7087);
and U9267 (N_9267,N_7491,N_7053);
xnor U9268 (N_9268,N_7521,N_6673);
nand U9269 (N_9269,N_6716,N_7242);
xnor U9270 (N_9270,N_7615,N_6437);
nor U9271 (N_9271,N_6712,N_6174);
and U9272 (N_9272,N_6879,N_6079);
and U9273 (N_9273,N_6512,N_7450);
xnor U9274 (N_9274,N_6236,N_6602);
nand U9275 (N_9275,N_7658,N_6515);
and U9276 (N_9276,N_6395,N_6401);
nor U9277 (N_9277,N_7708,N_7808);
and U9278 (N_9278,N_6561,N_7904);
xnor U9279 (N_9279,N_7651,N_7259);
nand U9280 (N_9280,N_6009,N_6014);
xor U9281 (N_9281,N_6507,N_6077);
or U9282 (N_9282,N_6541,N_6018);
nand U9283 (N_9283,N_6317,N_7847);
or U9284 (N_9284,N_7179,N_7654);
or U9285 (N_9285,N_7685,N_6534);
nor U9286 (N_9286,N_6856,N_7003);
xor U9287 (N_9287,N_7507,N_6108);
nand U9288 (N_9288,N_7414,N_6906);
nand U9289 (N_9289,N_7663,N_7463);
and U9290 (N_9290,N_6772,N_7351);
nor U9291 (N_9291,N_7046,N_7827);
and U9292 (N_9292,N_6486,N_6237);
or U9293 (N_9293,N_7979,N_7152);
nor U9294 (N_9294,N_7249,N_6615);
and U9295 (N_9295,N_7064,N_6768);
nand U9296 (N_9296,N_6224,N_6686);
xnor U9297 (N_9297,N_7977,N_6271);
nand U9298 (N_9298,N_6381,N_6716);
or U9299 (N_9299,N_6943,N_6008);
and U9300 (N_9300,N_6315,N_7841);
nor U9301 (N_9301,N_7773,N_7622);
xor U9302 (N_9302,N_7564,N_6062);
nor U9303 (N_9303,N_6256,N_7849);
and U9304 (N_9304,N_7571,N_7025);
and U9305 (N_9305,N_6145,N_6278);
xnor U9306 (N_9306,N_7999,N_6189);
and U9307 (N_9307,N_7016,N_7514);
nand U9308 (N_9308,N_7601,N_7047);
nor U9309 (N_9309,N_7764,N_7984);
and U9310 (N_9310,N_7473,N_6439);
xnor U9311 (N_9311,N_6478,N_7972);
or U9312 (N_9312,N_7358,N_7775);
or U9313 (N_9313,N_7761,N_6315);
xor U9314 (N_9314,N_6842,N_7762);
nor U9315 (N_9315,N_6518,N_7468);
nand U9316 (N_9316,N_7944,N_7956);
and U9317 (N_9317,N_7259,N_7264);
or U9318 (N_9318,N_7074,N_6386);
nand U9319 (N_9319,N_7224,N_7666);
or U9320 (N_9320,N_7258,N_7314);
or U9321 (N_9321,N_6135,N_7713);
nand U9322 (N_9322,N_6534,N_6554);
and U9323 (N_9323,N_6799,N_6686);
and U9324 (N_9324,N_7780,N_6383);
and U9325 (N_9325,N_7073,N_7414);
nand U9326 (N_9326,N_7380,N_7315);
nor U9327 (N_9327,N_7205,N_6483);
xnor U9328 (N_9328,N_7404,N_6466);
nand U9329 (N_9329,N_6179,N_7347);
and U9330 (N_9330,N_6203,N_7933);
and U9331 (N_9331,N_7143,N_6794);
and U9332 (N_9332,N_6394,N_7413);
and U9333 (N_9333,N_6833,N_6080);
or U9334 (N_9334,N_7503,N_7728);
xor U9335 (N_9335,N_6479,N_6728);
or U9336 (N_9336,N_7316,N_6970);
nor U9337 (N_9337,N_7339,N_6157);
nand U9338 (N_9338,N_7339,N_7025);
nand U9339 (N_9339,N_6975,N_7195);
nor U9340 (N_9340,N_6683,N_7828);
nand U9341 (N_9341,N_7619,N_6927);
nand U9342 (N_9342,N_7482,N_7012);
and U9343 (N_9343,N_7107,N_7120);
nand U9344 (N_9344,N_7576,N_7829);
and U9345 (N_9345,N_7901,N_6474);
and U9346 (N_9346,N_7640,N_7963);
and U9347 (N_9347,N_6701,N_7118);
or U9348 (N_9348,N_6605,N_7713);
nand U9349 (N_9349,N_7320,N_7864);
nor U9350 (N_9350,N_7606,N_6858);
xor U9351 (N_9351,N_7380,N_7213);
xor U9352 (N_9352,N_6618,N_6359);
nor U9353 (N_9353,N_6601,N_6909);
and U9354 (N_9354,N_6378,N_7188);
or U9355 (N_9355,N_7328,N_6264);
and U9356 (N_9356,N_7735,N_6579);
xor U9357 (N_9357,N_6173,N_7804);
nand U9358 (N_9358,N_7489,N_7424);
and U9359 (N_9359,N_7462,N_7609);
and U9360 (N_9360,N_6828,N_7311);
nor U9361 (N_9361,N_6368,N_6724);
and U9362 (N_9362,N_6473,N_6502);
xor U9363 (N_9363,N_6799,N_6485);
nand U9364 (N_9364,N_7010,N_7989);
nand U9365 (N_9365,N_7059,N_6081);
nor U9366 (N_9366,N_7248,N_6232);
or U9367 (N_9367,N_6429,N_7848);
or U9368 (N_9368,N_7188,N_7269);
or U9369 (N_9369,N_6048,N_7884);
xnor U9370 (N_9370,N_7150,N_6443);
nand U9371 (N_9371,N_7017,N_6338);
xor U9372 (N_9372,N_6297,N_6030);
xnor U9373 (N_9373,N_6023,N_6455);
and U9374 (N_9374,N_7101,N_7823);
and U9375 (N_9375,N_7740,N_7928);
xnor U9376 (N_9376,N_7477,N_6844);
or U9377 (N_9377,N_6179,N_6669);
nand U9378 (N_9378,N_7734,N_7140);
and U9379 (N_9379,N_7316,N_7193);
nor U9380 (N_9380,N_7508,N_7843);
nor U9381 (N_9381,N_7419,N_6955);
nand U9382 (N_9382,N_6828,N_7914);
xnor U9383 (N_9383,N_7827,N_6200);
nand U9384 (N_9384,N_7462,N_7090);
or U9385 (N_9385,N_6797,N_6071);
and U9386 (N_9386,N_6174,N_7227);
nor U9387 (N_9387,N_6628,N_6750);
or U9388 (N_9388,N_6620,N_7240);
nor U9389 (N_9389,N_7041,N_7161);
nor U9390 (N_9390,N_6839,N_7056);
and U9391 (N_9391,N_7075,N_7383);
nor U9392 (N_9392,N_7116,N_7346);
nand U9393 (N_9393,N_7626,N_6446);
xnor U9394 (N_9394,N_7911,N_7894);
nand U9395 (N_9395,N_7320,N_6190);
or U9396 (N_9396,N_6658,N_7543);
nand U9397 (N_9397,N_6596,N_6936);
or U9398 (N_9398,N_7717,N_7843);
xor U9399 (N_9399,N_7883,N_6964);
nand U9400 (N_9400,N_6196,N_6124);
nand U9401 (N_9401,N_7426,N_6358);
nor U9402 (N_9402,N_6655,N_6749);
xor U9403 (N_9403,N_7463,N_6952);
nand U9404 (N_9404,N_7520,N_6261);
nand U9405 (N_9405,N_7721,N_6463);
xor U9406 (N_9406,N_7270,N_6270);
xor U9407 (N_9407,N_7807,N_7605);
and U9408 (N_9408,N_6892,N_7402);
and U9409 (N_9409,N_7653,N_6212);
and U9410 (N_9410,N_6147,N_7387);
xnor U9411 (N_9411,N_7583,N_7273);
or U9412 (N_9412,N_6020,N_6423);
nand U9413 (N_9413,N_7301,N_7647);
xor U9414 (N_9414,N_6258,N_6957);
xor U9415 (N_9415,N_6600,N_6250);
or U9416 (N_9416,N_6819,N_7319);
nor U9417 (N_9417,N_7925,N_6529);
xnor U9418 (N_9418,N_6552,N_6994);
and U9419 (N_9419,N_6975,N_7397);
or U9420 (N_9420,N_7593,N_6712);
and U9421 (N_9421,N_6973,N_6332);
or U9422 (N_9422,N_6250,N_6335);
or U9423 (N_9423,N_7041,N_7252);
and U9424 (N_9424,N_7976,N_7503);
or U9425 (N_9425,N_6528,N_7148);
and U9426 (N_9426,N_7596,N_7733);
nand U9427 (N_9427,N_6895,N_7088);
nand U9428 (N_9428,N_6041,N_6142);
xnor U9429 (N_9429,N_7752,N_6986);
xor U9430 (N_9430,N_7831,N_6081);
xor U9431 (N_9431,N_6190,N_7038);
xor U9432 (N_9432,N_7572,N_6672);
or U9433 (N_9433,N_6393,N_7381);
xnor U9434 (N_9434,N_7951,N_7162);
and U9435 (N_9435,N_7981,N_7758);
or U9436 (N_9436,N_6326,N_6951);
and U9437 (N_9437,N_7147,N_7619);
xnor U9438 (N_9438,N_7741,N_6221);
nor U9439 (N_9439,N_7059,N_6857);
nor U9440 (N_9440,N_6921,N_7620);
xor U9441 (N_9441,N_7638,N_7042);
or U9442 (N_9442,N_7317,N_6290);
nor U9443 (N_9443,N_7438,N_7306);
nand U9444 (N_9444,N_7981,N_7149);
and U9445 (N_9445,N_7590,N_7218);
xnor U9446 (N_9446,N_7757,N_6523);
or U9447 (N_9447,N_6666,N_6428);
nor U9448 (N_9448,N_6291,N_7299);
and U9449 (N_9449,N_7528,N_7095);
nor U9450 (N_9450,N_7414,N_7147);
nand U9451 (N_9451,N_7075,N_6316);
nand U9452 (N_9452,N_7580,N_7858);
nor U9453 (N_9453,N_7814,N_6880);
or U9454 (N_9454,N_6651,N_6282);
and U9455 (N_9455,N_6166,N_7191);
or U9456 (N_9456,N_7944,N_7806);
nand U9457 (N_9457,N_7383,N_6648);
nor U9458 (N_9458,N_7101,N_6739);
and U9459 (N_9459,N_7459,N_7621);
xnor U9460 (N_9460,N_7194,N_6718);
nand U9461 (N_9461,N_6515,N_7379);
xnor U9462 (N_9462,N_7550,N_6307);
xor U9463 (N_9463,N_6563,N_6251);
nand U9464 (N_9464,N_7377,N_6062);
xor U9465 (N_9465,N_7517,N_6619);
nand U9466 (N_9466,N_7423,N_6991);
nand U9467 (N_9467,N_6761,N_7908);
nand U9468 (N_9468,N_7493,N_7505);
and U9469 (N_9469,N_6251,N_7233);
nor U9470 (N_9470,N_7042,N_7391);
or U9471 (N_9471,N_6844,N_6803);
or U9472 (N_9472,N_6279,N_6889);
and U9473 (N_9473,N_7563,N_7050);
xnor U9474 (N_9474,N_7943,N_7677);
or U9475 (N_9475,N_7860,N_7474);
or U9476 (N_9476,N_7578,N_6989);
or U9477 (N_9477,N_6353,N_7061);
and U9478 (N_9478,N_6311,N_6962);
nor U9479 (N_9479,N_6903,N_6017);
nand U9480 (N_9480,N_7692,N_6916);
nor U9481 (N_9481,N_6874,N_6964);
and U9482 (N_9482,N_6921,N_7069);
nand U9483 (N_9483,N_6813,N_6134);
nor U9484 (N_9484,N_6323,N_7354);
and U9485 (N_9485,N_7144,N_6241);
xor U9486 (N_9486,N_7252,N_6343);
xnor U9487 (N_9487,N_6110,N_6353);
xor U9488 (N_9488,N_6930,N_6226);
xor U9489 (N_9489,N_7021,N_7901);
and U9490 (N_9490,N_6946,N_6480);
nor U9491 (N_9491,N_7958,N_6958);
nor U9492 (N_9492,N_7065,N_7781);
and U9493 (N_9493,N_6593,N_7683);
nor U9494 (N_9494,N_6176,N_7606);
or U9495 (N_9495,N_7368,N_7017);
xor U9496 (N_9496,N_7336,N_6347);
nor U9497 (N_9497,N_7330,N_6467);
and U9498 (N_9498,N_7638,N_7754);
and U9499 (N_9499,N_7479,N_7444);
nor U9500 (N_9500,N_6095,N_7347);
or U9501 (N_9501,N_7673,N_7392);
and U9502 (N_9502,N_6691,N_6221);
and U9503 (N_9503,N_7704,N_6504);
nand U9504 (N_9504,N_6155,N_7477);
and U9505 (N_9505,N_7463,N_6322);
or U9506 (N_9506,N_7212,N_7039);
and U9507 (N_9507,N_6161,N_7542);
xor U9508 (N_9508,N_6053,N_6891);
or U9509 (N_9509,N_7441,N_6501);
xor U9510 (N_9510,N_7279,N_6096);
or U9511 (N_9511,N_7522,N_7350);
xnor U9512 (N_9512,N_7123,N_6687);
or U9513 (N_9513,N_6481,N_6523);
and U9514 (N_9514,N_6981,N_6416);
nor U9515 (N_9515,N_7180,N_6807);
or U9516 (N_9516,N_7010,N_6017);
nor U9517 (N_9517,N_6418,N_7507);
and U9518 (N_9518,N_7859,N_6337);
xnor U9519 (N_9519,N_6461,N_7818);
nand U9520 (N_9520,N_6332,N_6435);
nand U9521 (N_9521,N_7596,N_6820);
nor U9522 (N_9522,N_6787,N_6049);
xnor U9523 (N_9523,N_7093,N_7736);
or U9524 (N_9524,N_6356,N_7492);
nand U9525 (N_9525,N_7932,N_7540);
xnor U9526 (N_9526,N_7717,N_6470);
nor U9527 (N_9527,N_7408,N_6455);
and U9528 (N_9528,N_6808,N_7042);
and U9529 (N_9529,N_6133,N_6684);
or U9530 (N_9530,N_6500,N_6416);
nor U9531 (N_9531,N_6603,N_6362);
nor U9532 (N_9532,N_7537,N_6504);
or U9533 (N_9533,N_6508,N_6967);
xnor U9534 (N_9534,N_6802,N_6635);
nor U9535 (N_9535,N_7427,N_7130);
nor U9536 (N_9536,N_6420,N_7801);
nor U9537 (N_9537,N_6077,N_6927);
nand U9538 (N_9538,N_6062,N_6486);
or U9539 (N_9539,N_6532,N_7433);
and U9540 (N_9540,N_6167,N_6169);
or U9541 (N_9541,N_6490,N_6115);
and U9542 (N_9542,N_6814,N_7611);
and U9543 (N_9543,N_7307,N_6052);
xor U9544 (N_9544,N_7710,N_6379);
nand U9545 (N_9545,N_7794,N_7695);
xnor U9546 (N_9546,N_6061,N_7029);
xor U9547 (N_9547,N_6525,N_6230);
xnor U9548 (N_9548,N_7601,N_6959);
and U9549 (N_9549,N_6392,N_6503);
and U9550 (N_9550,N_7319,N_7413);
and U9551 (N_9551,N_7283,N_6854);
and U9552 (N_9552,N_7367,N_7594);
and U9553 (N_9553,N_7954,N_7854);
nand U9554 (N_9554,N_7067,N_6133);
and U9555 (N_9555,N_6437,N_7898);
nor U9556 (N_9556,N_7751,N_7798);
nand U9557 (N_9557,N_7600,N_6904);
or U9558 (N_9558,N_6927,N_6014);
or U9559 (N_9559,N_6179,N_6029);
nand U9560 (N_9560,N_7314,N_6563);
xnor U9561 (N_9561,N_6193,N_6291);
xor U9562 (N_9562,N_7502,N_7351);
nor U9563 (N_9563,N_6518,N_7053);
or U9564 (N_9564,N_7935,N_6381);
or U9565 (N_9565,N_6548,N_7981);
nand U9566 (N_9566,N_6668,N_7919);
and U9567 (N_9567,N_7668,N_7281);
and U9568 (N_9568,N_7919,N_6871);
nor U9569 (N_9569,N_7857,N_7501);
nand U9570 (N_9570,N_6596,N_7459);
xor U9571 (N_9571,N_6445,N_6603);
or U9572 (N_9572,N_6438,N_6555);
and U9573 (N_9573,N_7069,N_6711);
nand U9574 (N_9574,N_7828,N_6638);
or U9575 (N_9575,N_6259,N_6027);
nand U9576 (N_9576,N_6740,N_6828);
nor U9577 (N_9577,N_7441,N_7499);
nand U9578 (N_9578,N_6292,N_7251);
or U9579 (N_9579,N_6794,N_6540);
and U9580 (N_9580,N_7730,N_7108);
nor U9581 (N_9581,N_6485,N_6672);
and U9582 (N_9582,N_6848,N_7668);
xnor U9583 (N_9583,N_7670,N_6041);
nand U9584 (N_9584,N_6134,N_7275);
nor U9585 (N_9585,N_6835,N_6550);
nor U9586 (N_9586,N_6426,N_7449);
or U9587 (N_9587,N_6610,N_6265);
and U9588 (N_9588,N_6980,N_6547);
and U9589 (N_9589,N_7917,N_6447);
xor U9590 (N_9590,N_7064,N_6703);
nand U9591 (N_9591,N_6456,N_7575);
nor U9592 (N_9592,N_6955,N_7727);
xnor U9593 (N_9593,N_7998,N_7226);
or U9594 (N_9594,N_7748,N_7890);
nor U9595 (N_9595,N_6940,N_6045);
nand U9596 (N_9596,N_6130,N_6552);
xnor U9597 (N_9597,N_6496,N_6993);
nor U9598 (N_9598,N_6467,N_7622);
or U9599 (N_9599,N_6592,N_7164);
and U9600 (N_9600,N_6312,N_7616);
nor U9601 (N_9601,N_7469,N_7316);
or U9602 (N_9602,N_6944,N_6705);
nor U9603 (N_9603,N_6333,N_7874);
nor U9604 (N_9604,N_7996,N_6274);
and U9605 (N_9605,N_6843,N_6368);
xor U9606 (N_9606,N_6154,N_7819);
and U9607 (N_9607,N_6239,N_7031);
xor U9608 (N_9608,N_6030,N_6655);
or U9609 (N_9609,N_6864,N_6971);
nand U9610 (N_9610,N_6855,N_7488);
nand U9611 (N_9611,N_6175,N_7026);
nand U9612 (N_9612,N_7087,N_7515);
nor U9613 (N_9613,N_6382,N_7840);
xnor U9614 (N_9614,N_6286,N_7833);
xnor U9615 (N_9615,N_7334,N_7591);
nand U9616 (N_9616,N_6659,N_6821);
or U9617 (N_9617,N_6859,N_6329);
nand U9618 (N_9618,N_7945,N_7237);
xor U9619 (N_9619,N_7713,N_7206);
and U9620 (N_9620,N_6402,N_6767);
or U9621 (N_9621,N_6794,N_6552);
xor U9622 (N_9622,N_7300,N_7969);
nand U9623 (N_9623,N_7501,N_7080);
or U9624 (N_9624,N_6694,N_7900);
and U9625 (N_9625,N_7622,N_6312);
nand U9626 (N_9626,N_7135,N_7062);
and U9627 (N_9627,N_6374,N_7774);
xnor U9628 (N_9628,N_6972,N_7020);
nor U9629 (N_9629,N_6301,N_7352);
nor U9630 (N_9630,N_6079,N_6402);
xor U9631 (N_9631,N_7378,N_7724);
nor U9632 (N_9632,N_7609,N_7793);
xor U9633 (N_9633,N_6794,N_7210);
and U9634 (N_9634,N_6380,N_6585);
nand U9635 (N_9635,N_7572,N_7145);
and U9636 (N_9636,N_6376,N_6193);
or U9637 (N_9637,N_7400,N_6832);
or U9638 (N_9638,N_6323,N_6024);
nor U9639 (N_9639,N_7991,N_7328);
xor U9640 (N_9640,N_7162,N_6668);
xor U9641 (N_9641,N_6640,N_7667);
and U9642 (N_9642,N_6309,N_7328);
and U9643 (N_9643,N_7908,N_7544);
and U9644 (N_9644,N_7983,N_6690);
and U9645 (N_9645,N_6336,N_7783);
nand U9646 (N_9646,N_6289,N_7134);
and U9647 (N_9647,N_6112,N_6355);
and U9648 (N_9648,N_6473,N_7825);
nor U9649 (N_9649,N_7450,N_7389);
xor U9650 (N_9650,N_6984,N_6830);
and U9651 (N_9651,N_6768,N_7048);
xnor U9652 (N_9652,N_7077,N_7403);
or U9653 (N_9653,N_6100,N_6185);
and U9654 (N_9654,N_6103,N_7959);
nor U9655 (N_9655,N_6560,N_7826);
or U9656 (N_9656,N_6800,N_6452);
or U9657 (N_9657,N_7100,N_6635);
xnor U9658 (N_9658,N_6671,N_6154);
and U9659 (N_9659,N_6406,N_7185);
xnor U9660 (N_9660,N_7867,N_6949);
nor U9661 (N_9661,N_6226,N_6089);
xnor U9662 (N_9662,N_6794,N_7372);
nor U9663 (N_9663,N_7596,N_6372);
and U9664 (N_9664,N_7455,N_6109);
xnor U9665 (N_9665,N_7204,N_7265);
and U9666 (N_9666,N_6006,N_7579);
nand U9667 (N_9667,N_6328,N_6882);
or U9668 (N_9668,N_7041,N_6963);
or U9669 (N_9669,N_7814,N_6524);
or U9670 (N_9670,N_7057,N_6332);
and U9671 (N_9671,N_7365,N_7170);
nand U9672 (N_9672,N_6235,N_7232);
and U9673 (N_9673,N_6302,N_7402);
and U9674 (N_9674,N_7058,N_7924);
or U9675 (N_9675,N_6968,N_6190);
nand U9676 (N_9676,N_7235,N_7945);
and U9677 (N_9677,N_6370,N_7665);
xnor U9678 (N_9678,N_7575,N_6180);
xnor U9679 (N_9679,N_7108,N_6977);
xor U9680 (N_9680,N_6707,N_6585);
nand U9681 (N_9681,N_6809,N_6431);
nor U9682 (N_9682,N_7450,N_6338);
nand U9683 (N_9683,N_7107,N_7476);
or U9684 (N_9684,N_7553,N_7322);
nor U9685 (N_9685,N_7103,N_7101);
xnor U9686 (N_9686,N_6817,N_7940);
nand U9687 (N_9687,N_6578,N_6217);
and U9688 (N_9688,N_6871,N_6666);
or U9689 (N_9689,N_6184,N_7711);
nand U9690 (N_9690,N_7547,N_7844);
nand U9691 (N_9691,N_6225,N_6871);
or U9692 (N_9692,N_6310,N_6364);
nor U9693 (N_9693,N_7226,N_7973);
or U9694 (N_9694,N_7043,N_6934);
nand U9695 (N_9695,N_6205,N_7114);
nand U9696 (N_9696,N_6060,N_6600);
nor U9697 (N_9697,N_7098,N_7255);
xor U9698 (N_9698,N_6014,N_6685);
nor U9699 (N_9699,N_7730,N_6040);
nand U9700 (N_9700,N_6311,N_7300);
nand U9701 (N_9701,N_6240,N_6621);
or U9702 (N_9702,N_6623,N_6230);
or U9703 (N_9703,N_7980,N_7486);
nand U9704 (N_9704,N_6577,N_6403);
and U9705 (N_9705,N_7508,N_7129);
or U9706 (N_9706,N_7053,N_6573);
xnor U9707 (N_9707,N_6585,N_6163);
xor U9708 (N_9708,N_7522,N_7882);
or U9709 (N_9709,N_6038,N_6676);
nand U9710 (N_9710,N_7411,N_6609);
nor U9711 (N_9711,N_7974,N_6500);
and U9712 (N_9712,N_6618,N_7645);
xnor U9713 (N_9713,N_7063,N_7813);
or U9714 (N_9714,N_7672,N_7062);
and U9715 (N_9715,N_7485,N_6900);
nand U9716 (N_9716,N_7824,N_6566);
and U9717 (N_9717,N_6104,N_6078);
nand U9718 (N_9718,N_6368,N_7545);
nor U9719 (N_9719,N_6664,N_7404);
or U9720 (N_9720,N_7765,N_6278);
nand U9721 (N_9721,N_6372,N_6419);
or U9722 (N_9722,N_7720,N_7695);
xor U9723 (N_9723,N_6874,N_6406);
nor U9724 (N_9724,N_7186,N_6107);
and U9725 (N_9725,N_7948,N_7587);
nor U9726 (N_9726,N_6668,N_6357);
nor U9727 (N_9727,N_7783,N_6787);
and U9728 (N_9728,N_7111,N_7574);
nor U9729 (N_9729,N_7941,N_6193);
nor U9730 (N_9730,N_7233,N_6600);
xnor U9731 (N_9731,N_6666,N_7740);
nor U9732 (N_9732,N_6252,N_7409);
nand U9733 (N_9733,N_7986,N_6463);
xnor U9734 (N_9734,N_6025,N_7428);
xnor U9735 (N_9735,N_7154,N_6267);
nand U9736 (N_9736,N_6018,N_7749);
xnor U9737 (N_9737,N_7590,N_7072);
nand U9738 (N_9738,N_7013,N_7528);
and U9739 (N_9739,N_7776,N_6436);
or U9740 (N_9740,N_6206,N_7571);
nor U9741 (N_9741,N_6686,N_6979);
nand U9742 (N_9742,N_6878,N_6968);
nand U9743 (N_9743,N_6135,N_6826);
nor U9744 (N_9744,N_7898,N_6817);
or U9745 (N_9745,N_7356,N_6349);
nor U9746 (N_9746,N_7039,N_6027);
xnor U9747 (N_9747,N_6547,N_6619);
nand U9748 (N_9748,N_6948,N_6944);
nor U9749 (N_9749,N_7728,N_6987);
nand U9750 (N_9750,N_7425,N_7073);
nand U9751 (N_9751,N_7087,N_6539);
nand U9752 (N_9752,N_6083,N_7468);
or U9753 (N_9753,N_6260,N_6298);
xor U9754 (N_9754,N_7135,N_7436);
nand U9755 (N_9755,N_6904,N_6696);
nor U9756 (N_9756,N_7183,N_7217);
nand U9757 (N_9757,N_7663,N_7937);
and U9758 (N_9758,N_7026,N_6690);
nand U9759 (N_9759,N_6287,N_6666);
or U9760 (N_9760,N_6168,N_6861);
nand U9761 (N_9761,N_6585,N_6355);
and U9762 (N_9762,N_6871,N_6233);
and U9763 (N_9763,N_7267,N_7357);
or U9764 (N_9764,N_6441,N_7524);
nand U9765 (N_9765,N_7841,N_6745);
xnor U9766 (N_9766,N_6365,N_6024);
or U9767 (N_9767,N_6609,N_7689);
and U9768 (N_9768,N_6319,N_7933);
and U9769 (N_9769,N_6972,N_7869);
xnor U9770 (N_9770,N_7401,N_7452);
nand U9771 (N_9771,N_6396,N_6806);
nor U9772 (N_9772,N_6585,N_7154);
nor U9773 (N_9773,N_6020,N_7744);
or U9774 (N_9774,N_7476,N_6781);
or U9775 (N_9775,N_6078,N_6458);
xnor U9776 (N_9776,N_6583,N_7087);
nand U9777 (N_9777,N_6336,N_6022);
xnor U9778 (N_9778,N_6959,N_7654);
nand U9779 (N_9779,N_6578,N_7711);
or U9780 (N_9780,N_6021,N_6700);
xnor U9781 (N_9781,N_6811,N_6600);
and U9782 (N_9782,N_6944,N_6069);
and U9783 (N_9783,N_6392,N_7326);
nand U9784 (N_9784,N_7991,N_6181);
xnor U9785 (N_9785,N_6921,N_6549);
nand U9786 (N_9786,N_7074,N_7755);
nor U9787 (N_9787,N_6354,N_6266);
nor U9788 (N_9788,N_7433,N_7392);
nor U9789 (N_9789,N_7329,N_7426);
nor U9790 (N_9790,N_6560,N_7564);
nand U9791 (N_9791,N_7695,N_7383);
nor U9792 (N_9792,N_6375,N_6808);
nand U9793 (N_9793,N_7950,N_6668);
xor U9794 (N_9794,N_6991,N_7045);
nor U9795 (N_9795,N_6412,N_6680);
xnor U9796 (N_9796,N_7311,N_6365);
or U9797 (N_9797,N_6319,N_7781);
and U9798 (N_9798,N_7742,N_7357);
nand U9799 (N_9799,N_6486,N_7009);
and U9800 (N_9800,N_7622,N_6880);
nor U9801 (N_9801,N_6557,N_6167);
nor U9802 (N_9802,N_6431,N_6773);
nand U9803 (N_9803,N_6235,N_7427);
or U9804 (N_9804,N_7036,N_7512);
xnor U9805 (N_9805,N_6258,N_7117);
xnor U9806 (N_9806,N_7099,N_6673);
and U9807 (N_9807,N_7382,N_7649);
or U9808 (N_9808,N_7826,N_7339);
and U9809 (N_9809,N_6060,N_6145);
nor U9810 (N_9810,N_7622,N_6867);
nor U9811 (N_9811,N_6613,N_6135);
and U9812 (N_9812,N_7938,N_6103);
and U9813 (N_9813,N_6103,N_6107);
and U9814 (N_9814,N_7861,N_6011);
or U9815 (N_9815,N_6599,N_7232);
xnor U9816 (N_9816,N_7327,N_7528);
xor U9817 (N_9817,N_7961,N_6409);
or U9818 (N_9818,N_7030,N_7502);
and U9819 (N_9819,N_7626,N_7062);
nand U9820 (N_9820,N_7881,N_6110);
nand U9821 (N_9821,N_6699,N_6669);
nor U9822 (N_9822,N_7476,N_7665);
or U9823 (N_9823,N_7124,N_6569);
and U9824 (N_9824,N_7059,N_6800);
nor U9825 (N_9825,N_6095,N_7520);
or U9826 (N_9826,N_6916,N_7235);
nor U9827 (N_9827,N_7643,N_6114);
xor U9828 (N_9828,N_7034,N_6609);
xor U9829 (N_9829,N_6910,N_7603);
xor U9830 (N_9830,N_7101,N_7471);
nor U9831 (N_9831,N_7285,N_6038);
and U9832 (N_9832,N_6700,N_6045);
nand U9833 (N_9833,N_7581,N_6942);
xnor U9834 (N_9834,N_7603,N_7425);
or U9835 (N_9835,N_7768,N_7454);
and U9836 (N_9836,N_7620,N_7591);
and U9837 (N_9837,N_6418,N_6599);
or U9838 (N_9838,N_6642,N_7877);
and U9839 (N_9839,N_7436,N_7775);
nor U9840 (N_9840,N_7390,N_7309);
nand U9841 (N_9841,N_7059,N_7851);
xnor U9842 (N_9842,N_6285,N_6141);
nor U9843 (N_9843,N_7938,N_6768);
xor U9844 (N_9844,N_6992,N_6895);
xor U9845 (N_9845,N_6522,N_7537);
nor U9846 (N_9846,N_6324,N_6540);
xnor U9847 (N_9847,N_7318,N_7761);
nor U9848 (N_9848,N_6491,N_6456);
nand U9849 (N_9849,N_6164,N_6480);
nand U9850 (N_9850,N_7161,N_6019);
nand U9851 (N_9851,N_6876,N_6234);
and U9852 (N_9852,N_7282,N_6044);
or U9853 (N_9853,N_7439,N_6034);
and U9854 (N_9854,N_6565,N_6879);
nand U9855 (N_9855,N_7232,N_6045);
nand U9856 (N_9856,N_7634,N_7432);
xnor U9857 (N_9857,N_6834,N_6335);
xnor U9858 (N_9858,N_6867,N_6193);
or U9859 (N_9859,N_6464,N_6737);
xnor U9860 (N_9860,N_7298,N_6994);
nand U9861 (N_9861,N_6332,N_7714);
xor U9862 (N_9862,N_7808,N_7590);
xnor U9863 (N_9863,N_7861,N_6022);
nor U9864 (N_9864,N_6990,N_7945);
nand U9865 (N_9865,N_6388,N_7212);
and U9866 (N_9866,N_7771,N_6148);
and U9867 (N_9867,N_6331,N_6089);
or U9868 (N_9868,N_6030,N_6885);
xor U9869 (N_9869,N_6375,N_7384);
nor U9870 (N_9870,N_7182,N_6602);
and U9871 (N_9871,N_6680,N_7934);
nand U9872 (N_9872,N_7877,N_6307);
and U9873 (N_9873,N_7267,N_6137);
nand U9874 (N_9874,N_7616,N_6728);
nor U9875 (N_9875,N_7053,N_7598);
xnor U9876 (N_9876,N_6359,N_7232);
and U9877 (N_9877,N_6106,N_7192);
or U9878 (N_9878,N_7625,N_6878);
nand U9879 (N_9879,N_7302,N_7745);
nor U9880 (N_9880,N_6858,N_6736);
xnor U9881 (N_9881,N_6689,N_7041);
or U9882 (N_9882,N_6174,N_7152);
xnor U9883 (N_9883,N_6409,N_6663);
nor U9884 (N_9884,N_6173,N_7202);
xnor U9885 (N_9885,N_7179,N_6484);
nor U9886 (N_9886,N_7304,N_7668);
or U9887 (N_9887,N_7204,N_6556);
xor U9888 (N_9888,N_7513,N_6146);
or U9889 (N_9889,N_7567,N_6344);
and U9890 (N_9890,N_6198,N_6974);
nor U9891 (N_9891,N_7867,N_6582);
nand U9892 (N_9892,N_7984,N_7905);
and U9893 (N_9893,N_6315,N_6036);
or U9894 (N_9894,N_7958,N_6336);
nor U9895 (N_9895,N_7214,N_6004);
and U9896 (N_9896,N_7949,N_6297);
or U9897 (N_9897,N_7193,N_6198);
or U9898 (N_9898,N_6948,N_7104);
nand U9899 (N_9899,N_7765,N_7467);
nor U9900 (N_9900,N_7326,N_6382);
xnor U9901 (N_9901,N_6063,N_7062);
or U9902 (N_9902,N_7030,N_7690);
or U9903 (N_9903,N_7847,N_7609);
nor U9904 (N_9904,N_6405,N_7702);
xnor U9905 (N_9905,N_7986,N_6160);
and U9906 (N_9906,N_6768,N_7757);
nor U9907 (N_9907,N_6019,N_7520);
nor U9908 (N_9908,N_6508,N_7794);
xor U9909 (N_9909,N_7151,N_6625);
xnor U9910 (N_9910,N_6396,N_7716);
and U9911 (N_9911,N_7446,N_7556);
nand U9912 (N_9912,N_6643,N_7782);
or U9913 (N_9913,N_6856,N_7112);
or U9914 (N_9914,N_6073,N_7532);
and U9915 (N_9915,N_6280,N_6434);
or U9916 (N_9916,N_6315,N_6972);
or U9917 (N_9917,N_6306,N_7178);
xor U9918 (N_9918,N_7465,N_7012);
nor U9919 (N_9919,N_6720,N_7532);
xnor U9920 (N_9920,N_7267,N_7781);
xor U9921 (N_9921,N_7451,N_6099);
xor U9922 (N_9922,N_7779,N_7592);
nor U9923 (N_9923,N_7091,N_6869);
nand U9924 (N_9924,N_7406,N_6073);
nand U9925 (N_9925,N_6327,N_7098);
or U9926 (N_9926,N_6219,N_7367);
nor U9927 (N_9927,N_7513,N_6169);
and U9928 (N_9928,N_7500,N_6676);
or U9929 (N_9929,N_6824,N_6677);
nand U9930 (N_9930,N_6324,N_6993);
nand U9931 (N_9931,N_6489,N_7418);
and U9932 (N_9932,N_7859,N_7135);
and U9933 (N_9933,N_6432,N_6535);
nand U9934 (N_9934,N_6526,N_6956);
and U9935 (N_9935,N_7363,N_6775);
xnor U9936 (N_9936,N_7483,N_6404);
nor U9937 (N_9937,N_6900,N_7535);
nand U9938 (N_9938,N_7895,N_6914);
xnor U9939 (N_9939,N_6003,N_7353);
nor U9940 (N_9940,N_6247,N_6181);
or U9941 (N_9941,N_6912,N_6400);
nand U9942 (N_9942,N_7104,N_6509);
nand U9943 (N_9943,N_7927,N_6773);
nand U9944 (N_9944,N_6803,N_7848);
xor U9945 (N_9945,N_7311,N_6765);
or U9946 (N_9946,N_6330,N_7931);
nand U9947 (N_9947,N_6777,N_7918);
xor U9948 (N_9948,N_7510,N_6688);
nor U9949 (N_9949,N_6994,N_7638);
or U9950 (N_9950,N_7666,N_6595);
and U9951 (N_9951,N_6075,N_6901);
nor U9952 (N_9952,N_6247,N_6998);
nor U9953 (N_9953,N_7147,N_7652);
nand U9954 (N_9954,N_7264,N_6998);
or U9955 (N_9955,N_7651,N_7726);
xnor U9956 (N_9956,N_6236,N_7632);
nor U9957 (N_9957,N_7309,N_7769);
xnor U9958 (N_9958,N_7716,N_6250);
xnor U9959 (N_9959,N_6483,N_6142);
nor U9960 (N_9960,N_7673,N_7793);
and U9961 (N_9961,N_7978,N_7937);
nand U9962 (N_9962,N_6785,N_7151);
nand U9963 (N_9963,N_7753,N_6111);
nand U9964 (N_9964,N_7889,N_6817);
or U9965 (N_9965,N_6562,N_6148);
xnor U9966 (N_9966,N_7962,N_6562);
and U9967 (N_9967,N_6271,N_7195);
nand U9968 (N_9968,N_7424,N_7832);
or U9969 (N_9969,N_6706,N_7450);
nor U9970 (N_9970,N_6325,N_7706);
or U9971 (N_9971,N_6891,N_6586);
xor U9972 (N_9972,N_6367,N_6192);
or U9973 (N_9973,N_7707,N_6896);
or U9974 (N_9974,N_6731,N_6000);
nor U9975 (N_9975,N_7937,N_6267);
xor U9976 (N_9976,N_7394,N_7525);
nor U9977 (N_9977,N_7979,N_7976);
and U9978 (N_9978,N_7287,N_7351);
nor U9979 (N_9979,N_6003,N_6204);
nand U9980 (N_9980,N_6629,N_7497);
xnor U9981 (N_9981,N_7455,N_7992);
or U9982 (N_9982,N_7572,N_7465);
nor U9983 (N_9983,N_7977,N_7252);
or U9984 (N_9984,N_7386,N_7475);
or U9985 (N_9985,N_7084,N_6362);
nand U9986 (N_9986,N_6897,N_7175);
nand U9987 (N_9987,N_7129,N_7108);
nand U9988 (N_9988,N_6594,N_6595);
xor U9989 (N_9989,N_7961,N_6301);
nor U9990 (N_9990,N_6281,N_6368);
and U9991 (N_9991,N_6633,N_6418);
or U9992 (N_9992,N_6680,N_7720);
and U9993 (N_9993,N_6688,N_7145);
nor U9994 (N_9994,N_6703,N_7376);
and U9995 (N_9995,N_6303,N_7150);
xnor U9996 (N_9996,N_6674,N_6756);
xor U9997 (N_9997,N_7970,N_7047);
or U9998 (N_9998,N_6000,N_6206);
nand U9999 (N_9999,N_7312,N_6572);
and U10000 (N_10000,N_9951,N_9866);
or U10001 (N_10001,N_8286,N_8300);
and U10002 (N_10002,N_9145,N_8293);
nor U10003 (N_10003,N_8511,N_9012);
or U10004 (N_10004,N_8119,N_9739);
nor U10005 (N_10005,N_8120,N_9035);
nand U10006 (N_10006,N_8464,N_8797);
or U10007 (N_10007,N_9728,N_8156);
and U10008 (N_10008,N_8658,N_8834);
and U10009 (N_10009,N_9000,N_9967);
nor U10010 (N_10010,N_8446,N_8673);
nand U10011 (N_10011,N_9124,N_9348);
xor U10012 (N_10012,N_8984,N_8266);
and U10013 (N_10013,N_9864,N_9171);
xnor U10014 (N_10014,N_9977,N_9989);
and U10015 (N_10015,N_8296,N_9644);
nand U10016 (N_10016,N_8486,N_9935);
and U10017 (N_10017,N_8132,N_9328);
or U10018 (N_10018,N_8155,N_9112);
or U10019 (N_10019,N_9815,N_8488);
xnor U10020 (N_10020,N_8198,N_9104);
and U10021 (N_10021,N_9660,N_8543);
xor U10022 (N_10022,N_9257,N_9220);
xor U10023 (N_10023,N_9318,N_8302);
and U10024 (N_10024,N_8659,N_9811);
xor U10025 (N_10025,N_8676,N_8416);
nor U10026 (N_10026,N_9006,N_9478);
or U10027 (N_10027,N_9261,N_9139);
nand U10028 (N_10028,N_8480,N_9681);
xor U10029 (N_10029,N_9835,N_8079);
xnor U10030 (N_10030,N_9201,N_9309);
and U10031 (N_10031,N_9673,N_9441);
or U10032 (N_10032,N_9380,N_8831);
nor U10033 (N_10033,N_8711,N_8474);
and U10034 (N_10034,N_8310,N_9860);
and U10035 (N_10035,N_8648,N_9926);
and U10036 (N_10036,N_9600,N_9718);
nand U10037 (N_10037,N_9232,N_8779);
xor U10038 (N_10038,N_8569,N_9507);
nand U10039 (N_10039,N_9493,N_8023);
xnor U10040 (N_10040,N_8548,N_9604);
nor U10041 (N_10041,N_8072,N_9900);
xor U10042 (N_10042,N_9912,N_9529);
and U10043 (N_10043,N_9253,N_8083);
nor U10044 (N_10044,N_9639,N_8895);
or U10045 (N_10045,N_9931,N_8517);
or U10046 (N_10046,N_8759,N_8894);
or U10047 (N_10047,N_9239,N_9704);
nand U10048 (N_10048,N_9160,N_8228);
nor U10049 (N_10049,N_8448,N_9762);
and U10050 (N_10050,N_9522,N_9980);
nor U10051 (N_10051,N_8458,N_9116);
or U10052 (N_10052,N_9668,N_8267);
nor U10053 (N_10053,N_9975,N_9260);
and U10054 (N_10054,N_9636,N_9455);
xnor U10055 (N_10055,N_9939,N_9616);
nor U10056 (N_10056,N_8399,N_9126);
and U10057 (N_10057,N_9407,N_8269);
and U10058 (N_10058,N_8146,N_9779);
nand U10059 (N_10059,N_8563,N_8104);
and U10060 (N_10060,N_8793,N_9483);
or U10061 (N_10061,N_8046,N_9898);
and U10062 (N_10062,N_8504,N_9674);
and U10063 (N_10063,N_9504,N_9712);
nor U10064 (N_10064,N_8145,N_9786);
nor U10065 (N_10065,N_8126,N_8655);
or U10066 (N_10066,N_8394,N_9008);
xnor U10067 (N_10067,N_9894,N_9468);
xor U10068 (N_10068,N_8103,N_9439);
and U10069 (N_10069,N_9254,N_8249);
nand U10070 (N_10070,N_8647,N_9375);
nand U10071 (N_10071,N_8827,N_9320);
nand U10072 (N_10072,N_8964,N_9177);
nor U10073 (N_10073,N_8945,N_9958);
and U10074 (N_10074,N_9875,N_8348);
nor U10075 (N_10075,N_9885,N_8116);
and U10076 (N_10076,N_8304,N_9621);
or U10077 (N_10077,N_8874,N_8843);
nand U10078 (N_10078,N_8076,N_8953);
nand U10079 (N_10079,N_8439,N_8508);
nand U10080 (N_10080,N_9515,N_9047);
or U10081 (N_10081,N_9530,N_8096);
xnor U10082 (N_10082,N_8883,N_8541);
and U10083 (N_10083,N_8067,N_9999);
nand U10084 (N_10084,N_9060,N_8520);
nor U10085 (N_10085,N_8477,N_8966);
xor U10086 (N_10086,N_9776,N_9783);
nand U10087 (N_10087,N_8778,N_9358);
nor U10088 (N_10088,N_9959,N_8705);
and U10089 (N_10089,N_8333,N_9542);
and U10090 (N_10090,N_9315,N_9852);
xor U10091 (N_10091,N_8396,N_8173);
xnor U10092 (N_10092,N_8929,N_8913);
xor U10093 (N_10093,N_8846,N_9151);
xnor U10094 (N_10094,N_9297,N_9284);
and U10095 (N_10095,N_8581,N_8959);
nor U10096 (N_10096,N_9357,N_8727);
nand U10097 (N_10097,N_8932,N_9577);
or U10098 (N_10098,N_8652,N_9250);
nand U10099 (N_10099,N_9453,N_9140);
and U10100 (N_10100,N_9196,N_8558);
or U10101 (N_10101,N_9136,N_9765);
and U10102 (N_10102,N_9998,N_8789);
and U10103 (N_10103,N_8224,N_8197);
nand U10104 (N_10104,N_8250,N_9994);
and U10105 (N_10105,N_8426,N_8366);
and U10106 (N_10106,N_9859,N_9552);
xnor U10107 (N_10107,N_8958,N_8766);
nor U10108 (N_10108,N_8259,N_9854);
xor U10109 (N_10109,N_9186,N_9606);
or U10110 (N_10110,N_8842,N_9321);
and U10111 (N_10111,N_8899,N_9591);
nand U10112 (N_10112,N_8178,N_8127);
xnor U10113 (N_10113,N_9426,N_9554);
and U10114 (N_10114,N_9856,N_9784);
and U10115 (N_10115,N_9929,N_9043);
xor U10116 (N_10116,N_8395,N_9678);
and U10117 (N_10117,N_9039,N_9509);
and U10118 (N_10118,N_8410,N_9755);
nand U10119 (N_10119,N_8599,N_8080);
nor U10120 (N_10120,N_9170,N_8334);
or U10121 (N_10121,N_8704,N_8926);
or U10122 (N_10122,N_9661,N_8923);
or U10123 (N_10123,N_9026,N_9524);
nor U10124 (N_10124,N_8176,N_9518);
xnor U10125 (N_10125,N_9411,N_9448);
nand U10126 (N_10126,N_8876,N_9608);
xnor U10127 (N_10127,N_8890,N_8358);
or U10128 (N_10128,N_8280,N_9467);
and U10129 (N_10129,N_9569,N_9570);
nand U10130 (N_10130,N_8376,N_9602);
nand U10131 (N_10131,N_8552,N_9651);
or U10132 (N_10132,N_9212,N_8775);
nor U10133 (N_10133,N_8559,N_9079);
or U10134 (N_10134,N_9174,N_9816);
xor U10135 (N_10135,N_8963,N_8449);
nor U10136 (N_10136,N_8615,N_9512);
nor U10137 (N_10137,N_8089,N_9390);
nor U10138 (N_10138,N_8368,N_9848);
and U10139 (N_10139,N_8755,N_9155);
xnor U10140 (N_10140,N_9027,N_9785);
and U10141 (N_10141,N_9846,N_9323);
xnor U10142 (N_10142,N_8974,N_9858);
nor U10143 (N_10143,N_9832,N_8007);
nor U10144 (N_10144,N_9156,N_8382);
and U10145 (N_10145,N_8037,N_9218);
and U10146 (N_10146,N_8812,N_8716);
xor U10147 (N_10147,N_8062,N_9022);
xor U10148 (N_10148,N_9640,N_9495);
and U10149 (N_10149,N_8768,N_8671);
xnor U10150 (N_10150,N_8459,N_8896);
nor U10151 (N_10151,N_9396,N_9995);
and U10152 (N_10152,N_8139,N_9625);
nand U10153 (N_10153,N_9557,N_9833);
xor U10154 (N_10154,N_8022,N_9839);
xnor U10155 (N_10155,N_8186,N_8568);
xor U10156 (N_10156,N_8586,N_8030);
xor U10157 (N_10157,N_8408,N_8175);
nor U10158 (N_10158,N_8624,N_8814);
xor U10159 (N_10159,N_8108,N_8445);
nor U10160 (N_10160,N_8816,N_9695);
and U10161 (N_10161,N_8038,N_9029);
nand U10162 (N_10162,N_9275,N_8684);
nand U10163 (N_10163,N_9389,N_9325);
nand U10164 (N_10164,N_8940,N_8740);
nor U10165 (N_10165,N_8373,N_8193);
xnor U10166 (N_10166,N_8493,N_8109);
nand U10167 (N_10167,N_9751,N_8743);
nor U10168 (N_10168,N_8747,N_8646);
and U10169 (N_10169,N_8004,N_9419);
xnor U10170 (N_10170,N_8950,N_9298);
and U10171 (N_10171,N_9295,N_8774);
and U10172 (N_10172,N_8035,N_8528);
and U10173 (N_10173,N_9282,N_9161);
xnor U10174 (N_10174,N_9773,N_8582);
nand U10175 (N_10175,N_9222,N_9986);
or U10176 (N_10176,N_8554,N_8318);
nor U10177 (N_10177,N_8125,N_9133);
xor U10178 (N_10178,N_9702,N_9756);
nor U10179 (N_10179,N_8041,N_9682);
xor U10180 (N_10180,N_8245,N_9292);
nand U10181 (N_10181,N_8536,N_8979);
and U10182 (N_10182,N_8235,N_8463);
or U10183 (N_10183,N_9603,N_8687);
or U10184 (N_10184,N_8593,N_9761);
nand U10185 (N_10185,N_8131,N_9760);
and U10186 (N_10186,N_9586,N_9451);
nor U10187 (N_10187,N_9664,N_9184);
nor U10188 (N_10188,N_8147,N_8380);
or U10189 (N_10189,N_9537,N_8000);
or U10190 (N_10190,N_8858,N_8886);
xor U10191 (N_10191,N_9410,N_9534);
or U10192 (N_10192,N_8393,N_8608);
or U10193 (N_10193,N_8623,N_9662);
xnor U10194 (N_10194,N_9683,N_8203);
nand U10195 (N_10195,N_8326,N_9742);
nand U10196 (N_10196,N_9709,N_8996);
nor U10197 (N_10197,N_8044,N_8353);
nand U10198 (N_10198,N_9023,N_9217);
and U10199 (N_10199,N_8026,N_9412);
nand U10200 (N_10200,N_9965,N_9204);
nor U10201 (N_10201,N_8534,N_8758);
nand U10202 (N_10202,N_8935,N_9107);
xor U10203 (N_10203,N_8330,N_9115);
or U10204 (N_10204,N_8248,N_8595);
or U10205 (N_10205,N_8532,N_9422);
xor U10206 (N_10206,N_9802,N_8028);
nor U10207 (N_10207,N_8164,N_8725);
or U10208 (N_10208,N_8881,N_9893);
and U10209 (N_10209,N_9423,N_8021);
and U10210 (N_10210,N_9111,N_8994);
nand U10211 (N_10211,N_9219,N_8675);
and U10212 (N_10212,N_9082,N_8815);
xnor U10213 (N_10213,N_9091,N_8682);
and U10214 (N_10214,N_8140,N_9906);
and U10215 (N_10215,N_8009,N_9937);
nor U10216 (N_10216,N_8356,N_9098);
or U10217 (N_10217,N_8268,N_8664);
or U10218 (N_10218,N_8482,N_8257);
xnor U10219 (N_10219,N_9032,N_9233);
and U10220 (N_10220,N_8010,N_8202);
or U10221 (N_10221,N_9214,N_8731);
xnor U10222 (N_10222,N_8644,N_8696);
and U10223 (N_10223,N_8430,N_9656);
nand U10224 (N_10224,N_8830,N_9633);
nand U10225 (N_10225,N_8053,N_8437);
or U10226 (N_10226,N_8391,N_9795);
nand U10227 (N_10227,N_8765,N_8183);
nand U10228 (N_10228,N_8471,N_9655);
nand U10229 (N_10229,N_9304,N_8875);
or U10230 (N_10230,N_9734,N_9236);
and U10231 (N_10231,N_9265,N_9064);
and U10232 (N_10232,N_8314,N_9988);
nor U10233 (N_10233,N_8002,N_9895);
and U10234 (N_10234,N_9560,N_8506);
xor U10235 (N_10235,N_9452,N_8859);
nand U10236 (N_10236,N_8435,N_9094);
nand U10237 (N_10237,N_9149,N_9470);
xor U10238 (N_10238,N_9401,N_8311);
nand U10239 (N_10239,N_9805,N_9883);
or U10240 (N_10240,N_8533,N_9120);
nand U10241 (N_10241,N_8538,N_8383);
xor U10242 (N_10242,N_8732,N_8736);
and U10243 (N_10243,N_8355,N_9844);
and U10244 (N_10244,N_9889,N_9163);
nand U10245 (N_10245,N_9888,N_8605);
and U10246 (N_10246,N_9436,N_9465);
nor U10247 (N_10247,N_9574,N_8260);
xor U10248 (N_10248,N_8699,N_8162);
nand U10249 (N_10249,N_9782,N_8901);
xnor U10250 (N_10250,N_9631,N_8639);
or U10251 (N_10251,N_8045,N_8931);
or U10252 (N_10252,N_9305,N_8211);
nor U10253 (N_10253,N_8189,N_9724);
and U10254 (N_10254,N_9356,N_8828);
or U10255 (N_10255,N_8888,N_8171);
xnor U10256 (N_10256,N_8871,N_8161);
nand U10257 (N_10257,N_9244,N_8502);
nor U10258 (N_10258,N_9652,N_9425);
xnor U10259 (N_10259,N_8485,N_8360);
and U10260 (N_10260,N_8167,N_9141);
and U10261 (N_10261,N_8291,N_9164);
nand U10262 (N_10262,N_9413,N_8346);
and U10263 (N_10263,N_9287,N_9658);
nor U10264 (N_10264,N_8823,N_9367);
or U10265 (N_10265,N_9264,N_9580);
nand U10266 (N_10266,N_8349,N_8195);
xnor U10267 (N_10267,N_8357,N_9281);
or U10268 (N_10268,N_8625,N_8184);
nand U10269 (N_10269,N_8254,N_8866);
nor U10270 (N_10270,N_9211,N_8637);
or U10271 (N_10271,N_9421,N_9538);
and U10272 (N_10272,N_8436,N_8479);
nor U10273 (N_10273,N_9477,N_9242);
nor U10274 (N_10274,N_9696,N_8230);
xnor U10275 (N_10275,N_9238,N_9223);
or U10276 (N_10276,N_9376,N_9581);
or U10277 (N_10277,N_9824,N_9273);
and U10278 (N_10278,N_9240,N_8078);
xor U10279 (N_10279,N_8200,N_9052);
nand U10280 (N_10280,N_8272,N_8872);
and U10281 (N_10281,N_8729,N_9645);
xor U10282 (N_10282,N_8181,N_9523);
nor U10283 (N_10283,N_8606,N_9166);
nand U10284 (N_10284,N_8452,N_8453);
or U10285 (N_10285,N_9469,N_8916);
xnor U10286 (N_10286,N_9373,N_9159);
or U10287 (N_10287,N_8848,N_8723);
xor U10288 (N_10288,N_8631,N_9982);
or U10289 (N_10289,N_9378,N_8961);
xor U10290 (N_10290,N_9209,N_8345);
nand U10291 (N_10291,N_8634,N_9248);
nand U10292 (N_10292,N_8472,N_9927);
and U10293 (N_10293,N_8135,N_9377);
xnor U10294 (N_10294,N_8043,N_9772);
xnor U10295 (N_10295,N_9350,N_9733);
and U10296 (N_10296,N_8255,N_9293);
and U10297 (N_10297,N_8813,N_9391);
nor U10298 (N_10298,N_9178,N_8635);
and U10299 (N_10299,N_9228,N_9371);
or U10300 (N_10300,N_9096,N_8281);
or U10301 (N_10301,N_8320,N_8102);
and U10302 (N_10302,N_8492,N_8077);
and U10303 (N_10303,N_8434,N_8903);
or U10304 (N_10304,N_8802,N_9550);
xnor U10305 (N_10305,N_9830,N_9545);
or U10306 (N_10306,N_9583,N_8402);
nand U10307 (N_10307,N_8385,N_8042);
xnor U10308 (N_10308,N_9985,N_8651);
nand U10309 (N_10309,N_8274,N_9601);
nor U10310 (N_10310,N_9970,N_9018);
or U10311 (N_10311,N_8243,N_8837);
nor U10312 (N_10312,N_8934,N_9482);
and U10313 (N_10313,N_8168,N_8930);
nand U10314 (N_10314,N_8772,N_8075);
xor U10315 (N_10315,N_8851,N_8036);
nor U10316 (N_10316,N_8040,N_9194);
nor U10317 (N_10317,N_9622,N_8516);
xor U10318 (N_10318,N_8438,N_8978);
nor U10319 (N_10319,N_9270,N_8719);
and U10320 (N_10320,N_8414,N_9987);
and U10321 (N_10321,N_8390,N_9118);
or U10322 (N_10322,N_9774,N_9919);
nand U10323 (N_10323,N_8407,N_8570);
nor U10324 (N_10324,N_8667,N_9940);
xor U10325 (N_10325,N_8397,N_9647);
or U10326 (N_10326,N_9767,N_8751);
or U10327 (N_10327,N_9311,N_9387);
xnor U10328 (N_10328,N_9122,N_8187);
nand U10329 (N_10329,N_8617,N_9381);
xnor U10330 (N_10330,N_8838,N_8339);
nor U10331 (N_10331,N_8422,N_8997);
or U10332 (N_10332,N_8902,N_9263);
or U10333 (N_10333,N_9517,N_9113);
nor U10334 (N_10334,N_9546,N_9925);
nand U10335 (N_10335,N_9245,N_8019);
nand U10336 (N_10336,N_9716,N_9942);
xor U10337 (N_10337,N_8404,N_8764);
or U10338 (N_10338,N_8642,N_8347);
or U10339 (N_10339,N_8371,N_8303);
and U10340 (N_10340,N_8656,N_8622);
and U10341 (N_10341,N_9624,N_9961);
xor U10342 (N_10342,N_8316,N_9370);
or U10343 (N_10343,N_9333,N_8885);
or U10344 (N_10344,N_8064,N_8327);
xnor U10345 (N_10345,N_8873,N_8577);
nor U10346 (N_10346,N_9137,N_8588);
nand U10347 (N_10347,N_8082,N_9650);
nand U10348 (N_10348,N_9641,N_9344);
nand U10349 (N_10349,N_9769,N_8094);
and U10350 (N_10350,N_9936,N_8527);
nor U10351 (N_10351,N_8565,N_9078);
or U10352 (N_10352,N_8968,N_9341);
and U10353 (N_10353,N_8722,N_9338);
nor U10354 (N_10354,N_8367,N_8956);
nor U10355 (N_10355,N_8524,N_9665);
or U10356 (N_10356,N_8014,N_8553);
nor U10357 (N_10357,N_9234,N_9729);
or U10358 (N_10358,N_9775,N_8223);
and U10359 (N_10359,N_9715,N_8680);
nor U10360 (N_10360,N_8419,N_8008);
or U10361 (N_10361,N_9913,N_9582);
and U10362 (N_10362,N_8201,N_9612);
nor U10363 (N_10363,N_8549,N_8972);
xor U10364 (N_10364,N_9978,N_9933);
nor U10365 (N_10365,N_8865,N_8460);
or U10366 (N_10366,N_8522,N_9092);
xnor U10367 (N_10367,N_8803,N_9365);
and U10368 (N_10368,N_9901,N_8491);
nor U10369 (N_10369,N_9819,N_9001);
xor U10370 (N_10370,N_9067,N_9599);
xor U10371 (N_10371,N_8672,N_8498);
or U10372 (N_10372,N_8388,N_8417);
or U10373 (N_10373,N_9246,N_9831);
or U10374 (N_10374,N_8362,N_9890);
nor U10375 (N_10375,N_9267,N_8566);
nand U10376 (N_10376,N_9463,N_9764);
and U10377 (N_10377,N_9167,N_9471);
and U10378 (N_10378,N_9154,N_9649);
and U10379 (N_10379,N_8134,N_9123);
nor U10380 (N_10380,N_8596,N_9481);
xor U10381 (N_10381,N_8279,N_9713);
nand U10382 (N_10382,N_9634,N_8800);
nor U10383 (N_10383,N_9867,N_9181);
nand U10384 (N_10384,N_9814,N_8970);
xor U10385 (N_10385,N_9229,N_9457);
or U10386 (N_10386,N_8985,N_9521);
nand U10387 (N_10387,N_9404,N_9553);
and U10388 (N_10388,N_9085,N_8579);
and U10389 (N_10389,N_9458,N_9974);
or U10390 (N_10390,N_9009,N_9886);
nand U10391 (N_10391,N_8336,N_9374);
and U10392 (N_10392,N_9200,N_9252);
nor U10393 (N_10393,N_9654,N_9207);
or U10394 (N_10394,N_8746,N_8443);
and U10395 (N_10395,N_9024,N_9700);
or U10396 (N_10396,N_8610,N_8071);
and U10397 (N_10397,N_9105,N_8713);
nor U10398 (N_10398,N_8868,N_8454);
and U10399 (N_10399,N_8199,N_9313);
or U10400 (N_10400,N_8483,N_8805);
or U10401 (N_10401,N_9853,N_9884);
nor U10402 (N_10402,N_9617,N_8425);
or U10403 (N_10403,N_8212,N_9849);
and U10404 (N_10404,N_9191,N_8822);
xnor U10405 (N_10405,N_8324,N_8106);
xor U10406 (N_10406,N_8061,N_8246);
nand U10407 (N_10407,N_9578,N_8572);
and U10408 (N_10408,N_9964,N_9828);
xor U10409 (N_10409,N_8006,N_8451);
or U10410 (N_10410,N_8661,N_9500);
and U10411 (N_10411,N_8507,N_8537);
xor U10412 (N_10412,N_9005,N_8191);
nand U10413 (N_10413,N_8811,N_8820);
xnor U10414 (N_10414,N_8880,N_9498);
xnor U10415 (N_10415,N_9036,N_8048);
nor U10416 (N_10416,N_8335,N_8401);
and U10417 (N_10417,N_9271,N_9677);
xor U10418 (N_10418,N_9444,N_8289);
or U10419 (N_10419,N_8239,N_9754);
nand U10420 (N_10420,N_8188,N_9555);
xnor U10421 (N_10421,N_8403,N_9619);
nand U10422 (N_10422,N_9450,N_8323);
or U10423 (N_10423,N_8091,N_9508);
xnor U10424 (N_10424,N_9566,N_8580);
nand U10425 (N_10425,N_8332,N_8059);
and U10426 (N_10426,N_9258,N_9923);
nor U10427 (N_10427,N_8887,N_8295);
nand U10428 (N_10428,N_9629,N_9347);
and U10429 (N_10429,N_9594,N_9635);
nand U10430 (N_10430,N_9213,N_9692);
or U10431 (N_10431,N_8341,N_8653);
or U10432 (N_10432,N_9345,N_9561);
nor U10433 (N_10433,N_9334,N_8817);
xnor U10434 (N_10434,N_8216,N_8133);
nor U10435 (N_10435,N_8495,N_9763);
or U10436 (N_10436,N_9675,N_9968);
xor U10437 (N_10437,N_9033,N_9168);
or U10438 (N_10438,N_9195,N_9598);
nand U10439 (N_10439,N_8757,N_9717);
nor U10440 (N_10440,N_9648,N_8911);
xnor U10441 (N_10441,N_8431,N_9506);
and U10442 (N_10442,N_9991,N_9235);
nor U10443 (N_10443,N_9676,N_8056);
nor U10444 (N_10444,N_8669,N_8703);
or U10445 (N_10445,N_9409,N_9869);
or U10446 (N_10446,N_8551,N_8897);
and U10447 (N_10447,N_8850,N_9585);
or U10448 (N_10448,N_8475,N_9745);
nor U10449 (N_10449,N_9372,N_8938);
xor U10450 (N_10450,N_9902,N_8238);
and U10451 (N_10451,N_9097,N_8735);
or U10452 (N_10452,N_9300,N_9630);
and U10453 (N_10453,N_8949,N_9801);
or U10454 (N_10454,N_8649,N_8179);
xnor U10455 (N_10455,N_8290,N_9723);
or U10456 (N_10456,N_9567,N_8379);
or U10457 (N_10457,N_8905,N_9153);
nand U10458 (N_10458,N_9687,N_9659);
and U10459 (N_10459,N_9799,N_9984);
xor U10460 (N_10460,N_8594,N_8790);
xnor U10461 (N_10461,N_8619,N_8744);
or U10462 (N_10462,N_9921,N_9949);
or U10463 (N_10463,N_8231,N_8750);
and U10464 (N_10464,N_8708,N_9564);
xor U10465 (N_10465,N_9368,N_9056);
nand U10466 (N_10466,N_8616,N_9803);
nor U10467 (N_10467,N_9778,N_9225);
or U10468 (N_10468,N_9904,N_8465);
nor U10469 (N_10469,N_9397,N_8798);
and U10470 (N_10470,N_9479,N_8900);
nor U10471 (N_10471,N_9266,N_8251);
or U10472 (N_10472,N_9972,N_9918);
or U10473 (N_10473,N_8143,N_8697);
nor U10474 (N_10474,N_8282,N_8636);
or U10475 (N_10475,N_8400,N_8763);
nor U10476 (N_10476,N_9494,N_8180);
nand U10477 (N_10477,N_9416,N_9331);
xnor U10478 (N_10478,N_9473,N_9593);
and U10479 (N_10479,N_9541,N_8954);
and U10480 (N_10480,N_8989,N_9903);
nor U10481 (N_10481,N_8627,N_9924);
xnor U10482 (N_10482,N_8057,N_8157);
or U10483 (N_10483,N_8392,N_8093);
xor U10484 (N_10484,N_8114,N_9237);
or U10485 (N_10485,N_8470,N_9420);
and U10486 (N_10486,N_9584,N_9596);
or U10487 (N_10487,N_9464,N_8988);
or U10488 (N_10488,N_8450,N_9335);
or U10489 (N_10489,N_8922,N_9771);
or U10490 (N_10490,N_9806,N_9993);
xnor U10491 (N_10491,N_9976,N_9822);
nand U10492 (N_10492,N_9443,N_9189);
and U10493 (N_10493,N_8182,N_8128);
or U10494 (N_10494,N_9003,N_9462);
nor U10495 (N_10495,N_9106,N_8879);
xnor U10496 (N_10496,N_8287,N_8361);
or U10497 (N_10497,N_8264,N_8794);
and U10498 (N_10498,N_9938,N_9059);
or U10499 (N_10499,N_9071,N_8234);
xnor U10500 (N_10500,N_8971,N_9487);
nand U10501 (N_10501,N_8845,N_8726);
or U10502 (N_10502,N_8149,N_8073);
xnor U10503 (N_10503,N_8378,N_9354);
and U10504 (N_10504,N_9289,N_9548);
or U10505 (N_10505,N_8208,N_9827);
or U10506 (N_10506,N_8284,N_9953);
and U10507 (N_10507,N_9736,N_8070);
xnor U10508 (N_10508,N_9040,N_8993);
xor U10509 (N_10509,N_8177,N_8777);
and U10510 (N_10510,N_9908,N_9807);
nand U10511 (N_10511,N_8384,N_9053);
xnor U10512 (N_10512,N_9607,N_9353);
or U10513 (N_10513,N_8597,N_9456);
and U10514 (N_10514,N_9428,N_8307);
nand U10515 (N_10515,N_8690,N_9069);
xor U10516 (N_10516,N_8919,N_8169);
xnor U10517 (N_10517,N_9007,N_9221);
nand U10518 (N_10518,N_8991,N_9058);
nor U10519 (N_10519,N_8564,N_9680);
nand U10520 (N_10520,N_9892,N_9710);
nor U10521 (N_10521,N_8039,N_8309);
xor U10522 (N_10522,N_9862,N_8152);
or U10523 (N_10523,N_9547,N_9917);
or U10524 (N_10524,N_8276,N_9996);
or U10525 (N_10525,N_9326,N_9336);
nor U10526 (N_10526,N_8468,N_8981);
and U10527 (N_10527,N_9572,N_8626);
xor U10528 (N_10528,N_8085,N_8665);
and U10529 (N_10529,N_8484,N_8456);
nand U10530 (N_10530,N_8518,N_9488);
and U10531 (N_10531,N_9130,N_9330);
or U10532 (N_10532,N_8869,N_8965);
nor U10533 (N_10533,N_8692,N_9626);
nand U10534 (N_10534,N_8515,N_8592);
or U10535 (N_10535,N_8535,N_8792);
nand U10536 (N_10536,N_9502,N_9398);
or U10537 (N_10537,N_9632,N_9131);
xor U10538 (N_10538,N_9306,N_8607);
xnor U10539 (N_10539,N_8337,N_9671);
or U10540 (N_10540,N_8262,N_8317);
nor U10541 (N_10541,N_9180,N_8469);
xnor U10542 (N_10542,N_9366,N_9614);
and U10543 (N_10543,N_9535,N_8707);
or U10544 (N_10544,N_9544,N_9708);
and U10545 (N_10545,N_8165,N_8826);
and U10546 (N_10546,N_9531,N_9089);
nor U10547 (N_10547,N_8645,N_9162);
nand U10548 (N_10548,N_9726,N_9017);
nand U10549 (N_10549,N_9016,N_9101);
nor U10550 (N_10550,N_8090,N_8578);
nor U10551 (N_10551,N_8587,N_8657);
xor U10552 (N_10552,N_8236,N_8017);
or U10553 (N_10553,N_9255,N_8745);
xnor U10554 (N_10554,N_9794,N_9355);
nand U10555 (N_10555,N_9990,N_9691);
nor U10556 (N_10556,N_9046,N_9914);
or U10557 (N_10557,N_8222,N_9013);
nand U10558 (N_10558,N_9272,N_9247);
or U10559 (N_10559,N_9610,N_9277);
xnor U10560 (N_10560,N_9780,N_8771);
or U10561 (N_10561,N_8918,N_8921);
nor U10562 (N_10562,N_8297,N_9400);
nor U10563 (N_10563,N_8912,N_9100);
nand U10564 (N_10564,N_9346,N_9301);
or U10565 (N_10565,N_8205,N_8788);
nand U10566 (N_10566,N_8663,N_9956);
xnor U10567 (N_10567,N_8051,N_8947);
nor U10568 (N_10568,N_8427,N_9851);
nand U10569 (N_10569,N_9408,N_8769);
or U10570 (N_10570,N_9510,N_9699);
nor U10571 (N_10571,N_9836,N_8804);
or U10572 (N_10572,N_8050,N_9820);
nand U10573 (N_10573,N_9646,N_8441);
or U10574 (N_10574,N_8529,N_9727);
xnor U10575 (N_10575,N_9399,N_9262);
xor U10576 (N_10576,N_8904,N_9431);
xor U10577 (N_10577,N_8748,N_8069);
or U10578 (N_10578,N_9759,N_9768);
xnor U10579 (N_10579,N_9302,N_9628);
and U10580 (N_10580,N_9480,N_9590);
xnor U10581 (N_10581,N_8862,N_9870);
xor U10582 (N_10582,N_8629,N_9857);
nor U10583 (N_10583,N_8691,N_9922);
nor U10584 (N_10584,N_9707,N_8312);
nand U10585 (N_10585,N_8514,N_9520);
nand U10586 (N_10586,N_8832,N_9132);
nor U10587 (N_10587,N_9948,N_8807);
or U10588 (N_10588,N_9010,N_9798);
and U10589 (N_10589,N_9747,N_9615);
or U10590 (N_10590,N_9823,N_8752);
and U10591 (N_10591,N_8298,N_9057);
and U10592 (N_10592,N_8909,N_8001);
and U10593 (N_10593,N_8677,N_8914);
or U10594 (N_10594,N_9847,N_8322);
and U10595 (N_10595,N_8018,N_8638);
nand U10596 (N_10596,N_9296,N_8455);
nand U10597 (N_10597,N_8967,N_8060);
nand U10598 (N_10598,N_8261,N_8944);
or U10599 (N_10599,N_8547,N_8560);
and U10600 (N_10600,N_9643,N_8466);
xnor U10601 (N_10601,N_8825,N_8783);
and U10602 (N_10602,N_8153,N_9789);
and U10603 (N_10603,N_8097,N_9573);
and U10604 (N_10604,N_8003,N_8863);
xnor U10605 (N_10605,N_9442,N_9693);
nand U10606 (N_10606,N_9087,N_9004);
xor U10607 (N_10607,N_8503,N_8013);
nand U10608 (N_10608,N_9514,N_9362);
xnor U10609 (N_10609,N_8387,N_9015);
xor U10610 (N_10610,N_9427,N_8305);
nor U10611 (N_10611,N_9511,N_8363);
and U10612 (N_10612,N_8760,N_8123);
or U10613 (N_10613,N_9028,N_8688);
and U10614 (N_10614,N_8686,N_9251);
or U10615 (N_10615,N_9073,N_8782);
nor U10616 (N_10616,N_9663,N_9711);
nand U10617 (N_10617,N_8590,N_9491);
nand U10618 (N_10618,N_9743,N_8100);
and U10619 (N_10619,N_8689,N_9241);
and U10620 (N_10620,N_8365,N_8462);
xnor U10621 (N_10621,N_8185,N_8130);
nor U10622 (N_10622,N_8217,N_9226);
nor U10623 (N_10623,N_9486,N_8150);
or U10624 (N_10624,N_8105,N_8562);
nand U10625 (N_10625,N_9539,N_9369);
or U10626 (N_10626,N_9280,N_8948);
xnor U10627 (N_10627,N_8992,N_8854);
and U10628 (N_10628,N_8561,N_9386);
nand U10629 (N_10629,N_8342,N_9796);
nor U10630 (N_10630,N_9672,N_8720);
xor U10631 (N_10631,N_9571,N_9910);
or U10632 (N_10632,N_8785,N_9020);
or U10633 (N_10633,N_8343,N_9383);
or U10634 (N_10634,N_9689,N_9299);
and U10635 (N_10635,N_8159,N_8095);
nor U10636 (N_10636,N_8531,N_8776);
nand U10637 (N_10637,N_8306,N_8983);
nand U10638 (N_10638,N_8893,N_8215);
nand U10639 (N_10639,N_9329,N_8550);
nor U10640 (N_10640,N_8166,N_9045);
and U10641 (N_10641,N_8841,N_9623);
and U10642 (N_10642,N_9414,N_8121);
or U10643 (N_10643,N_8233,N_8074);
nor U10644 (N_10644,N_9109,N_9620);
or U10645 (N_10645,N_9074,N_9735);
or U10646 (N_10646,N_8092,N_8099);
or U10647 (N_10647,N_9840,N_8192);
and U10648 (N_10648,N_8232,N_9125);
nand U10649 (N_10649,N_9749,N_8406);
xnor U10650 (N_10650,N_8271,N_8519);
nand U10651 (N_10651,N_9882,N_8247);
or U10652 (N_10652,N_8601,N_8718);
nand U10653 (N_10653,N_9099,N_9911);
nor U10654 (N_10654,N_9288,N_8292);
xnor U10655 (N_10655,N_8476,N_9084);
nand U10656 (N_10656,N_8660,N_8325);
nor U10657 (N_10657,N_9719,N_9960);
nor U10658 (N_10658,N_9190,N_8389);
nor U10659 (N_10659,N_8278,N_8544);
xnor U10660 (N_10660,N_8115,N_8398);
xor U10661 (N_10661,N_8252,N_9138);
xnor U10662 (N_10662,N_9283,N_9916);
nor U10663 (N_10663,N_8328,N_9278);
xnor U10664 (N_10664,N_9791,N_9014);
nand U10665 (N_10665,N_9434,N_9424);
xnor U10666 (N_10666,N_9563,N_9874);
nor U10667 (N_10667,N_8494,N_8065);
and U10668 (N_10668,N_9268,N_8674);
or U10669 (N_10669,N_8136,N_8509);
nor U10670 (N_10670,N_8810,N_9187);
nand U10671 (N_10671,N_8668,N_9188);
nor U10672 (N_10672,N_8241,N_9714);
and U10673 (N_10673,N_8025,N_8172);
xor U10674 (N_10674,N_9405,N_9215);
xor U10675 (N_10675,N_8315,N_9838);
xnor U10676 (N_10676,N_9793,N_9034);
nor U10677 (N_10677,N_8721,N_9030);
nor U10678 (N_10678,N_8420,N_9134);
and U10679 (N_10679,N_9418,N_8489);
or U10680 (N_10680,N_8294,N_9750);
nor U10681 (N_10681,N_8068,N_9597);
nor U10682 (N_10682,N_8490,N_9722);
or U10683 (N_10683,N_8882,N_8542);
nand U10684 (N_10684,N_8749,N_8521);
xor U10685 (N_10685,N_8975,N_9088);
or U10686 (N_10686,N_9528,N_8943);
or U10687 (N_10687,N_8210,N_9351);
or U10688 (N_10688,N_9395,N_8609);
xnor U10689 (N_10689,N_9896,N_8107);
xnor U10690 (N_10690,N_8052,N_8024);
or U10691 (N_10691,N_8939,N_9038);
and U10692 (N_10692,N_9360,N_9135);
nand U10693 (N_10693,N_8818,N_8329);
and U10694 (N_10694,N_9737,N_8762);
nor U10695 (N_10695,N_9385,N_8352);
nor U10696 (N_10696,N_8032,N_8301);
nand U10697 (N_10697,N_9706,N_9144);
and U10698 (N_10698,N_8917,N_8602);
xnor U10699 (N_10699,N_8209,N_9308);
xor U10700 (N_10700,N_9954,N_8824);
or U10701 (N_10701,N_9962,N_8029);
nor U10702 (N_10702,N_8695,N_8941);
xnor U10703 (N_10703,N_9364,N_8808);
xor U10704 (N_10704,N_9446,N_8447);
nor U10705 (N_10705,N_9834,N_9216);
or U10706 (N_10706,N_9152,N_9979);
nor U10707 (N_10707,N_8864,N_9559);
nor U10708 (N_10708,N_9666,N_8194);
or U10709 (N_10709,N_8374,N_9950);
xnor U10710 (N_10710,N_8999,N_9496);
or U10711 (N_10711,N_8087,N_8148);
nor U10712 (N_10712,N_9128,N_8928);
nand U10713 (N_10713,N_9945,N_9766);
nor U10714 (N_10714,N_8780,N_8849);
xnor U10715 (N_10715,N_8611,N_9992);
xor U10716 (N_10716,N_9657,N_8728);
or U10717 (N_10717,N_9291,N_9332);
or U10718 (N_10718,N_9720,N_9061);
nand U10719 (N_10719,N_8375,N_9025);
or U10720 (N_10720,N_8204,N_9172);
xnor U10721 (N_10721,N_9361,N_9359);
and U10722 (N_10722,N_8319,N_8867);
nand U10723 (N_10723,N_8556,N_8283);
or U10724 (N_10724,N_8962,N_9192);
or U10725 (N_10725,N_8258,N_8781);
nor U10726 (N_10726,N_9705,N_8288);
or U10727 (N_10727,N_8101,N_9489);
xnor U10728 (N_10728,N_9878,N_8005);
and U10729 (N_10729,N_8936,N_8058);
and U10730 (N_10730,N_9957,N_9568);
nor U10731 (N_10731,N_8063,N_8612);
nor U10732 (N_10732,N_9206,N_8158);
or U10733 (N_10733,N_8457,N_8016);
xor U10734 (N_10734,N_8557,N_9698);
xnor U10735 (N_10735,N_9415,N_8990);
xor U10736 (N_10736,N_9314,N_9829);
and U10737 (N_10737,N_8122,N_8510);
nor U10738 (N_10738,N_9147,N_8423);
nand U10739 (N_10739,N_9589,N_8821);
xnor U10740 (N_10740,N_9905,N_9684);
or U10741 (N_10741,N_8937,N_9558);
xor U10742 (N_10742,N_9501,N_9454);
or U10743 (N_10743,N_9800,N_8377);
xnor U10744 (N_10744,N_9503,N_9943);
xor U10745 (N_10745,N_8112,N_9611);
and U10746 (N_10746,N_9740,N_9947);
or U10747 (N_10747,N_8603,N_8724);
nand U10748 (N_10748,N_8898,N_8142);
nand U10749 (N_10749,N_9474,N_9516);
nor U10750 (N_10750,N_9579,N_8986);
nor U10751 (N_10751,N_9080,N_9158);
nor U10752 (N_10752,N_9813,N_9179);
xnor U10753 (N_10753,N_8226,N_9746);
or U10754 (N_10754,N_8237,N_8784);
and U10755 (N_10755,N_8839,N_9066);
nand U10756 (N_10756,N_8737,N_9055);
or U10757 (N_10757,N_9432,N_8976);
xnor U10758 (N_10758,N_9440,N_8256);
or U10759 (N_10759,N_9703,N_8015);
xnor U10760 (N_10760,N_8681,N_8712);
xor U10761 (N_10761,N_9103,N_8227);
and U10762 (N_10762,N_8229,N_8786);
nor U10763 (N_10763,N_9231,N_8946);
nand U10764 (N_10764,N_9505,N_9543);
or U10765 (N_10765,N_9757,N_8047);
and U10766 (N_10766,N_8643,N_8584);
nand U10767 (N_10767,N_9997,N_9438);
and U10768 (N_10768,N_8117,N_9199);
or U10769 (N_10769,N_9817,N_8666);
nand U10770 (N_10770,N_9932,N_8621);
and U10771 (N_10771,N_8835,N_8641);
nor U10772 (N_10772,N_8925,N_9322);
and U10773 (N_10773,N_8600,N_8020);
and U10774 (N_10774,N_8889,N_8933);
and U10775 (N_10775,N_9070,N_9679);
and U10776 (N_10776,N_9777,N_9183);
or U10777 (N_10777,N_9871,N_8370);
nor U10778 (N_10778,N_9176,N_8411);
or U10779 (N_10779,N_8331,N_8049);
and U10780 (N_10780,N_9821,N_9382);
xnor U10781 (N_10781,N_9449,N_9792);
or U10782 (N_10782,N_8840,N_8987);
nand U10783 (N_10783,N_9303,N_8613);
nor U10784 (N_10784,N_8220,N_9127);
and U10785 (N_10785,N_8801,N_9788);
xnor U10786 (N_10786,N_8787,N_8273);
xnor U10787 (N_10787,N_9394,N_8571);
nor U10788 (N_10788,N_8567,N_9525);
nor U10789 (N_10789,N_8861,N_8742);
and U10790 (N_10790,N_9392,N_9907);
and U10791 (N_10791,N_9732,N_9294);
nand U10792 (N_10792,N_9129,N_9119);
xnor U10793 (N_10793,N_9618,N_9460);
or U10794 (N_10794,N_9044,N_8338);
nand U10795 (N_10795,N_8413,N_8539);
nor U10796 (N_10796,N_9143,N_8214);
xnor U10797 (N_10797,N_9062,N_8853);
and U10798 (N_10798,N_8359,N_9447);
nor U10799 (N_10799,N_8770,N_9290);
or U10800 (N_10800,N_9208,N_9256);
nor U10801 (N_10801,N_9165,N_8806);
and U10802 (N_10802,N_8878,N_8372);
and U10803 (N_10803,N_9891,N_9810);
and U10804 (N_10804,N_8221,N_9259);
and U10805 (N_10805,N_8715,N_9388);
xor U10806 (N_10806,N_8086,N_8678);
nor U10807 (N_10807,N_9193,N_9753);
or U10808 (N_10808,N_9669,N_9286);
or U10809 (N_10809,N_9797,N_9316);
nor U10810 (N_10810,N_9276,N_9685);
or U10811 (N_10811,N_9845,N_9499);
nor U10812 (N_10812,N_8847,N_8920);
or U10813 (N_10813,N_9050,N_9093);
nand U10814 (N_10814,N_8526,N_9887);
or U10815 (N_10815,N_8977,N_9279);
and U10816 (N_10816,N_9688,N_8701);
or U10817 (N_10817,N_9973,N_9429);
or U10818 (N_10818,N_9095,N_8650);
nand U10819 (N_10819,N_9551,N_9946);
nor U10820 (N_10820,N_8170,N_9384);
and U10821 (N_10821,N_8084,N_8415);
and U10822 (N_10822,N_9540,N_9587);
nand U10823 (N_10823,N_8907,N_8055);
or U10824 (N_10824,N_8154,N_8369);
nor U10825 (N_10825,N_8836,N_9565);
xnor U10826 (N_10826,N_9484,N_8574);
nor U10827 (N_10827,N_9877,N_8421);
or U10828 (N_10828,N_8513,N_9533);
or U10829 (N_10829,N_9575,N_8540);
nor U10830 (N_10830,N_8027,N_9075);
xor U10831 (N_10831,N_9349,N_9342);
nor U10832 (N_10832,N_9576,N_9363);
and U10833 (N_10833,N_9317,N_9417);
or U10834 (N_10834,N_8891,N_9781);
or U10835 (N_10835,N_8364,N_8952);
nor U10836 (N_10836,N_9041,N_9230);
and U10837 (N_10837,N_9808,N_8011);
or U10838 (N_10838,N_8555,N_8710);
or U10839 (N_10839,N_8405,N_8433);
and U10840 (N_10840,N_8299,N_9307);
xor U10841 (N_10841,N_8118,N_8844);
or U10842 (N_10842,N_9210,N_9076);
nand U10843 (N_10843,N_9731,N_9758);
or U10844 (N_10844,N_9475,N_9197);
or U10845 (N_10845,N_9920,N_9002);
or U10846 (N_10846,N_8031,N_8951);
nand U10847 (N_10847,N_8124,N_9865);
nand U10848 (N_10848,N_9653,N_8190);
xor U10849 (N_10849,N_9403,N_8225);
nand U10850 (N_10850,N_9185,N_9202);
or U10851 (N_10851,N_9748,N_8218);
nand U10852 (N_10852,N_9402,N_9108);
nand U10853 (N_10853,N_9146,N_9274);
nor U10854 (N_10854,N_8855,N_9642);
and U10855 (N_10855,N_9588,N_9876);
nor U10856 (N_10856,N_9437,N_9863);
nor U10857 (N_10857,N_8478,N_9048);
nand U10858 (N_10858,N_9285,N_9430);
nor U10859 (N_10859,N_9472,N_8739);
nand U10860 (N_10860,N_8791,N_8754);
and U10861 (N_10861,N_9243,N_8693);
xnor U10862 (N_10862,N_9701,N_8819);
and U10863 (N_10863,N_9855,N_8113);
nand U10864 (N_10864,N_8906,N_9941);
nor U10865 (N_10865,N_8618,N_9667);
or U10866 (N_10866,N_9605,N_9339);
nand U10867 (N_10867,N_8497,N_9818);
nor U10868 (N_10868,N_9804,N_8444);
and U10869 (N_10869,N_9868,N_8525);
xor U10870 (N_10870,N_8110,N_8589);
nor U10871 (N_10871,N_8717,N_9556);
nor U10872 (N_10872,N_9637,N_8213);
and U10873 (N_10873,N_8995,N_8809);
xnor U10874 (N_10874,N_9686,N_9627);
and U10875 (N_10875,N_9744,N_8098);
and U10876 (N_10876,N_9072,N_8354);
and U10877 (N_10877,N_9842,N_9324);
or U10878 (N_10878,N_8683,N_9536);
xnor U10879 (N_10879,N_8054,N_8892);
nand U10880 (N_10880,N_9049,N_9873);
xor U10881 (N_10881,N_9490,N_8499);
and U10882 (N_10882,N_8285,N_9466);
and U10883 (N_10883,N_8344,N_8138);
xnor U10884 (N_10884,N_9741,N_9340);
or U10885 (N_10885,N_8263,N_9909);
nand U10886 (N_10886,N_8033,N_9613);
and U10887 (N_10887,N_9406,N_9086);
nand U10888 (N_10888,N_8694,N_9433);
or U10889 (N_10889,N_8955,N_9738);
nor U10890 (N_10890,N_8163,N_9343);
and U10891 (N_10891,N_9476,N_9861);
nor U10892 (N_10892,N_8829,N_9173);
nand U10893 (N_10893,N_8340,N_9203);
nor U10894 (N_10894,N_8505,N_8685);
or U10895 (N_10895,N_8265,N_8129);
xor U10896 (N_10896,N_9983,N_9114);
and U10897 (N_10897,N_8481,N_9227);
nand U10898 (N_10898,N_8206,N_8730);
nand U10899 (N_10899,N_8585,N_8700);
nor U10900 (N_10900,N_8620,N_8270);
nor U10901 (N_10901,N_9393,N_8632);
or U10902 (N_10902,N_8756,N_9725);
xnor U10903 (N_10903,N_9198,N_9562);
or U10904 (N_10904,N_9526,N_9944);
or U10905 (N_10905,N_9850,N_8957);
and U10906 (N_10906,N_8523,N_9752);
or U10907 (N_10907,N_9021,N_9812);
nor U10908 (N_10908,N_8860,N_9930);
xor U10909 (N_10909,N_8141,N_9971);
nor U10910 (N_10910,N_8741,N_8432);
or U10911 (N_10911,N_9826,N_9981);
or U10912 (N_10912,N_8412,N_9011);
xnor U10913 (N_10913,N_9899,N_8662);
and U10914 (N_10914,N_8111,N_8767);
nand U10915 (N_10915,N_8910,N_9081);
and U10916 (N_10916,N_8277,N_9880);
nor U10917 (N_10917,N_8440,N_9148);
and U10918 (N_10918,N_9837,N_8321);
or U10919 (N_10919,N_9117,N_8982);
xnor U10920 (N_10920,N_8351,N_9031);
nand U10921 (N_10921,N_9694,N_9461);
xnor U10922 (N_10922,N_9249,N_8796);
nand U10923 (N_10923,N_8501,N_9595);
and U10924 (N_10924,N_8942,N_9881);
xor U10925 (N_10925,N_8308,N_9319);
nor U10926 (N_10926,N_8473,N_8240);
nor U10927 (N_10927,N_8242,N_9934);
and U10928 (N_10928,N_8545,N_9019);
nor U10929 (N_10929,N_9037,N_8640);
nand U10930 (N_10930,N_8409,N_8698);
or U10931 (N_10931,N_8381,N_9549);
xnor U10932 (N_10932,N_8196,N_8980);
nand U10933 (N_10933,N_8012,N_8573);
or U10934 (N_10934,N_9312,N_9459);
and U10935 (N_10935,N_9065,N_8424);
or U10936 (N_10936,N_8467,N_8761);
and U10937 (N_10937,N_8386,N_8856);
or U10938 (N_10938,N_8160,N_8733);
or U10939 (N_10939,N_9102,N_8833);
nor U10940 (N_10940,N_9609,N_9770);
and U10941 (N_10941,N_8799,N_9670);
and U10942 (N_10942,N_9809,N_8591);
and U10943 (N_10943,N_9352,N_9337);
nand U10944 (N_10944,N_8734,N_9157);
and U10945 (N_10945,N_9445,N_8628);
xor U10946 (N_10946,N_8852,N_8877);
and U10947 (N_10947,N_8244,N_8583);
and U10948 (N_10948,N_8088,N_9224);
nor U10949 (N_10949,N_8915,N_9121);
xor U10950 (N_10950,N_8442,N_9182);
xnor U10951 (N_10951,N_9042,N_8630);
xor U10952 (N_10952,N_8633,N_8960);
nor U10953 (N_10953,N_9841,N_8702);
or U10954 (N_10954,N_8034,N_9150);
and U10955 (N_10955,N_9963,N_9790);
and U10956 (N_10956,N_8598,N_8253);
nand U10957 (N_10957,N_8530,N_9843);
nor U10958 (N_10958,N_9532,N_9327);
nand U10959 (N_10959,N_9513,N_9969);
nand U10960 (N_10960,N_8418,N_8857);
xnor U10961 (N_10961,N_8496,N_9897);
nand U10962 (N_10962,N_8753,N_8927);
nor U10963 (N_10963,N_8207,N_8546);
and U10964 (N_10964,N_8614,N_9485);
and U10965 (N_10965,N_9090,N_8487);
xor U10966 (N_10966,N_9787,N_9077);
xor U10967 (N_10967,N_8795,N_9527);
nand U10968 (N_10968,N_8350,N_8576);
nand U10969 (N_10969,N_9169,N_8709);
and U10970 (N_10970,N_9638,N_9142);
xor U10971 (N_10971,N_9051,N_8066);
and U10972 (N_10972,N_8924,N_9872);
or U10973 (N_10973,N_9063,N_8870);
xnor U10974 (N_10974,N_8081,N_8969);
nor U10975 (N_10975,N_8313,N_8998);
and U10976 (N_10976,N_9175,N_9110);
and U10977 (N_10977,N_9952,N_8738);
and U10978 (N_10978,N_8512,N_9928);
nor U10979 (N_10979,N_9915,N_8174);
and U10980 (N_10980,N_8144,N_9697);
nand U10981 (N_10981,N_9205,N_8773);
nor U10982 (N_10982,N_8973,N_9966);
nand U10983 (N_10983,N_8654,N_8137);
and U10984 (N_10984,N_9068,N_9730);
nor U10985 (N_10985,N_9879,N_8575);
xnor U10986 (N_10986,N_9497,N_8428);
or U10987 (N_10987,N_9083,N_8884);
and U10988 (N_10988,N_9519,N_8461);
xor U10989 (N_10989,N_8275,N_9435);
nor U10990 (N_10990,N_8429,N_8604);
and U10991 (N_10991,N_9269,N_9690);
xor U10992 (N_10992,N_8670,N_9492);
xnor U10993 (N_10993,N_9721,N_8679);
xnor U10994 (N_10994,N_9379,N_9054);
xor U10995 (N_10995,N_9592,N_8219);
and U10996 (N_10996,N_9310,N_9955);
nand U10997 (N_10997,N_8151,N_8706);
or U10998 (N_10998,N_8500,N_9825);
nand U10999 (N_10999,N_8714,N_8908);
and U11000 (N_11000,N_9451,N_9725);
nand U11001 (N_11001,N_9637,N_9989);
nor U11002 (N_11002,N_9127,N_8121);
nand U11003 (N_11003,N_8953,N_8530);
or U11004 (N_11004,N_8387,N_9930);
nand U11005 (N_11005,N_8500,N_8275);
nor U11006 (N_11006,N_8986,N_9030);
and U11007 (N_11007,N_9901,N_9335);
xnor U11008 (N_11008,N_8014,N_9164);
and U11009 (N_11009,N_9988,N_8052);
or U11010 (N_11010,N_9330,N_9452);
nand U11011 (N_11011,N_8928,N_9179);
xor U11012 (N_11012,N_8022,N_8476);
nand U11013 (N_11013,N_8993,N_9579);
nor U11014 (N_11014,N_8758,N_8129);
and U11015 (N_11015,N_8404,N_9285);
or U11016 (N_11016,N_8530,N_9577);
and U11017 (N_11017,N_8834,N_9767);
nand U11018 (N_11018,N_9992,N_9656);
or U11019 (N_11019,N_8572,N_9665);
nor U11020 (N_11020,N_8400,N_9505);
nand U11021 (N_11021,N_9020,N_8324);
and U11022 (N_11022,N_9674,N_9745);
or U11023 (N_11023,N_8496,N_8950);
and U11024 (N_11024,N_9643,N_8238);
or U11025 (N_11025,N_9941,N_8226);
and U11026 (N_11026,N_8250,N_8155);
xor U11027 (N_11027,N_9206,N_8448);
nand U11028 (N_11028,N_9596,N_8554);
or U11029 (N_11029,N_9682,N_8305);
and U11030 (N_11030,N_8986,N_8369);
xnor U11031 (N_11031,N_8416,N_9374);
nand U11032 (N_11032,N_8779,N_9057);
nor U11033 (N_11033,N_9689,N_8958);
nor U11034 (N_11034,N_8678,N_9795);
and U11035 (N_11035,N_9871,N_9755);
xnor U11036 (N_11036,N_8155,N_9237);
nor U11037 (N_11037,N_8094,N_8335);
and U11038 (N_11038,N_8718,N_8462);
xor U11039 (N_11039,N_9015,N_9649);
nor U11040 (N_11040,N_8472,N_9415);
or U11041 (N_11041,N_8332,N_9772);
and U11042 (N_11042,N_8690,N_9354);
or U11043 (N_11043,N_8105,N_9575);
xor U11044 (N_11044,N_9512,N_8497);
xnor U11045 (N_11045,N_9607,N_9687);
xnor U11046 (N_11046,N_8207,N_8243);
nor U11047 (N_11047,N_9812,N_9196);
or U11048 (N_11048,N_9658,N_9954);
or U11049 (N_11049,N_8021,N_9215);
or U11050 (N_11050,N_8172,N_9137);
and U11051 (N_11051,N_8198,N_8256);
nand U11052 (N_11052,N_8533,N_9544);
or U11053 (N_11053,N_8357,N_9490);
or U11054 (N_11054,N_8815,N_8349);
xnor U11055 (N_11055,N_8706,N_9296);
and U11056 (N_11056,N_8742,N_8803);
xnor U11057 (N_11057,N_9540,N_9507);
xor U11058 (N_11058,N_9437,N_9603);
or U11059 (N_11059,N_8384,N_9528);
xnor U11060 (N_11060,N_9805,N_9453);
xnor U11061 (N_11061,N_9653,N_9423);
or U11062 (N_11062,N_9290,N_9596);
or U11063 (N_11063,N_8276,N_8650);
xor U11064 (N_11064,N_9435,N_9178);
nand U11065 (N_11065,N_9422,N_9818);
nand U11066 (N_11066,N_8717,N_8557);
nor U11067 (N_11067,N_8314,N_8494);
nand U11068 (N_11068,N_8780,N_9802);
nor U11069 (N_11069,N_8404,N_8189);
nor U11070 (N_11070,N_8362,N_9283);
xnor U11071 (N_11071,N_9748,N_8388);
and U11072 (N_11072,N_9190,N_9899);
xor U11073 (N_11073,N_9803,N_9137);
or U11074 (N_11074,N_9526,N_8359);
xnor U11075 (N_11075,N_8381,N_9103);
or U11076 (N_11076,N_9891,N_8661);
or U11077 (N_11077,N_8239,N_8820);
xnor U11078 (N_11078,N_8950,N_8085);
nand U11079 (N_11079,N_9198,N_9405);
or U11080 (N_11080,N_8758,N_8941);
and U11081 (N_11081,N_8687,N_9901);
xor U11082 (N_11082,N_8077,N_8957);
xnor U11083 (N_11083,N_9366,N_9245);
and U11084 (N_11084,N_9363,N_9176);
and U11085 (N_11085,N_8380,N_9657);
xnor U11086 (N_11086,N_9785,N_8808);
and U11087 (N_11087,N_8890,N_9982);
nand U11088 (N_11088,N_8560,N_8982);
and U11089 (N_11089,N_9333,N_8349);
or U11090 (N_11090,N_8634,N_8785);
xor U11091 (N_11091,N_9381,N_8650);
nand U11092 (N_11092,N_8191,N_9779);
and U11093 (N_11093,N_9601,N_8527);
nor U11094 (N_11094,N_9781,N_9236);
nand U11095 (N_11095,N_9619,N_8793);
or U11096 (N_11096,N_9253,N_9339);
and U11097 (N_11097,N_9476,N_8871);
nor U11098 (N_11098,N_9727,N_9613);
and U11099 (N_11099,N_9011,N_9865);
or U11100 (N_11100,N_9974,N_9212);
nand U11101 (N_11101,N_9020,N_9918);
nor U11102 (N_11102,N_8333,N_9870);
xor U11103 (N_11103,N_8477,N_9994);
nand U11104 (N_11104,N_8888,N_8827);
or U11105 (N_11105,N_8149,N_9838);
nand U11106 (N_11106,N_9386,N_8459);
or U11107 (N_11107,N_9088,N_8364);
or U11108 (N_11108,N_9160,N_9723);
nand U11109 (N_11109,N_8079,N_8676);
nor U11110 (N_11110,N_9758,N_8306);
nand U11111 (N_11111,N_8211,N_9315);
nor U11112 (N_11112,N_9310,N_9945);
xor U11113 (N_11113,N_9879,N_9110);
xnor U11114 (N_11114,N_9975,N_8526);
and U11115 (N_11115,N_9301,N_8676);
or U11116 (N_11116,N_9772,N_9260);
and U11117 (N_11117,N_9678,N_8627);
and U11118 (N_11118,N_9489,N_8739);
and U11119 (N_11119,N_9952,N_9981);
xor U11120 (N_11120,N_8908,N_9025);
xnor U11121 (N_11121,N_8280,N_8547);
nand U11122 (N_11122,N_8158,N_8611);
nand U11123 (N_11123,N_8797,N_8964);
nand U11124 (N_11124,N_8488,N_8545);
xnor U11125 (N_11125,N_9227,N_8784);
nor U11126 (N_11126,N_9163,N_8427);
and U11127 (N_11127,N_8665,N_9748);
nand U11128 (N_11128,N_8492,N_9573);
nand U11129 (N_11129,N_9616,N_8560);
nor U11130 (N_11130,N_8296,N_8666);
and U11131 (N_11131,N_8149,N_9852);
or U11132 (N_11132,N_8588,N_9403);
and U11133 (N_11133,N_8149,N_8185);
or U11134 (N_11134,N_9923,N_8602);
nand U11135 (N_11135,N_9176,N_9879);
or U11136 (N_11136,N_8138,N_8235);
and U11137 (N_11137,N_8008,N_8690);
nor U11138 (N_11138,N_8272,N_8057);
or U11139 (N_11139,N_9577,N_9758);
xor U11140 (N_11140,N_8008,N_8563);
or U11141 (N_11141,N_8435,N_9346);
or U11142 (N_11142,N_8826,N_9844);
and U11143 (N_11143,N_8327,N_9872);
or U11144 (N_11144,N_8667,N_9776);
nand U11145 (N_11145,N_8903,N_8551);
or U11146 (N_11146,N_9457,N_9164);
nand U11147 (N_11147,N_8234,N_9082);
nor U11148 (N_11148,N_8446,N_8094);
or U11149 (N_11149,N_9616,N_9309);
and U11150 (N_11150,N_8345,N_9523);
or U11151 (N_11151,N_9248,N_8149);
nor U11152 (N_11152,N_9513,N_8418);
and U11153 (N_11153,N_9106,N_9683);
xnor U11154 (N_11154,N_9277,N_9238);
nor U11155 (N_11155,N_8113,N_9053);
xnor U11156 (N_11156,N_8927,N_8540);
or U11157 (N_11157,N_9152,N_9082);
or U11158 (N_11158,N_9866,N_8123);
nor U11159 (N_11159,N_9365,N_9685);
nand U11160 (N_11160,N_8416,N_9647);
nor U11161 (N_11161,N_9202,N_9589);
xor U11162 (N_11162,N_9510,N_9451);
xor U11163 (N_11163,N_8308,N_8780);
and U11164 (N_11164,N_9011,N_9272);
and U11165 (N_11165,N_8851,N_8814);
nand U11166 (N_11166,N_8941,N_9198);
and U11167 (N_11167,N_9521,N_9492);
nor U11168 (N_11168,N_9570,N_8268);
or U11169 (N_11169,N_9943,N_8661);
and U11170 (N_11170,N_9738,N_8886);
or U11171 (N_11171,N_8053,N_8987);
and U11172 (N_11172,N_9673,N_8672);
or U11173 (N_11173,N_9608,N_8715);
nor U11174 (N_11174,N_8116,N_9417);
and U11175 (N_11175,N_9884,N_8506);
and U11176 (N_11176,N_8074,N_8304);
nor U11177 (N_11177,N_9641,N_8896);
or U11178 (N_11178,N_8600,N_8207);
and U11179 (N_11179,N_8267,N_8669);
or U11180 (N_11180,N_8463,N_8306);
or U11181 (N_11181,N_8722,N_8502);
xor U11182 (N_11182,N_9343,N_8673);
nor U11183 (N_11183,N_9572,N_9485);
nor U11184 (N_11184,N_9934,N_8660);
and U11185 (N_11185,N_9358,N_8381);
nand U11186 (N_11186,N_9256,N_9950);
xor U11187 (N_11187,N_8838,N_8456);
nand U11188 (N_11188,N_9778,N_9584);
or U11189 (N_11189,N_8124,N_9965);
xnor U11190 (N_11190,N_8853,N_8846);
xor U11191 (N_11191,N_8485,N_9970);
nor U11192 (N_11192,N_8796,N_8381);
nor U11193 (N_11193,N_8536,N_9914);
and U11194 (N_11194,N_8210,N_9495);
or U11195 (N_11195,N_9563,N_9146);
xnor U11196 (N_11196,N_9492,N_9362);
nor U11197 (N_11197,N_8839,N_8364);
and U11198 (N_11198,N_9360,N_9298);
nor U11199 (N_11199,N_8259,N_8708);
nand U11200 (N_11200,N_8675,N_9105);
nor U11201 (N_11201,N_9273,N_8265);
nand U11202 (N_11202,N_8745,N_9807);
xnor U11203 (N_11203,N_9813,N_8858);
xnor U11204 (N_11204,N_8746,N_9477);
xnor U11205 (N_11205,N_8062,N_8667);
nand U11206 (N_11206,N_8967,N_9809);
nand U11207 (N_11207,N_8508,N_9215);
nor U11208 (N_11208,N_9910,N_9247);
nor U11209 (N_11209,N_8105,N_8232);
nand U11210 (N_11210,N_8406,N_8945);
and U11211 (N_11211,N_8896,N_8726);
nand U11212 (N_11212,N_9628,N_8111);
nand U11213 (N_11213,N_9878,N_9213);
nand U11214 (N_11214,N_8888,N_9177);
xor U11215 (N_11215,N_9076,N_9867);
nand U11216 (N_11216,N_9022,N_8602);
and U11217 (N_11217,N_9545,N_9879);
nand U11218 (N_11218,N_8211,N_9605);
nor U11219 (N_11219,N_8255,N_9586);
xnor U11220 (N_11220,N_8074,N_8422);
xnor U11221 (N_11221,N_8888,N_8622);
or U11222 (N_11222,N_8979,N_9154);
and U11223 (N_11223,N_9401,N_8652);
and U11224 (N_11224,N_8542,N_8234);
nand U11225 (N_11225,N_8754,N_9401);
or U11226 (N_11226,N_8145,N_9056);
or U11227 (N_11227,N_8204,N_8974);
nand U11228 (N_11228,N_8376,N_8161);
nand U11229 (N_11229,N_8651,N_8182);
xnor U11230 (N_11230,N_8686,N_8627);
or U11231 (N_11231,N_9405,N_9100);
and U11232 (N_11232,N_8042,N_8672);
or U11233 (N_11233,N_8695,N_8684);
xnor U11234 (N_11234,N_9071,N_9131);
and U11235 (N_11235,N_8379,N_8495);
nor U11236 (N_11236,N_8189,N_8452);
and U11237 (N_11237,N_8798,N_9418);
nand U11238 (N_11238,N_8080,N_9649);
and U11239 (N_11239,N_9518,N_8600);
and U11240 (N_11240,N_9393,N_9524);
and U11241 (N_11241,N_8300,N_9438);
or U11242 (N_11242,N_8891,N_9159);
nand U11243 (N_11243,N_8376,N_8273);
nand U11244 (N_11244,N_9795,N_9127);
nand U11245 (N_11245,N_8928,N_8620);
nand U11246 (N_11246,N_9462,N_8593);
or U11247 (N_11247,N_8023,N_8461);
and U11248 (N_11248,N_9317,N_9183);
or U11249 (N_11249,N_8142,N_9185);
and U11250 (N_11250,N_8220,N_9839);
nor U11251 (N_11251,N_9738,N_9952);
or U11252 (N_11252,N_8148,N_9093);
nand U11253 (N_11253,N_9259,N_9286);
nand U11254 (N_11254,N_9516,N_8772);
or U11255 (N_11255,N_9872,N_8016);
and U11256 (N_11256,N_9396,N_9075);
and U11257 (N_11257,N_8860,N_8866);
xor U11258 (N_11258,N_8530,N_8829);
and U11259 (N_11259,N_9902,N_9522);
and U11260 (N_11260,N_9560,N_9120);
nand U11261 (N_11261,N_9319,N_9112);
xnor U11262 (N_11262,N_8296,N_8965);
nand U11263 (N_11263,N_8783,N_8288);
or U11264 (N_11264,N_8534,N_9502);
nand U11265 (N_11265,N_9749,N_8113);
nor U11266 (N_11266,N_9250,N_9559);
nor U11267 (N_11267,N_8053,N_8182);
xor U11268 (N_11268,N_9724,N_8262);
nand U11269 (N_11269,N_8178,N_9250);
or U11270 (N_11270,N_9192,N_9359);
nand U11271 (N_11271,N_9436,N_9648);
nand U11272 (N_11272,N_8034,N_8081);
or U11273 (N_11273,N_9696,N_8677);
nor U11274 (N_11274,N_8691,N_9815);
nor U11275 (N_11275,N_9271,N_9088);
and U11276 (N_11276,N_9791,N_8038);
or U11277 (N_11277,N_8037,N_9615);
xnor U11278 (N_11278,N_9275,N_8893);
xor U11279 (N_11279,N_9917,N_9084);
nand U11280 (N_11280,N_9767,N_8011);
and U11281 (N_11281,N_9852,N_8632);
nor U11282 (N_11282,N_9670,N_9288);
or U11283 (N_11283,N_9573,N_8621);
nor U11284 (N_11284,N_9921,N_9127);
or U11285 (N_11285,N_9070,N_8319);
and U11286 (N_11286,N_9882,N_9771);
and U11287 (N_11287,N_9646,N_8736);
or U11288 (N_11288,N_8584,N_9162);
and U11289 (N_11289,N_9078,N_8063);
or U11290 (N_11290,N_8810,N_8579);
nor U11291 (N_11291,N_9232,N_8254);
and U11292 (N_11292,N_8145,N_8403);
nor U11293 (N_11293,N_8084,N_8645);
nor U11294 (N_11294,N_8689,N_8686);
nand U11295 (N_11295,N_9747,N_9554);
nand U11296 (N_11296,N_9584,N_8331);
nand U11297 (N_11297,N_8832,N_9393);
or U11298 (N_11298,N_9973,N_9219);
nor U11299 (N_11299,N_8083,N_9600);
nor U11300 (N_11300,N_8030,N_9796);
xnor U11301 (N_11301,N_8913,N_8411);
or U11302 (N_11302,N_9137,N_9760);
or U11303 (N_11303,N_9602,N_8537);
nor U11304 (N_11304,N_8581,N_8466);
nor U11305 (N_11305,N_8936,N_9614);
nor U11306 (N_11306,N_9132,N_8076);
xnor U11307 (N_11307,N_9009,N_9725);
and U11308 (N_11308,N_9475,N_9263);
nand U11309 (N_11309,N_9181,N_9153);
or U11310 (N_11310,N_8537,N_8919);
and U11311 (N_11311,N_8042,N_9073);
and U11312 (N_11312,N_9345,N_9952);
nor U11313 (N_11313,N_8654,N_8252);
nor U11314 (N_11314,N_9679,N_9532);
nand U11315 (N_11315,N_9198,N_8836);
nand U11316 (N_11316,N_8976,N_8177);
or U11317 (N_11317,N_9245,N_9297);
nand U11318 (N_11318,N_9607,N_9469);
or U11319 (N_11319,N_8182,N_9466);
xnor U11320 (N_11320,N_8454,N_8600);
nor U11321 (N_11321,N_9448,N_9933);
nand U11322 (N_11322,N_9782,N_8662);
nor U11323 (N_11323,N_9008,N_9689);
and U11324 (N_11324,N_9290,N_9801);
nand U11325 (N_11325,N_9861,N_9367);
or U11326 (N_11326,N_9031,N_9351);
xor U11327 (N_11327,N_9249,N_8456);
or U11328 (N_11328,N_9399,N_8184);
or U11329 (N_11329,N_9141,N_9556);
nand U11330 (N_11330,N_9085,N_9416);
and U11331 (N_11331,N_8495,N_8355);
xor U11332 (N_11332,N_9608,N_8570);
xnor U11333 (N_11333,N_8267,N_9981);
and U11334 (N_11334,N_8293,N_9762);
nor U11335 (N_11335,N_8922,N_9473);
or U11336 (N_11336,N_9189,N_8929);
xnor U11337 (N_11337,N_8460,N_9508);
or U11338 (N_11338,N_9525,N_8101);
nand U11339 (N_11339,N_8387,N_9159);
and U11340 (N_11340,N_9677,N_9057);
nor U11341 (N_11341,N_9866,N_9705);
and U11342 (N_11342,N_8608,N_9646);
and U11343 (N_11343,N_9205,N_8196);
nor U11344 (N_11344,N_9721,N_9662);
nand U11345 (N_11345,N_9364,N_8455);
nor U11346 (N_11346,N_8993,N_8888);
and U11347 (N_11347,N_8651,N_9006);
nand U11348 (N_11348,N_9675,N_9646);
nor U11349 (N_11349,N_8512,N_8381);
or U11350 (N_11350,N_9876,N_9323);
or U11351 (N_11351,N_9016,N_9803);
and U11352 (N_11352,N_9793,N_8176);
xnor U11353 (N_11353,N_9516,N_8844);
xnor U11354 (N_11354,N_9126,N_8467);
nand U11355 (N_11355,N_9404,N_9429);
and U11356 (N_11356,N_9551,N_9321);
xnor U11357 (N_11357,N_8988,N_8322);
and U11358 (N_11358,N_8175,N_9110);
or U11359 (N_11359,N_9306,N_8546);
nand U11360 (N_11360,N_8114,N_8960);
and U11361 (N_11361,N_9693,N_8095);
and U11362 (N_11362,N_8356,N_9431);
xnor U11363 (N_11363,N_9390,N_9227);
and U11364 (N_11364,N_8265,N_8633);
xor U11365 (N_11365,N_9121,N_9648);
nor U11366 (N_11366,N_9095,N_8069);
nor U11367 (N_11367,N_9201,N_9248);
and U11368 (N_11368,N_8249,N_8550);
nor U11369 (N_11369,N_9550,N_9645);
and U11370 (N_11370,N_9825,N_8017);
and U11371 (N_11371,N_8268,N_8497);
and U11372 (N_11372,N_9980,N_9804);
or U11373 (N_11373,N_9603,N_8838);
or U11374 (N_11374,N_8945,N_9321);
nand U11375 (N_11375,N_8857,N_8029);
and U11376 (N_11376,N_9578,N_9810);
nor U11377 (N_11377,N_9738,N_8342);
or U11378 (N_11378,N_8205,N_8869);
nand U11379 (N_11379,N_9105,N_8011);
and U11380 (N_11380,N_9620,N_9398);
nor U11381 (N_11381,N_9346,N_9952);
or U11382 (N_11382,N_9415,N_8207);
nand U11383 (N_11383,N_9433,N_9637);
xnor U11384 (N_11384,N_8102,N_8567);
or U11385 (N_11385,N_8015,N_8245);
nand U11386 (N_11386,N_8317,N_9167);
nor U11387 (N_11387,N_8576,N_9365);
or U11388 (N_11388,N_8110,N_9755);
or U11389 (N_11389,N_8958,N_9100);
and U11390 (N_11390,N_9105,N_8913);
or U11391 (N_11391,N_9099,N_8785);
and U11392 (N_11392,N_8528,N_8507);
xnor U11393 (N_11393,N_9745,N_9860);
nor U11394 (N_11394,N_9888,N_8342);
nor U11395 (N_11395,N_9418,N_8556);
nor U11396 (N_11396,N_9780,N_9195);
and U11397 (N_11397,N_8718,N_8960);
nor U11398 (N_11398,N_9000,N_9061);
or U11399 (N_11399,N_9401,N_9085);
or U11400 (N_11400,N_8495,N_9102);
nand U11401 (N_11401,N_9101,N_8334);
xnor U11402 (N_11402,N_8494,N_8261);
and U11403 (N_11403,N_8466,N_8315);
nor U11404 (N_11404,N_8775,N_8449);
nor U11405 (N_11405,N_9595,N_9636);
and U11406 (N_11406,N_9806,N_9364);
nand U11407 (N_11407,N_8029,N_9911);
nor U11408 (N_11408,N_9148,N_8741);
nor U11409 (N_11409,N_9863,N_9993);
or U11410 (N_11410,N_8324,N_9502);
and U11411 (N_11411,N_9168,N_8971);
nand U11412 (N_11412,N_9914,N_9264);
nor U11413 (N_11413,N_8784,N_9360);
or U11414 (N_11414,N_9363,N_9385);
nand U11415 (N_11415,N_8033,N_9119);
or U11416 (N_11416,N_8083,N_8689);
or U11417 (N_11417,N_8911,N_8256);
or U11418 (N_11418,N_8278,N_9671);
xor U11419 (N_11419,N_8599,N_8778);
xnor U11420 (N_11420,N_8216,N_9716);
nor U11421 (N_11421,N_8479,N_8557);
nor U11422 (N_11422,N_9173,N_9420);
or U11423 (N_11423,N_8115,N_8439);
nand U11424 (N_11424,N_9371,N_8766);
and U11425 (N_11425,N_9639,N_8419);
nor U11426 (N_11426,N_9022,N_8084);
or U11427 (N_11427,N_9586,N_8011);
nor U11428 (N_11428,N_9873,N_9635);
and U11429 (N_11429,N_9321,N_8276);
nand U11430 (N_11430,N_8358,N_8624);
and U11431 (N_11431,N_8525,N_8316);
or U11432 (N_11432,N_9302,N_9157);
nand U11433 (N_11433,N_9566,N_9889);
or U11434 (N_11434,N_8094,N_8671);
or U11435 (N_11435,N_8980,N_8340);
xnor U11436 (N_11436,N_8448,N_8918);
or U11437 (N_11437,N_8194,N_9230);
and U11438 (N_11438,N_8400,N_9400);
xnor U11439 (N_11439,N_9691,N_9818);
and U11440 (N_11440,N_8028,N_9448);
xnor U11441 (N_11441,N_8841,N_9536);
xnor U11442 (N_11442,N_8444,N_9795);
and U11443 (N_11443,N_8903,N_9578);
nor U11444 (N_11444,N_8565,N_8338);
and U11445 (N_11445,N_8280,N_9590);
or U11446 (N_11446,N_9670,N_9960);
or U11447 (N_11447,N_9555,N_9260);
or U11448 (N_11448,N_9336,N_8373);
nor U11449 (N_11449,N_8452,N_9434);
xnor U11450 (N_11450,N_8045,N_9846);
xor U11451 (N_11451,N_9588,N_9722);
xnor U11452 (N_11452,N_9025,N_8933);
nand U11453 (N_11453,N_9352,N_9467);
nand U11454 (N_11454,N_9769,N_9708);
nor U11455 (N_11455,N_8606,N_8964);
nor U11456 (N_11456,N_8429,N_8171);
nand U11457 (N_11457,N_9068,N_9413);
and U11458 (N_11458,N_9002,N_9610);
nor U11459 (N_11459,N_8258,N_9356);
and U11460 (N_11460,N_9938,N_9334);
and U11461 (N_11461,N_8153,N_9893);
and U11462 (N_11462,N_8755,N_9300);
or U11463 (N_11463,N_9054,N_9006);
nor U11464 (N_11464,N_9887,N_8507);
and U11465 (N_11465,N_9582,N_9580);
and U11466 (N_11466,N_9449,N_8290);
nor U11467 (N_11467,N_9199,N_9618);
nor U11468 (N_11468,N_9062,N_8054);
and U11469 (N_11469,N_8970,N_8969);
nand U11470 (N_11470,N_8952,N_8187);
nor U11471 (N_11471,N_8688,N_9006);
xor U11472 (N_11472,N_8174,N_9811);
and U11473 (N_11473,N_9043,N_8961);
and U11474 (N_11474,N_9578,N_8897);
xnor U11475 (N_11475,N_9298,N_8690);
and U11476 (N_11476,N_9160,N_8690);
nand U11477 (N_11477,N_9058,N_8035);
or U11478 (N_11478,N_9469,N_8861);
nor U11479 (N_11479,N_8200,N_9876);
and U11480 (N_11480,N_8754,N_8350);
nor U11481 (N_11481,N_9754,N_9183);
or U11482 (N_11482,N_9316,N_8995);
and U11483 (N_11483,N_9257,N_9505);
nand U11484 (N_11484,N_9130,N_8607);
xor U11485 (N_11485,N_8918,N_8209);
or U11486 (N_11486,N_9187,N_8373);
nand U11487 (N_11487,N_8197,N_8595);
nand U11488 (N_11488,N_8658,N_8031);
xor U11489 (N_11489,N_9772,N_9447);
nand U11490 (N_11490,N_9828,N_8644);
and U11491 (N_11491,N_9715,N_8258);
or U11492 (N_11492,N_9643,N_8692);
or U11493 (N_11493,N_8554,N_8521);
nand U11494 (N_11494,N_8482,N_9493);
nand U11495 (N_11495,N_8174,N_9613);
xnor U11496 (N_11496,N_8283,N_8944);
and U11497 (N_11497,N_9228,N_9264);
or U11498 (N_11498,N_9985,N_8933);
and U11499 (N_11499,N_8994,N_8794);
and U11500 (N_11500,N_8392,N_9067);
nand U11501 (N_11501,N_8733,N_9634);
and U11502 (N_11502,N_9571,N_8981);
nor U11503 (N_11503,N_9791,N_9847);
xnor U11504 (N_11504,N_8411,N_9437);
nor U11505 (N_11505,N_8215,N_8323);
nor U11506 (N_11506,N_9181,N_9480);
xnor U11507 (N_11507,N_9552,N_8130);
xnor U11508 (N_11508,N_9417,N_8731);
or U11509 (N_11509,N_8487,N_8608);
nor U11510 (N_11510,N_9876,N_8155);
or U11511 (N_11511,N_9076,N_8521);
and U11512 (N_11512,N_9995,N_8784);
or U11513 (N_11513,N_8867,N_8659);
nor U11514 (N_11514,N_8815,N_9705);
nor U11515 (N_11515,N_8680,N_8045);
and U11516 (N_11516,N_8942,N_9122);
nand U11517 (N_11517,N_8837,N_8676);
nand U11518 (N_11518,N_9507,N_9033);
xor U11519 (N_11519,N_9373,N_9682);
nor U11520 (N_11520,N_9544,N_9128);
nor U11521 (N_11521,N_8808,N_8050);
or U11522 (N_11522,N_8005,N_8014);
nor U11523 (N_11523,N_9955,N_9740);
nand U11524 (N_11524,N_9838,N_9442);
and U11525 (N_11525,N_8131,N_8254);
or U11526 (N_11526,N_8172,N_8563);
and U11527 (N_11527,N_8003,N_9710);
nand U11528 (N_11528,N_9437,N_9818);
nor U11529 (N_11529,N_9183,N_8326);
nor U11530 (N_11530,N_8326,N_8960);
nand U11531 (N_11531,N_9001,N_8898);
xnor U11532 (N_11532,N_8609,N_8849);
nand U11533 (N_11533,N_8565,N_9077);
or U11534 (N_11534,N_8186,N_9224);
xor U11535 (N_11535,N_8642,N_8430);
nor U11536 (N_11536,N_8009,N_9023);
nand U11537 (N_11537,N_8776,N_9986);
or U11538 (N_11538,N_8735,N_9550);
nand U11539 (N_11539,N_9124,N_9525);
nand U11540 (N_11540,N_8146,N_9039);
and U11541 (N_11541,N_9995,N_9690);
xor U11542 (N_11542,N_9218,N_8298);
xnor U11543 (N_11543,N_9219,N_8324);
nand U11544 (N_11544,N_8307,N_9082);
or U11545 (N_11545,N_9293,N_9997);
and U11546 (N_11546,N_9017,N_9930);
xor U11547 (N_11547,N_8086,N_8834);
or U11548 (N_11548,N_8445,N_9028);
nand U11549 (N_11549,N_9693,N_9536);
and U11550 (N_11550,N_8199,N_8086);
nor U11551 (N_11551,N_8837,N_9454);
xor U11552 (N_11552,N_8794,N_9044);
nand U11553 (N_11553,N_9020,N_8952);
nand U11554 (N_11554,N_9577,N_9472);
and U11555 (N_11555,N_8463,N_8457);
xor U11556 (N_11556,N_8800,N_9648);
nand U11557 (N_11557,N_9862,N_8549);
or U11558 (N_11558,N_8646,N_9338);
nor U11559 (N_11559,N_9601,N_8177);
nor U11560 (N_11560,N_8154,N_8940);
nand U11561 (N_11561,N_8813,N_9652);
nand U11562 (N_11562,N_8558,N_9616);
and U11563 (N_11563,N_8624,N_9361);
nand U11564 (N_11564,N_9392,N_9193);
xnor U11565 (N_11565,N_9663,N_8867);
nor U11566 (N_11566,N_8020,N_9944);
or U11567 (N_11567,N_8048,N_9652);
nand U11568 (N_11568,N_9478,N_9416);
or U11569 (N_11569,N_9908,N_8465);
nor U11570 (N_11570,N_9238,N_8547);
nor U11571 (N_11571,N_8100,N_8932);
and U11572 (N_11572,N_9153,N_9113);
and U11573 (N_11573,N_8189,N_9652);
nand U11574 (N_11574,N_8922,N_8622);
xor U11575 (N_11575,N_9947,N_8308);
and U11576 (N_11576,N_8119,N_9762);
xnor U11577 (N_11577,N_8492,N_9391);
nor U11578 (N_11578,N_9993,N_8609);
or U11579 (N_11579,N_8232,N_8428);
and U11580 (N_11580,N_8758,N_9335);
or U11581 (N_11581,N_8841,N_9921);
or U11582 (N_11582,N_8799,N_8643);
nor U11583 (N_11583,N_9895,N_9994);
nand U11584 (N_11584,N_8610,N_9348);
and U11585 (N_11585,N_9034,N_8485);
or U11586 (N_11586,N_8665,N_8423);
xnor U11587 (N_11587,N_8494,N_9659);
and U11588 (N_11588,N_9565,N_8362);
or U11589 (N_11589,N_9401,N_8858);
xor U11590 (N_11590,N_9757,N_9990);
nand U11591 (N_11591,N_8629,N_9229);
nor U11592 (N_11592,N_9571,N_8989);
nor U11593 (N_11593,N_8013,N_9004);
nor U11594 (N_11594,N_9679,N_8388);
or U11595 (N_11595,N_9162,N_8209);
or U11596 (N_11596,N_8252,N_8343);
nand U11597 (N_11597,N_9996,N_8524);
or U11598 (N_11598,N_9394,N_9089);
nor U11599 (N_11599,N_8824,N_8246);
or U11600 (N_11600,N_9357,N_9799);
and U11601 (N_11601,N_8762,N_8614);
or U11602 (N_11602,N_8520,N_9525);
nor U11603 (N_11603,N_8514,N_9123);
nand U11604 (N_11604,N_8084,N_8218);
nor U11605 (N_11605,N_9499,N_8951);
xor U11606 (N_11606,N_9780,N_9996);
nor U11607 (N_11607,N_9016,N_8812);
or U11608 (N_11608,N_8085,N_9061);
or U11609 (N_11609,N_8942,N_8710);
or U11610 (N_11610,N_8126,N_8531);
nand U11611 (N_11611,N_9371,N_8941);
or U11612 (N_11612,N_8703,N_9836);
nor U11613 (N_11613,N_9777,N_9372);
xor U11614 (N_11614,N_8275,N_9014);
or U11615 (N_11615,N_9800,N_8696);
nand U11616 (N_11616,N_8076,N_8838);
nor U11617 (N_11617,N_8623,N_8457);
and U11618 (N_11618,N_9259,N_9442);
and U11619 (N_11619,N_8142,N_8416);
nand U11620 (N_11620,N_8940,N_9850);
nand U11621 (N_11621,N_8724,N_9400);
nand U11622 (N_11622,N_8505,N_8269);
xor U11623 (N_11623,N_9720,N_9488);
or U11624 (N_11624,N_8269,N_8428);
nand U11625 (N_11625,N_9198,N_8102);
or U11626 (N_11626,N_9302,N_8748);
or U11627 (N_11627,N_9565,N_9955);
nand U11628 (N_11628,N_9192,N_9893);
xnor U11629 (N_11629,N_9182,N_8509);
nand U11630 (N_11630,N_9564,N_8341);
or U11631 (N_11631,N_8932,N_9275);
xor U11632 (N_11632,N_8199,N_9764);
nand U11633 (N_11633,N_8951,N_9851);
xnor U11634 (N_11634,N_8917,N_9197);
xnor U11635 (N_11635,N_8786,N_8393);
xnor U11636 (N_11636,N_8013,N_9585);
nor U11637 (N_11637,N_8529,N_9928);
and U11638 (N_11638,N_9221,N_9463);
xnor U11639 (N_11639,N_8233,N_9327);
nand U11640 (N_11640,N_9427,N_8593);
or U11641 (N_11641,N_9429,N_8762);
nand U11642 (N_11642,N_8678,N_9735);
or U11643 (N_11643,N_9281,N_9878);
nor U11644 (N_11644,N_9326,N_9952);
nor U11645 (N_11645,N_9518,N_8059);
xnor U11646 (N_11646,N_8606,N_9622);
nor U11647 (N_11647,N_8447,N_8798);
nand U11648 (N_11648,N_9165,N_8883);
or U11649 (N_11649,N_8270,N_8858);
nor U11650 (N_11650,N_8957,N_9127);
nand U11651 (N_11651,N_8258,N_8247);
xnor U11652 (N_11652,N_8618,N_8158);
and U11653 (N_11653,N_8747,N_8507);
and U11654 (N_11654,N_9252,N_8915);
xnor U11655 (N_11655,N_9331,N_9095);
xnor U11656 (N_11656,N_9804,N_8728);
or U11657 (N_11657,N_8697,N_9339);
and U11658 (N_11658,N_8532,N_8384);
xor U11659 (N_11659,N_8768,N_9953);
or U11660 (N_11660,N_8894,N_8909);
or U11661 (N_11661,N_9814,N_8314);
or U11662 (N_11662,N_9522,N_9613);
nor U11663 (N_11663,N_8261,N_8491);
xor U11664 (N_11664,N_8302,N_9895);
nor U11665 (N_11665,N_9245,N_8964);
xor U11666 (N_11666,N_9928,N_9251);
nor U11667 (N_11667,N_8192,N_9397);
nand U11668 (N_11668,N_9823,N_8986);
and U11669 (N_11669,N_9973,N_8859);
xnor U11670 (N_11670,N_8785,N_9030);
xor U11671 (N_11671,N_9473,N_8322);
and U11672 (N_11672,N_8867,N_9442);
nor U11673 (N_11673,N_8870,N_9264);
or U11674 (N_11674,N_8474,N_8924);
and U11675 (N_11675,N_8327,N_9789);
or U11676 (N_11676,N_8361,N_9571);
and U11677 (N_11677,N_9872,N_8558);
nor U11678 (N_11678,N_9528,N_9668);
xor U11679 (N_11679,N_9713,N_9156);
or U11680 (N_11680,N_8878,N_9694);
and U11681 (N_11681,N_9236,N_8606);
xor U11682 (N_11682,N_8943,N_9651);
xnor U11683 (N_11683,N_9560,N_9470);
or U11684 (N_11684,N_9767,N_8135);
nor U11685 (N_11685,N_9194,N_9709);
xnor U11686 (N_11686,N_8173,N_8979);
nand U11687 (N_11687,N_9576,N_9954);
xor U11688 (N_11688,N_9622,N_8077);
or U11689 (N_11689,N_9473,N_8345);
or U11690 (N_11690,N_9047,N_8709);
or U11691 (N_11691,N_8313,N_9372);
nand U11692 (N_11692,N_8083,N_8847);
or U11693 (N_11693,N_8008,N_8278);
or U11694 (N_11694,N_8825,N_8162);
and U11695 (N_11695,N_8226,N_9141);
nor U11696 (N_11696,N_8175,N_9870);
and U11697 (N_11697,N_8649,N_9101);
nand U11698 (N_11698,N_8306,N_8422);
nand U11699 (N_11699,N_8366,N_9583);
or U11700 (N_11700,N_8534,N_9252);
xor U11701 (N_11701,N_9304,N_9971);
or U11702 (N_11702,N_9809,N_8775);
nor U11703 (N_11703,N_8826,N_8179);
nand U11704 (N_11704,N_8551,N_8523);
or U11705 (N_11705,N_8356,N_8690);
or U11706 (N_11706,N_8934,N_8659);
or U11707 (N_11707,N_9871,N_8206);
nand U11708 (N_11708,N_8744,N_9754);
and U11709 (N_11709,N_8388,N_9862);
xnor U11710 (N_11710,N_9904,N_8818);
xor U11711 (N_11711,N_8742,N_9585);
or U11712 (N_11712,N_9776,N_8162);
or U11713 (N_11713,N_8168,N_9355);
nand U11714 (N_11714,N_9350,N_8262);
nand U11715 (N_11715,N_9398,N_8158);
or U11716 (N_11716,N_8548,N_9161);
nand U11717 (N_11717,N_9337,N_8270);
or U11718 (N_11718,N_9755,N_9863);
nand U11719 (N_11719,N_9176,N_9464);
xnor U11720 (N_11720,N_8085,N_9732);
nor U11721 (N_11721,N_9339,N_9481);
and U11722 (N_11722,N_8129,N_9985);
and U11723 (N_11723,N_8545,N_8417);
xor U11724 (N_11724,N_8892,N_8937);
or U11725 (N_11725,N_8282,N_9870);
nand U11726 (N_11726,N_8681,N_8812);
and U11727 (N_11727,N_8947,N_9630);
and U11728 (N_11728,N_9791,N_8969);
nand U11729 (N_11729,N_9435,N_9982);
nor U11730 (N_11730,N_8363,N_9095);
xor U11731 (N_11731,N_8024,N_9770);
nor U11732 (N_11732,N_9731,N_8005);
nor U11733 (N_11733,N_8668,N_9316);
xnor U11734 (N_11734,N_9278,N_8661);
nor U11735 (N_11735,N_9561,N_8945);
nand U11736 (N_11736,N_9149,N_9821);
xnor U11737 (N_11737,N_8790,N_9565);
xor U11738 (N_11738,N_9308,N_9947);
nor U11739 (N_11739,N_8830,N_9509);
nand U11740 (N_11740,N_8505,N_8517);
nand U11741 (N_11741,N_8140,N_8486);
and U11742 (N_11742,N_8387,N_8524);
or U11743 (N_11743,N_8817,N_8394);
and U11744 (N_11744,N_9739,N_8326);
xnor U11745 (N_11745,N_8134,N_9958);
or U11746 (N_11746,N_8863,N_8751);
nor U11747 (N_11747,N_8225,N_8158);
or U11748 (N_11748,N_8922,N_9767);
nor U11749 (N_11749,N_8522,N_9883);
and U11750 (N_11750,N_9826,N_9295);
nor U11751 (N_11751,N_8453,N_8220);
and U11752 (N_11752,N_9119,N_9516);
nor U11753 (N_11753,N_9395,N_9810);
nand U11754 (N_11754,N_8666,N_8617);
and U11755 (N_11755,N_8004,N_9754);
nand U11756 (N_11756,N_8647,N_9859);
nor U11757 (N_11757,N_9821,N_8516);
nor U11758 (N_11758,N_8292,N_8864);
xor U11759 (N_11759,N_8675,N_9857);
nand U11760 (N_11760,N_9442,N_8918);
or U11761 (N_11761,N_8745,N_8999);
nand U11762 (N_11762,N_9959,N_9359);
or U11763 (N_11763,N_9132,N_8511);
or U11764 (N_11764,N_8148,N_9265);
nand U11765 (N_11765,N_9322,N_9999);
xnor U11766 (N_11766,N_9001,N_8179);
or U11767 (N_11767,N_8683,N_9569);
or U11768 (N_11768,N_9201,N_8971);
nand U11769 (N_11769,N_8107,N_8195);
nor U11770 (N_11770,N_8000,N_8481);
and U11771 (N_11771,N_8763,N_9600);
nand U11772 (N_11772,N_8137,N_8433);
nand U11773 (N_11773,N_8578,N_9729);
nand U11774 (N_11774,N_9063,N_9844);
xnor U11775 (N_11775,N_9698,N_8238);
and U11776 (N_11776,N_8376,N_8259);
nand U11777 (N_11777,N_8822,N_8189);
xnor U11778 (N_11778,N_9814,N_9838);
nand U11779 (N_11779,N_9734,N_8818);
or U11780 (N_11780,N_8762,N_8863);
nor U11781 (N_11781,N_9438,N_9596);
nand U11782 (N_11782,N_9064,N_9629);
or U11783 (N_11783,N_8438,N_9107);
nand U11784 (N_11784,N_9178,N_9216);
nor U11785 (N_11785,N_9334,N_8362);
nor U11786 (N_11786,N_8415,N_9520);
and U11787 (N_11787,N_9753,N_9183);
or U11788 (N_11788,N_9053,N_8975);
or U11789 (N_11789,N_9566,N_8553);
nor U11790 (N_11790,N_8053,N_9327);
nand U11791 (N_11791,N_9942,N_8153);
or U11792 (N_11792,N_8804,N_9364);
and U11793 (N_11793,N_9121,N_8663);
or U11794 (N_11794,N_9572,N_9751);
nand U11795 (N_11795,N_9309,N_8225);
nand U11796 (N_11796,N_9670,N_8902);
or U11797 (N_11797,N_8338,N_9641);
or U11798 (N_11798,N_8987,N_8231);
nor U11799 (N_11799,N_8804,N_8376);
and U11800 (N_11800,N_9010,N_9255);
xnor U11801 (N_11801,N_8110,N_8359);
or U11802 (N_11802,N_8960,N_9282);
nand U11803 (N_11803,N_9562,N_8599);
or U11804 (N_11804,N_8561,N_9284);
nor U11805 (N_11805,N_9650,N_8282);
nor U11806 (N_11806,N_9461,N_8826);
nor U11807 (N_11807,N_8529,N_8760);
nand U11808 (N_11808,N_9448,N_8412);
xnor U11809 (N_11809,N_9882,N_8795);
or U11810 (N_11810,N_9671,N_9987);
and U11811 (N_11811,N_9870,N_8368);
nor U11812 (N_11812,N_9205,N_8635);
nand U11813 (N_11813,N_9630,N_8350);
nand U11814 (N_11814,N_8071,N_8110);
nand U11815 (N_11815,N_8438,N_9119);
nand U11816 (N_11816,N_8036,N_9133);
nor U11817 (N_11817,N_8769,N_9476);
nor U11818 (N_11818,N_8284,N_9190);
nor U11819 (N_11819,N_9354,N_9534);
or U11820 (N_11820,N_9863,N_8429);
or U11821 (N_11821,N_9414,N_8306);
and U11822 (N_11822,N_9678,N_9208);
nand U11823 (N_11823,N_9985,N_9838);
xor U11824 (N_11824,N_9465,N_9544);
nor U11825 (N_11825,N_9481,N_9492);
and U11826 (N_11826,N_9003,N_8745);
nor U11827 (N_11827,N_8250,N_8605);
xnor U11828 (N_11828,N_8628,N_8510);
and U11829 (N_11829,N_9928,N_8077);
xor U11830 (N_11830,N_8572,N_9868);
and U11831 (N_11831,N_9056,N_9400);
xor U11832 (N_11832,N_8414,N_9522);
nand U11833 (N_11833,N_8705,N_9470);
or U11834 (N_11834,N_8519,N_9657);
xnor U11835 (N_11835,N_8716,N_9365);
nand U11836 (N_11836,N_8073,N_9916);
and U11837 (N_11837,N_9774,N_9188);
and U11838 (N_11838,N_8966,N_9277);
nand U11839 (N_11839,N_9742,N_9262);
nor U11840 (N_11840,N_8764,N_8305);
nor U11841 (N_11841,N_8072,N_9766);
xnor U11842 (N_11842,N_8698,N_9935);
nor U11843 (N_11843,N_9355,N_8343);
and U11844 (N_11844,N_8253,N_8982);
or U11845 (N_11845,N_8997,N_8724);
nor U11846 (N_11846,N_8316,N_8449);
or U11847 (N_11847,N_9720,N_9626);
xnor U11848 (N_11848,N_8366,N_9993);
and U11849 (N_11849,N_9172,N_9442);
or U11850 (N_11850,N_9333,N_9441);
nand U11851 (N_11851,N_9576,N_9728);
nand U11852 (N_11852,N_8814,N_9056);
and U11853 (N_11853,N_8287,N_9300);
nand U11854 (N_11854,N_9781,N_9116);
or U11855 (N_11855,N_9323,N_8020);
and U11856 (N_11856,N_8666,N_8145);
nand U11857 (N_11857,N_9544,N_9734);
nand U11858 (N_11858,N_9919,N_8567);
xnor U11859 (N_11859,N_8611,N_9110);
and U11860 (N_11860,N_8681,N_8092);
or U11861 (N_11861,N_9246,N_8467);
and U11862 (N_11862,N_8427,N_9373);
or U11863 (N_11863,N_8084,N_9896);
nor U11864 (N_11864,N_8920,N_8003);
and U11865 (N_11865,N_8527,N_9769);
xnor U11866 (N_11866,N_8274,N_9967);
or U11867 (N_11867,N_9929,N_9685);
xnor U11868 (N_11868,N_9707,N_8327);
nand U11869 (N_11869,N_8352,N_8770);
and U11870 (N_11870,N_9714,N_9847);
nor U11871 (N_11871,N_8233,N_8177);
and U11872 (N_11872,N_8286,N_9830);
or U11873 (N_11873,N_9354,N_9313);
and U11874 (N_11874,N_8190,N_8845);
nand U11875 (N_11875,N_9354,N_8195);
or U11876 (N_11876,N_8048,N_9339);
xnor U11877 (N_11877,N_8593,N_8825);
nand U11878 (N_11878,N_9074,N_9323);
or U11879 (N_11879,N_8644,N_8521);
nor U11880 (N_11880,N_9836,N_8712);
nor U11881 (N_11881,N_9982,N_8265);
and U11882 (N_11882,N_9671,N_9878);
nand U11883 (N_11883,N_8335,N_8684);
and U11884 (N_11884,N_9617,N_8053);
nand U11885 (N_11885,N_8178,N_9192);
or U11886 (N_11886,N_9998,N_8867);
nand U11887 (N_11887,N_8865,N_8276);
or U11888 (N_11888,N_9320,N_9281);
or U11889 (N_11889,N_8215,N_8896);
nand U11890 (N_11890,N_9580,N_9191);
xnor U11891 (N_11891,N_8461,N_8714);
and U11892 (N_11892,N_8365,N_9787);
nor U11893 (N_11893,N_9828,N_9983);
nor U11894 (N_11894,N_8513,N_8496);
nor U11895 (N_11895,N_9610,N_8277);
and U11896 (N_11896,N_9544,N_9321);
nand U11897 (N_11897,N_9674,N_9151);
xnor U11898 (N_11898,N_9258,N_8464);
and U11899 (N_11899,N_8034,N_9677);
nor U11900 (N_11900,N_9756,N_8526);
and U11901 (N_11901,N_8470,N_8495);
nor U11902 (N_11902,N_9450,N_9804);
or U11903 (N_11903,N_8691,N_9653);
nor U11904 (N_11904,N_8102,N_8394);
or U11905 (N_11905,N_8297,N_8175);
nand U11906 (N_11906,N_9692,N_8603);
nor U11907 (N_11907,N_9777,N_9046);
or U11908 (N_11908,N_8675,N_8487);
xor U11909 (N_11909,N_9221,N_9284);
nor U11910 (N_11910,N_9115,N_9978);
nand U11911 (N_11911,N_8704,N_8798);
xor U11912 (N_11912,N_8547,N_9207);
nand U11913 (N_11913,N_9890,N_8452);
xnor U11914 (N_11914,N_8262,N_8185);
or U11915 (N_11915,N_9436,N_9033);
and U11916 (N_11916,N_8809,N_8591);
or U11917 (N_11917,N_9139,N_8867);
nand U11918 (N_11918,N_8235,N_8087);
nor U11919 (N_11919,N_8916,N_8231);
nor U11920 (N_11920,N_8258,N_9358);
nor U11921 (N_11921,N_9254,N_8124);
and U11922 (N_11922,N_9671,N_8760);
xor U11923 (N_11923,N_9128,N_9984);
nor U11924 (N_11924,N_8974,N_8658);
and U11925 (N_11925,N_9448,N_8083);
nor U11926 (N_11926,N_8833,N_8658);
nand U11927 (N_11927,N_8046,N_9188);
nand U11928 (N_11928,N_9280,N_8067);
xnor U11929 (N_11929,N_8063,N_9648);
xor U11930 (N_11930,N_8641,N_9449);
or U11931 (N_11931,N_9686,N_9326);
or U11932 (N_11932,N_8317,N_8341);
and U11933 (N_11933,N_8636,N_9033);
and U11934 (N_11934,N_8253,N_8409);
and U11935 (N_11935,N_9291,N_9567);
nor U11936 (N_11936,N_9699,N_8941);
or U11937 (N_11937,N_8698,N_8332);
xnor U11938 (N_11938,N_9371,N_8080);
or U11939 (N_11939,N_9599,N_9549);
xnor U11940 (N_11940,N_9939,N_9346);
xnor U11941 (N_11941,N_9870,N_8976);
and U11942 (N_11942,N_8469,N_9295);
and U11943 (N_11943,N_8978,N_8737);
xnor U11944 (N_11944,N_8864,N_9502);
or U11945 (N_11945,N_8861,N_9118);
nor U11946 (N_11946,N_9370,N_8335);
nand U11947 (N_11947,N_9301,N_9118);
or U11948 (N_11948,N_8911,N_8796);
or U11949 (N_11949,N_8246,N_9185);
nor U11950 (N_11950,N_9241,N_9676);
nor U11951 (N_11951,N_9788,N_8444);
xor U11952 (N_11952,N_9704,N_8610);
nor U11953 (N_11953,N_8173,N_9372);
nor U11954 (N_11954,N_8998,N_8504);
or U11955 (N_11955,N_9742,N_9940);
or U11956 (N_11956,N_9014,N_9291);
and U11957 (N_11957,N_8462,N_9089);
nand U11958 (N_11958,N_8407,N_9067);
xor U11959 (N_11959,N_8030,N_9152);
nor U11960 (N_11960,N_9049,N_9639);
nor U11961 (N_11961,N_8403,N_9396);
nand U11962 (N_11962,N_8664,N_8239);
nand U11963 (N_11963,N_8395,N_9412);
nor U11964 (N_11964,N_9213,N_8586);
nand U11965 (N_11965,N_9412,N_9705);
xor U11966 (N_11966,N_8237,N_9822);
nor U11967 (N_11967,N_9435,N_8104);
and U11968 (N_11968,N_9861,N_8701);
and U11969 (N_11969,N_8725,N_9259);
nor U11970 (N_11970,N_9906,N_9606);
or U11971 (N_11971,N_9775,N_9527);
and U11972 (N_11972,N_9839,N_8271);
xnor U11973 (N_11973,N_8246,N_8058);
and U11974 (N_11974,N_8393,N_8514);
nand U11975 (N_11975,N_9961,N_8435);
or U11976 (N_11976,N_8005,N_8682);
nor U11977 (N_11977,N_9109,N_9694);
or U11978 (N_11978,N_8156,N_9752);
xnor U11979 (N_11979,N_9647,N_8612);
or U11980 (N_11980,N_9410,N_9109);
and U11981 (N_11981,N_9228,N_9709);
xnor U11982 (N_11982,N_9216,N_9185);
or U11983 (N_11983,N_9466,N_8704);
xnor U11984 (N_11984,N_8331,N_9774);
or U11985 (N_11985,N_9681,N_9746);
nand U11986 (N_11986,N_8953,N_8911);
nor U11987 (N_11987,N_8201,N_8405);
xnor U11988 (N_11988,N_9259,N_8373);
nand U11989 (N_11989,N_8728,N_9598);
xnor U11990 (N_11990,N_8915,N_8867);
or U11991 (N_11991,N_8216,N_8406);
xnor U11992 (N_11992,N_9759,N_9499);
nand U11993 (N_11993,N_8168,N_9538);
or U11994 (N_11994,N_9477,N_9143);
xnor U11995 (N_11995,N_9739,N_8543);
nor U11996 (N_11996,N_9053,N_8611);
or U11997 (N_11997,N_9864,N_8854);
or U11998 (N_11998,N_9858,N_8029);
or U11999 (N_11999,N_8519,N_8742);
or U12000 (N_12000,N_11046,N_10391);
xor U12001 (N_12001,N_11073,N_11319);
and U12002 (N_12002,N_10101,N_11437);
nand U12003 (N_12003,N_10687,N_10916);
and U12004 (N_12004,N_10668,N_10670);
and U12005 (N_12005,N_10225,N_11756);
xnor U12006 (N_12006,N_10015,N_10021);
nor U12007 (N_12007,N_10199,N_11485);
nor U12008 (N_12008,N_11725,N_10580);
nor U12009 (N_12009,N_11406,N_11938);
xor U12010 (N_12010,N_10809,N_10691);
xor U12011 (N_12011,N_11116,N_10406);
nand U12012 (N_12012,N_10781,N_11313);
nor U12013 (N_12013,N_11977,N_11642);
and U12014 (N_12014,N_11509,N_11267);
nor U12015 (N_12015,N_11692,N_10060);
nor U12016 (N_12016,N_10073,N_10362);
or U12017 (N_12017,N_11742,N_11235);
or U12018 (N_12018,N_11015,N_11654);
and U12019 (N_12019,N_10645,N_10657);
or U12020 (N_12020,N_11576,N_10495);
nand U12021 (N_12021,N_11214,N_11338);
or U12022 (N_12022,N_10742,N_10539);
or U12023 (N_12023,N_10681,N_11249);
and U12024 (N_12024,N_11035,N_11841);
nor U12025 (N_12025,N_11131,N_10125);
or U12026 (N_12026,N_10690,N_11113);
nand U12027 (N_12027,N_11278,N_10948);
and U12028 (N_12028,N_10925,N_10014);
and U12029 (N_12029,N_11252,N_11499);
nand U12030 (N_12030,N_11829,N_10148);
nand U12031 (N_12031,N_10924,N_10266);
xnor U12032 (N_12032,N_10595,N_11306);
xor U12033 (N_12033,N_10052,N_10956);
and U12034 (N_12034,N_11102,N_11143);
nor U12035 (N_12035,N_11592,N_11473);
and U12036 (N_12036,N_11611,N_11813);
or U12037 (N_12037,N_10984,N_10335);
nand U12038 (N_12038,N_10200,N_11582);
and U12039 (N_12039,N_10336,N_10233);
nand U12040 (N_12040,N_10591,N_10864);
or U12041 (N_12041,N_10971,N_11285);
nand U12042 (N_12042,N_11453,N_11491);
or U12043 (N_12043,N_11941,N_10585);
nand U12044 (N_12044,N_11699,N_10597);
or U12045 (N_12045,N_11626,N_10277);
nor U12046 (N_12046,N_11401,N_11939);
nand U12047 (N_12047,N_11641,N_10483);
and U12048 (N_12048,N_10557,N_10902);
and U12049 (N_12049,N_10800,N_10538);
xnor U12050 (N_12050,N_11317,N_10083);
xor U12051 (N_12051,N_11442,N_10805);
nor U12052 (N_12052,N_11812,N_10001);
nor U12053 (N_12053,N_10959,N_10556);
or U12054 (N_12054,N_10491,N_10622);
xnor U12055 (N_12055,N_10744,N_10222);
nor U12056 (N_12056,N_11649,N_11365);
or U12057 (N_12057,N_11480,N_10050);
xnor U12058 (N_12058,N_11470,N_10067);
or U12059 (N_12059,N_10772,N_10770);
xor U12060 (N_12060,N_10150,N_10260);
or U12061 (N_12061,N_10082,N_10127);
nor U12062 (N_12062,N_10636,N_11221);
nand U12063 (N_12063,N_11656,N_11281);
nor U12064 (N_12064,N_10875,N_10341);
nor U12065 (N_12065,N_10940,N_10903);
nor U12066 (N_12066,N_10117,N_10288);
or U12067 (N_12067,N_10129,N_11018);
and U12068 (N_12068,N_10255,N_10510);
nor U12069 (N_12069,N_10671,N_10347);
and U12070 (N_12070,N_11684,N_11662);
nor U12071 (N_12071,N_11447,N_10138);
nand U12072 (N_12072,N_11646,N_10416);
nor U12073 (N_12073,N_10504,N_10996);
and U12074 (N_12074,N_11392,N_11346);
nand U12075 (N_12075,N_10434,N_11661);
xor U12076 (N_12076,N_11802,N_11976);
nor U12077 (N_12077,N_10814,N_10968);
or U12078 (N_12078,N_10316,N_11227);
or U12079 (N_12079,N_11651,N_10787);
or U12080 (N_12080,N_10618,N_11198);
or U12081 (N_12081,N_11922,N_11593);
nand U12082 (N_12082,N_11157,N_10145);
and U12083 (N_12083,N_11492,N_11905);
or U12084 (N_12084,N_10040,N_11872);
and U12085 (N_12085,N_10766,N_11153);
and U12086 (N_12086,N_11632,N_10477);
or U12087 (N_12087,N_10066,N_10221);
and U12088 (N_12088,N_11417,N_11605);
nor U12089 (N_12089,N_10723,N_11533);
and U12090 (N_12090,N_10323,N_11248);
nand U12091 (N_12091,N_11388,N_11712);
nor U12092 (N_12092,N_11121,N_10782);
or U12093 (N_12093,N_11541,N_10802);
and U12094 (N_12094,N_10081,N_11151);
nor U12095 (N_12095,N_10149,N_10880);
nand U12096 (N_12096,N_11849,N_10536);
xnor U12097 (N_12097,N_10778,N_10877);
or U12098 (N_12098,N_11530,N_10686);
nor U12099 (N_12099,N_10895,N_10216);
nor U12100 (N_12100,N_10540,N_11929);
and U12101 (N_12101,N_10793,N_10534);
and U12102 (N_12102,N_10115,N_10286);
xnor U12103 (N_12103,N_11482,N_11867);
and U12104 (N_12104,N_10166,N_11142);
nor U12105 (N_12105,N_11347,N_10408);
and U12106 (N_12106,N_10227,N_10048);
or U12107 (N_12107,N_11122,N_11820);
or U12108 (N_12108,N_10301,N_11586);
nor U12109 (N_12109,N_11280,N_11061);
xnor U12110 (N_12110,N_11192,N_11964);
or U12111 (N_12111,N_10649,N_10777);
or U12112 (N_12112,N_11109,N_11033);
nand U12113 (N_12113,N_10454,N_10063);
or U12114 (N_12114,N_11924,N_10685);
and U12115 (N_12115,N_10946,N_10709);
and U12116 (N_12116,N_11194,N_11856);
nor U12117 (N_12117,N_10547,N_10569);
xnor U12118 (N_12118,N_11718,N_10939);
nor U12119 (N_12119,N_10708,N_10741);
xor U12120 (N_12120,N_11047,N_10244);
nor U12121 (N_12121,N_10771,N_11567);
nor U12122 (N_12122,N_10969,N_11197);
or U12123 (N_12123,N_10624,N_10695);
and U12124 (N_12124,N_10724,N_10384);
or U12125 (N_12125,N_11776,N_11980);
xor U12126 (N_12126,N_11665,N_10185);
xnor U12127 (N_12127,N_10499,N_10300);
xnor U12128 (N_12128,N_10905,N_11495);
and U12129 (N_12129,N_10355,N_11629);
nor U12130 (N_12130,N_10816,N_11778);
xor U12131 (N_12131,N_10480,N_11393);
nand U12132 (N_12132,N_11445,N_10870);
xor U12133 (N_12133,N_10195,N_11390);
and U12134 (N_12134,N_10628,N_11022);
nand U12135 (N_12135,N_10057,N_10620);
or U12136 (N_12136,N_11009,N_11225);
or U12137 (N_12137,N_11126,N_10059);
and U12138 (N_12138,N_10158,N_11570);
nand U12139 (N_12139,N_10289,N_11387);
and U12140 (N_12140,N_10998,N_11246);
and U12141 (N_12141,N_11244,N_10731);
and U12142 (N_12142,N_11762,N_10560);
xor U12143 (N_12143,N_10721,N_11412);
and U12144 (N_12144,N_11222,N_10604);
xor U12145 (N_12145,N_11655,N_11298);
xnor U12146 (N_12146,N_10352,N_11483);
nor U12147 (N_12147,N_11430,N_10364);
and U12148 (N_12148,N_10209,N_10737);
nor U12149 (N_12149,N_11374,N_11024);
and U12150 (N_12150,N_10826,N_10562);
and U12151 (N_12151,N_11765,N_10938);
nor U12152 (N_12152,N_11761,N_11077);
nand U12153 (N_12153,N_11339,N_11696);
nand U12154 (N_12154,N_10632,N_11023);
nor U12155 (N_12155,N_11734,N_11542);
and U12156 (N_12156,N_11880,N_10462);
and U12157 (N_12157,N_11769,N_11946);
nand U12158 (N_12158,N_10099,N_10134);
xor U12159 (N_12159,N_10997,N_10069);
xnor U12160 (N_12160,N_10854,N_10439);
xnor U12161 (N_12161,N_10400,N_11028);
nor U12162 (N_12162,N_11479,N_11352);
nor U12163 (N_12163,N_11261,N_10375);
nor U12164 (N_12164,N_10779,N_10531);
nor U12165 (N_12165,N_10614,N_11243);
xnor U12166 (N_12166,N_10677,N_11947);
nand U12167 (N_12167,N_10623,N_11270);
and U12168 (N_12168,N_10911,N_11054);
nor U12169 (N_12169,N_11963,N_10732);
nand U12170 (N_12170,N_10785,N_10047);
or U12171 (N_12171,N_11763,N_10000);
nand U12172 (N_12172,N_10763,N_10162);
nand U12173 (N_12173,N_11477,N_11784);
xor U12174 (N_12174,N_10193,N_10239);
and U12175 (N_12175,N_10934,N_11408);
nor U12176 (N_12176,N_11139,N_11367);
and U12177 (N_12177,N_10789,N_11361);
xor U12178 (N_12178,N_10589,N_10501);
xnor U12179 (N_12179,N_10603,N_10310);
nand U12180 (N_12180,N_10697,N_11177);
xor U12181 (N_12181,N_11726,N_11606);
nand U12182 (N_12182,N_11386,N_11609);
and U12183 (N_12183,N_10643,N_11522);
xor U12184 (N_12184,N_10119,N_10706);
or U12185 (N_12185,N_10542,N_11103);
and U12186 (N_12186,N_11962,N_10043);
nand U12187 (N_12187,N_11195,N_11773);
or U12188 (N_12188,N_11695,N_11217);
nor U12189 (N_12189,N_11932,N_10071);
or U12190 (N_12190,N_10461,N_10088);
and U12191 (N_12191,N_10563,N_10422);
nor U12192 (N_12192,N_11004,N_11764);
or U12193 (N_12193,N_10906,N_11808);
or U12194 (N_12194,N_11580,N_10273);
xor U12195 (N_12195,N_11897,N_10985);
and U12196 (N_12196,N_10022,N_10937);
and U12197 (N_12197,N_10530,N_10374);
nand U12198 (N_12198,N_10463,N_11254);
nand U12199 (N_12199,N_11970,N_10153);
or U12200 (N_12200,N_10836,N_11272);
nand U12201 (N_12201,N_11057,N_11643);
and U12202 (N_12202,N_11071,N_10009);
nand U12203 (N_12203,N_10342,N_11155);
or U12204 (N_12204,N_10447,N_11241);
nor U12205 (N_12205,N_11096,N_11326);
or U12206 (N_12206,N_10629,N_11832);
and U12207 (N_12207,N_11613,N_11276);
and U12208 (N_12208,N_11729,N_10258);
or U12209 (N_12209,N_10329,N_10188);
nand U12210 (N_12210,N_11760,N_10498);
xnor U12211 (N_12211,N_11968,N_11353);
xor U12212 (N_12212,N_10835,N_11169);
xor U12213 (N_12213,N_11998,N_10656);
and U12214 (N_12214,N_11163,N_10904);
or U12215 (N_12215,N_10860,N_11511);
nand U12216 (N_12216,N_11916,N_10449);
or U12217 (N_12217,N_11721,N_10516);
xnor U12218 (N_12218,N_11637,N_10172);
or U12219 (N_12219,N_11100,N_10550);
xor U12220 (N_12220,N_11150,N_10062);
xor U12221 (N_12221,N_10314,N_10428);
xnor U12222 (N_12222,N_11119,N_11749);
xor U12223 (N_12223,N_11134,N_11830);
or U12224 (N_12224,N_10320,N_11603);
and U12225 (N_12225,N_11147,N_11926);
nand U12226 (N_12226,N_10960,N_10298);
nor U12227 (N_12227,N_11800,N_10927);
nand U12228 (N_12228,N_10928,N_11336);
nand U12229 (N_12229,N_11951,N_10752);
xor U12230 (N_12230,N_11239,N_10058);
nand U12231 (N_12231,N_10068,N_10727);
xor U12232 (N_12232,N_11099,N_10443);
xnor U12233 (N_12233,N_11870,N_11310);
and U12234 (N_12234,N_10907,N_10315);
and U12235 (N_12235,N_10935,N_10285);
or U12236 (N_12236,N_10248,N_10806);
nand U12237 (N_12237,N_11474,N_10437);
and U12238 (N_12238,N_10372,N_11332);
nor U12239 (N_12239,N_11379,N_10646);
or U12240 (N_12240,N_10481,N_10363);
nor U12241 (N_12241,N_10955,N_11253);
nor U12242 (N_12242,N_10198,N_10871);
and U12243 (N_12243,N_11173,N_11578);
nor U12244 (N_12244,N_11698,N_11790);
nand U12245 (N_12245,N_10759,N_11436);
nor U12246 (N_12246,N_10028,N_10505);
nand U12247 (N_12247,N_11788,N_10033);
and U12248 (N_12248,N_11209,N_11465);
xor U12249 (N_12249,N_10346,N_11263);
xor U12250 (N_12250,N_11208,N_10988);
nand U12251 (N_12251,N_11616,N_10947);
xor U12252 (N_12252,N_10212,N_10941);
xnor U12253 (N_12253,N_10665,N_11438);
or U12254 (N_12254,N_10160,N_11959);
or U12255 (N_12255,N_10466,N_10745);
or U12256 (N_12256,N_10526,N_11888);
nor U12257 (N_12257,N_11051,N_11913);
xnor U12258 (N_12258,N_11891,N_11991);
nand U12259 (N_12259,N_10476,N_10652);
or U12260 (N_12260,N_10251,N_10576);
or U12261 (N_12261,N_11215,N_10007);
nand U12262 (N_12262,N_10942,N_10719);
or U12263 (N_12263,N_10559,N_10858);
nand U12264 (N_12264,N_10159,N_10278);
or U12265 (N_12265,N_10855,N_11823);
nand U12266 (N_12266,N_10673,N_11440);
xor U12267 (N_12267,N_10598,N_10219);
or U12268 (N_12268,N_11958,N_11628);
and U12269 (N_12269,N_11451,N_11572);
nand U12270 (N_12270,N_11159,N_10856);
nor U12271 (N_12271,N_11219,N_11428);
nor U12272 (N_12272,N_10360,N_10850);
and U12273 (N_12273,N_10223,N_11389);
nand U12274 (N_12274,N_11536,N_10885);
or U12275 (N_12275,N_10581,N_10901);
or U12276 (N_12276,N_11385,N_11552);
or U12277 (N_12277,N_10549,N_11889);
or U12278 (N_12278,N_10249,N_11847);
nor U12279 (N_12279,N_11799,N_10511);
xnor U12280 (N_12280,N_10201,N_10133);
and U12281 (N_12281,N_11551,N_11011);
nor U12282 (N_12282,N_10820,N_10993);
and U12283 (N_12283,N_10775,N_10573);
nand U12284 (N_12284,N_11282,N_11462);
nor U12285 (N_12285,N_10366,N_11648);
nor U12286 (N_12286,N_10173,N_11638);
xnor U12287 (N_12287,N_10259,N_11988);
or U12288 (N_12288,N_11260,N_11098);
and U12289 (N_12289,N_11848,N_11064);
nand U12290 (N_12290,N_10368,N_10541);
xor U12291 (N_12291,N_10736,N_11952);
nand U12292 (N_12292,N_11550,N_11021);
xor U12293 (N_12293,N_10163,N_10566);
nand U12294 (N_12294,N_10650,N_10171);
or U12295 (N_12295,N_10458,N_10943);
xnor U12296 (N_12296,N_11316,N_10290);
xnor U12297 (N_12297,N_11171,N_11797);
nor U12298 (N_12298,N_11325,N_11783);
and U12299 (N_12299,N_11358,N_11660);
nand U12300 (N_12300,N_11469,N_10507);
nor U12301 (N_12301,N_10207,N_10100);
xor U12302 (N_12302,N_11943,N_11434);
nand U12303 (N_12303,N_11454,N_11052);
or U12304 (N_12304,N_10896,N_11266);
and U12305 (N_12305,N_10819,N_10813);
or U12306 (N_12306,N_10553,N_11657);
or U12307 (N_12307,N_10197,N_11031);
and U12308 (N_12308,N_11376,N_10699);
nor U12309 (N_12309,N_10508,N_10568);
and U12310 (N_12310,N_10867,N_10002);
nor U12311 (N_12311,N_11187,N_11344);
xnor U12312 (N_12312,N_10302,N_10883);
nand U12313 (N_12313,N_10036,N_10420);
or U12314 (N_12314,N_10210,N_10882);
and U12315 (N_12315,N_11036,N_11433);
nor U12316 (N_12316,N_10235,N_10647);
xor U12317 (N_12317,N_10349,N_10236);
or U12318 (N_12318,N_11443,N_11521);
nor U12319 (N_12319,N_11918,N_10799);
nor U12320 (N_12320,N_11074,N_10999);
and U12321 (N_12321,N_10654,N_11703);
xor U12322 (N_12322,N_10552,N_11597);
nand U12323 (N_12323,N_10817,N_10610);
xor U12324 (N_12324,N_11141,N_10831);
and U12325 (N_12325,N_11183,N_10839);
xor U12326 (N_12326,N_11457,N_11329);
or U12327 (N_12327,N_11405,N_10423);
xnor U12328 (N_12328,N_11546,N_11826);
xor U12329 (N_12329,N_10373,N_11420);
or U12330 (N_12330,N_10274,N_11682);
nor U12331 (N_12331,N_10812,N_11132);
nand U12332 (N_12332,N_11810,N_11312);
nor U12333 (N_12333,N_11982,N_10293);
nand U12334 (N_12334,N_11311,N_10967);
xor U12335 (N_12335,N_11238,N_10913);
or U12336 (N_12336,N_10108,N_11748);
nor U12337 (N_12337,N_11708,N_10204);
or U12338 (N_12338,N_10915,N_11568);
nor U12339 (N_12339,N_10684,N_11391);
and U12340 (N_12340,N_10484,N_11577);
and U12341 (N_12341,N_11149,N_10593);
xor U12342 (N_12342,N_11954,N_10308);
or U12343 (N_12343,N_11111,N_11744);
and U12344 (N_12344,N_10672,N_11138);
or U12345 (N_12345,N_11758,N_10433);
nand U12346 (N_12346,N_10945,N_11581);
nand U12347 (N_12347,N_11921,N_10011);
and U12348 (N_12348,N_11753,N_11295);
xnor U12349 (N_12349,N_11908,N_10792);
xor U12350 (N_12350,N_10205,N_10804);
xor U12351 (N_12351,N_11893,N_10010);
or U12352 (N_12352,N_10045,N_10111);
nor U12353 (N_12353,N_10253,N_11679);
nor U12354 (N_12354,N_11912,N_11730);
and U12355 (N_12355,N_11415,N_10154);
nand U12356 (N_12356,N_11600,N_11328);
nor U12357 (N_12357,N_10730,N_10863);
nor U12358 (N_12358,N_10740,N_10280);
nand U12359 (N_12359,N_10502,N_11513);
and U12360 (N_12360,N_10324,N_10371);
or U12361 (N_12361,N_11294,N_11409);
or U12362 (N_12362,N_10348,N_11005);
xor U12363 (N_12363,N_10203,N_10004);
nor U12364 (N_12364,N_11997,N_11565);
xnor U12365 (N_12365,N_11727,N_11191);
xnor U12366 (N_12366,N_10811,N_11123);
xnor U12367 (N_12367,N_10444,N_11446);
nand U12368 (N_12368,N_11432,N_11514);
xnor U12369 (N_12369,N_11633,N_11670);
nand U12370 (N_12370,N_11548,N_10440);
xnor U12371 (N_12371,N_10151,N_10178);
or U12372 (N_12372,N_11416,N_11531);
or U12373 (N_12373,N_11357,N_11145);
nor U12374 (N_12374,N_11569,N_11640);
and U12375 (N_12375,N_11224,N_10257);
nor U12376 (N_12376,N_10046,N_10523);
or U12377 (N_12377,N_11907,N_10768);
nand U12378 (N_12378,N_11402,N_11092);
nand U12379 (N_12379,N_11088,N_11291);
or U12380 (N_12380,N_11400,N_10733);
nand U12381 (N_12381,N_11965,N_11302);
nand U12382 (N_12382,N_10165,N_11579);
or U12383 (N_12383,N_10098,N_11685);
and U12384 (N_12384,N_10294,N_10184);
nor U12385 (N_12385,N_10013,N_11199);
nand U12386 (N_12386,N_11618,N_11639);
xor U12387 (N_12387,N_11337,N_10990);
nor U12388 (N_12388,N_11287,N_10532);
and U12389 (N_12389,N_11614,N_10268);
nand U12390 (N_12390,N_10729,N_11429);
nor U12391 (N_12391,N_10753,N_11162);
and U12392 (N_12392,N_10910,N_10750);
and U12393 (N_12393,N_11481,N_11558);
nand U12394 (N_12394,N_10696,N_11961);
nand U12395 (N_12395,N_10426,N_11240);
xnor U12396 (N_12396,N_10633,N_10242);
nor U12397 (N_12397,N_10535,N_10754);
and U12398 (N_12398,N_10613,N_11720);
nor U12399 (N_12399,N_10761,N_10735);
or U12400 (N_12400,N_10388,N_10520);
xor U12401 (N_12401,N_10626,N_10702);
nand U12402 (N_12402,N_11403,N_10472);
nor U12403 (N_12403,N_10359,N_11494);
xnor U12404 (N_12404,N_10261,N_10417);
and U12405 (N_12405,N_11647,N_10079);
xor U12406 (N_12406,N_11527,N_10704);
nand U12407 (N_12407,N_11075,N_11590);
xor U12408 (N_12408,N_10714,N_11452);
nand U12409 (N_12409,N_11002,N_11852);
nor U12410 (N_12410,N_10972,N_11067);
xor U12411 (N_12411,N_10287,N_10339);
xor U12412 (N_12412,N_10031,N_11879);
and U12413 (N_12413,N_11256,N_11923);
nor U12414 (N_12414,N_10232,N_10431);
nand U12415 (N_12415,N_11619,N_11274);
and U12416 (N_12416,N_11471,N_10179);
nor U12417 (N_12417,N_10884,N_11885);
and U12418 (N_12418,N_11324,N_11904);
and U12419 (N_12419,N_11269,N_11874);
nand U12420 (N_12420,N_10121,N_11168);
nor U12421 (N_12421,N_11320,N_11663);
xor U12422 (N_12422,N_10716,N_10411);
or U12423 (N_12423,N_11493,N_10297);
xnor U12424 (N_12424,N_10606,N_11082);
or U12425 (N_12425,N_11560,N_11296);
and U12426 (N_12426,N_11804,N_11375);
nor U12427 (N_12427,N_11711,N_11230);
and U12428 (N_12428,N_11012,N_10120);
nor U12429 (N_12429,N_11625,N_11101);
or U12430 (N_12430,N_10818,N_10381);
nand U12431 (N_12431,N_11843,N_11182);
and U12432 (N_12432,N_10829,N_11909);
nor U12433 (N_12433,N_11903,N_10515);
or U12434 (N_12434,N_10393,N_11079);
nor U12435 (N_12435,N_11059,N_11297);
xor U12436 (N_12436,N_10694,N_11944);
or U12437 (N_12437,N_10380,N_10634);
xor U12438 (N_12438,N_10965,N_10313);
nand U12439 (N_12439,N_10202,N_11026);
and U12440 (N_12440,N_10191,N_10131);
and U12441 (N_12441,N_11950,N_11259);
nor U12442 (N_12442,N_10521,N_11348);
xor U12443 (N_12443,N_10561,N_10106);
and U12444 (N_12444,N_11097,N_10387);
and U12445 (N_12445,N_10038,N_10144);
xnor U12446 (N_12446,N_10954,N_10514);
nor U12447 (N_12447,N_11475,N_10608);
xnor U12448 (N_12448,N_11608,N_11985);
and U12449 (N_12449,N_11937,N_11786);
nand U12450 (N_12450,N_10292,N_11978);
nand U12451 (N_12451,N_11309,N_11878);
nor U12452 (N_12452,N_10660,N_10485);
and U12453 (N_12453,N_11094,N_10586);
or U12454 (N_12454,N_10023,N_10438);
xor U12455 (N_12455,N_11724,N_11300);
nor U12456 (N_12456,N_10551,N_11086);
nand U12457 (N_12457,N_11359,N_10053);
or U12458 (N_12458,N_11770,N_11811);
and U12459 (N_12459,N_10078,N_11204);
or U12460 (N_12460,N_11264,N_11557);
or U12461 (N_12461,N_11936,N_10378);
and U12462 (N_12462,N_11321,N_10455);
and U12463 (N_12463,N_10086,N_11284);
nand U12464 (N_12464,N_11114,N_11752);
nor U12465 (N_12465,N_11019,N_11245);
nand U12466 (N_12466,N_11135,N_11896);
xnor U12467 (N_12467,N_11029,N_11652);
and U12468 (N_12468,N_11979,N_10857);
xor U12469 (N_12469,N_11419,N_10533);
or U12470 (N_12470,N_11688,N_11677);
nor U12471 (N_12471,N_10717,N_11421);
nand U12472 (N_12472,N_11915,N_10427);
nand U12473 (N_12473,N_10847,N_11427);
or U12474 (N_12474,N_10487,N_11540);
and U12475 (N_12475,N_10676,N_11496);
nor U12476 (N_12476,N_10005,N_10072);
nor U12477 (N_12477,N_11910,N_11289);
and U12478 (N_12478,N_11265,N_10164);
or U12479 (N_12479,N_10669,N_10140);
and U12480 (N_12480,N_10074,N_10575);
or U12481 (N_12481,N_10424,N_11612);
nand U12482 (N_12482,N_11710,N_11973);
nand U12483 (N_12483,N_10571,N_10361);
nor U12484 (N_12484,N_10054,N_11207);
nor U12485 (N_12485,N_11771,N_10037);
nor U12486 (N_12486,N_10030,N_11747);
and U12487 (N_12487,N_10252,N_11627);
nand U12488 (N_12488,N_11062,N_10126);
and U12489 (N_12489,N_11425,N_10311);
xnor U12490 (N_12490,N_10044,N_11884);
nand U12491 (N_12491,N_10177,N_11584);
and U12492 (N_12492,N_11136,N_11855);
nand U12493 (N_12493,N_10966,N_11439);
or U12494 (N_12494,N_10141,N_11414);
xnor U12495 (N_12495,N_11030,N_11886);
xor U12496 (N_12496,N_11805,N_11032);
nor U12497 (N_12497,N_10155,N_10246);
or U12498 (N_12498,N_10748,N_10648);
or U12499 (N_12499,N_11397,N_10658);
xor U12500 (N_12500,N_10478,N_11706);
nor U12501 (N_12501,N_11591,N_11411);
or U12502 (N_12502,N_10627,N_10852);
nor U12503 (N_12503,N_11366,N_11719);
and U12504 (N_12504,N_11304,N_11831);
nand U12505 (N_12505,N_10784,N_11396);
or U12506 (N_12506,N_11701,N_10304);
nor U12507 (N_12507,N_10611,N_10386);
nor U12508 (N_12508,N_11356,N_10157);
and U12509 (N_12509,N_11065,N_10356);
nor U12510 (N_12510,N_11362,N_10572);
nor U12511 (N_12511,N_10061,N_10116);
xor U12512 (N_12512,N_10827,N_10096);
and U12513 (N_12513,N_10087,N_10869);
nor U12514 (N_12514,N_11842,N_11288);
nand U12515 (N_12515,N_10621,N_11056);
nand U12516 (N_12516,N_11589,N_11839);
xnor U12517 (N_12517,N_11863,N_10228);
nor U12518 (N_12518,N_10332,N_11404);
xnor U12519 (N_12519,N_11084,N_10849);
nand U12520 (N_12520,N_11112,N_10113);
nor U12521 (N_12521,N_10345,N_10281);
xnor U12522 (N_12522,N_10020,N_10464);
or U12523 (N_12523,N_11486,N_11156);
xor U12524 (N_12524,N_11299,N_10441);
or U12525 (N_12525,N_11250,N_10776);
nand U12526 (N_12526,N_11060,N_10307);
xnor U12527 (N_12527,N_10263,N_11172);
and U12528 (N_12528,N_11524,N_10230);
and U12529 (N_12529,N_11315,N_10599);
nor U12530 (N_12530,N_10080,N_10951);
nand U12531 (N_12531,N_11602,N_10110);
or U12532 (N_12532,N_11461,N_10545);
nand U12533 (N_12533,N_10003,N_10987);
nand U12534 (N_12534,N_10174,N_11667);
or U12535 (N_12535,N_10490,N_11206);
or U12536 (N_12536,N_11732,N_10952);
and U12537 (N_12537,N_11468,N_11877);
nor U12538 (N_12538,N_11426,N_10012);
xor U12539 (N_12539,N_11722,N_11972);
or U12540 (N_12540,N_10607,N_11775);
xor U12541 (N_12541,N_11650,N_10338);
nor U12542 (N_12542,N_11450,N_10897);
or U12543 (N_12543,N_11331,N_10977);
nand U12544 (N_12544,N_10389,N_11003);
and U12545 (N_12545,N_11573,N_11520);
and U12546 (N_12546,N_10773,N_11330);
nand U12547 (N_12547,N_10392,N_11620);
xnor U12548 (N_12548,N_10584,N_10963);
nor U12549 (N_12549,N_11717,N_11571);
nor U12550 (N_12550,N_10722,N_10453);
or U12551 (N_12551,N_11875,N_11838);
and U12552 (N_12552,N_10834,N_10588);
or U12553 (N_12553,N_11981,N_11423);
nor U12554 (N_12554,N_11069,N_10467);
and U12555 (N_12555,N_11538,N_10326);
xnor U12556 (N_12556,N_11283,N_11516);
and U12557 (N_12557,N_11038,N_11049);
nand U12558 (N_12558,N_10094,N_11822);
nor U12559 (N_12559,N_10651,N_11738);
or U12560 (N_12560,N_11883,N_10625);
nor U12561 (N_12561,N_10042,N_10105);
nand U12562 (N_12562,N_10312,N_11598);
and U12563 (N_12563,N_11928,N_11301);
nor U12564 (N_12564,N_10112,N_11464);
and U12565 (N_12565,N_10774,N_11040);
or U12566 (N_12566,N_11817,N_11824);
or U12567 (N_12567,N_11399,N_11942);
or U12568 (N_12568,N_11467,N_11906);
nand U12569 (N_12569,N_10325,N_10077);
nor U12570 (N_12570,N_10932,N_10208);
nor U12571 (N_12571,N_10964,N_10565);
nor U12572 (N_12572,N_10616,N_10385);
and U12573 (N_12573,N_10457,N_10524);
and U12574 (N_12574,N_10786,N_10482);
or U12575 (N_12575,N_10630,N_11107);
nand U12576 (N_12576,N_10838,N_10284);
nand U12577 (N_12577,N_11993,N_11745);
nor U12578 (N_12578,N_11994,N_10486);
and U12579 (N_12579,N_11574,N_11683);
and U12580 (N_12580,N_11739,N_11078);
xnor U12581 (N_12581,N_10936,N_11549);
xor U12582 (N_12582,N_11341,N_10653);
nand U12583 (N_12583,N_10218,N_11242);
xor U12584 (N_12584,N_11037,N_10180);
nor U12585 (N_12585,N_10612,N_11372);
nor U12586 (N_12586,N_10796,N_11636);
nor U12587 (N_12587,N_10851,N_10846);
nor U12588 (N_12588,N_11292,N_11407);
or U12589 (N_12589,N_10262,N_10868);
xnor U12590 (N_12590,N_10309,N_11193);
xor U12591 (N_12591,N_10412,N_10525);
and U12592 (N_12592,N_10139,N_11890);
or U12593 (N_12593,N_11125,N_10409);
nand U12594 (N_12594,N_10830,N_11892);
nor U12595 (N_12595,N_11791,N_10032);
xnor U12596 (N_12596,N_11216,N_10639);
nand U12597 (N_12597,N_10496,N_10700);
and U12598 (N_12598,N_10751,N_10680);
nor U12599 (N_12599,N_11179,N_11435);
nand U12600 (N_12600,N_10922,N_11165);
and U12601 (N_12601,N_11833,N_10452);
and U12602 (N_12602,N_11006,N_10953);
or U12603 (N_12603,N_10892,N_11448);
nor U12604 (N_12604,N_11723,N_10635);
and U12605 (N_12605,N_10544,N_10637);
and U12606 (N_12606,N_11599,N_10473);
and U12607 (N_12607,N_10918,N_10543);
and U12608 (N_12608,N_11161,N_11894);
xor U12609 (N_12609,N_10760,N_11203);
xor U12610 (N_12610,N_11774,N_10234);
and U12611 (N_12611,N_10056,N_11999);
and U12612 (N_12612,N_11792,N_11129);
xor U12613 (N_12613,N_10136,N_10919);
or U12614 (N_12614,N_11676,N_10728);
nor U12615 (N_12615,N_11034,N_10644);
nand U12616 (N_12616,N_10196,N_10888);
nand U12617 (N_12617,N_10828,N_11345);
and U12618 (N_12618,N_10794,N_10147);
or U12619 (N_12619,N_11691,N_11690);
nor U12620 (N_12620,N_11085,N_11307);
nor U12621 (N_12621,N_11277,N_10189);
or U12622 (N_12622,N_10343,N_10394);
and U12623 (N_12623,N_11213,N_11463);
nor U12624 (N_12624,N_11675,N_10241);
nor U12625 (N_12625,N_10414,N_10837);
nand U12626 (N_12626,N_10995,N_10026);
or U12627 (N_12627,N_10041,N_11681);
and U12628 (N_12628,N_11969,N_10889);
nor U12629 (N_12629,N_11526,N_10275);
or U12630 (N_12630,N_10803,N_11525);
or U12631 (N_12631,N_10582,N_11507);
xor U12632 (N_12632,N_11045,N_11777);
or U12633 (N_12633,N_10103,N_11068);
nand U12634 (N_12634,N_11705,N_10034);
nand U12635 (N_12635,N_10845,N_11455);
nand U12636 (N_12636,N_10152,N_10469);
nor U12637 (N_12637,N_11501,N_11354);
nor U12638 (N_12638,N_10353,N_11176);
xor U12639 (N_12639,N_11919,N_11873);
or U12640 (N_12640,N_11202,N_11793);
or U12641 (N_12641,N_11271,N_10186);
xnor U12642 (N_12642,N_11547,N_11158);
nand U12643 (N_12643,N_10247,N_10674);
xnor U12644 (N_12644,N_10479,N_10291);
xnor U12645 (N_12645,N_10790,N_10224);
or U12646 (N_12646,N_11081,N_10450);
or U12647 (N_12647,N_10451,N_10711);
or U12648 (N_12648,N_10592,N_11816);
nand U12649 (N_12649,N_11058,N_10642);
xnor U12650 (N_12650,N_10430,N_10833);
nor U12651 (N_12651,N_11806,N_10276);
xnor U12652 (N_12652,N_10407,N_11911);
and U12653 (N_12653,N_10659,N_10707);
nor U12654 (N_12654,N_11860,N_10862);
and U12655 (N_12655,N_10421,N_10666);
or U12656 (N_12656,N_10930,N_10570);
nor U12657 (N_12657,N_10548,N_11895);
nor U12658 (N_12658,N_10170,N_10425);
nor U12659 (N_12659,N_11990,N_11837);
xor U12660 (N_12660,N_11343,N_10279);
xor U12661 (N_12661,N_10471,N_11866);
xor U12662 (N_12662,N_11743,N_11363);
and U12663 (N_12663,N_10878,N_11704);
nand U12664 (N_12664,N_10705,N_10240);
nand U12665 (N_12665,N_11234,N_10853);
xor U12666 (N_12666,N_10764,N_10950);
nand U12667 (N_12667,N_10333,N_10970);
nand U12668 (N_12668,N_10317,N_10395);
nand U12669 (N_12669,N_11497,N_10076);
nor U12670 (N_12670,N_11106,N_11715);
xor U12671 (N_12671,N_11110,N_10306);
and U12672 (N_12672,N_10554,N_10397);
and U12673 (N_12673,N_10893,N_10128);
nand U12674 (N_12674,N_10703,N_11373);
or U12675 (N_12675,N_10564,N_11914);
nand U12676 (N_12676,N_10340,N_10084);
xor U12677 (N_12677,N_11128,N_10305);
or U12678 (N_12678,N_11042,N_11917);
xnor U12679 (N_12679,N_10866,N_10456);
nor U12680 (N_12680,N_11459,N_11787);
xor U12681 (N_12681,N_10879,N_11766);
xor U12682 (N_12682,N_11555,N_11898);
nor U12683 (N_12683,N_11413,N_11955);
or U12684 (N_12684,N_10980,N_11072);
or U12685 (N_12685,N_11095,N_11821);
and U12686 (N_12686,N_11382,N_10619);
nor U12687 (N_12687,N_11148,N_10376);
nand U12688 (N_12688,N_10269,N_11133);
xor U12689 (N_12689,N_10176,N_10841);
xnor U12690 (N_12690,N_10206,N_10555);
nand U12691 (N_12691,N_10747,N_11535);
nand U12692 (N_12692,N_11010,N_11566);
nand U12693 (N_12693,N_11562,N_11255);
nor U12694 (N_12694,N_11105,N_10746);
nand U12695 (N_12695,N_11953,N_11305);
and U12696 (N_12696,N_11740,N_10810);
or U12697 (N_12697,N_10107,N_11779);
nand U12698 (N_12698,N_11622,N_10698);
nor U12699 (N_12699,N_10978,N_11251);
xor U12700 (N_12700,N_11001,N_10085);
nor U12701 (N_12701,N_11940,N_11957);
nor U12702 (N_12702,N_11043,N_11528);
nand U12703 (N_12703,N_10460,N_10114);
and U12704 (N_12704,N_10981,N_11554);
nor U12705 (N_12705,N_10825,N_10390);
nand U12706 (N_12706,N_10917,N_11181);
xnor U12707 (N_12707,N_10404,N_10587);
nand U12708 (N_12708,N_10874,N_10567);
or U12709 (N_12709,N_11152,N_10881);
nor U12710 (N_12710,N_10493,N_10328);
xor U12711 (N_12711,N_11635,N_11925);
xnor U12712 (N_12712,N_11621,N_11184);
xnor U12713 (N_12713,N_11671,N_10492);
and U12714 (N_12714,N_10436,N_10093);
xor U12715 (N_12715,N_10419,N_11610);
and U12716 (N_12716,N_10923,N_11381);
or U12717 (N_12717,N_11190,N_10016);
xor U12718 (N_12718,N_11458,N_11472);
and U12719 (N_12719,N_11564,N_10876);
and U12720 (N_12720,N_10459,N_10749);
or U12721 (N_12721,N_10413,N_11449);
nand U12722 (N_12722,N_11956,N_10143);
or U12723 (N_12723,N_10135,N_11137);
xor U12724 (N_12724,N_11583,N_10519);
and U12725 (N_12725,N_10738,N_11000);
xor U12726 (N_12726,N_10350,N_10908);
nand U12727 (N_12727,N_10055,N_10843);
and U12728 (N_12728,N_10962,N_10720);
xnor U12729 (N_12729,N_10756,N_11899);
and U12730 (N_12730,N_11882,N_11757);
xnor U12731 (N_12731,N_10758,N_10182);
or U12732 (N_12732,N_10090,N_10823);
or U12733 (N_12733,N_11871,N_11160);
or U12734 (N_12734,N_11124,N_10265);
or U12735 (N_12735,N_11927,N_11490);
nor U12736 (N_12736,N_10824,N_10912);
nand U12737 (N_12737,N_10442,N_11960);
or U12738 (N_12738,N_11934,N_10006);
nor U12739 (N_12739,N_10104,N_11851);
nand U12740 (N_12740,N_11167,N_11751);
or U12741 (N_12741,N_10398,N_11063);
nand U12742 (N_12742,N_11876,N_11201);
nor U12743 (N_12743,N_10602,N_10415);
xor U12744 (N_12744,N_10991,N_10019);
and U12745 (N_12745,N_11900,N_10282);
nor U12746 (N_12746,N_11728,N_11226);
nor U12747 (N_12747,N_11083,N_11117);
or U12748 (N_12748,N_11818,N_11519);
xnor U12749 (N_12749,N_11933,N_10992);
or U12750 (N_12750,N_10780,N_10064);
xor U12751 (N_12751,N_10370,N_11601);
and U12752 (N_12752,N_11360,N_10641);
and U12753 (N_12753,N_11115,N_11733);
nor U12754 (N_12754,N_11016,N_11700);
and U12755 (N_12755,N_11205,N_10734);
or U12756 (N_12756,N_11055,N_11355);
xnor U12757 (N_12757,N_11754,N_10894);
nor U12758 (N_12758,N_11441,N_10445);
nand U12759 (N_12759,N_10303,N_11901);
xnor U12760 (N_12760,N_11967,N_11624);
and U12761 (N_12761,N_11864,N_11975);
or U12762 (N_12762,N_10583,N_11869);
xor U12763 (N_12763,N_11707,N_11862);
and U12764 (N_12764,N_11410,N_11746);
nor U12765 (N_12765,N_11575,N_11500);
nor U12766 (N_12766,N_10283,N_10008);
nor U12767 (N_12767,N_10410,N_10574);
nand U12768 (N_12768,N_10215,N_11834);
nor U12769 (N_12769,N_10900,N_11798);
xnor U12770 (N_12770,N_11127,N_10921);
and U12771 (N_12771,N_10399,N_11984);
xnor U12772 (N_12772,N_11185,N_10238);
xor U12773 (N_12773,N_10365,N_10726);
or U12774 (N_12774,N_10788,N_10049);
nor U12775 (N_12775,N_10319,N_11476);
xnor U12776 (N_12776,N_10891,N_11537);
nor U12777 (N_12777,N_10840,N_11803);
nor U12778 (N_12778,N_10795,N_11273);
nand U12779 (N_12779,N_10909,N_11634);
nor U12780 (N_12780,N_11333,N_10682);
or U12781 (N_12781,N_10403,N_11759);
and U12782 (N_12782,N_11840,N_10590);
or U12783 (N_12783,N_11789,N_11076);
or U12784 (N_12784,N_11587,N_11782);
or U12785 (N_12785,N_10506,N_11090);
and U12786 (N_12786,N_11796,N_11286);
and U12787 (N_12787,N_10640,N_11080);
or U12788 (N_12788,N_10661,N_11750);
xnor U12789 (N_12789,N_11247,N_11370);
and U12790 (N_12790,N_10220,N_10383);
nor U12791 (N_12791,N_10986,N_11992);
or U12792 (N_12792,N_11017,N_10245);
nand U12793 (N_12793,N_10529,N_10264);
nand U12794 (N_12794,N_10367,N_11174);
nor U12795 (N_12795,N_10156,N_11971);
nor U12796 (N_12796,N_10609,N_11220);
nand U12797 (N_12797,N_11418,N_10865);
and U12798 (N_12798,N_11920,N_11053);
nor U12799 (N_12799,N_11518,N_10018);
and U12800 (N_12800,N_11368,N_10214);
and U12801 (N_12801,N_11819,N_10982);
nand U12802 (N_12802,N_10027,N_11529);
or U12803 (N_12803,N_11314,N_10330);
and U12804 (N_12804,N_10822,N_10663);
or U12805 (N_12805,N_10832,N_11484);
xor U12806 (N_12806,N_10405,N_11488);
nand U12807 (N_12807,N_10757,N_11666);
nor U12808 (N_12808,N_10024,N_11515);
xnor U12809 (N_12809,N_10092,N_10807);
or U12810 (N_12810,N_11858,N_10091);
nand U12811 (N_12811,N_11737,N_10097);
or U12812 (N_12812,N_10194,N_11279);
or U12813 (N_12813,N_11140,N_10801);
or U12814 (N_12814,N_11258,N_10675);
nor U12815 (N_12815,N_10429,N_10983);
nand U12816 (N_12816,N_11422,N_10710);
xor U12817 (N_12817,N_10712,N_11709);
nor U12818 (N_12818,N_10369,N_11595);
nor U12819 (N_12819,N_10254,N_11630);
nor U12820 (N_12820,N_11007,N_11478);
or U12821 (N_12821,N_10861,N_11398);
and U12822 (N_12822,N_10075,N_10522);
or U12823 (N_12823,N_11850,N_10693);
nor U12824 (N_12824,N_11303,N_11008);
nor U12825 (N_12825,N_11680,N_11322);
or U12826 (N_12826,N_10494,N_10181);
xor U12827 (N_12827,N_11563,N_10692);
or U12828 (N_12828,N_11857,N_11801);
nand U12829 (N_12829,N_11861,N_10678);
or U12830 (N_12830,N_10161,N_11539);
xor U12831 (N_12831,N_10528,N_11070);
nor U12832 (N_12832,N_10142,N_11814);
nor U12833 (N_12833,N_11966,N_11146);
xnor U12834 (N_12834,N_10334,N_11694);
xor U12835 (N_12835,N_10931,N_10468);
and U12836 (N_12836,N_11659,N_11487);
xor U12837 (N_12837,N_10890,N_11093);
nand U12838 (N_12838,N_10169,N_11702);
xor U12839 (N_12839,N_10418,N_10821);
nand U12840 (N_12840,N_11377,N_11532);
nor U12841 (N_12841,N_11713,N_11233);
or U12842 (N_12842,N_10979,N_10130);
and U12843 (N_12843,N_11673,N_11859);
nand U12844 (N_12844,N_10944,N_10994);
and U12845 (N_12845,N_10920,N_11604);
and U12846 (N_12846,N_10167,N_11118);
nor U12847 (N_12847,N_11229,N_10512);
nor U12848 (N_12848,N_11809,N_11534);
nor U12849 (N_12849,N_10183,N_10579);
or U12850 (N_12850,N_10500,N_10237);
and U12851 (N_12851,N_10631,N_11553);
xnor U12852 (N_12852,N_11556,N_11902);
and U12853 (N_12853,N_10465,N_10844);
or U12854 (N_12854,N_11334,N_10743);
xnor U12855 (N_12855,N_11931,N_10815);
or U12856 (N_12856,N_10102,N_11678);
nand U12857 (N_12857,N_11188,N_10396);
and U12858 (N_12858,N_10808,N_11369);
nor U12859 (N_12859,N_10600,N_10226);
or U12860 (N_12860,N_10272,N_11154);
xor U12861 (N_12861,N_10243,N_11020);
and U12862 (N_12862,N_10187,N_10231);
or U12863 (N_12863,N_11543,N_11989);
nand U12864 (N_12864,N_11949,N_10546);
nor U12865 (N_12865,N_11506,N_11846);
or U12866 (N_12866,N_11275,N_10957);
or U12867 (N_12867,N_11218,N_10488);
or U12868 (N_12868,N_10594,N_11523);
or U12869 (N_12869,N_11510,N_10762);
xor U12870 (N_12870,N_10229,N_11854);
xor U12871 (N_12871,N_10327,N_11668);
nor U12872 (N_12872,N_10089,N_10124);
nand U12873 (N_12873,N_10596,N_10344);
or U12874 (N_12874,N_11835,N_10605);
xnor U12875 (N_12875,N_11180,N_11544);
nor U12876 (N_12876,N_10432,N_10267);
xor U12877 (N_12877,N_10168,N_10132);
nor U12878 (N_12878,N_10035,N_11027);
nand U12879 (N_12879,N_10558,N_10382);
and U12880 (N_12880,N_10791,N_10331);
nand U12881 (N_12881,N_11164,N_11120);
xnor U12882 (N_12882,N_11384,N_11394);
or U12883 (N_12883,N_11795,N_11089);
and U12884 (N_12884,N_11815,N_11785);
nand U12885 (N_12885,N_11170,N_10537);
nor U12886 (N_12886,N_10713,N_11351);
nand U12887 (N_12887,N_10211,N_11996);
nor U12888 (N_12888,N_11930,N_11505);
xor U12889 (N_12889,N_11987,N_11262);
or U12890 (N_12890,N_11232,N_11689);
xor U12891 (N_12891,N_11489,N_11130);
nor U12892 (N_12892,N_10250,N_11364);
xor U12893 (N_12893,N_10872,N_11588);
xor U12894 (N_12894,N_11504,N_10448);
and U12895 (N_12895,N_10192,N_11664);
xnor U12896 (N_12896,N_11228,N_11512);
or U12897 (N_12897,N_11781,N_10949);
or U12898 (N_12898,N_11594,N_11175);
and U12899 (N_12899,N_10688,N_10065);
nor U12900 (N_12900,N_11144,N_10354);
or U12901 (N_12901,N_11669,N_10527);
nand U12902 (N_12902,N_10638,N_10217);
xnor U12903 (N_12903,N_11559,N_11825);
and U12904 (N_12904,N_10783,N_11460);
and U12905 (N_12905,N_11091,N_11935);
nor U12906 (N_12906,N_11383,N_11395);
or U12907 (N_12907,N_11644,N_10474);
nor U12908 (N_12908,N_11466,N_11293);
nor U12909 (N_12909,N_11186,N_11050);
or U12910 (N_12910,N_10929,N_11887);
and U12911 (N_12911,N_11731,N_11048);
nand U12912 (N_12912,N_10489,N_11041);
nand U12913 (N_12913,N_10322,N_10887);
or U12914 (N_12914,N_10715,N_11503);
and U12915 (N_12915,N_10933,N_10039);
nor U12916 (N_12916,N_10518,N_10679);
or U12917 (N_12917,N_10577,N_10318);
nor U12918 (N_12918,N_11674,N_11517);
nand U12919 (N_12919,N_11716,N_11868);
or U12920 (N_12920,N_10351,N_11257);
nand U12921 (N_12921,N_10859,N_10299);
xor U12922 (N_12922,N_11025,N_11014);
nor U12923 (N_12923,N_10070,N_10798);
and U12924 (N_12924,N_10683,N_10765);
xnor U12925 (N_12925,N_11290,N_10337);
nor U12926 (N_12926,N_10146,N_11166);
xnor U12927 (N_12927,N_11735,N_10615);
or U12928 (N_12928,N_11844,N_10976);
xor U12929 (N_12929,N_11211,N_11498);
and U12930 (N_12930,N_10213,N_11431);
nand U12931 (N_12931,N_11615,N_10898);
nand U12932 (N_12932,N_10667,N_10617);
nor U12933 (N_12933,N_10961,N_10470);
nand U12934 (N_12934,N_11349,N_11456);
xnor U12935 (N_12935,N_11066,N_11108);
nor U12936 (N_12936,N_10379,N_11617);
xor U12937 (N_12937,N_11741,N_10122);
and U12938 (N_12938,N_10095,N_10664);
nor U12939 (N_12939,N_10357,N_11828);
nand U12940 (N_12940,N_11378,N_10377);
nor U12941 (N_12941,N_10886,N_11687);
and U12942 (N_12942,N_11767,N_11236);
and U12943 (N_12943,N_11087,N_11200);
and U12944 (N_12944,N_11697,N_11212);
nand U12945 (N_12945,N_11631,N_11237);
nand U12946 (N_12946,N_11335,N_10958);
or U12947 (N_12947,N_10842,N_10725);
nor U12948 (N_12948,N_10109,N_11865);
and U12949 (N_12949,N_11342,N_10873);
nor U12950 (N_12950,N_11794,N_11827);
xnor U12951 (N_12951,N_11585,N_11645);
nand U12952 (N_12952,N_11561,N_10701);
nand U12953 (N_12953,N_10175,N_10739);
xnor U12954 (N_12954,N_11350,N_10256);
xnor U12955 (N_12955,N_11340,N_11686);
nor U12956 (N_12956,N_10755,N_11502);
xnor U12957 (N_12957,N_11327,N_10051);
and U12958 (N_12958,N_10497,N_10689);
and U12959 (N_12959,N_10435,N_11044);
and U12960 (N_12960,N_10848,N_10989);
xor U12961 (N_12961,N_10118,N_10926);
xnor U12962 (N_12962,N_10358,N_11945);
and U12963 (N_12963,N_10296,N_11995);
and U12964 (N_12964,N_11380,N_10475);
and U12965 (N_12965,N_11545,N_11772);
nor U12966 (N_12966,N_10899,N_10509);
xor U12967 (N_12967,N_11104,N_11231);
or U12968 (N_12968,N_11323,N_11807);
nand U12969 (N_12969,N_10769,N_10503);
nor U12970 (N_12970,N_10973,N_11768);
and U12971 (N_12971,N_11013,N_11693);
nor U12972 (N_12972,N_10401,N_10517);
and U12973 (N_12973,N_11658,N_11881);
or U12974 (N_12974,N_11607,N_11986);
xnor U12975 (N_12975,N_11424,N_10662);
nand U12976 (N_12976,N_11196,N_11983);
or U12977 (N_12977,N_11444,N_10513);
or U12978 (N_12978,N_10601,N_11845);
or U12979 (N_12979,N_10295,N_10270);
and U12980 (N_12980,N_10655,N_10578);
nand U12981 (N_12981,N_10137,N_11948);
nor U12982 (N_12982,N_11755,N_11853);
nor U12983 (N_12983,N_11653,N_11836);
or U12984 (N_12984,N_10767,N_10446);
nand U12985 (N_12985,N_11189,N_11178);
xor U12986 (N_12986,N_11623,N_10190);
xor U12987 (N_12987,N_10797,N_11974);
nand U12988 (N_12988,N_10974,N_10123);
xnor U12989 (N_12989,N_11210,N_11223);
xnor U12990 (N_12990,N_11318,N_10718);
nand U12991 (N_12991,N_11508,N_11736);
nand U12992 (N_12992,N_10017,N_10321);
nand U12993 (N_12993,N_11672,N_11268);
or U12994 (N_12994,N_11308,N_10025);
and U12995 (N_12995,N_11371,N_10271);
nand U12996 (N_12996,N_10914,N_11596);
and U12997 (N_12997,N_11780,N_10975);
or U12998 (N_12998,N_10029,N_11039);
and U12999 (N_12999,N_11714,N_10402);
nor U13000 (N_13000,N_11277,N_10731);
and U13001 (N_13001,N_11277,N_10101);
and U13002 (N_13002,N_10582,N_11715);
or U13003 (N_13003,N_11089,N_10509);
and U13004 (N_13004,N_11085,N_11973);
and U13005 (N_13005,N_10555,N_11153);
nand U13006 (N_13006,N_10358,N_10871);
xnor U13007 (N_13007,N_10552,N_10167);
or U13008 (N_13008,N_10048,N_11425);
xnor U13009 (N_13009,N_10127,N_11087);
nand U13010 (N_13010,N_10935,N_11473);
nand U13011 (N_13011,N_10209,N_11844);
nor U13012 (N_13012,N_11953,N_11939);
nand U13013 (N_13013,N_10987,N_11421);
nor U13014 (N_13014,N_10411,N_10576);
xor U13015 (N_13015,N_11634,N_11837);
and U13016 (N_13016,N_11330,N_11646);
nand U13017 (N_13017,N_11213,N_10574);
xnor U13018 (N_13018,N_11807,N_11914);
xor U13019 (N_13019,N_11219,N_11030);
nand U13020 (N_13020,N_10811,N_11436);
or U13021 (N_13021,N_11364,N_11816);
xnor U13022 (N_13022,N_10390,N_11674);
and U13023 (N_13023,N_11166,N_10308);
and U13024 (N_13024,N_11876,N_10329);
xnor U13025 (N_13025,N_10776,N_10872);
xor U13026 (N_13026,N_10715,N_10580);
xnor U13027 (N_13027,N_10070,N_11413);
or U13028 (N_13028,N_10681,N_10733);
nand U13029 (N_13029,N_10477,N_10414);
and U13030 (N_13030,N_10290,N_11620);
and U13031 (N_13031,N_11015,N_11603);
and U13032 (N_13032,N_11029,N_11910);
and U13033 (N_13033,N_10588,N_10250);
or U13034 (N_13034,N_10402,N_11895);
and U13035 (N_13035,N_10188,N_11174);
nor U13036 (N_13036,N_10264,N_10002);
nand U13037 (N_13037,N_10161,N_10232);
nor U13038 (N_13038,N_11735,N_11175);
and U13039 (N_13039,N_10631,N_10132);
nand U13040 (N_13040,N_11556,N_11885);
or U13041 (N_13041,N_11987,N_11261);
xor U13042 (N_13042,N_10780,N_10346);
and U13043 (N_13043,N_10448,N_10105);
and U13044 (N_13044,N_10618,N_11714);
nand U13045 (N_13045,N_10778,N_11709);
nor U13046 (N_13046,N_10719,N_11802);
or U13047 (N_13047,N_11000,N_10268);
xor U13048 (N_13048,N_10262,N_11421);
nand U13049 (N_13049,N_10468,N_10698);
or U13050 (N_13050,N_11765,N_10022);
xnor U13051 (N_13051,N_11083,N_11329);
xor U13052 (N_13052,N_10000,N_11153);
and U13053 (N_13053,N_10912,N_11424);
and U13054 (N_13054,N_11728,N_11912);
nor U13055 (N_13055,N_11313,N_10385);
nor U13056 (N_13056,N_10775,N_11817);
nand U13057 (N_13057,N_11281,N_10199);
or U13058 (N_13058,N_11658,N_11740);
nand U13059 (N_13059,N_11050,N_10128);
nand U13060 (N_13060,N_11752,N_10567);
and U13061 (N_13061,N_11565,N_10298);
or U13062 (N_13062,N_11691,N_10265);
xor U13063 (N_13063,N_10914,N_10377);
and U13064 (N_13064,N_10439,N_10001);
or U13065 (N_13065,N_11931,N_11941);
nor U13066 (N_13066,N_10726,N_11514);
or U13067 (N_13067,N_10837,N_11404);
and U13068 (N_13068,N_10666,N_10879);
and U13069 (N_13069,N_11362,N_10310);
nor U13070 (N_13070,N_10249,N_10282);
nor U13071 (N_13071,N_11277,N_10606);
nand U13072 (N_13072,N_11487,N_10294);
or U13073 (N_13073,N_11373,N_10728);
or U13074 (N_13074,N_11371,N_11692);
nor U13075 (N_13075,N_11974,N_11133);
nor U13076 (N_13076,N_10530,N_11097);
nor U13077 (N_13077,N_10719,N_11957);
or U13078 (N_13078,N_10437,N_11531);
nand U13079 (N_13079,N_10744,N_11487);
nand U13080 (N_13080,N_11304,N_11820);
or U13081 (N_13081,N_11993,N_10184);
nor U13082 (N_13082,N_10362,N_10357);
nand U13083 (N_13083,N_10961,N_10726);
nand U13084 (N_13084,N_10622,N_11648);
xnor U13085 (N_13085,N_10538,N_10641);
nand U13086 (N_13086,N_11396,N_10289);
or U13087 (N_13087,N_10675,N_10732);
and U13088 (N_13088,N_10922,N_10239);
nand U13089 (N_13089,N_11586,N_11123);
or U13090 (N_13090,N_10734,N_10927);
and U13091 (N_13091,N_11105,N_11828);
or U13092 (N_13092,N_10449,N_11003);
nor U13093 (N_13093,N_10808,N_11092);
nor U13094 (N_13094,N_11903,N_11512);
or U13095 (N_13095,N_10377,N_10667);
or U13096 (N_13096,N_11120,N_11489);
nor U13097 (N_13097,N_11158,N_11152);
xor U13098 (N_13098,N_11286,N_11945);
and U13099 (N_13099,N_10364,N_11605);
nor U13100 (N_13100,N_11428,N_10184);
nor U13101 (N_13101,N_10257,N_10190);
or U13102 (N_13102,N_10866,N_11041);
and U13103 (N_13103,N_10746,N_11692);
or U13104 (N_13104,N_11382,N_10452);
and U13105 (N_13105,N_10191,N_11310);
nor U13106 (N_13106,N_10520,N_11334);
or U13107 (N_13107,N_11281,N_11365);
or U13108 (N_13108,N_10725,N_10853);
nand U13109 (N_13109,N_11029,N_10084);
and U13110 (N_13110,N_10932,N_11489);
nand U13111 (N_13111,N_11826,N_11326);
nand U13112 (N_13112,N_11661,N_11200);
or U13113 (N_13113,N_11783,N_10765);
xnor U13114 (N_13114,N_10178,N_10779);
nand U13115 (N_13115,N_11233,N_10702);
and U13116 (N_13116,N_10036,N_11312);
nand U13117 (N_13117,N_10817,N_10250);
or U13118 (N_13118,N_11669,N_10409);
or U13119 (N_13119,N_10890,N_11933);
or U13120 (N_13120,N_10718,N_11415);
or U13121 (N_13121,N_10890,N_10733);
nand U13122 (N_13122,N_11255,N_10569);
nor U13123 (N_13123,N_10580,N_11368);
xor U13124 (N_13124,N_11710,N_10393);
nor U13125 (N_13125,N_10269,N_10936);
nor U13126 (N_13126,N_11287,N_11490);
nor U13127 (N_13127,N_10333,N_10753);
or U13128 (N_13128,N_11164,N_11073);
xor U13129 (N_13129,N_11460,N_10854);
xor U13130 (N_13130,N_10624,N_11172);
or U13131 (N_13131,N_11283,N_11052);
and U13132 (N_13132,N_11138,N_11715);
xnor U13133 (N_13133,N_11269,N_11214);
and U13134 (N_13134,N_11570,N_11754);
xnor U13135 (N_13135,N_11196,N_11369);
nand U13136 (N_13136,N_11959,N_10646);
nor U13137 (N_13137,N_10562,N_10426);
and U13138 (N_13138,N_10683,N_11581);
nor U13139 (N_13139,N_11298,N_10585);
and U13140 (N_13140,N_11630,N_10367);
and U13141 (N_13141,N_10890,N_10793);
nor U13142 (N_13142,N_10276,N_11668);
or U13143 (N_13143,N_10018,N_10942);
nor U13144 (N_13144,N_11779,N_11705);
nand U13145 (N_13145,N_11386,N_10407);
or U13146 (N_13146,N_10798,N_10698);
and U13147 (N_13147,N_10326,N_11556);
xor U13148 (N_13148,N_10650,N_10750);
and U13149 (N_13149,N_10037,N_10114);
or U13150 (N_13150,N_10913,N_10993);
or U13151 (N_13151,N_10935,N_10724);
xnor U13152 (N_13152,N_10135,N_11980);
or U13153 (N_13153,N_11760,N_11977);
nor U13154 (N_13154,N_11566,N_11280);
xor U13155 (N_13155,N_10702,N_10573);
nor U13156 (N_13156,N_11418,N_10075);
nor U13157 (N_13157,N_10009,N_11475);
nand U13158 (N_13158,N_11407,N_11659);
nor U13159 (N_13159,N_10026,N_11647);
or U13160 (N_13160,N_10282,N_10727);
and U13161 (N_13161,N_11038,N_10096);
xor U13162 (N_13162,N_11547,N_10830);
or U13163 (N_13163,N_11177,N_10850);
nor U13164 (N_13164,N_11204,N_10427);
or U13165 (N_13165,N_10407,N_11465);
nand U13166 (N_13166,N_11749,N_10215);
xnor U13167 (N_13167,N_11817,N_11807);
and U13168 (N_13168,N_11993,N_11305);
nand U13169 (N_13169,N_10375,N_11218);
xor U13170 (N_13170,N_11081,N_10454);
nor U13171 (N_13171,N_10605,N_10166);
nor U13172 (N_13172,N_10681,N_10617);
nand U13173 (N_13173,N_10958,N_11120);
and U13174 (N_13174,N_10376,N_11704);
nand U13175 (N_13175,N_11463,N_10021);
nor U13176 (N_13176,N_10277,N_11432);
nor U13177 (N_13177,N_10009,N_10769);
nor U13178 (N_13178,N_10330,N_10518);
or U13179 (N_13179,N_10797,N_10473);
xnor U13180 (N_13180,N_10177,N_11630);
nor U13181 (N_13181,N_10137,N_10617);
nand U13182 (N_13182,N_10377,N_10219);
nor U13183 (N_13183,N_10917,N_11801);
nand U13184 (N_13184,N_10574,N_11684);
nand U13185 (N_13185,N_10508,N_11927);
nand U13186 (N_13186,N_10060,N_10189);
xnor U13187 (N_13187,N_11804,N_11646);
xnor U13188 (N_13188,N_10051,N_11000);
nand U13189 (N_13189,N_10993,N_11796);
xnor U13190 (N_13190,N_10064,N_11045);
and U13191 (N_13191,N_10113,N_11186);
nand U13192 (N_13192,N_11837,N_10718);
or U13193 (N_13193,N_11748,N_11933);
nand U13194 (N_13194,N_10347,N_10644);
nand U13195 (N_13195,N_10033,N_11027);
nand U13196 (N_13196,N_11727,N_11175);
or U13197 (N_13197,N_11409,N_10727);
and U13198 (N_13198,N_10779,N_10408);
nor U13199 (N_13199,N_11672,N_10659);
nor U13200 (N_13200,N_10390,N_11228);
or U13201 (N_13201,N_10803,N_11713);
nand U13202 (N_13202,N_10558,N_11663);
or U13203 (N_13203,N_10196,N_11036);
and U13204 (N_13204,N_11494,N_11768);
or U13205 (N_13205,N_10833,N_10032);
and U13206 (N_13206,N_10356,N_10881);
nand U13207 (N_13207,N_11576,N_10486);
and U13208 (N_13208,N_11543,N_10869);
nor U13209 (N_13209,N_11827,N_10264);
xor U13210 (N_13210,N_10515,N_10774);
nand U13211 (N_13211,N_10386,N_11457);
nand U13212 (N_13212,N_10694,N_11616);
and U13213 (N_13213,N_11415,N_11468);
or U13214 (N_13214,N_10557,N_11574);
and U13215 (N_13215,N_11640,N_11036);
xor U13216 (N_13216,N_11984,N_11174);
or U13217 (N_13217,N_11265,N_10074);
or U13218 (N_13218,N_11782,N_10049);
or U13219 (N_13219,N_10438,N_11892);
nor U13220 (N_13220,N_10595,N_10766);
and U13221 (N_13221,N_11901,N_11447);
xor U13222 (N_13222,N_10049,N_11097);
xor U13223 (N_13223,N_10774,N_11669);
and U13224 (N_13224,N_10640,N_11734);
nor U13225 (N_13225,N_11613,N_11679);
or U13226 (N_13226,N_11866,N_10810);
xor U13227 (N_13227,N_10964,N_11403);
nand U13228 (N_13228,N_11436,N_10040);
xnor U13229 (N_13229,N_10549,N_10425);
and U13230 (N_13230,N_11466,N_11610);
or U13231 (N_13231,N_11442,N_11546);
xnor U13232 (N_13232,N_11754,N_11911);
nor U13233 (N_13233,N_10053,N_10709);
nand U13234 (N_13234,N_11455,N_10094);
and U13235 (N_13235,N_11983,N_11990);
nand U13236 (N_13236,N_10978,N_10966);
nand U13237 (N_13237,N_10982,N_11161);
and U13238 (N_13238,N_10295,N_11023);
or U13239 (N_13239,N_10488,N_10020);
nor U13240 (N_13240,N_10696,N_10441);
or U13241 (N_13241,N_11481,N_10222);
and U13242 (N_13242,N_10034,N_11818);
nand U13243 (N_13243,N_10771,N_10679);
nor U13244 (N_13244,N_10024,N_10632);
nor U13245 (N_13245,N_10348,N_11694);
and U13246 (N_13246,N_11371,N_10441);
or U13247 (N_13247,N_11639,N_11731);
nor U13248 (N_13248,N_10864,N_10917);
nand U13249 (N_13249,N_10304,N_10690);
nor U13250 (N_13250,N_10864,N_10837);
nand U13251 (N_13251,N_10514,N_11448);
nor U13252 (N_13252,N_10230,N_11699);
and U13253 (N_13253,N_10005,N_11171);
nor U13254 (N_13254,N_10262,N_10207);
or U13255 (N_13255,N_10713,N_10779);
nand U13256 (N_13256,N_11107,N_10321);
xor U13257 (N_13257,N_10495,N_11111);
or U13258 (N_13258,N_10147,N_11336);
nor U13259 (N_13259,N_11375,N_11556);
nor U13260 (N_13260,N_11003,N_11406);
nor U13261 (N_13261,N_11266,N_11987);
nand U13262 (N_13262,N_11242,N_11685);
or U13263 (N_13263,N_11383,N_11627);
nand U13264 (N_13264,N_11930,N_10321);
xor U13265 (N_13265,N_11664,N_10032);
xnor U13266 (N_13266,N_10701,N_11152);
and U13267 (N_13267,N_11933,N_11523);
nand U13268 (N_13268,N_10124,N_10901);
nor U13269 (N_13269,N_11478,N_10275);
and U13270 (N_13270,N_10755,N_11189);
and U13271 (N_13271,N_10015,N_11529);
nor U13272 (N_13272,N_10024,N_11892);
xor U13273 (N_13273,N_11934,N_10698);
or U13274 (N_13274,N_11223,N_10631);
nand U13275 (N_13275,N_10729,N_11513);
or U13276 (N_13276,N_10649,N_10666);
or U13277 (N_13277,N_10441,N_10122);
or U13278 (N_13278,N_11065,N_11259);
or U13279 (N_13279,N_11613,N_10325);
and U13280 (N_13280,N_10593,N_11576);
nand U13281 (N_13281,N_11929,N_11623);
xor U13282 (N_13282,N_10817,N_11068);
or U13283 (N_13283,N_11734,N_11495);
nand U13284 (N_13284,N_10291,N_11017);
nand U13285 (N_13285,N_10543,N_10629);
or U13286 (N_13286,N_10152,N_11165);
or U13287 (N_13287,N_10245,N_11826);
nor U13288 (N_13288,N_10719,N_10481);
nand U13289 (N_13289,N_10296,N_11849);
or U13290 (N_13290,N_10308,N_11186);
or U13291 (N_13291,N_11217,N_11912);
xor U13292 (N_13292,N_11719,N_10902);
nand U13293 (N_13293,N_10175,N_11822);
nor U13294 (N_13294,N_11233,N_10584);
xor U13295 (N_13295,N_10615,N_10542);
xor U13296 (N_13296,N_11090,N_10889);
and U13297 (N_13297,N_11426,N_10429);
and U13298 (N_13298,N_11180,N_10191);
or U13299 (N_13299,N_11084,N_10195);
or U13300 (N_13300,N_10740,N_11164);
nand U13301 (N_13301,N_11242,N_10871);
or U13302 (N_13302,N_10380,N_10429);
or U13303 (N_13303,N_10586,N_10523);
and U13304 (N_13304,N_10567,N_11912);
nand U13305 (N_13305,N_10704,N_10871);
nand U13306 (N_13306,N_11375,N_10323);
or U13307 (N_13307,N_10651,N_10561);
and U13308 (N_13308,N_11731,N_11075);
nor U13309 (N_13309,N_10749,N_10132);
xor U13310 (N_13310,N_11096,N_10087);
xnor U13311 (N_13311,N_10393,N_11966);
or U13312 (N_13312,N_11882,N_11145);
nor U13313 (N_13313,N_11937,N_11105);
nor U13314 (N_13314,N_10508,N_11990);
and U13315 (N_13315,N_10460,N_11447);
and U13316 (N_13316,N_10212,N_11415);
xor U13317 (N_13317,N_10640,N_10805);
and U13318 (N_13318,N_10163,N_11626);
xor U13319 (N_13319,N_10773,N_11139);
nand U13320 (N_13320,N_10311,N_10556);
nand U13321 (N_13321,N_10142,N_11068);
nand U13322 (N_13322,N_11815,N_10370);
xnor U13323 (N_13323,N_10321,N_10831);
nand U13324 (N_13324,N_10824,N_10661);
or U13325 (N_13325,N_11053,N_11807);
nor U13326 (N_13326,N_10956,N_10753);
nor U13327 (N_13327,N_10863,N_11645);
or U13328 (N_13328,N_11367,N_10847);
or U13329 (N_13329,N_10059,N_10766);
nand U13330 (N_13330,N_11706,N_11459);
nand U13331 (N_13331,N_10297,N_11957);
xnor U13332 (N_13332,N_11149,N_10776);
xnor U13333 (N_13333,N_10005,N_10982);
nor U13334 (N_13334,N_11063,N_11799);
and U13335 (N_13335,N_11172,N_10749);
xor U13336 (N_13336,N_10951,N_10645);
or U13337 (N_13337,N_10697,N_10579);
nand U13338 (N_13338,N_10411,N_10820);
and U13339 (N_13339,N_10542,N_10314);
and U13340 (N_13340,N_10909,N_10004);
xor U13341 (N_13341,N_11862,N_11310);
and U13342 (N_13342,N_11878,N_11983);
nor U13343 (N_13343,N_10807,N_11008);
or U13344 (N_13344,N_10449,N_11041);
nand U13345 (N_13345,N_11327,N_11469);
xor U13346 (N_13346,N_10042,N_10837);
nand U13347 (N_13347,N_11723,N_10204);
and U13348 (N_13348,N_11814,N_10513);
xnor U13349 (N_13349,N_11890,N_10829);
nor U13350 (N_13350,N_11458,N_10357);
and U13351 (N_13351,N_10160,N_10089);
nand U13352 (N_13352,N_10285,N_11980);
nand U13353 (N_13353,N_10749,N_11073);
nor U13354 (N_13354,N_11569,N_11884);
or U13355 (N_13355,N_10680,N_10977);
xor U13356 (N_13356,N_10237,N_10771);
nand U13357 (N_13357,N_10524,N_10029);
or U13358 (N_13358,N_10976,N_11816);
nor U13359 (N_13359,N_11787,N_10853);
xnor U13360 (N_13360,N_11014,N_10677);
or U13361 (N_13361,N_11472,N_11861);
and U13362 (N_13362,N_11253,N_10929);
or U13363 (N_13363,N_10717,N_10708);
nor U13364 (N_13364,N_10784,N_11697);
xor U13365 (N_13365,N_10734,N_11326);
nor U13366 (N_13366,N_10703,N_11348);
nand U13367 (N_13367,N_10473,N_11883);
nand U13368 (N_13368,N_10209,N_11633);
nand U13369 (N_13369,N_11961,N_10848);
nor U13370 (N_13370,N_11537,N_11414);
nand U13371 (N_13371,N_11033,N_10155);
nor U13372 (N_13372,N_11997,N_11899);
xnor U13373 (N_13373,N_10431,N_10756);
and U13374 (N_13374,N_11920,N_10452);
nor U13375 (N_13375,N_11075,N_10539);
or U13376 (N_13376,N_10638,N_11316);
nor U13377 (N_13377,N_10735,N_11635);
xnor U13378 (N_13378,N_11629,N_10590);
and U13379 (N_13379,N_11517,N_10660);
nand U13380 (N_13380,N_11249,N_10972);
nor U13381 (N_13381,N_11094,N_11751);
nand U13382 (N_13382,N_10627,N_11406);
nand U13383 (N_13383,N_10290,N_11154);
xnor U13384 (N_13384,N_11046,N_10357);
nor U13385 (N_13385,N_10683,N_10645);
and U13386 (N_13386,N_11763,N_11350);
or U13387 (N_13387,N_10241,N_11966);
and U13388 (N_13388,N_11055,N_10582);
or U13389 (N_13389,N_11144,N_11667);
nor U13390 (N_13390,N_11795,N_10806);
nand U13391 (N_13391,N_10550,N_10010);
nor U13392 (N_13392,N_11094,N_11812);
xnor U13393 (N_13393,N_10233,N_10523);
nand U13394 (N_13394,N_10430,N_10463);
or U13395 (N_13395,N_11542,N_11059);
nand U13396 (N_13396,N_11579,N_11997);
xnor U13397 (N_13397,N_10037,N_11024);
xor U13398 (N_13398,N_11666,N_10144);
nor U13399 (N_13399,N_11079,N_11970);
nand U13400 (N_13400,N_11096,N_10805);
and U13401 (N_13401,N_10458,N_10875);
nand U13402 (N_13402,N_11628,N_10936);
nor U13403 (N_13403,N_10086,N_11787);
or U13404 (N_13404,N_10441,N_10281);
or U13405 (N_13405,N_11818,N_11939);
or U13406 (N_13406,N_10842,N_10969);
and U13407 (N_13407,N_10982,N_11471);
or U13408 (N_13408,N_11838,N_11882);
and U13409 (N_13409,N_10759,N_10906);
and U13410 (N_13410,N_11233,N_11589);
xor U13411 (N_13411,N_10266,N_10732);
or U13412 (N_13412,N_11538,N_11598);
and U13413 (N_13413,N_10532,N_10075);
nor U13414 (N_13414,N_11263,N_10757);
xor U13415 (N_13415,N_11752,N_11606);
nor U13416 (N_13416,N_11427,N_11935);
nand U13417 (N_13417,N_10960,N_11767);
nand U13418 (N_13418,N_11156,N_10118);
and U13419 (N_13419,N_10643,N_10769);
or U13420 (N_13420,N_10664,N_10073);
or U13421 (N_13421,N_11358,N_10352);
nor U13422 (N_13422,N_10293,N_11998);
xnor U13423 (N_13423,N_11365,N_11669);
nand U13424 (N_13424,N_11227,N_10975);
xor U13425 (N_13425,N_10809,N_10399);
and U13426 (N_13426,N_10203,N_11445);
xor U13427 (N_13427,N_11096,N_10926);
nor U13428 (N_13428,N_11905,N_10164);
xor U13429 (N_13429,N_11649,N_11476);
xnor U13430 (N_13430,N_11082,N_10351);
or U13431 (N_13431,N_10626,N_11076);
xnor U13432 (N_13432,N_11020,N_11145);
and U13433 (N_13433,N_11459,N_10425);
and U13434 (N_13434,N_10105,N_10877);
nor U13435 (N_13435,N_10849,N_10608);
and U13436 (N_13436,N_10029,N_11268);
and U13437 (N_13437,N_10386,N_11880);
nor U13438 (N_13438,N_11007,N_10969);
nand U13439 (N_13439,N_10930,N_10329);
nor U13440 (N_13440,N_11575,N_10258);
xor U13441 (N_13441,N_11069,N_11988);
nand U13442 (N_13442,N_10896,N_11969);
nand U13443 (N_13443,N_10450,N_11220);
xnor U13444 (N_13444,N_10605,N_10868);
or U13445 (N_13445,N_11843,N_10981);
or U13446 (N_13446,N_10591,N_11604);
xnor U13447 (N_13447,N_10134,N_10823);
xor U13448 (N_13448,N_10321,N_11618);
xor U13449 (N_13449,N_11139,N_10368);
nor U13450 (N_13450,N_11667,N_11964);
nand U13451 (N_13451,N_11957,N_10063);
or U13452 (N_13452,N_10684,N_11332);
nand U13453 (N_13453,N_10299,N_11822);
and U13454 (N_13454,N_11497,N_10158);
nor U13455 (N_13455,N_11731,N_10411);
and U13456 (N_13456,N_11924,N_11010);
and U13457 (N_13457,N_10808,N_11810);
xor U13458 (N_13458,N_10727,N_10676);
nor U13459 (N_13459,N_11536,N_11915);
and U13460 (N_13460,N_11161,N_10743);
nand U13461 (N_13461,N_10617,N_11302);
xor U13462 (N_13462,N_10372,N_11448);
or U13463 (N_13463,N_11479,N_10138);
xnor U13464 (N_13464,N_10709,N_11059);
or U13465 (N_13465,N_10993,N_10873);
or U13466 (N_13466,N_10387,N_11570);
nor U13467 (N_13467,N_10610,N_10852);
nand U13468 (N_13468,N_10407,N_10604);
nand U13469 (N_13469,N_10450,N_11789);
nor U13470 (N_13470,N_10551,N_11032);
xnor U13471 (N_13471,N_11573,N_11899);
and U13472 (N_13472,N_11527,N_10998);
nand U13473 (N_13473,N_11843,N_11769);
nor U13474 (N_13474,N_10307,N_11975);
xnor U13475 (N_13475,N_11144,N_11615);
nor U13476 (N_13476,N_10406,N_11728);
nand U13477 (N_13477,N_10170,N_10553);
nand U13478 (N_13478,N_10824,N_11304);
or U13479 (N_13479,N_11620,N_11318);
nor U13480 (N_13480,N_10309,N_10134);
xnor U13481 (N_13481,N_10216,N_10341);
nand U13482 (N_13482,N_10064,N_11342);
nor U13483 (N_13483,N_10030,N_11444);
nor U13484 (N_13484,N_10084,N_11407);
xnor U13485 (N_13485,N_10222,N_11616);
or U13486 (N_13486,N_10575,N_11062);
or U13487 (N_13487,N_10326,N_10055);
nor U13488 (N_13488,N_11671,N_10513);
nand U13489 (N_13489,N_11126,N_10721);
nand U13490 (N_13490,N_10389,N_10863);
or U13491 (N_13491,N_11664,N_11794);
nand U13492 (N_13492,N_10558,N_10959);
nand U13493 (N_13493,N_11054,N_10199);
and U13494 (N_13494,N_10810,N_10011);
and U13495 (N_13495,N_10938,N_11344);
nand U13496 (N_13496,N_10424,N_11103);
nor U13497 (N_13497,N_11284,N_10920);
nor U13498 (N_13498,N_11972,N_11686);
xor U13499 (N_13499,N_10215,N_11766);
and U13500 (N_13500,N_10421,N_11288);
nand U13501 (N_13501,N_10324,N_11583);
xor U13502 (N_13502,N_10592,N_10315);
or U13503 (N_13503,N_11157,N_10780);
nor U13504 (N_13504,N_10322,N_11597);
and U13505 (N_13505,N_11090,N_11391);
nor U13506 (N_13506,N_11766,N_11093);
nor U13507 (N_13507,N_11410,N_11466);
or U13508 (N_13508,N_10348,N_11798);
or U13509 (N_13509,N_11900,N_10862);
xor U13510 (N_13510,N_10595,N_11064);
nand U13511 (N_13511,N_10183,N_10220);
and U13512 (N_13512,N_11018,N_11161);
and U13513 (N_13513,N_10374,N_10793);
nor U13514 (N_13514,N_10530,N_11115);
nand U13515 (N_13515,N_11377,N_10241);
and U13516 (N_13516,N_11813,N_10402);
xor U13517 (N_13517,N_10617,N_10689);
nor U13518 (N_13518,N_10784,N_11949);
and U13519 (N_13519,N_10048,N_11830);
xnor U13520 (N_13520,N_11949,N_10755);
nor U13521 (N_13521,N_10990,N_10200);
xor U13522 (N_13522,N_10223,N_10290);
nand U13523 (N_13523,N_11695,N_10934);
or U13524 (N_13524,N_11344,N_11040);
xor U13525 (N_13525,N_11341,N_11520);
or U13526 (N_13526,N_11344,N_10775);
or U13527 (N_13527,N_11133,N_10511);
xnor U13528 (N_13528,N_11429,N_10438);
or U13529 (N_13529,N_11903,N_11080);
or U13530 (N_13530,N_11829,N_10399);
nand U13531 (N_13531,N_10310,N_10201);
or U13532 (N_13532,N_11883,N_11114);
xor U13533 (N_13533,N_11277,N_11687);
nand U13534 (N_13534,N_11725,N_11274);
nor U13535 (N_13535,N_11655,N_10347);
xnor U13536 (N_13536,N_11719,N_11414);
xor U13537 (N_13537,N_10621,N_11843);
xor U13538 (N_13538,N_10918,N_11724);
and U13539 (N_13539,N_11676,N_11630);
and U13540 (N_13540,N_10604,N_10630);
and U13541 (N_13541,N_11453,N_10357);
xnor U13542 (N_13542,N_11544,N_11385);
or U13543 (N_13543,N_11222,N_10377);
nand U13544 (N_13544,N_11128,N_10744);
nand U13545 (N_13545,N_11572,N_11836);
xor U13546 (N_13546,N_11335,N_10007);
nor U13547 (N_13547,N_11255,N_11406);
and U13548 (N_13548,N_10021,N_11567);
nor U13549 (N_13549,N_11917,N_11486);
nand U13550 (N_13550,N_10065,N_10843);
or U13551 (N_13551,N_10489,N_10814);
nor U13552 (N_13552,N_10225,N_10374);
nand U13553 (N_13553,N_11507,N_11420);
xnor U13554 (N_13554,N_10796,N_11958);
or U13555 (N_13555,N_11603,N_11842);
xor U13556 (N_13556,N_10281,N_11077);
nand U13557 (N_13557,N_10655,N_10709);
nand U13558 (N_13558,N_11905,N_11834);
nor U13559 (N_13559,N_10446,N_10914);
nand U13560 (N_13560,N_11274,N_10210);
or U13561 (N_13561,N_11277,N_11105);
nand U13562 (N_13562,N_10387,N_10557);
xor U13563 (N_13563,N_10501,N_10406);
or U13564 (N_13564,N_10658,N_10609);
nor U13565 (N_13565,N_10733,N_11978);
nor U13566 (N_13566,N_11062,N_11033);
nand U13567 (N_13567,N_11630,N_10779);
nand U13568 (N_13568,N_11281,N_10651);
xor U13569 (N_13569,N_10679,N_11666);
nor U13570 (N_13570,N_10529,N_10241);
nand U13571 (N_13571,N_10753,N_10708);
or U13572 (N_13572,N_11767,N_11472);
and U13573 (N_13573,N_11053,N_11770);
xor U13574 (N_13574,N_10581,N_10878);
xor U13575 (N_13575,N_11807,N_10417);
nand U13576 (N_13576,N_11456,N_10149);
xnor U13577 (N_13577,N_11778,N_11273);
nand U13578 (N_13578,N_11506,N_11538);
and U13579 (N_13579,N_11492,N_10779);
and U13580 (N_13580,N_11952,N_11073);
xor U13581 (N_13581,N_10908,N_11698);
and U13582 (N_13582,N_11109,N_11307);
xor U13583 (N_13583,N_10087,N_10171);
and U13584 (N_13584,N_11286,N_10302);
nor U13585 (N_13585,N_11409,N_10926);
or U13586 (N_13586,N_10345,N_11446);
or U13587 (N_13587,N_10954,N_11083);
or U13588 (N_13588,N_11001,N_11115);
xor U13589 (N_13589,N_11775,N_10976);
xor U13590 (N_13590,N_10243,N_10801);
nand U13591 (N_13591,N_10588,N_10420);
xnor U13592 (N_13592,N_10167,N_11670);
xnor U13593 (N_13593,N_11801,N_10243);
or U13594 (N_13594,N_10658,N_10186);
and U13595 (N_13595,N_11159,N_11093);
xor U13596 (N_13596,N_10504,N_11469);
and U13597 (N_13597,N_10372,N_10416);
nor U13598 (N_13598,N_11847,N_10731);
xnor U13599 (N_13599,N_11129,N_10813);
nor U13600 (N_13600,N_10886,N_11526);
xnor U13601 (N_13601,N_10972,N_11684);
xor U13602 (N_13602,N_10581,N_10297);
nor U13603 (N_13603,N_10661,N_11828);
xnor U13604 (N_13604,N_11047,N_11383);
nand U13605 (N_13605,N_10881,N_10771);
and U13606 (N_13606,N_11657,N_11803);
xnor U13607 (N_13607,N_10450,N_11792);
nand U13608 (N_13608,N_10053,N_10346);
nand U13609 (N_13609,N_11049,N_11930);
xor U13610 (N_13610,N_11322,N_11062);
and U13611 (N_13611,N_11166,N_11435);
and U13612 (N_13612,N_11167,N_11789);
nor U13613 (N_13613,N_11606,N_10587);
nand U13614 (N_13614,N_11265,N_11315);
xnor U13615 (N_13615,N_11727,N_11527);
or U13616 (N_13616,N_10437,N_10124);
nand U13617 (N_13617,N_10541,N_10640);
nand U13618 (N_13618,N_10102,N_10636);
nor U13619 (N_13619,N_11332,N_10769);
nor U13620 (N_13620,N_11506,N_10443);
xnor U13621 (N_13621,N_11581,N_11320);
and U13622 (N_13622,N_10382,N_11244);
nor U13623 (N_13623,N_10589,N_10936);
or U13624 (N_13624,N_10494,N_10182);
or U13625 (N_13625,N_11480,N_10666);
nand U13626 (N_13626,N_10481,N_11560);
nor U13627 (N_13627,N_10199,N_10163);
nor U13628 (N_13628,N_10771,N_10555);
and U13629 (N_13629,N_10964,N_11853);
and U13630 (N_13630,N_10588,N_10776);
and U13631 (N_13631,N_11942,N_11976);
nand U13632 (N_13632,N_11517,N_11177);
xnor U13633 (N_13633,N_10342,N_10883);
xor U13634 (N_13634,N_11534,N_11846);
or U13635 (N_13635,N_10477,N_11340);
or U13636 (N_13636,N_11263,N_11866);
nand U13637 (N_13637,N_11616,N_11592);
and U13638 (N_13638,N_11826,N_10053);
xor U13639 (N_13639,N_10508,N_10757);
xnor U13640 (N_13640,N_11008,N_10713);
or U13641 (N_13641,N_11800,N_10166);
xnor U13642 (N_13642,N_10906,N_11972);
xor U13643 (N_13643,N_10620,N_10996);
nor U13644 (N_13644,N_11690,N_11314);
or U13645 (N_13645,N_11161,N_11865);
nand U13646 (N_13646,N_11747,N_10745);
nor U13647 (N_13647,N_10441,N_10389);
and U13648 (N_13648,N_10048,N_10424);
or U13649 (N_13649,N_11243,N_10212);
xnor U13650 (N_13650,N_10559,N_11307);
nand U13651 (N_13651,N_10799,N_11478);
or U13652 (N_13652,N_10158,N_10073);
nor U13653 (N_13653,N_10938,N_10099);
xor U13654 (N_13654,N_10517,N_11087);
and U13655 (N_13655,N_10458,N_11443);
or U13656 (N_13656,N_11396,N_10408);
xor U13657 (N_13657,N_10064,N_11155);
and U13658 (N_13658,N_11941,N_11045);
nor U13659 (N_13659,N_11043,N_11721);
or U13660 (N_13660,N_10358,N_11062);
xnor U13661 (N_13661,N_10715,N_10511);
or U13662 (N_13662,N_10589,N_10509);
nand U13663 (N_13663,N_10469,N_10557);
xor U13664 (N_13664,N_11368,N_11042);
and U13665 (N_13665,N_10246,N_11306);
nor U13666 (N_13666,N_11455,N_10367);
nor U13667 (N_13667,N_10049,N_10819);
nor U13668 (N_13668,N_10235,N_10840);
or U13669 (N_13669,N_11817,N_11503);
xnor U13670 (N_13670,N_11738,N_11963);
nor U13671 (N_13671,N_10460,N_10364);
nor U13672 (N_13672,N_11764,N_10274);
xnor U13673 (N_13673,N_10594,N_10700);
or U13674 (N_13674,N_11166,N_10101);
nand U13675 (N_13675,N_10810,N_10885);
or U13676 (N_13676,N_11802,N_11134);
nor U13677 (N_13677,N_11507,N_11486);
xnor U13678 (N_13678,N_11728,N_10537);
nor U13679 (N_13679,N_10615,N_11549);
xnor U13680 (N_13680,N_10331,N_11139);
xor U13681 (N_13681,N_11096,N_10577);
xnor U13682 (N_13682,N_10210,N_10850);
nor U13683 (N_13683,N_10481,N_10478);
nor U13684 (N_13684,N_11443,N_11076);
or U13685 (N_13685,N_10506,N_10061);
xnor U13686 (N_13686,N_11685,N_10459);
and U13687 (N_13687,N_10506,N_11878);
xor U13688 (N_13688,N_11384,N_10618);
or U13689 (N_13689,N_11559,N_10104);
nand U13690 (N_13690,N_10170,N_10672);
nand U13691 (N_13691,N_11974,N_11220);
or U13692 (N_13692,N_11183,N_10895);
or U13693 (N_13693,N_11033,N_11216);
or U13694 (N_13694,N_10990,N_10415);
nor U13695 (N_13695,N_10551,N_10614);
or U13696 (N_13696,N_10579,N_11459);
xor U13697 (N_13697,N_10640,N_10268);
nand U13698 (N_13698,N_10373,N_11003);
xnor U13699 (N_13699,N_10927,N_11444);
xnor U13700 (N_13700,N_11117,N_11332);
nor U13701 (N_13701,N_11704,N_11505);
or U13702 (N_13702,N_10139,N_10741);
nor U13703 (N_13703,N_11784,N_11692);
nor U13704 (N_13704,N_11139,N_10736);
or U13705 (N_13705,N_11113,N_10253);
and U13706 (N_13706,N_10326,N_10247);
and U13707 (N_13707,N_11909,N_11282);
nor U13708 (N_13708,N_11685,N_11915);
or U13709 (N_13709,N_10877,N_10355);
and U13710 (N_13710,N_10539,N_11948);
nand U13711 (N_13711,N_11562,N_11462);
xor U13712 (N_13712,N_10327,N_10497);
or U13713 (N_13713,N_10306,N_11778);
nand U13714 (N_13714,N_11492,N_11398);
xor U13715 (N_13715,N_11915,N_10386);
xor U13716 (N_13716,N_11292,N_11497);
and U13717 (N_13717,N_10091,N_11252);
and U13718 (N_13718,N_10339,N_10902);
or U13719 (N_13719,N_10432,N_10697);
nor U13720 (N_13720,N_11941,N_11086);
and U13721 (N_13721,N_10840,N_11139);
and U13722 (N_13722,N_10494,N_10395);
and U13723 (N_13723,N_10746,N_11904);
nand U13724 (N_13724,N_11153,N_10234);
nand U13725 (N_13725,N_11317,N_11623);
and U13726 (N_13726,N_11318,N_11996);
or U13727 (N_13727,N_11101,N_11760);
nor U13728 (N_13728,N_10712,N_10467);
or U13729 (N_13729,N_10336,N_10653);
and U13730 (N_13730,N_11240,N_11458);
xor U13731 (N_13731,N_11804,N_11829);
and U13732 (N_13732,N_11202,N_11718);
xor U13733 (N_13733,N_11265,N_10981);
nand U13734 (N_13734,N_10248,N_10268);
and U13735 (N_13735,N_11185,N_11286);
nand U13736 (N_13736,N_11018,N_10387);
xnor U13737 (N_13737,N_10924,N_10425);
nand U13738 (N_13738,N_10957,N_11535);
nor U13739 (N_13739,N_11825,N_11945);
and U13740 (N_13740,N_10175,N_11009);
and U13741 (N_13741,N_10714,N_11190);
nor U13742 (N_13742,N_11964,N_10268);
and U13743 (N_13743,N_11310,N_11920);
and U13744 (N_13744,N_11706,N_11965);
or U13745 (N_13745,N_11812,N_11521);
and U13746 (N_13746,N_11079,N_11502);
or U13747 (N_13747,N_10379,N_11040);
nand U13748 (N_13748,N_10632,N_10215);
nand U13749 (N_13749,N_10079,N_11356);
nand U13750 (N_13750,N_10505,N_11457);
nor U13751 (N_13751,N_11741,N_10994);
nor U13752 (N_13752,N_11513,N_11437);
xor U13753 (N_13753,N_11665,N_10686);
xor U13754 (N_13754,N_11640,N_11688);
xor U13755 (N_13755,N_10320,N_11210);
nor U13756 (N_13756,N_10390,N_11687);
and U13757 (N_13757,N_10613,N_10710);
nand U13758 (N_13758,N_11084,N_10019);
nor U13759 (N_13759,N_10756,N_10367);
nand U13760 (N_13760,N_11785,N_10094);
or U13761 (N_13761,N_10912,N_11954);
xor U13762 (N_13762,N_11714,N_11448);
and U13763 (N_13763,N_10005,N_11726);
or U13764 (N_13764,N_11507,N_10673);
nor U13765 (N_13765,N_11627,N_11112);
nor U13766 (N_13766,N_11136,N_10646);
xnor U13767 (N_13767,N_11937,N_10004);
or U13768 (N_13768,N_11318,N_11108);
and U13769 (N_13769,N_11890,N_10178);
nand U13770 (N_13770,N_10344,N_11637);
or U13771 (N_13771,N_11318,N_10083);
or U13772 (N_13772,N_11439,N_11662);
and U13773 (N_13773,N_10598,N_10994);
nor U13774 (N_13774,N_10011,N_11864);
or U13775 (N_13775,N_10216,N_11060);
or U13776 (N_13776,N_10152,N_11593);
nor U13777 (N_13777,N_11598,N_10473);
xnor U13778 (N_13778,N_10702,N_10796);
xor U13779 (N_13779,N_11527,N_10589);
and U13780 (N_13780,N_11258,N_11478);
and U13781 (N_13781,N_11435,N_10789);
nor U13782 (N_13782,N_10713,N_10656);
nand U13783 (N_13783,N_10938,N_10243);
or U13784 (N_13784,N_10910,N_11926);
nor U13785 (N_13785,N_11423,N_10076);
xor U13786 (N_13786,N_11285,N_11007);
or U13787 (N_13787,N_10583,N_11027);
or U13788 (N_13788,N_10989,N_10928);
xor U13789 (N_13789,N_10559,N_10756);
or U13790 (N_13790,N_11131,N_10138);
nor U13791 (N_13791,N_11261,N_11720);
xor U13792 (N_13792,N_10553,N_10960);
nand U13793 (N_13793,N_11682,N_10915);
xnor U13794 (N_13794,N_11627,N_10859);
or U13795 (N_13795,N_11587,N_11370);
nor U13796 (N_13796,N_11272,N_10663);
xnor U13797 (N_13797,N_10895,N_10064);
nor U13798 (N_13798,N_11245,N_11530);
or U13799 (N_13799,N_11886,N_10888);
xor U13800 (N_13800,N_10469,N_10515);
or U13801 (N_13801,N_10847,N_11618);
nor U13802 (N_13802,N_10837,N_11750);
or U13803 (N_13803,N_11522,N_11893);
nor U13804 (N_13804,N_10715,N_11466);
nand U13805 (N_13805,N_11869,N_11558);
nor U13806 (N_13806,N_10543,N_10225);
nor U13807 (N_13807,N_11414,N_11650);
nand U13808 (N_13808,N_11423,N_10706);
or U13809 (N_13809,N_10087,N_10663);
and U13810 (N_13810,N_11356,N_11620);
nor U13811 (N_13811,N_10873,N_11954);
or U13812 (N_13812,N_11617,N_11062);
or U13813 (N_13813,N_11732,N_11461);
nand U13814 (N_13814,N_11107,N_10980);
xnor U13815 (N_13815,N_10848,N_10219);
or U13816 (N_13816,N_11168,N_11309);
nand U13817 (N_13817,N_10936,N_10404);
nand U13818 (N_13818,N_10715,N_11112);
nor U13819 (N_13819,N_11050,N_10733);
nand U13820 (N_13820,N_11629,N_10939);
xor U13821 (N_13821,N_11309,N_11891);
xor U13822 (N_13822,N_10438,N_11483);
and U13823 (N_13823,N_10188,N_10904);
nand U13824 (N_13824,N_11125,N_10072);
and U13825 (N_13825,N_11071,N_10362);
xor U13826 (N_13826,N_11278,N_10866);
or U13827 (N_13827,N_10415,N_10023);
and U13828 (N_13828,N_10474,N_10347);
xor U13829 (N_13829,N_10015,N_11723);
and U13830 (N_13830,N_11301,N_10528);
nand U13831 (N_13831,N_11980,N_10536);
xnor U13832 (N_13832,N_10103,N_10638);
nor U13833 (N_13833,N_11199,N_10157);
or U13834 (N_13834,N_11256,N_10550);
and U13835 (N_13835,N_11064,N_11745);
and U13836 (N_13836,N_10107,N_10821);
xnor U13837 (N_13837,N_11099,N_11009);
nor U13838 (N_13838,N_10217,N_11053);
or U13839 (N_13839,N_11208,N_10144);
or U13840 (N_13840,N_11101,N_11242);
or U13841 (N_13841,N_11024,N_11603);
and U13842 (N_13842,N_11562,N_10296);
nand U13843 (N_13843,N_11489,N_11510);
nor U13844 (N_13844,N_11409,N_11181);
or U13845 (N_13845,N_10783,N_11742);
or U13846 (N_13846,N_10802,N_11826);
and U13847 (N_13847,N_10665,N_11961);
or U13848 (N_13848,N_10173,N_10592);
nand U13849 (N_13849,N_11087,N_11523);
nand U13850 (N_13850,N_11689,N_10685);
xor U13851 (N_13851,N_10557,N_10981);
nor U13852 (N_13852,N_10379,N_10640);
nand U13853 (N_13853,N_11495,N_11252);
nand U13854 (N_13854,N_11765,N_11285);
xnor U13855 (N_13855,N_10011,N_11673);
or U13856 (N_13856,N_10951,N_11212);
xnor U13857 (N_13857,N_11066,N_10723);
nor U13858 (N_13858,N_11017,N_10049);
and U13859 (N_13859,N_11245,N_10169);
or U13860 (N_13860,N_10276,N_10487);
and U13861 (N_13861,N_11554,N_10640);
and U13862 (N_13862,N_10999,N_11070);
or U13863 (N_13863,N_10065,N_10214);
or U13864 (N_13864,N_10419,N_10136);
nor U13865 (N_13865,N_11324,N_10263);
nand U13866 (N_13866,N_10446,N_11364);
xnor U13867 (N_13867,N_10929,N_11014);
xor U13868 (N_13868,N_10514,N_10543);
and U13869 (N_13869,N_10733,N_11642);
xnor U13870 (N_13870,N_11601,N_11091);
nor U13871 (N_13871,N_11237,N_11700);
nand U13872 (N_13872,N_11722,N_10171);
nand U13873 (N_13873,N_10717,N_11364);
nor U13874 (N_13874,N_10669,N_11187);
nand U13875 (N_13875,N_11823,N_10663);
and U13876 (N_13876,N_10002,N_10174);
and U13877 (N_13877,N_10940,N_10858);
or U13878 (N_13878,N_10457,N_10143);
nand U13879 (N_13879,N_10248,N_11924);
nand U13880 (N_13880,N_10535,N_10744);
or U13881 (N_13881,N_11970,N_11634);
and U13882 (N_13882,N_11377,N_10221);
or U13883 (N_13883,N_11356,N_10446);
nor U13884 (N_13884,N_10644,N_10612);
nor U13885 (N_13885,N_10106,N_10185);
or U13886 (N_13886,N_11094,N_11818);
and U13887 (N_13887,N_11098,N_11367);
and U13888 (N_13888,N_10522,N_10173);
nor U13889 (N_13889,N_11290,N_10701);
nor U13890 (N_13890,N_10622,N_11621);
nor U13891 (N_13891,N_10164,N_11094);
xnor U13892 (N_13892,N_11722,N_11519);
and U13893 (N_13893,N_11667,N_11581);
or U13894 (N_13894,N_11418,N_10935);
xor U13895 (N_13895,N_10258,N_10468);
nand U13896 (N_13896,N_11235,N_10165);
xor U13897 (N_13897,N_11425,N_10310);
and U13898 (N_13898,N_11632,N_11113);
nand U13899 (N_13899,N_11870,N_10601);
and U13900 (N_13900,N_10957,N_11202);
nand U13901 (N_13901,N_11170,N_10375);
or U13902 (N_13902,N_11239,N_11920);
xnor U13903 (N_13903,N_10653,N_11219);
and U13904 (N_13904,N_11117,N_11445);
nor U13905 (N_13905,N_11796,N_11023);
and U13906 (N_13906,N_10859,N_10825);
and U13907 (N_13907,N_11685,N_10975);
nor U13908 (N_13908,N_11667,N_11600);
xor U13909 (N_13909,N_10518,N_11338);
nand U13910 (N_13910,N_11031,N_10764);
or U13911 (N_13911,N_10861,N_10279);
xor U13912 (N_13912,N_11752,N_11112);
or U13913 (N_13913,N_11218,N_11360);
nand U13914 (N_13914,N_10456,N_10757);
nor U13915 (N_13915,N_10003,N_11315);
and U13916 (N_13916,N_10067,N_10063);
or U13917 (N_13917,N_10121,N_10584);
nor U13918 (N_13918,N_10285,N_11649);
and U13919 (N_13919,N_11142,N_11217);
xor U13920 (N_13920,N_10731,N_11307);
or U13921 (N_13921,N_11797,N_11950);
xor U13922 (N_13922,N_11206,N_10307);
and U13923 (N_13923,N_10657,N_11758);
and U13924 (N_13924,N_11736,N_10093);
xor U13925 (N_13925,N_11535,N_10027);
xnor U13926 (N_13926,N_11834,N_10336);
or U13927 (N_13927,N_11188,N_11653);
or U13928 (N_13928,N_10773,N_10373);
and U13929 (N_13929,N_11311,N_11331);
nor U13930 (N_13930,N_10174,N_11550);
nand U13931 (N_13931,N_10374,N_11494);
xor U13932 (N_13932,N_10985,N_11490);
nand U13933 (N_13933,N_11399,N_10754);
nand U13934 (N_13934,N_10091,N_10840);
xor U13935 (N_13935,N_11007,N_10366);
or U13936 (N_13936,N_10094,N_10888);
and U13937 (N_13937,N_10105,N_10258);
nor U13938 (N_13938,N_10339,N_10766);
and U13939 (N_13939,N_11561,N_11600);
xor U13940 (N_13940,N_11359,N_11414);
and U13941 (N_13941,N_11618,N_11307);
and U13942 (N_13942,N_11164,N_10379);
and U13943 (N_13943,N_10553,N_10111);
and U13944 (N_13944,N_11984,N_10086);
nand U13945 (N_13945,N_11155,N_10727);
xnor U13946 (N_13946,N_11163,N_11430);
nand U13947 (N_13947,N_10704,N_10329);
nand U13948 (N_13948,N_10538,N_11373);
xnor U13949 (N_13949,N_11507,N_11126);
xor U13950 (N_13950,N_10161,N_10537);
and U13951 (N_13951,N_10668,N_10822);
nand U13952 (N_13952,N_10519,N_11754);
xor U13953 (N_13953,N_10552,N_10714);
or U13954 (N_13954,N_10172,N_10232);
nor U13955 (N_13955,N_10371,N_11422);
or U13956 (N_13956,N_10185,N_11997);
and U13957 (N_13957,N_11662,N_10844);
or U13958 (N_13958,N_11347,N_11579);
nand U13959 (N_13959,N_11683,N_11726);
or U13960 (N_13960,N_10343,N_11939);
nand U13961 (N_13961,N_11698,N_11303);
nor U13962 (N_13962,N_10057,N_11112);
nand U13963 (N_13963,N_11441,N_11640);
xnor U13964 (N_13964,N_11127,N_10346);
or U13965 (N_13965,N_10681,N_11260);
and U13966 (N_13966,N_10638,N_10002);
or U13967 (N_13967,N_10876,N_10632);
and U13968 (N_13968,N_11239,N_10665);
nand U13969 (N_13969,N_10626,N_11763);
or U13970 (N_13970,N_11170,N_10068);
xnor U13971 (N_13971,N_10716,N_11157);
or U13972 (N_13972,N_11996,N_11449);
nor U13973 (N_13973,N_10097,N_10317);
nor U13974 (N_13974,N_10123,N_11255);
nor U13975 (N_13975,N_10448,N_10208);
xor U13976 (N_13976,N_10425,N_11258);
or U13977 (N_13977,N_10919,N_11564);
and U13978 (N_13978,N_11799,N_11358);
or U13979 (N_13979,N_10979,N_10128);
and U13980 (N_13980,N_10680,N_10887);
xnor U13981 (N_13981,N_11938,N_10099);
xnor U13982 (N_13982,N_11516,N_10689);
xnor U13983 (N_13983,N_10384,N_11199);
xor U13984 (N_13984,N_11153,N_10739);
nor U13985 (N_13985,N_10068,N_10281);
or U13986 (N_13986,N_11588,N_10025);
nor U13987 (N_13987,N_10648,N_11881);
nor U13988 (N_13988,N_11230,N_10886);
and U13989 (N_13989,N_11644,N_11346);
and U13990 (N_13990,N_10310,N_10766);
nor U13991 (N_13991,N_11007,N_11766);
and U13992 (N_13992,N_11768,N_10017);
and U13993 (N_13993,N_11875,N_11054);
and U13994 (N_13994,N_10458,N_11315);
and U13995 (N_13995,N_10251,N_10781);
or U13996 (N_13996,N_10731,N_10179);
nand U13997 (N_13997,N_10180,N_10514);
xnor U13998 (N_13998,N_11045,N_10875);
and U13999 (N_13999,N_10536,N_11892);
and U14000 (N_14000,N_13605,N_12604);
and U14001 (N_14001,N_13785,N_13089);
or U14002 (N_14002,N_13245,N_13853);
xnor U14003 (N_14003,N_13370,N_13517);
and U14004 (N_14004,N_13112,N_12670);
and U14005 (N_14005,N_12873,N_13889);
or U14006 (N_14006,N_13279,N_13304);
and U14007 (N_14007,N_13477,N_12933);
and U14008 (N_14008,N_12851,N_13412);
nor U14009 (N_14009,N_13638,N_12720);
nor U14010 (N_14010,N_13585,N_13914);
and U14011 (N_14011,N_12066,N_12689);
nor U14012 (N_14012,N_12448,N_12141);
and U14013 (N_14013,N_12554,N_13482);
or U14014 (N_14014,N_13437,N_13678);
nor U14015 (N_14015,N_12455,N_13149);
and U14016 (N_14016,N_13064,N_12775);
xnor U14017 (N_14017,N_13184,N_13784);
xor U14018 (N_14018,N_12312,N_13818);
or U14019 (N_14019,N_12633,N_12621);
nor U14020 (N_14020,N_13132,N_13713);
or U14021 (N_14021,N_12167,N_12279);
or U14022 (N_14022,N_12155,N_13364);
or U14023 (N_14023,N_12702,N_12516);
nand U14024 (N_14024,N_13580,N_12493);
nand U14025 (N_14025,N_13087,N_12449);
and U14026 (N_14026,N_13121,N_12630);
and U14027 (N_14027,N_13221,N_12246);
nor U14028 (N_14028,N_12238,N_12972);
and U14029 (N_14029,N_12602,N_12081);
nand U14030 (N_14030,N_13310,N_12294);
xnor U14031 (N_14031,N_13211,N_12926);
or U14032 (N_14032,N_13986,N_12645);
nor U14033 (N_14033,N_12548,N_13977);
nand U14034 (N_14034,N_13410,N_12491);
or U14035 (N_14035,N_12817,N_12408);
xnor U14036 (N_14036,N_12919,N_13990);
and U14037 (N_14037,N_12901,N_12747);
nor U14038 (N_14038,N_13242,N_12531);
or U14039 (N_14039,N_12121,N_12757);
or U14040 (N_14040,N_12570,N_12407);
nand U14041 (N_14041,N_12502,N_13062);
or U14042 (N_14042,N_13476,N_13207);
or U14043 (N_14043,N_13483,N_13396);
and U14044 (N_14044,N_12115,N_12084);
nand U14045 (N_14045,N_13057,N_13674);
and U14046 (N_14046,N_13694,N_13208);
xor U14047 (N_14047,N_12792,N_12158);
nor U14048 (N_14048,N_13265,N_13652);
nor U14049 (N_14049,N_13401,N_13009);
xor U14050 (N_14050,N_12831,N_13071);
nor U14051 (N_14051,N_12613,N_13416);
nor U14052 (N_14052,N_13948,N_13447);
and U14053 (N_14053,N_12587,N_12423);
and U14054 (N_14054,N_13692,N_13204);
nor U14055 (N_14055,N_13332,N_12827);
nand U14056 (N_14056,N_13540,N_12459);
nor U14057 (N_14057,N_12654,N_12674);
nor U14058 (N_14058,N_12788,N_12023);
or U14059 (N_14059,N_12850,N_12481);
nor U14060 (N_14060,N_13884,N_13442);
nand U14061 (N_14061,N_12242,N_13543);
xor U14062 (N_14062,N_13193,N_13180);
nand U14063 (N_14063,N_13969,N_13160);
or U14064 (N_14064,N_12403,N_13849);
nor U14065 (N_14065,N_13759,N_13533);
xor U14066 (N_14066,N_13766,N_13863);
xnor U14067 (N_14067,N_13272,N_12910);
nand U14068 (N_14068,N_12145,N_13937);
nor U14069 (N_14069,N_12194,N_12805);
and U14070 (N_14070,N_13925,N_12691);
xnor U14071 (N_14071,N_12639,N_13491);
xor U14072 (N_14072,N_12371,N_13308);
xor U14073 (N_14073,N_13197,N_13851);
nor U14074 (N_14074,N_13756,N_13343);
nand U14075 (N_14075,N_13455,N_12983);
nand U14076 (N_14076,N_12405,N_12632);
xor U14077 (N_14077,N_12551,N_13811);
or U14078 (N_14078,N_13649,N_13562);
nand U14079 (N_14079,N_13943,N_13873);
or U14080 (N_14080,N_12657,N_12483);
nor U14081 (N_14081,N_12681,N_13203);
xor U14082 (N_14082,N_12909,N_12787);
nor U14083 (N_14083,N_12785,N_12385);
nor U14084 (N_14084,N_13407,N_12024);
nor U14085 (N_14085,N_12903,N_12881);
or U14086 (N_14086,N_13994,N_12686);
xnor U14087 (N_14087,N_13190,N_13901);
and U14088 (N_14088,N_13838,N_13904);
nor U14089 (N_14089,N_13687,N_12037);
nor U14090 (N_14090,N_13258,N_13590);
xnor U14091 (N_14091,N_13913,N_12259);
and U14092 (N_14092,N_12107,N_13307);
nand U14093 (N_14093,N_12998,N_12964);
and U14094 (N_14094,N_12510,N_13708);
xor U14095 (N_14095,N_13338,N_12065);
nor U14096 (N_14096,N_12004,N_13353);
nand U14097 (N_14097,N_12537,N_13518);
xor U14098 (N_14098,N_13110,N_12966);
xnor U14099 (N_14099,N_12628,N_12303);
nor U14100 (N_14100,N_13519,N_12178);
or U14101 (N_14101,N_13438,N_12469);
or U14102 (N_14102,N_13892,N_12197);
nand U14103 (N_14103,N_12376,N_12116);
or U14104 (N_14104,N_12914,N_12588);
nand U14105 (N_14105,N_13806,N_13752);
xor U14106 (N_14106,N_13052,N_13557);
nand U14107 (N_14107,N_13825,N_12542);
xnor U14108 (N_14108,N_13701,N_13117);
nand U14109 (N_14109,N_12022,N_13252);
xnor U14110 (N_14110,N_12624,N_12383);
nand U14111 (N_14111,N_12798,N_12233);
and U14112 (N_14112,N_13929,N_13225);
xnor U14113 (N_14113,N_12927,N_12027);
nand U14114 (N_14114,N_12234,N_12090);
and U14115 (N_14115,N_12801,N_12348);
nand U14116 (N_14116,N_13340,N_13963);
or U14117 (N_14117,N_13363,N_13256);
and U14118 (N_14118,N_12756,N_13249);
nand U14119 (N_14119,N_12976,N_12036);
and U14120 (N_14120,N_12637,N_13191);
nand U14121 (N_14121,N_12853,N_13541);
nand U14122 (N_14122,N_12617,N_12653);
xnor U14123 (N_14123,N_13726,N_13226);
xnor U14124 (N_14124,N_12620,N_13885);
nor U14125 (N_14125,N_12350,N_12500);
nand U14126 (N_14126,N_12451,N_13781);
and U14127 (N_14127,N_12048,N_12422);
nand U14128 (N_14128,N_13022,N_13246);
nand U14129 (N_14129,N_13115,N_13228);
nand U14130 (N_14130,N_13457,N_12665);
nand U14131 (N_14131,N_13431,N_13951);
or U14132 (N_14132,N_13730,N_13615);
nand U14133 (N_14133,N_13799,N_12104);
or U14134 (N_14134,N_12466,N_12687);
nor U14135 (N_14135,N_12077,N_12339);
xor U14136 (N_14136,N_12997,N_12395);
or U14137 (N_14137,N_12390,N_12000);
nor U14138 (N_14138,N_12800,N_12487);
nand U14139 (N_14139,N_12213,N_13633);
or U14140 (N_14140,N_12230,N_12330);
nand U14141 (N_14141,N_12547,N_13871);
nand U14142 (N_14142,N_12867,N_13425);
nor U14143 (N_14143,N_13096,N_13324);
and U14144 (N_14144,N_12143,N_12492);
nand U14145 (N_14145,N_13496,N_12341);
nand U14146 (N_14146,N_13031,N_13976);
and U14147 (N_14147,N_12638,N_13097);
nand U14148 (N_14148,N_12270,N_13761);
or U14149 (N_14149,N_13887,N_13715);
or U14150 (N_14150,N_12778,N_12241);
nand U14151 (N_14151,N_12297,N_12047);
nand U14152 (N_14152,N_12461,N_13143);
and U14153 (N_14153,N_13306,N_13059);
xnor U14154 (N_14154,N_12506,N_13597);
or U14155 (N_14155,N_12532,N_12298);
nor U14156 (N_14156,N_13280,N_13586);
nand U14157 (N_14157,N_13934,N_13141);
xor U14158 (N_14158,N_12345,N_12535);
xor U14159 (N_14159,N_12969,N_12967);
nor U14160 (N_14160,N_12030,N_13460);
nand U14161 (N_14161,N_12699,N_12679);
nand U14162 (N_14162,N_13802,N_13840);
xor U14163 (N_14163,N_12735,N_13981);
or U14164 (N_14164,N_12877,N_12227);
nand U14165 (N_14165,N_12418,N_12404);
nand U14166 (N_14166,N_13041,N_13801);
nand U14167 (N_14167,N_13899,N_12454);
or U14168 (N_14168,N_13151,N_13333);
xor U14169 (N_14169,N_12274,N_12095);
and U14170 (N_14170,N_13594,N_12748);
and U14171 (N_14171,N_13625,N_12737);
nand U14172 (N_14172,N_12007,N_12988);
nor U14173 (N_14173,N_12954,N_12252);
or U14174 (N_14174,N_13985,N_13247);
or U14175 (N_14175,N_13008,N_12057);
xor U14176 (N_14176,N_12716,N_13738);
or U14177 (N_14177,N_13685,N_13152);
nand U14178 (N_14178,N_13268,N_13065);
nor U14179 (N_14179,N_12533,N_13828);
xor U14180 (N_14180,N_13375,N_13769);
nand U14181 (N_14181,N_12283,N_12006);
nor U14182 (N_14182,N_12753,N_13800);
nand U14183 (N_14183,N_13956,N_13138);
or U14184 (N_14184,N_12021,N_12507);
or U14185 (N_14185,N_12728,N_13660);
xor U14186 (N_14186,N_12684,N_12783);
and U14187 (N_14187,N_13101,N_12123);
nor U14188 (N_14188,N_13917,N_13419);
xnor U14189 (N_14189,N_12203,N_13911);
nand U14190 (N_14190,N_13485,N_12321);
nand U14191 (N_14191,N_12878,N_13961);
nor U14192 (N_14192,N_12437,N_12056);
or U14193 (N_14193,N_12369,N_13636);
or U14194 (N_14194,N_12412,N_13171);
nand U14195 (N_14195,N_13627,N_13217);
and U14196 (N_14196,N_12368,N_13923);
or U14197 (N_14197,N_12773,N_13076);
and U14198 (N_14198,N_12049,N_13592);
and U14199 (N_14199,N_13045,N_13706);
nor U14200 (N_14200,N_13376,N_13857);
nand U14201 (N_14201,N_13804,N_12237);
nand U14202 (N_14202,N_12595,N_13218);
nor U14203 (N_14203,N_13821,N_12782);
nor U14204 (N_14204,N_13720,N_12215);
or U14205 (N_14205,N_13305,N_12635);
nor U14206 (N_14206,N_13150,N_12002);
and U14207 (N_14207,N_12603,N_13409);
and U14208 (N_14208,N_13704,N_12411);
nor U14209 (N_14209,N_12565,N_13408);
nand U14210 (N_14210,N_12068,N_13001);
xor U14211 (N_14211,N_13525,N_12069);
xnor U14212 (N_14212,N_12485,N_12094);
nand U14213 (N_14213,N_12916,N_12925);
nor U14214 (N_14214,N_13005,N_12396);
nor U14215 (N_14215,N_12338,N_13803);
or U14216 (N_14216,N_12228,N_12025);
or U14217 (N_14217,N_13182,N_12401);
nor U14218 (N_14218,N_12690,N_12320);
or U14219 (N_14219,N_13843,N_12111);
or U14220 (N_14220,N_13921,N_13047);
xor U14221 (N_14221,N_12307,N_13133);
xnor U14222 (N_14222,N_12184,N_13100);
nand U14223 (N_14223,N_12634,N_13861);
or U14224 (N_14224,N_12680,N_13329);
nor U14225 (N_14225,N_13063,N_13582);
and U14226 (N_14226,N_12247,N_13631);
nor U14227 (N_14227,N_12999,N_13366);
or U14228 (N_14228,N_12709,N_13516);
nor U14229 (N_14229,N_13789,N_12475);
or U14230 (N_14230,N_12172,N_13458);
nor U14231 (N_14231,N_12764,N_12585);
nor U14232 (N_14232,N_13142,N_12193);
and U14233 (N_14233,N_13910,N_12417);
or U14234 (N_14234,N_13697,N_12505);
nor U14235 (N_14235,N_12908,N_13168);
nand U14236 (N_14236,N_12271,N_13946);
nor U14237 (N_14237,N_12103,N_13710);
or U14238 (N_14238,N_12682,N_12807);
or U14239 (N_14239,N_12770,N_12351);
or U14240 (N_14240,N_12384,N_13548);
xnor U14241 (N_14241,N_13507,N_12708);
xnor U14242 (N_14242,N_13188,N_12629);
nor U14243 (N_14243,N_13588,N_12947);
nand U14244 (N_14244,N_13847,N_13405);
nand U14245 (N_14245,N_12923,N_12540);
nor U14246 (N_14246,N_12488,N_12362);
nor U14247 (N_14247,N_12110,N_12696);
nor U14248 (N_14248,N_13979,N_12079);
or U14249 (N_14249,N_12833,N_12568);
nor U14250 (N_14250,N_13102,N_13350);
nor U14251 (N_14251,N_12059,N_13373);
and U14252 (N_14252,N_12062,N_13161);
nor U14253 (N_14253,N_12694,N_12573);
nor U14254 (N_14254,N_12353,N_13155);
nor U14255 (N_14255,N_12991,N_13116);
or U14256 (N_14256,N_12743,N_12832);
or U14257 (N_14257,N_12344,N_12122);
or U14258 (N_14258,N_13935,N_12290);
or U14259 (N_14259,N_12476,N_12912);
or U14260 (N_14260,N_13655,N_13259);
or U14261 (N_14261,N_12519,N_12352);
xor U14262 (N_14262,N_12758,N_12140);
nand U14263 (N_14263,N_12599,N_13289);
nand U14264 (N_14264,N_12127,N_13081);
nor U14265 (N_14265,N_13068,N_12484);
or U14266 (N_14266,N_12426,N_13426);
nand U14267 (N_14267,N_12114,N_13122);
xnor U14268 (N_14268,N_13842,N_12882);
nor U14269 (N_14269,N_13947,N_13967);
nor U14270 (N_14270,N_13779,N_13058);
xor U14271 (N_14271,N_12965,N_13090);
or U14272 (N_14272,N_12734,N_12443);
and U14273 (N_14273,N_12836,N_12142);
xor U14274 (N_14274,N_13606,N_12078);
xnor U14275 (N_14275,N_12326,N_12631);
xnor U14276 (N_14276,N_12462,N_12165);
nor U14277 (N_14277,N_13154,N_12661);
xor U14278 (N_14278,N_12161,N_13916);
or U14279 (N_14279,N_13523,N_13912);
or U14280 (N_14280,N_12772,N_13679);
or U14281 (N_14281,N_13119,N_13888);
or U14282 (N_14282,N_13732,N_12678);
and U14283 (N_14283,N_12131,N_12486);
nand U14284 (N_14284,N_13470,N_13144);
nand U14285 (N_14285,N_13695,N_13107);
or U14286 (N_14286,N_13183,N_12175);
or U14287 (N_14287,N_12074,N_13607);
or U14288 (N_14288,N_13462,N_13998);
xnor U14289 (N_14289,N_13378,N_12360);
nand U14290 (N_14290,N_12073,N_12300);
nand U14291 (N_14291,N_13468,N_12672);
xnor U14292 (N_14292,N_12526,N_13814);
nor U14293 (N_14293,N_12387,N_12730);
or U14294 (N_14294,N_12545,N_13841);
and U14295 (N_14295,N_13290,N_12164);
or U14296 (N_14296,N_12655,N_12789);
nand U14297 (N_14297,N_12340,N_12211);
or U14298 (N_14298,N_13328,N_13538);
nand U14299 (N_14299,N_12306,N_12497);
xor U14300 (N_14300,N_12922,N_12472);
nand U14301 (N_14301,N_12740,N_13984);
nor U14302 (N_14302,N_12996,N_12393);
nand U14303 (N_14303,N_13475,N_12317);
nor U14304 (N_14304,N_13093,N_12216);
and U14305 (N_14305,N_12465,N_13479);
or U14306 (N_14306,N_13729,N_13369);
nand U14307 (N_14307,N_12567,N_12821);
xor U14308 (N_14308,N_13365,N_13267);
xor U14309 (N_14309,N_13284,N_12605);
xor U14310 (N_14310,N_13750,N_13770);
xor U14311 (N_14311,N_13866,N_12174);
nand U14312 (N_14312,N_13839,N_13080);
xnor U14313 (N_14313,N_12425,N_12610);
nand U14314 (N_14314,N_13711,N_13326);
nand U14315 (N_14315,N_13812,N_13025);
nand U14316 (N_14316,N_12780,N_12314);
nand U14317 (N_14317,N_13647,N_13212);
nor U14318 (N_14318,N_12399,N_12198);
and U14319 (N_14319,N_13240,N_13648);
nand U14320 (N_14320,N_12051,N_12529);
or U14321 (N_14321,N_13399,N_12170);
nor U14322 (N_14322,N_13616,N_13415);
or U14323 (N_14323,N_12139,N_12210);
nand U14324 (N_14324,N_13665,N_13398);
xor U14325 (N_14325,N_13167,N_12538);
xor U14326 (N_14326,N_13868,N_12153);
xor U14327 (N_14327,N_13422,N_13300);
nor U14328 (N_14328,N_13114,N_13535);
and U14329 (N_14329,N_12082,N_13509);
nor U14330 (N_14330,N_12264,N_12377);
or U14331 (N_14331,N_13675,N_12275);
nor U14332 (N_14332,N_13229,N_13354);
and U14333 (N_14333,N_12880,N_12668);
and U14334 (N_14334,N_12961,N_13091);
and U14335 (N_14335,N_12128,N_13325);
nor U14336 (N_14336,N_13344,N_13424);
and U14337 (N_14337,N_12931,N_13048);
nor U14338 (N_14338,N_13949,N_12612);
xor U14339 (N_14339,N_12192,N_12618);
nor U14340 (N_14340,N_13508,N_12895);
and U14341 (N_14341,N_13493,N_13077);
xnor U14342 (N_14342,N_13795,N_12265);
nor U14343 (N_14343,N_12424,N_12117);
nor U14344 (N_14344,N_13510,N_12189);
nor U14345 (N_14345,N_12669,N_12660);
or U14346 (N_14346,N_12700,N_13270);
nor U14347 (N_14347,N_12287,N_12200);
and U14348 (N_14348,N_12349,N_12869);
xor U14349 (N_14349,N_13745,N_12844);
xor U14350 (N_14350,N_13312,N_12266);
or U14351 (N_14351,N_12316,N_13805);
nor U14352 (N_14352,N_13807,N_12989);
and U14353 (N_14353,N_13587,N_12614);
nor U14354 (N_14354,N_12951,N_13362);
xnor U14355 (N_14355,N_13469,N_12962);
and U14356 (N_14356,N_12572,N_13854);
or U14357 (N_14357,N_13124,N_13176);
xor U14358 (N_14358,N_13753,N_13512);
nand U14359 (N_14359,N_13954,N_13833);
nor U14360 (N_14360,N_13021,N_12781);
xor U14361 (N_14361,N_13567,N_12796);
and U14362 (N_14362,N_13875,N_12101);
xnor U14363 (N_14363,N_13744,N_13007);
nor U14364 (N_14364,N_13233,N_12035);
or U14365 (N_14365,N_12248,N_12366);
nor U14366 (N_14366,N_12712,N_12291);
nor U14367 (N_14367,N_13235,N_13560);
xnor U14368 (N_14368,N_12984,N_13536);
and U14369 (N_14369,N_13922,N_13776);
or U14370 (N_14370,N_12892,N_12790);
and U14371 (N_14371,N_13846,N_12406);
or U14372 (N_14372,N_13680,N_13236);
or U14373 (N_14373,N_13351,N_13563);
nand U14374 (N_14374,N_13734,N_12898);
or U14375 (N_14375,N_13032,N_12470);
xor U14376 (N_14376,N_13178,N_12732);
nand U14377 (N_14377,N_13530,N_13822);
nand U14378 (N_14378,N_13645,N_13945);
xnor U14379 (N_14379,N_12400,N_13224);
xnor U14380 (N_14380,N_13069,N_13359);
or U14381 (N_14381,N_12093,N_13886);
nor U14382 (N_14382,N_13443,N_12956);
nor U14383 (N_14383,N_12693,N_12640);
nand U14384 (N_14384,N_13900,N_13931);
and U14385 (N_14385,N_12324,N_12692);
or U14386 (N_14386,N_12119,N_13264);
nand U14387 (N_14387,N_13672,N_13860);
and U14388 (N_14388,N_12202,N_12935);
nor U14389 (N_14389,N_12957,N_12040);
or U14390 (N_14390,N_12218,N_12755);
nor U14391 (N_14391,N_12724,N_12808);
or U14392 (N_14392,N_13239,N_12251);
or U14393 (N_14393,N_12017,N_13668);
or U14394 (N_14394,N_13819,N_13372);
or U14395 (N_14395,N_13944,N_13978);
nand U14396 (N_14396,N_13646,N_12196);
nor U14397 (N_14397,N_13004,N_13712);
or U14398 (N_14398,N_12176,N_12917);
or U14399 (N_14399,N_12135,N_12651);
nand U14400 (N_14400,N_13663,N_12380);
or U14401 (N_14401,N_13737,N_13958);
xor U14402 (N_14402,N_13794,N_13282);
nand U14403 (N_14403,N_12530,N_13617);
nor U14404 (N_14404,N_12489,N_12409);
nand U14405 (N_14405,N_12508,N_12058);
xor U14406 (N_14406,N_13198,N_13880);
or U14407 (N_14407,N_12856,N_13628);
nor U14408 (N_14408,N_12235,N_12190);
xnor U14409 (N_14409,N_12955,N_12154);
and U14410 (N_14410,N_13698,N_12226);
and U14411 (N_14411,N_13195,N_13384);
xnor U14412 (N_14412,N_13699,N_13445);
xnor U14413 (N_14413,N_12315,N_13968);
nor U14414 (N_14414,N_13497,N_13971);
xnor U14415 (N_14415,N_12221,N_13552);
and U14416 (N_14416,N_12705,N_12342);
or U14417 (N_14417,N_12864,N_13164);
and U14418 (N_14418,N_13686,N_12091);
nor U14419 (N_14419,N_12289,N_13792);
xor U14420 (N_14420,N_13526,N_13589);
xnor U14421 (N_14421,N_12391,N_12843);
nor U14422 (N_14422,N_13050,N_12125);
nand U14423 (N_14423,N_12803,N_12296);
xor U14424 (N_14424,N_13128,N_13681);
xor U14425 (N_14425,N_13844,N_12029);
or U14426 (N_14426,N_12420,N_12372);
or U14427 (N_14427,N_13214,N_12813);
nor U14428 (N_14428,N_12332,N_12828);
nor U14429 (N_14429,N_13850,N_13894);
nor U14430 (N_14430,N_12163,N_12549);
nor U14431 (N_14431,N_13169,N_13767);
and U14432 (N_14432,N_13514,N_13137);
nand U14433 (N_14433,N_12034,N_13932);
nor U14434 (N_14434,N_13054,N_12906);
nor U14435 (N_14435,N_12656,N_12896);
and U14436 (N_14436,N_13952,N_13953);
nor U14437 (N_14437,N_12994,N_13539);
or U14438 (N_14438,N_13650,N_12075);
xor U14439 (N_14439,N_13404,N_12611);
or U14440 (N_14440,N_13276,N_13599);
nor U14441 (N_14441,N_13158,N_13573);
nor U14442 (N_14442,N_12766,N_13200);
or U14443 (N_14443,N_13816,N_12597);
and U14444 (N_14444,N_13965,N_12625);
and U14445 (N_14445,N_12685,N_12858);
xor U14446 (N_14446,N_13690,N_12421);
nand U14447 (N_14447,N_12607,N_13034);
nand U14448 (N_14448,N_13908,N_12835);
nand U14449 (N_14449,N_13286,N_12137);
nand U14450 (N_14450,N_12008,N_13577);
and U14451 (N_14451,N_13867,N_13347);
xnor U14452 (N_14452,N_12089,N_13432);
xnor U14453 (N_14453,N_13484,N_13322);
xnor U14454 (N_14454,N_12581,N_13046);
xor U14455 (N_14455,N_13696,N_12722);
nor U14456 (N_14456,N_12677,N_13388);
and U14457 (N_14457,N_12849,N_12032);
or U14458 (N_14458,N_12126,N_13988);
nand U14459 (N_14459,N_13827,N_13011);
or U14460 (N_14460,N_13583,N_12150);
nor U14461 (N_14461,N_12992,N_12038);
nor U14462 (N_14462,N_13126,N_12427);
xnor U14463 (N_14463,N_13400,N_12206);
xnor U14464 (N_14464,N_12286,N_12325);
and U14465 (N_14465,N_13749,N_12811);
nand U14466 (N_14466,N_12441,N_12473);
or U14467 (N_14467,N_13478,N_13189);
or U14468 (N_14468,N_13368,N_13848);
or U14469 (N_14469,N_13620,N_12891);
and U14470 (N_14470,N_13296,N_12707);
nand U14471 (N_14471,N_12667,N_12897);
nand U14472 (N_14472,N_12105,N_13836);
or U14473 (N_14473,N_13383,N_13623);
and U14474 (N_14474,N_12151,N_13336);
nand U14475 (N_14475,N_13078,N_13016);
and U14476 (N_14476,N_13676,N_13859);
nor U14477 (N_14477,N_12852,N_12566);
nor U14478 (N_14478,N_13664,N_13394);
and U14479 (N_14479,N_12571,N_13575);
xor U14480 (N_14480,N_12839,N_13601);
and U14481 (N_14481,N_12845,N_13755);
or U14482 (N_14482,N_12162,N_13241);
or U14483 (N_14483,N_13129,N_12765);
and U14484 (N_14484,N_12958,N_12943);
or U14485 (N_14485,N_13070,N_12249);
or U14486 (N_14486,N_13635,N_13210);
and U14487 (N_14487,N_12179,N_13830);
nand U14488 (N_14488,N_13495,N_13056);
xor U14489 (N_14489,N_13315,N_13654);
or U14490 (N_14490,N_13473,N_13966);
nand U14491 (N_14491,N_13382,N_13074);
or U14492 (N_14492,N_13831,N_13780);
and U14493 (N_14493,N_13015,N_13657);
xor U14494 (N_14494,N_13834,N_13385);
nand U14495 (N_14495,N_12053,N_13716);
and U14496 (N_14496,N_12795,N_13153);
nand U14497 (N_14497,N_13618,N_12802);
nor U14498 (N_14498,N_12930,N_13626);
xor U14499 (N_14499,N_13722,N_13260);
nor U14500 (N_14500,N_13996,N_12592);
nor U14501 (N_14501,N_13318,N_13751);
nor U14502 (N_14502,N_12292,N_13919);
xor U14503 (N_14503,N_13823,N_12650);
xor U14504 (N_14504,N_12061,N_12367);
or U14505 (N_14505,N_12239,N_13970);
and U14506 (N_14506,N_13174,N_12745);
and U14507 (N_14507,N_13380,N_12866);
nor U14508 (N_14508,N_12695,N_12460);
or U14509 (N_14509,N_13377,N_12829);
xor U14510 (N_14510,N_13316,N_12759);
xnor U14511 (N_14511,N_12181,N_12842);
and U14512 (N_14512,N_13283,N_13196);
and U14513 (N_14513,N_12562,N_13106);
and U14514 (N_14514,N_13345,N_13731);
nand U14515 (N_14515,N_13231,N_12430);
xor U14516 (N_14516,N_12509,N_12382);
or U14517 (N_14517,N_12511,N_12622);
xor U14518 (N_14518,N_13768,N_13186);
xor U14519 (N_14519,N_13317,N_13725);
xor U14520 (N_14520,N_13824,N_12050);
xor U14521 (N_14521,N_12598,N_13550);
or U14522 (N_14522,N_13856,N_13902);
or U14523 (N_14523,N_13459,N_12711);
nand U14524 (N_14524,N_12060,N_13471);
xor U14525 (N_14525,N_12723,N_13492);
nand U14526 (N_14526,N_13000,N_12857);
or U14527 (N_14527,N_12381,N_13578);
and U14528 (N_14528,N_12014,N_13598);
and U14529 (N_14529,N_13146,N_13179);
nor U14530 (N_14530,N_12793,N_13251);
or U14531 (N_14531,N_13234,N_13983);
nand U14532 (N_14532,N_13295,N_12990);
and U14533 (N_14533,N_13817,N_13547);
nor U14534 (N_14534,N_12977,N_13992);
xnor U14535 (N_14535,N_12729,N_12544);
xor U14536 (N_14536,N_13689,N_12262);
nor U14537 (N_14537,N_13624,N_12440);
xnor U14538 (N_14538,N_13933,N_12337);
nor U14539 (N_14539,N_13130,N_12392);
xnor U14540 (N_14540,N_12386,N_12941);
nor U14541 (N_14541,N_13735,N_13262);
nor U14542 (N_14542,N_13778,N_12953);
nand U14543 (N_14543,N_13870,N_13465);
nor U14544 (N_14544,N_12222,N_13504);
nor U14545 (N_14545,N_12741,N_13746);
nor U14546 (N_14546,N_13837,N_12363);
or U14547 (N_14547,N_12948,N_13271);
nor U14548 (N_14548,N_12229,N_12706);
nor U14549 (N_14549,N_12763,N_13136);
nand U14550 (N_14550,N_13758,N_13060);
nor U14551 (N_14551,N_12480,N_13309);
xnor U14552 (N_14552,N_12028,N_13044);
or U14553 (N_14553,N_12295,N_13263);
nand U14554 (N_14554,N_13278,N_13505);
or U14555 (N_14555,N_13553,N_13441);
xor U14556 (N_14556,N_13320,N_13574);
and U14557 (N_14557,N_12899,N_12993);
xor U14558 (N_14558,N_12648,N_13556);
and U14559 (N_14559,N_12446,N_12550);
or U14560 (N_14560,N_13162,N_12183);
and U14561 (N_14561,N_13611,N_12168);
and U14562 (N_14562,N_13602,N_13783);
nand U14563 (N_14563,N_13747,N_12477);
nand U14564 (N_14564,N_12968,N_13003);
or U14565 (N_14565,N_12861,N_12494);
and U14566 (N_14566,N_13565,N_13604);
or U14567 (N_14567,N_12940,N_12092);
nor U14568 (N_14568,N_12946,N_13237);
and U14569 (N_14569,N_12245,N_13643);
nand U14570 (N_14570,N_13614,N_12177);
or U14571 (N_14571,N_13030,N_13542);
nand U14572 (N_14572,N_13012,N_13748);
nor U14573 (N_14573,N_12288,N_12985);
xnor U14574 (N_14574,N_13927,N_12318);
nand U14575 (N_14575,N_13619,N_12171);
and U14576 (N_14576,N_13499,N_13754);
nor U14577 (N_14577,N_12447,N_12883);
nand U14578 (N_14578,N_12335,N_12085);
nor U14579 (N_14579,N_13942,N_13466);
xnor U14580 (N_14580,N_13724,N_12261);
xnor U14581 (N_14581,N_13327,N_13334);
and U14582 (N_14582,N_13808,N_13040);
nand U14583 (N_14583,N_13600,N_12591);
nor U14584 (N_14584,N_12322,N_13337);
xor U14585 (N_14585,N_12428,N_12365);
or U14586 (N_14586,N_13703,N_12662);
or U14587 (N_14587,N_13346,N_13895);
nand U14588 (N_14588,N_13987,N_13170);
and U14589 (N_14589,N_13498,N_13702);
and U14590 (N_14590,N_12136,N_13177);
and U14591 (N_14591,N_13544,N_13793);
and U14592 (N_14592,N_13879,N_13786);
or U14593 (N_14593,N_12688,N_12555);
nor U14594 (N_14594,N_13464,N_12358);
nand U14595 (N_14595,N_13709,N_13406);
and U14596 (N_14596,N_12714,N_12872);
nor U14597 (N_14597,N_13835,N_13348);
nor U14598 (N_14598,N_12671,N_12911);
and U14599 (N_14599,N_13255,N_12003);
xnor U14600 (N_14600,N_12055,N_13250);
xor U14601 (N_14601,N_12995,N_13829);
nand U14602 (N_14602,N_13314,N_13430);
or U14603 (N_14603,N_13973,N_13435);
nand U14604 (N_14604,N_12044,N_13773);
nand U14605 (N_14605,N_12863,N_13593);
nand U14606 (N_14606,N_12209,N_12016);
xnor U14607 (N_14607,N_13630,N_13414);
xnor U14608 (N_14608,N_13997,N_13683);
and U14609 (N_14609,N_13311,N_13254);
xnor U14610 (N_14610,N_13222,N_13342);
nand U14611 (N_14611,N_12479,N_12416);
and U14612 (N_14612,N_12774,N_12945);
nand U14613 (N_14613,N_13936,N_13569);
nand U14614 (N_14614,N_13909,N_12838);
xor U14615 (N_14615,N_12979,N_13855);
nand U14616 (N_14616,N_13244,N_12579);
and U14617 (N_14617,N_13039,N_12559);
or U14618 (N_14618,N_13531,N_12503);
nand U14619 (N_14619,N_13511,N_12370);
xnor U14620 (N_14620,N_12018,N_12973);
and U14621 (N_14621,N_13740,N_12536);
and U14622 (N_14622,N_13094,N_13298);
nand U14623 (N_14623,N_12214,N_12713);
nand U14624 (N_14624,N_12963,N_12847);
xnor U14625 (N_14625,N_12478,N_12515);
nor U14626 (N_14626,N_12582,N_13449);
and U14627 (N_14627,N_12005,N_13002);
xor U14628 (N_14628,N_12936,N_12496);
and U14629 (N_14629,N_13386,N_12504);
or U14630 (N_14630,N_13528,N_12578);
nor U14631 (N_14631,N_13413,N_13073);
nand U14632 (N_14632,N_12525,N_12333);
nand U14633 (N_14633,N_12388,N_13907);
nand U14634 (N_14634,N_12815,N_12596);
and U14635 (N_14635,N_12072,N_13165);
nand U14636 (N_14636,N_12626,N_12433);
and U14637 (N_14637,N_13872,N_13223);
nand U14638 (N_14638,N_12419,N_13940);
and U14639 (N_14639,N_13637,N_13760);
nand U14640 (N_14640,N_13662,N_13420);
or U14641 (N_14641,N_13639,N_12187);
and U14642 (N_14642,N_12173,N_12981);
or U14643 (N_14643,N_13632,N_12601);
and U14644 (N_14644,N_12169,N_12900);
xnor U14645 (N_14645,N_12088,N_13782);
and U14646 (N_14646,N_12375,N_13974);
nor U14647 (N_14647,N_12108,N_12915);
nand U14648 (N_14648,N_12830,N_13104);
or U14649 (N_14649,N_13513,N_12942);
xnor U14650 (N_14650,N_12133,N_13157);
xnor U14651 (N_14651,N_13739,N_13453);
nor U14652 (N_14652,N_13938,N_13356);
or U14653 (N_14653,N_13815,N_12471);
xor U14654 (N_14654,N_12086,N_13020);
xnor U14655 (N_14655,N_13467,N_12738);
or U14656 (N_14656,N_13173,N_13736);
nor U14657 (N_14657,N_12099,N_12310);
xor U14658 (N_14658,N_12354,N_12697);
xnor U14659 (N_14659,N_13395,N_13551);
nand U14660 (N_14660,N_13905,N_13075);
and U14661 (N_14661,N_13294,N_13232);
or U14662 (N_14662,N_13502,N_13930);
nor U14663 (N_14663,N_12453,N_13024);
nand U14664 (N_14664,N_12894,N_12939);
and U14665 (N_14665,N_12499,N_12456);
nand U14666 (N_14666,N_12282,N_12166);
nand U14667 (N_14667,N_13878,N_12336);
and U14668 (N_14668,N_12243,N_12586);
and U14669 (N_14669,N_13813,N_12301);
xnor U14670 (N_14670,N_12130,N_13733);
nor U14671 (N_14671,N_12809,N_13147);
xor U14672 (N_14672,N_12464,N_13371);
xnor U14673 (N_14673,N_13564,N_12762);
and U14674 (N_14674,N_12641,N_13926);
xnor U14675 (N_14675,N_13451,N_13500);
xor U14676 (N_14676,N_12106,N_13055);
xnor U14677 (N_14677,N_12299,N_12812);
nor U14678 (N_14678,N_13417,N_12450);
and U14679 (N_14679,N_12254,N_12147);
or U14680 (N_14680,N_13448,N_12518);
and U14681 (N_14681,N_13201,N_12949);
and U14682 (N_14682,N_12583,N_13293);
and U14683 (N_14683,N_13135,N_12552);
or U14684 (N_14684,N_12546,N_13603);
or U14685 (N_14685,N_12937,N_13277);
and U14686 (N_14686,N_13893,N_13436);
xor U14687 (N_14687,N_13881,N_12276);
nand U14688 (N_14688,N_13666,N_12201);
and U14689 (N_14689,N_12733,N_12825);
and U14690 (N_14690,N_13527,N_12974);
and U14691 (N_14691,N_13199,N_13439);
nor U14692 (N_14692,N_12822,N_13810);
nand U14693 (N_14693,N_12468,N_13127);
and U14694 (N_14694,N_13521,N_13890);
or U14695 (N_14695,N_13608,N_12557);
or U14696 (N_14696,N_13028,N_12804);
xnor U14697 (N_14697,N_12952,N_13506);
and U14698 (N_14698,N_12258,N_12717);
xnor U14699 (N_14699,N_13389,N_13651);
nor U14700 (N_14700,N_13489,N_12054);
or U14701 (N_14701,N_12144,N_13113);
nand U14702 (N_14702,N_13450,N_12810);
nor U14703 (N_14703,N_13898,N_12594);
and U14704 (N_14704,N_13920,N_13010);
or U14705 (N_14705,N_13285,N_12268);
xor U14706 (N_14706,N_13243,N_13721);
and U14707 (N_14707,N_12432,N_13790);
and U14708 (N_14708,N_12590,N_12149);
and U14709 (N_14709,N_13862,N_13037);
nor U14710 (N_14710,N_13018,N_13960);
nor U14711 (N_14711,N_12960,N_12837);
and U14712 (N_14712,N_13480,N_12097);
or U14713 (N_14713,N_13134,N_13123);
nand U14714 (N_14714,N_12232,N_13051);
nand U14715 (N_14715,N_13494,N_13275);
and U14716 (N_14716,N_12816,N_13791);
nor U14717 (N_14717,N_12498,N_13140);
nand U14718 (N_14718,N_12015,N_12260);
and U14719 (N_14719,N_12731,N_13669);
nand U14720 (N_14720,N_12627,N_12742);
and U14721 (N_14721,N_13796,N_13049);
nand U14722 (N_14722,N_12308,N_13105);
nand U14723 (N_14723,N_13219,N_12950);
or U14724 (N_14724,N_13595,N_13248);
and U14725 (N_14725,N_12666,N_13172);
nand U14726 (N_14726,N_13017,N_13705);
nor U14727 (N_14727,N_13192,N_13490);
or U14728 (N_14728,N_12619,N_13185);
nand U14729 (N_14729,N_12256,N_12520);
xor U14730 (N_14730,N_12285,N_12938);
and U14731 (N_14731,N_12495,N_12779);
nand U14732 (N_14732,N_13299,N_13906);
nand U14733 (N_14733,N_12284,N_12195);
or U14734 (N_14734,N_12199,N_12944);
nand U14735 (N_14735,N_12806,N_13014);
and U14736 (N_14736,N_12124,N_13391);
xnor U14737 (N_14737,N_13472,N_12721);
or U14738 (N_14738,N_12769,N_13454);
and U14739 (N_14739,N_12255,N_12818);
or U14740 (N_14740,N_13896,N_13095);
nor U14741 (N_14741,N_12309,N_13897);
and U14742 (N_14742,N_12726,N_12379);
and U14743 (N_14743,N_12577,N_12100);
xor U14744 (N_14744,N_13982,N_12076);
nor U14745 (N_14745,N_12739,N_12364);
xor U14746 (N_14746,N_12267,N_13520);
nand U14747 (N_14747,N_12558,N_12727);
nand U14748 (N_14748,N_13313,N_13718);
nor U14749 (N_14749,N_13653,N_13741);
nand U14750 (N_14750,N_13423,N_13891);
and U14751 (N_14751,N_13341,N_13714);
nand U14752 (N_14752,N_13098,N_13109);
nand U14753 (N_14753,N_12304,N_13883);
xnor U14754 (N_14754,N_12361,N_12971);
nand U14755 (N_14755,N_12281,N_12553);
nand U14756 (N_14756,N_13086,N_12652);
or U14757 (N_14757,N_13033,N_13673);
and U14758 (N_14758,N_12576,N_13765);
xor U14759 (N_14759,N_12096,N_12563);
xor U14760 (N_14760,N_12220,N_12980);
and U14761 (N_14761,N_13555,N_13656);
or U14762 (N_14762,N_13440,N_12580);
or U14763 (N_14763,N_12715,N_13288);
nor U14764 (N_14764,N_13869,N_12767);
nand U14765 (N_14765,N_13529,N_12157);
nand U14766 (N_14766,N_13719,N_12205);
or U14767 (N_14767,N_13390,N_13501);
or U14768 (N_14768,N_13266,N_12884);
xor U14769 (N_14769,N_13216,N_13962);
nand U14770 (N_14770,N_12543,N_12280);
nand U14771 (N_14771,N_12272,N_12987);
xnor U14772 (N_14772,N_13957,N_13584);
or U14773 (N_14773,N_12865,N_12305);
nand U14774 (N_14774,N_13707,N_12208);
and U14775 (N_14775,N_13434,N_13321);
nor U14776 (N_14776,N_12098,N_13634);
or U14777 (N_14777,N_12904,N_12204);
xnor U14778 (N_14778,N_12834,N_13642);
nand U14779 (N_14779,N_12013,N_13777);
nor U14780 (N_14780,N_13131,N_13612);
nor U14781 (N_14781,N_12132,N_12207);
nand U14782 (N_14782,N_12429,N_13762);
and U14783 (N_14783,N_13554,N_13456);
and U14784 (N_14784,N_13175,N_13928);
nor U14785 (N_14785,N_13397,N_13085);
nor U14786 (N_14786,N_12436,N_13532);
or U14787 (N_14787,N_13877,N_12373);
nand U14788 (N_14788,N_13253,N_12616);
xor U14789 (N_14789,N_12710,N_12514);
or U14790 (N_14790,N_13579,N_13381);
or U14791 (N_14791,N_13392,N_12138);
nor U14792 (N_14792,N_13950,N_12071);
and U14793 (N_14793,N_12920,N_12442);
nand U14794 (N_14794,N_13139,N_12160);
nor U14795 (N_14795,N_13402,N_13013);
nand U14796 (N_14796,N_13545,N_13301);
and U14797 (N_14797,N_13524,N_13163);
or U14798 (N_14798,N_13488,N_13568);
or U14799 (N_14799,N_13622,N_12820);
and U14800 (N_14800,N_12064,N_12761);
or U14801 (N_14801,N_13303,N_12063);
or U14802 (N_14802,N_12019,N_12302);
nand U14803 (N_14803,N_12776,N_12786);
or U14804 (N_14804,N_12848,N_12327);
and U14805 (N_14805,N_13159,N_13558);
nor U14806 (N_14806,N_12664,N_13281);
or U14807 (N_14807,N_12534,N_12797);
and U14808 (N_14808,N_12278,N_12020);
or U14809 (N_14809,N_12148,N_12250);
and U14810 (N_14810,N_12589,N_13691);
nor U14811 (N_14811,N_13798,N_13066);
nor U14812 (N_14812,N_13742,N_13743);
and U14813 (N_14813,N_13522,N_13763);
or U14814 (N_14814,N_12134,N_13481);
nor U14815 (N_14815,N_12673,N_13181);
xor U14816 (N_14816,N_13205,N_13572);
and U14817 (N_14817,N_13989,N_13964);
nand U14818 (N_14818,N_13644,N_12888);
xnor U14819 (N_14819,N_12799,N_12676);
nor U14820 (N_14820,N_12754,N_13019);
xnor U14821 (N_14821,N_12885,N_12855);
and U14822 (N_14822,N_12791,N_13788);
xnor U14823 (N_14823,N_12152,N_12860);
xnor U14824 (N_14824,N_13213,N_12120);
nand U14825 (N_14825,N_13549,N_12263);
and U14826 (N_14826,N_13156,N_13027);
xor U14827 (N_14827,N_12879,N_13187);
or U14828 (N_14828,N_13688,N_13865);
or U14829 (N_14829,N_12760,N_12907);
or U14830 (N_14830,N_12823,N_12527);
or U14831 (N_14831,N_12609,N_12523);
xnor U14832 (N_14832,N_13367,N_12225);
nor U14833 (N_14833,N_12191,N_12959);
nor U14834 (N_14834,N_13319,N_13403);
nand U14835 (N_14835,N_12814,N_12182);
xor U14836 (N_14836,N_12001,N_12402);
and U14837 (N_14837,N_12874,N_12524);
and U14838 (N_14838,N_13991,N_13038);
or U14839 (N_14839,N_12644,N_12501);
or U14840 (N_14840,N_12356,N_12928);
or U14841 (N_14841,N_12905,N_12457);
and U14842 (N_14842,N_12313,N_12398);
or U14843 (N_14843,N_12052,N_12435);
or U14844 (N_14844,N_13428,N_12224);
or U14845 (N_14845,N_12841,N_12039);
nand U14846 (N_14846,N_13361,N_13220);
xor U14847 (N_14847,N_12180,N_13546);
and U14848 (N_14848,N_12982,N_13667);
and U14849 (N_14849,N_13658,N_12083);
nand U14850 (N_14850,N_13148,N_13995);
or U14851 (N_14851,N_13291,N_13446);
nand U14852 (N_14852,N_13924,N_13717);
nor U14853 (N_14853,N_12887,N_13082);
nor U14854 (N_14854,N_12868,N_12269);
nand U14855 (N_14855,N_13559,N_12042);
xnor U14856 (N_14856,N_13118,N_13515);
xnor U14857 (N_14857,N_12357,N_13084);
or U14858 (N_14858,N_13452,N_12431);
and U14859 (N_14859,N_12188,N_13330);
xnor U14860 (N_14860,N_13360,N_13809);
and U14861 (N_14861,N_13571,N_12704);
or U14862 (N_14862,N_12347,N_13903);
and U14863 (N_14863,N_12482,N_12698);
nand U14864 (N_14864,N_12129,N_13349);
xor U14865 (N_14865,N_13166,N_12784);
or U14866 (N_14866,N_12067,N_12608);
nand U14867 (N_14867,N_13576,N_13661);
nand U14868 (N_14868,N_12889,N_12918);
or U14869 (N_14869,N_13083,N_12569);
xnor U14870 (N_14870,N_13067,N_13023);
and U14871 (N_14871,N_12893,N_12438);
and U14872 (N_14872,N_12346,N_13772);
and U14873 (N_14873,N_13297,N_12675);
or U14874 (N_14874,N_13682,N_13797);
or U14875 (N_14875,N_12824,N_12045);
nand U14876 (N_14876,N_13125,N_12574);
nand U14877 (N_14877,N_12623,N_13596);
nor U14878 (N_14878,N_12219,N_12556);
xor U14879 (N_14879,N_12564,N_12768);
and U14880 (N_14880,N_12244,N_12541);
and U14881 (N_14881,N_12434,N_13486);
nand U14882 (N_14882,N_13787,N_13864);
and U14883 (N_14883,N_13757,N_13261);
or U14884 (N_14884,N_12862,N_13215);
xnor U14885 (N_14885,N_13876,N_13537);
xor U14886 (N_14886,N_13339,N_12584);
nor U14887 (N_14887,N_12986,N_12978);
xnor U14888 (N_14888,N_12870,N_12934);
nor U14889 (N_14889,N_13257,N_13609);
nand U14890 (N_14890,N_12902,N_12575);
xnor U14891 (N_14891,N_13874,N_13393);
xnor U14892 (N_14892,N_13727,N_12649);
or U14893 (N_14893,N_13641,N_12010);
xnor U14894 (N_14894,N_12718,N_12118);
xnor U14895 (N_14895,N_12439,N_12659);
or U14896 (N_14896,N_13269,N_13421);
nor U14897 (N_14897,N_13610,N_13659);
and U14898 (N_14898,N_12975,N_13352);
and U14899 (N_14899,N_13358,N_13581);
nor U14900 (N_14900,N_13640,N_12725);
or U14901 (N_14901,N_12331,N_13845);
and U14902 (N_14902,N_12185,N_12840);
nand U14903 (N_14903,N_12636,N_12328);
nand U14904 (N_14904,N_12374,N_13374);
and U14905 (N_14905,N_13972,N_12752);
nor U14906 (N_14906,N_12890,N_13826);
and U14907 (N_14907,N_12444,N_13993);
or U14908 (N_14908,N_13006,N_12240);
and U14909 (N_14909,N_12600,N_13570);
or U14910 (N_14910,N_12750,N_12413);
nor U14911 (N_14911,N_12871,N_13534);
nand U14912 (N_14912,N_12041,N_12031);
nor U14913 (N_14913,N_12593,N_12921);
nand U14914 (N_14914,N_12876,N_13099);
xor U14915 (N_14915,N_13433,N_13629);
nand U14916 (N_14916,N_12359,N_12463);
and U14917 (N_14917,N_13774,N_13613);
nand U14918 (N_14918,N_12512,N_13092);
or U14919 (N_14919,N_13053,N_13852);
or U14920 (N_14920,N_12794,N_12819);
nor U14921 (N_14921,N_13379,N_12109);
or U14922 (N_14922,N_13728,N_13036);
xor U14923 (N_14923,N_12846,N_13764);
xor U14924 (N_14924,N_12643,N_13463);
nor U14925 (N_14925,N_12924,N_13429);
and U14926 (N_14926,N_13882,N_13202);
or U14927 (N_14927,N_13061,N_12932);
nor U14928 (N_14928,N_12703,N_13043);
nor U14929 (N_14929,N_12156,N_13108);
xor U14930 (N_14930,N_12217,N_12970);
nor U14931 (N_14931,N_13444,N_12311);
xor U14932 (N_14932,N_13194,N_12011);
and U14933 (N_14933,N_12334,N_13671);
nor U14934 (N_14934,N_12751,N_12452);
or U14935 (N_14935,N_12012,N_13700);
xor U14936 (N_14936,N_13975,N_13693);
and U14937 (N_14937,N_13418,N_12560);
nor U14938 (N_14938,N_12647,N_12642);
nand U14939 (N_14939,N_13088,N_12397);
and U14940 (N_14940,N_12070,N_13684);
and U14941 (N_14941,N_12223,N_13120);
or U14942 (N_14942,N_13072,N_13918);
nand U14943 (N_14943,N_13287,N_12319);
nor U14944 (N_14944,N_13035,N_12646);
or U14945 (N_14945,N_12663,N_12236);
xor U14946 (N_14946,N_13227,N_12146);
xnor U14947 (N_14947,N_13079,N_12528);
xnor U14948 (N_14948,N_12293,N_12026);
nor U14949 (N_14949,N_12212,N_13832);
and U14950 (N_14950,N_13387,N_13103);
or U14951 (N_14951,N_12467,N_13230);
nor U14952 (N_14952,N_13980,N_13209);
xnor U14953 (N_14953,N_12658,N_13959);
nor U14954 (N_14954,N_12323,N_12517);
nor U14955 (N_14955,N_12826,N_13771);
or U14956 (N_14956,N_13292,N_12859);
nand U14957 (N_14957,N_12046,N_12606);
nand U14958 (N_14958,N_12378,N_12886);
nor U14959 (N_14959,N_12929,N_13487);
nor U14960 (N_14960,N_12445,N_13111);
nand U14961 (N_14961,N_12159,N_13427);
and U14962 (N_14962,N_12112,N_13026);
nor U14963 (N_14963,N_13723,N_13042);
and U14964 (N_14964,N_13941,N_13335);
xnor U14965 (N_14965,N_12561,N_12701);
or U14966 (N_14966,N_12719,N_12394);
nor U14967 (N_14967,N_13274,N_12277);
and U14968 (N_14968,N_13206,N_12253);
or U14969 (N_14969,N_13820,N_12033);
and U14970 (N_14970,N_13915,N_12777);
nor U14971 (N_14971,N_12458,N_12257);
xnor U14972 (N_14972,N_13323,N_13999);
xnor U14973 (N_14973,N_13273,N_13029);
and U14974 (N_14974,N_13411,N_13955);
nand U14975 (N_14975,N_13566,N_12513);
or U14976 (N_14976,N_12329,N_12474);
or U14977 (N_14977,N_12355,N_13561);
or U14978 (N_14978,N_12186,N_12854);
nor U14979 (N_14979,N_12102,N_12231);
or U14980 (N_14980,N_13331,N_12913);
nand U14981 (N_14981,N_13503,N_12539);
and U14982 (N_14982,N_13461,N_12683);
xor U14983 (N_14983,N_12736,N_12389);
and U14984 (N_14984,N_12490,N_13858);
and U14985 (N_14985,N_12521,N_13677);
xor U14986 (N_14986,N_12410,N_13621);
and U14987 (N_14987,N_13357,N_12522);
or U14988 (N_14988,N_13591,N_12273);
or U14989 (N_14989,N_13302,N_13145);
nand U14990 (N_14990,N_12343,N_12875);
nand U14991 (N_14991,N_12080,N_12087);
and U14992 (N_14992,N_12749,N_12615);
or U14993 (N_14993,N_13939,N_12744);
nand U14994 (N_14994,N_12415,N_12043);
and U14995 (N_14995,N_12746,N_12414);
or U14996 (N_14996,N_12009,N_12113);
xor U14997 (N_14997,N_13775,N_13670);
and U14998 (N_14998,N_12771,N_13238);
xor U14999 (N_14999,N_13355,N_13474);
and U15000 (N_15000,N_13333,N_12000);
and U15001 (N_15001,N_12209,N_12358);
or U15002 (N_15002,N_12553,N_13338);
nor U15003 (N_15003,N_13642,N_12966);
nor U15004 (N_15004,N_13597,N_13394);
nand U15005 (N_15005,N_13809,N_13007);
nor U15006 (N_15006,N_12358,N_13900);
and U15007 (N_15007,N_13631,N_12928);
and U15008 (N_15008,N_12618,N_13733);
or U15009 (N_15009,N_12013,N_13084);
nor U15010 (N_15010,N_12812,N_13297);
nand U15011 (N_15011,N_13662,N_13596);
or U15012 (N_15012,N_13969,N_13533);
nand U15013 (N_15013,N_12486,N_12261);
nor U15014 (N_15014,N_12661,N_13305);
and U15015 (N_15015,N_12815,N_12289);
nand U15016 (N_15016,N_13392,N_13842);
and U15017 (N_15017,N_12421,N_13720);
or U15018 (N_15018,N_12765,N_12055);
xnor U15019 (N_15019,N_13002,N_12370);
or U15020 (N_15020,N_13028,N_12042);
or U15021 (N_15021,N_13373,N_13312);
and U15022 (N_15022,N_12377,N_12066);
and U15023 (N_15023,N_13203,N_13855);
nand U15024 (N_15024,N_12737,N_13317);
nand U15025 (N_15025,N_12537,N_12265);
and U15026 (N_15026,N_12984,N_12294);
nand U15027 (N_15027,N_13915,N_13832);
nor U15028 (N_15028,N_13848,N_12986);
xnor U15029 (N_15029,N_13548,N_13289);
or U15030 (N_15030,N_12045,N_12614);
nand U15031 (N_15031,N_12150,N_13781);
nand U15032 (N_15032,N_13467,N_13021);
nor U15033 (N_15033,N_13512,N_13412);
nand U15034 (N_15034,N_12058,N_13181);
or U15035 (N_15035,N_13902,N_13666);
nor U15036 (N_15036,N_12768,N_12377);
and U15037 (N_15037,N_13206,N_13172);
nand U15038 (N_15038,N_13064,N_12376);
nand U15039 (N_15039,N_12822,N_12300);
xor U15040 (N_15040,N_13200,N_13918);
nand U15041 (N_15041,N_12946,N_13965);
and U15042 (N_15042,N_12470,N_12816);
and U15043 (N_15043,N_12569,N_13834);
or U15044 (N_15044,N_13460,N_13128);
nor U15045 (N_15045,N_12926,N_12847);
or U15046 (N_15046,N_13028,N_13122);
nand U15047 (N_15047,N_12015,N_13310);
or U15048 (N_15048,N_13801,N_13049);
and U15049 (N_15049,N_12365,N_12661);
xor U15050 (N_15050,N_13554,N_13583);
and U15051 (N_15051,N_12068,N_13243);
and U15052 (N_15052,N_13930,N_13361);
and U15053 (N_15053,N_13349,N_12579);
xnor U15054 (N_15054,N_12417,N_12273);
xor U15055 (N_15055,N_12223,N_13704);
nand U15056 (N_15056,N_13330,N_13527);
nand U15057 (N_15057,N_13779,N_13108);
nor U15058 (N_15058,N_12440,N_13608);
nor U15059 (N_15059,N_13355,N_13516);
xor U15060 (N_15060,N_13422,N_13918);
xnor U15061 (N_15061,N_12134,N_13002);
nand U15062 (N_15062,N_12590,N_13424);
nand U15063 (N_15063,N_13945,N_13890);
nor U15064 (N_15064,N_13562,N_13403);
and U15065 (N_15065,N_13859,N_13127);
nand U15066 (N_15066,N_12031,N_12288);
xor U15067 (N_15067,N_13964,N_13936);
nand U15068 (N_15068,N_13431,N_13767);
xnor U15069 (N_15069,N_12477,N_13900);
xnor U15070 (N_15070,N_12011,N_13273);
xor U15071 (N_15071,N_12967,N_13722);
nor U15072 (N_15072,N_12557,N_12040);
nor U15073 (N_15073,N_12336,N_13408);
or U15074 (N_15074,N_13779,N_12999);
and U15075 (N_15075,N_13123,N_12162);
or U15076 (N_15076,N_13786,N_13512);
nand U15077 (N_15077,N_13364,N_12182);
nor U15078 (N_15078,N_12446,N_12375);
nor U15079 (N_15079,N_12888,N_13454);
nand U15080 (N_15080,N_12595,N_13068);
nor U15081 (N_15081,N_13632,N_12036);
or U15082 (N_15082,N_12708,N_13226);
and U15083 (N_15083,N_13531,N_13505);
and U15084 (N_15084,N_12005,N_13892);
nand U15085 (N_15085,N_13489,N_12577);
nand U15086 (N_15086,N_12892,N_12769);
and U15087 (N_15087,N_12732,N_12554);
nand U15088 (N_15088,N_13920,N_13991);
or U15089 (N_15089,N_13552,N_13792);
and U15090 (N_15090,N_12517,N_12721);
xor U15091 (N_15091,N_13221,N_13943);
xnor U15092 (N_15092,N_12602,N_13696);
and U15093 (N_15093,N_12015,N_13918);
nor U15094 (N_15094,N_13750,N_13717);
and U15095 (N_15095,N_12176,N_13671);
or U15096 (N_15096,N_13647,N_13053);
xnor U15097 (N_15097,N_13751,N_13910);
or U15098 (N_15098,N_12137,N_13915);
and U15099 (N_15099,N_13966,N_12095);
xnor U15100 (N_15100,N_12729,N_12311);
nor U15101 (N_15101,N_13439,N_12600);
nor U15102 (N_15102,N_12067,N_13232);
and U15103 (N_15103,N_12851,N_12263);
or U15104 (N_15104,N_13245,N_12302);
xor U15105 (N_15105,N_12322,N_12119);
xnor U15106 (N_15106,N_13679,N_12697);
xnor U15107 (N_15107,N_12298,N_13197);
xnor U15108 (N_15108,N_13306,N_12170);
nand U15109 (N_15109,N_13461,N_12327);
nand U15110 (N_15110,N_12319,N_12535);
and U15111 (N_15111,N_12430,N_13298);
and U15112 (N_15112,N_13051,N_12429);
or U15113 (N_15113,N_13259,N_13156);
and U15114 (N_15114,N_13516,N_12859);
nor U15115 (N_15115,N_13004,N_12645);
nand U15116 (N_15116,N_13815,N_13770);
and U15117 (N_15117,N_12182,N_13705);
nand U15118 (N_15118,N_13287,N_13789);
nor U15119 (N_15119,N_12130,N_12076);
nand U15120 (N_15120,N_13120,N_12627);
xor U15121 (N_15121,N_13488,N_13936);
or U15122 (N_15122,N_12524,N_13393);
nand U15123 (N_15123,N_13886,N_12281);
and U15124 (N_15124,N_13004,N_13432);
and U15125 (N_15125,N_13887,N_13294);
xnor U15126 (N_15126,N_13582,N_12738);
nand U15127 (N_15127,N_12956,N_12816);
or U15128 (N_15128,N_12727,N_12941);
nand U15129 (N_15129,N_12362,N_12325);
and U15130 (N_15130,N_13655,N_13357);
and U15131 (N_15131,N_12105,N_12379);
or U15132 (N_15132,N_13490,N_12581);
and U15133 (N_15133,N_12279,N_12894);
nor U15134 (N_15134,N_12296,N_12355);
nor U15135 (N_15135,N_12589,N_13033);
nand U15136 (N_15136,N_12666,N_12142);
nand U15137 (N_15137,N_13102,N_13175);
nor U15138 (N_15138,N_13058,N_13923);
nand U15139 (N_15139,N_12276,N_13826);
or U15140 (N_15140,N_13465,N_13059);
nor U15141 (N_15141,N_12177,N_13789);
or U15142 (N_15142,N_12788,N_13512);
or U15143 (N_15143,N_13132,N_13700);
nor U15144 (N_15144,N_12791,N_13301);
nor U15145 (N_15145,N_13430,N_12274);
xor U15146 (N_15146,N_12422,N_13811);
xor U15147 (N_15147,N_12832,N_13909);
nand U15148 (N_15148,N_13803,N_12232);
nand U15149 (N_15149,N_13499,N_13727);
and U15150 (N_15150,N_12553,N_13938);
xnor U15151 (N_15151,N_13410,N_12356);
nor U15152 (N_15152,N_13755,N_13398);
nor U15153 (N_15153,N_12532,N_13762);
nor U15154 (N_15154,N_13632,N_12289);
or U15155 (N_15155,N_12224,N_13151);
nor U15156 (N_15156,N_12949,N_13406);
nand U15157 (N_15157,N_12410,N_13139);
or U15158 (N_15158,N_12495,N_13539);
xor U15159 (N_15159,N_12741,N_13129);
xnor U15160 (N_15160,N_13312,N_12734);
and U15161 (N_15161,N_12407,N_12612);
nor U15162 (N_15162,N_12512,N_13544);
or U15163 (N_15163,N_12460,N_13734);
xnor U15164 (N_15164,N_12121,N_13674);
xnor U15165 (N_15165,N_12960,N_12140);
and U15166 (N_15166,N_13091,N_12826);
nor U15167 (N_15167,N_12997,N_12541);
nand U15168 (N_15168,N_12141,N_12480);
and U15169 (N_15169,N_13705,N_13306);
nor U15170 (N_15170,N_13492,N_12331);
or U15171 (N_15171,N_13058,N_12657);
or U15172 (N_15172,N_13403,N_13658);
xor U15173 (N_15173,N_13196,N_12832);
xnor U15174 (N_15174,N_13542,N_13694);
nor U15175 (N_15175,N_12325,N_12763);
and U15176 (N_15176,N_13867,N_13625);
and U15177 (N_15177,N_13000,N_13580);
and U15178 (N_15178,N_12151,N_12322);
nor U15179 (N_15179,N_12272,N_12307);
and U15180 (N_15180,N_13554,N_12578);
xor U15181 (N_15181,N_12449,N_13312);
nor U15182 (N_15182,N_12703,N_13937);
or U15183 (N_15183,N_12042,N_12357);
xnor U15184 (N_15184,N_12695,N_12844);
xnor U15185 (N_15185,N_12865,N_13238);
nand U15186 (N_15186,N_13973,N_12672);
nand U15187 (N_15187,N_12429,N_12662);
or U15188 (N_15188,N_13248,N_12209);
or U15189 (N_15189,N_12210,N_12435);
and U15190 (N_15190,N_13851,N_13211);
nand U15191 (N_15191,N_13332,N_13684);
or U15192 (N_15192,N_12484,N_12881);
or U15193 (N_15193,N_13214,N_12533);
nor U15194 (N_15194,N_12375,N_12789);
xnor U15195 (N_15195,N_13806,N_13527);
nand U15196 (N_15196,N_12118,N_13494);
nand U15197 (N_15197,N_13303,N_13005);
nor U15198 (N_15198,N_13845,N_13954);
nor U15199 (N_15199,N_12477,N_12623);
xnor U15200 (N_15200,N_13075,N_13779);
nand U15201 (N_15201,N_13432,N_13716);
xor U15202 (N_15202,N_12341,N_12841);
nand U15203 (N_15203,N_13123,N_12758);
nor U15204 (N_15204,N_12638,N_12676);
nand U15205 (N_15205,N_13621,N_12189);
nor U15206 (N_15206,N_13405,N_13803);
nand U15207 (N_15207,N_12874,N_12715);
and U15208 (N_15208,N_13589,N_12058);
or U15209 (N_15209,N_12030,N_13276);
xnor U15210 (N_15210,N_13706,N_12308);
xnor U15211 (N_15211,N_12614,N_13414);
nor U15212 (N_15212,N_13680,N_12212);
xor U15213 (N_15213,N_12992,N_13030);
xnor U15214 (N_15214,N_13909,N_12418);
nand U15215 (N_15215,N_13336,N_13831);
or U15216 (N_15216,N_13315,N_13364);
nor U15217 (N_15217,N_13582,N_13182);
nor U15218 (N_15218,N_13776,N_12859);
nor U15219 (N_15219,N_12862,N_12442);
and U15220 (N_15220,N_13412,N_13396);
xor U15221 (N_15221,N_12263,N_12933);
and U15222 (N_15222,N_12124,N_12814);
nand U15223 (N_15223,N_13129,N_13773);
or U15224 (N_15224,N_12153,N_12840);
xnor U15225 (N_15225,N_12743,N_13931);
and U15226 (N_15226,N_12922,N_12957);
nand U15227 (N_15227,N_12162,N_12478);
and U15228 (N_15228,N_12905,N_12426);
nor U15229 (N_15229,N_13969,N_12937);
nor U15230 (N_15230,N_12890,N_13821);
xnor U15231 (N_15231,N_13713,N_12170);
and U15232 (N_15232,N_13871,N_12636);
nand U15233 (N_15233,N_12846,N_13600);
nor U15234 (N_15234,N_13138,N_12394);
or U15235 (N_15235,N_13490,N_13037);
nand U15236 (N_15236,N_12865,N_13990);
nand U15237 (N_15237,N_12923,N_12801);
xnor U15238 (N_15238,N_13398,N_12403);
and U15239 (N_15239,N_13322,N_12369);
nor U15240 (N_15240,N_13966,N_13589);
and U15241 (N_15241,N_12295,N_12691);
or U15242 (N_15242,N_12738,N_13881);
and U15243 (N_15243,N_12774,N_13298);
or U15244 (N_15244,N_13324,N_12939);
nor U15245 (N_15245,N_12764,N_13711);
nand U15246 (N_15246,N_12329,N_13915);
nand U15247 (N_15247,N_12159,N_13318);
nand U15248 (N_15248,N_13471,N_12727);
or U15249 (N_15249,N_12145,N_12627);
xnor U15250 (N_15250,N_12267,N_12675);
nor U15251 (N_15251,N_13906,N_12608);
or U15252 (N_15252,N_12669,N_12928);
nand U15253 (N_15253,N_13948,N_12846);
or U15254 (N_15254,N_13866,N_13220);
nand U15255 (N_15255,N_13379,N_12286);
nor U15256 (N_15256,N_13888,N_13296);
nor U15257 (N_15257,N_13147,N_12932);
and U15258 (N_15258,N_12503,N_13061);
or U15259 (N_15259,N_12457,N_12017);
and U15260 (N_15260,N_13621,N_13777);
nor U15261 (N_15261,N_13525,N_13324);
nand U15262 (N_15262,N_13978,N_13646);
xor U15263 (N_15263,N_13292,N_13068);
xnor U15264 (N_15264,N_12035,N_12707);
xor U15265 (N_15265,N_13925,N_12726);
nand U15266 (N_15266,N_12762,N_12681);
nand U15267 (N_15267,N_13154,N_13934);
or U15268 (N_15268,N_13408,N_13007);
nor U15269 (N_15269,N_13758,N_13440);
nand U15270 (N_15270,N_12467,N_12182);
or U15271 (N_15271,N_12127,N_12872);
or U15272 (N_15272,N_13930,N_13680);
xnor U15273 (N_15273,N_13109,N_12539);
nand U15274 (N_15274,N_13152,N_12464);
nand U15275 (N_15275,N_13755,N_12177);
nor U15276 (N_15276,N_13772,N_13721);
and U15277 (N_15277,N_13402,N_12322);
nor U15278 (N_15278,N_13858,N_13034);
nor U15279 (N_15279,N_13293,N_13662);
xor U15280 (N_15280,N_13203,N_13401);
nand U15281 (N_15281,N_13294,N_13412);
or U15282 (N_15282,N_12441,N_13231);
or U15283 (N_15283,N_12393,N_12664);
nand U15284 (N_15284,N_12396,N_12906);
and U15285 (N_15285,N_12937,N_12262);
xnor U15286 (N_15286,N_12297,N_13621);
nand U15287 (N_15287,N_12264,N_13157);
nor U15288 (N_15288,N_12733,N_13523);
nor U15289 (N_15289,N_12906,N_12117);
or U15290 (N_15290,N_13665,N_13015);
or U15291 (N_15291,N_12823,N_12011);
nor U15292 (N_15292,N_12387,N_13027);
or U15293 (N_15293,N_13809,N_13239);
xor U15294 (N_15294,N_12149,N_12493);
and U15295 (N_15295,N_13266,N_13008);
nand U15296 (N_15296,N_12328,N_13296);
and U15297 (N_15297,N_12583,N_13262);
or U15298 (N_15298,N_12441,N_12609);
xnor U15299 (N_15299,N_12176,N_13008);
nor U15300 (N_15300,N_13778,N_13178);
or U15301 (N_15301,N_13706,N_13767);
nor U15302 (N_15302,N_12046,N_13585);
nor U15303 (N_15303,N_13616,N_12847);
nor U15304 (N_15304,N_13170,N_12678);
nor U15305 (N_15305,N_12290,N_12096);
nand U15306 (N_15306,N_13464,N_13957);
and U15307 (N_15307,N_13037,N_13176);
or U15308 (N_15308,N_13840,N_12229);
and U15309 (N_15309,N_12386,N_13754);
xor U15310 (N_15310,N_13523,N_13748);
or U15311 (N_15311,N_12440,N_12436);
xor U15312 (N_15312,N_13688,N_13204);
and U15313 (N_15313,N_12822,N_13194);
nand U15314 (N_15314,N_13450,N_12174);
xnor U15315 (N_15315,N_12235,N_12059);
and U15316 (N_15316,N_13465,N_12334);
nor U15317 (N_15317,N_13045,N_13434);
nand U15318 (N_15318,N_13643,N_12887);
xor U15319 (N_15319,N_13568,N_13394);
nand U15320 (N_15320,N_12701,N_12360);
xor U15321 (N_15321,N_13253,N_12407);
or U15322 (N_15322,N_13120,N_12783);
nand U15323 (N_15323,N_13046,N_12711);
xor U15324 (N_15324,N_13969,N_13904);
nand U15325 (N_15325,N_13305,N_12605);
nor U15326 (N_15326,N_12981,N_13766);
and U15327 (N_15327,N_12295,N_12114);
or U15328 (N_15328,N_12953,N_13527);
nor U15329 (N_15329,N_13180,N_13289);
nor U15330 (N_15330,N_13766,N_13923);
and U15331 (N_15331,N_12172,N_13322);
or U15332 (N_15332,N_13098,N_13294);
nor U15333 (N_15333,N_13862,N_12440);
and U15334 (N_15334,N_12369,N_12791);
and U15335 (N_15335,N_12204,N_13009);
nor U15336 (N_15336,N_12345,N_12557);
or U15337 (N_15337,N_13167,N_13949);
and U15338 (N_15338,N_12173,N_12187);
and U15339 (N_15339,N_13690,N_13288);
nand U15340 (N_15340,N_12794,N_13569);
nor U15341 (N_15341,N_12163,N_13670);
or U15342 (N_15342,N_12616,N_12781);
nor U15343 (N_15343,N_13283,N_13850);
xor U15344 (N_15344,N_13786,N_13602);
xor U15345 (N_15345,N_13735,N_12398);
xor U15346 (N_15346,N_13486,N_12914);
xnor U15347 (N_15347,N_12209,N_13973);
nor U15348 (N_15348,N_12781,N_12632);
xor U15349 (N_15349,N_12726,N_13016);
or U15350 (N_15350,N_13335,N_13291);
or U15351 (N_15351,N_13783,N_13750);
and U15352 (N_15352,N_12683,N_12441);
or U15353 (N_15353,N_12908,N_12353);
nor U15354 (N_15354,N_13421,N_13174);
nand U15355 (N_15355,N_13528,N_13110);
or U15356 (N_15356,N_13088,N_13958);
xor U15357 (N_15357,N_13164,N_12709);
or U15358 (N_15358,N_12088,N_12876);
nand U15359 (N_15359,N_13638,N_12316);
and U15360 (N_15360,N_12059,N_12859);
nor U15361 (N_15361,N_13792,N_13906);
and U15362 (N_15362,N_12736,N_13281);
nor U15363 (N_15363,N_12143,N_13481);
and U15364 (N_15364,N_13436,N_12094);
nor U15365 (N_15365,N_12532,N_13737);
or U15366 (N_15366,N_13371,N_13309);
and U15367 (N_15367,N_13811,N_12237);
nor U15368 (N_15368,N_12378,N_13723);
xnor U15369 (N_15369,N_13087,N_13706);
nand U15370 (N_15370,N_12749,N_13871);
and U15371 (N_15371,N_12453,N_13905);
nand U15372 (N_15372,N_12065,N_13520);
nand U15373 (N_15373,N_12349,N_12357);
nand U15374 (N_15374,N_12427,N_12482);
and U15375 (N_15375,N_13375,N_13418);
nand U15376 (N_15376,N_12496,N_13557);
nor U15377 (N_15377,N_12450,N_13801);
xor U15378 (N_15378,N_12568,N_13673);
xor U15379 (N_15379,N_13761,N_12117);
nor U15380 (N_15380,N_12313,N_13337);
xnor U15381 (N_15381,N_12200,N_12831);
nand U15382 (N_15382,N_12872,N_12903);
nand U15383 (N_15383,N_13203,N_13746);
xnor U15384 (N_15384,N_12112,N_12988);
or U15385 (N_15385,N_13540,N_13779);
nand U15386 (N_15386,N_12882,N_13410);
or U15387 (N_15387,N_13667,N_13813);
and U15388 (N_15388,N_12760,N_12273);
or U15389 (N_15389,N_13368,N_13232);
or U15390 (N_15390,N_12041,N_13753);
or U15391 (N_15391,N_12549,N_13573);
nand U15392 (N_15392,N_12860,N_13150);
nand U15393 (N_15393,N_12176,N_12939);
nand U15394 (N_15394,N_12514,N_13330);
nand U15395 (N_15395,N_12952,N_13826);
nor U15396 (N_15396,N_13613,N_12207);
nor U15397 (N_15397,N_12152,N_13049);
or U15398 (N_15398,N_12095,N_13682);
xor U15399 (N_15399,N_13640,N_13642);
and U15400 (N_15400,N_13752,N_13061);
or U15401 (N_15401,N_13807,N_13787);
nand U15402 (N_15402,N_12868,N_12289);
nand U15403 (N_15403,N_13008,N_13313);
and U15404 (N_15404,N_12474,N_13793);
nor U15405 (N_15405,N_13543,N_12010);
and U15406 (N_15406,N_12183,N_13995);
or U15407 (N_15407,N_12466,N_13350);
nand U15408 (N_15408,N_13064,N_12526);
nor U15409 (N_15409,N_13408,N_13140);
or U15410 (N_15410,N_12884,N_12534);
and U15411 (N_15411,N_13154,N_12999);
nor U15412 (N_15412,N_13417,N_12677);
and U15413 (N_15413,N_12012,N_13998);
nand U15414 (N_15414,N_12993,N_12055);
nand U15415 (N_15415,N_12602,N_13819);
and U15416 (N_15416,N_12387,N_12051);
and U15417 (N_15417,N_12049,N_13135);
and U15418 (N_15418,N_13020,N_13712);
xor U15419 (N_15419,N_12212,N_13540);
nand U15420 (N_15420,N_13204,N_13332);
nand U15421 (N_15421,N_13831,N_12339);
or U15422 (N_15422,N_13694,N_13757);
nand U15423 (N_15423,N_13448,N_12097);
xnor U15424 (N_15424,N_12990,N_13736);
and U15425 (N_15425,N_12663,N_12350);
nor U15426 (N_15426,N_12464,N_13205);
nand U15427 (N_15427,N_12823,N_13067);
nand U15428 (N_15428,N_12510,N_12953);
nand U15429 (N_15429,N_12077,N_12985);
xor U15430 (N_15430,N_12794,N_12687);
nand U15431 (N_15431,N_13334,N_13623);
nand U15432 (N_15432,N_12322,N_13434);
xnor U15433 (N_15433,N_12654,N_13801);
xnor U15434 (N_15434,N_12125,N_12865);
xnor U15435 (N_15435,N_13701,N_13739);
or U15436 (N_15436,N_12483,N_13982);
or U15437 (N_15437,N_12264,N_12158);
nand U15438 (N_15438,N_12696,N_12473);
xor U15439 (N_15439,N_12133,N_12070);
nor U15440 (N_15440,N_13589,N_12721);
xnor U15441 (N_15441,N_13691,N_13172);
and U15442 (N_15442,N_13788,N_13434);
or U15443 (N_15443,N_12831,N_12451);
and U15444 (N_15444,N_12810,N_12101);
nor U15445 (N_15445,N_13489,N_12958);
or U15446 (N_15446,N_13072,N_12577);
xor U15447 (N_15447,N_13662,N_13363);
xnor U15448 (N_15448,N_13328,N_12601);
nand U15449 (N_15449,N_12102,N_12798);
nor U15450 (N_15450,N_12344,N_12310);
nand U15451 (N_15451,N_13972,N_12196);
or U15452 (N_15452,N_13404,N_12663);
or U15453 (N_15453,N_13526,N_12749);
or U15454 (N_15454,N_12039,N_12379);
and U15455 (N_15455,N_13337,N_12896);
and U15456 (N_15456,N_12902,N_12137);
nand U15457 (N_15457,N_13211,N_12765);
nor U15458 (N_15458,N_12287,N_13860);
and U15459 (N_15459,N_13511,N_12496);
nor U15460 (N_15460,N_12301,N_13750);
and U15461 (N_15461,N_12383,N_12743);
nor U15462 (N_15462,N_13902,N_12402);
and U15463 (N_15463,N_12915,N_12919);
xor U15464 (N_15464,N_13907,N_13353);
and U15465 (N_15465,N_13641,N_12833);
nor U15466 (N_15466,N_12866,N_13172);
or U15467 (N_15467,N_13226,N_13685);
or U15468 (N_15468,N_13995,N_12840);
nor U15469 (N_15469,N_13181,N_12379);
nor U15470 (N_15470,N_13807,N_12150);
nand U15471 (N_15471,N_12110,N_13521);
nor U15472 (N_15472,N_12484,N_13767);
and U15473 (N_15473,N_12048,N_12229);
and U15474 (N_15474,N_12272,N_13338);
nor U15475 (N_15475,N_12089,N_12146);
or U15476 (N_15476,N_13271,N_13246);
nand U15477 (N_15477,N_12018,N_12236);
and U15478 (N_15478,N_12920,N_13688);
or U15479 (N_15479,N_12875,N_12322);
or U15480 (N_15480,N_13478,N_13727);
or U15481 (N_15481,N_12692,N_13171);
xnor U15482 (N_15482,N_12520,N_13550);
or U15483 (N_15483,N_13911,N_13068);
xor U15484 (N_15484,N_13534,N_12483);
and U15485 (N_15485,N_12370,N_12375);
or U15486 (N_15486,N_12003,N_13987);
nor U15487 (N_15487,N_12502,N_13142);
xnor U15488 (N_15488,N_13194,N_12513);
and U15489 (N_15489,N_13174,N_12897);
nand U15490 (N_15490,N_12252,N_13653);
or U15491 (N_15491,N_12033,N_12876);
nand U15492 (N_15492,N_12461,N_12019);
and U15493 (N_15493,N_12540,N_13082);
nand U15494 (N_15494,N_13782,N_12634);
nor U15495 (N_15495,N_13268,N_13834);
xnor U15496 (N_15496,N_13362,N_13194);
or U15497 (N_15497,N_12102,N_13010);
and U15498 (N_15498,N_12656,N_12494);
or U15499 (N_15499,N_12050,N_12190);
xnor U15500 (N_15500,N_13668,N_13128);
and U15501 (N_15501,N_12170,N_12549);
and U15502 (N_15502,N_12044,N_13850);
nor U15503 (N_15503,N_12035,N_12452);
xor U15504 (N_15504,N_12940,N_12026);
or U15505 (N_15505,N_12327,N_12091);
xor U15506 (N_15506,N_13196,N_13539);
or U15507 (N_15507,N_13884,N_13358);
nand U15508 (N_15508,N_12565,N_13116);
nand U15509 (N_15509,N_12574,N_12997);
and U15510 (N_15510,N_13710,N_12280);
nor U15511 (N_15511,N_13816,N_12588);
xnor U15512 (N_15512,N_13632,N_12531);
nor U15513 (N_15513,N_12858,N_12690);
xor U15514 (N_15514,N_12888,N_12390);
nor U15515 (N_15515,N_13716,N_12153);
nor U15516 (N_15516,N_12124,N_12388);
nor U15517 (N_15517,N_13083,N_12033);
xnor U15518 (N_15518,N_12325,N_13143);
nand U15519 (N_15519,N_12156,N_12939);
xor U15520 (N_15520,N_13429,N_12759);
nand U15521 (N_15521,N_12004,N_12119);
or U15522 (N_15522,N_13933,N_12325);
and U15523 (N_15523,N_13619,N_12128);
xnor U15524 (N_15524,N_12522,N_13678);
or U15525 (N_15525,N_13965,N_12253);
xnor U15526 (N_15526,N_12750,N_12122);
xnor U15527 (N_15527,N_12983,N_13846);
xor U15528 (N_15528,N_13955,N_12237);
xor U15529 (N_15529,N_12895,N_13898);
and U15530 (N_15530,N_12188,N_12580);
or U15531 (N_15531,N_12736,N_13539);
nand U15532 (N_15532,N_12082,N_13792);
or U15533 (N_15533,N_13093,N_12269);
nor U15534 (N_15534,N_12343,N_12287);
xnor U15535 (N_15535,N_13954,N_12422);
xor U15536 (N_15536,N_13925,N_12517);
or U15537 (N_15537,N_12188,N_13391);
xor U15538 (N_15538,N_13121,N_13076);
nand U15539 (N_15539,N_13774,N_13056);
xor U15540 (N_15540,N_13736,N_13907);
nand U15541 (N_15541,N_13239,N_12387);
nor U15542 (N_15542,N_13245,N_12099);
or U15543 (N_15543,N_13256,N_12608);
and U15544 (N_15544,N_12597,N_12488);
xor U15545 (N_15545,N_13048,N_12447);
nor U15546 (N_15546,N_12270,N_13091);
xnor U15547 (N_15547,N_13755,N_13536);
or U15548 (N_15548,N_13084,N_12655);
nor U15549 (N_15549,N_12645,N_12532);
nand U15550 (N_15550,N_12782,N_13445);
nand U15551 (N_15551,N_12525,N_13038);
and U15552 (N_15552,N_13779,N_13486);
and U15553 (N_15553,N_13114,N_12497);
nand U15554 (N_15554,N_13219,N_12980);
or U15555 (N_15555,N_13381,N_12041);
or U15556 (N_15556,N_13496,N_13282);
nor U15557 (N_15557,N_12885,N_13428);
or U15558 (N_15558,N_13719,N_13731);
or U15559 (N_15559,N_12561,N_13199);
and U15560 (N_15560,N_13165,N_13492);
and U15561 (N_15561,N_13550,N_13303);
xor U15562 (N_15562,N_12246,N_12705);
xnor U15563 (N_15563,N_13075,N_12482);
or U15564 (N_15564,N_12922,N_13488);
xnor U15565 (N_15565,N_12096,N_13022);
and U15566 (N_15566,N_12100,N_12392);
or U15567 (N_15567,N_13582,N_13258);
xor U15568 (N_15568,N_13022,N_12345);
xnor U15569 (N_15569,N_13785,N_13533);
nand U15570 (N_15570,N_12505,N_13188);
nor U15571 (N_15571,N_12799,N_13970);
xnor U15572 (N_15572,N_12108,N_13284);
xor U15573 (N_15573,N_13864,N_12573);
or U15574 (N_15574,N_13324,N_12409);
nor U15575 (N_15575,N_13197,N_13802);
and U15576 (N_15576,N_12687,N_13212);
nand U15577 (N_15577,N_12266,N_13943);
nor U15578 (N_15578,N_12087,N_13639);
nand U15579 (N_15579,N_12977,N_12426);
nor U15580 (N_15580,N_13119,N_12071);
and U15581 (N_15581,N_12693,N_12383);
or U15582 (N_15582,N_13706,N_13664);
nand U15583 (N_15583,N_13553,N_12377);
nand U15584 (N_15584,N_13199,N_13184);
and U15585 (N_15585,N_13073,N_12192);
nand U15586 (N_15586,N_13909,N_13330);
or U15587 (N_15587,N_12543,N_12100);
and U15588 (N_15588,N_12890,N_12881);
nor U15589 (N_15589,N_12794,N_12836);
nor U15590 (N_15590,N_13097,N_12540);
nand U15591 (N_15591,N_12089,N_13155);
nand U15592 (N_15592,N_13226,N_12048);
and U15593 (N_15593,N_12008,N_13759);
or U15594 (N_15594,N_12355,N_13795);
nor U15595 (N_15595,N_12422,N_12806);
nor U15596 (N_15596,N_13654,N_12484);
nor U15597 (N_15597,N_13274,N_13311);
and U15598 (N_15598,N_12641,N_13156);
nand U15599 (N_15599,N_13135,N_12497);
and U15600 (N_15600,N_13056,N_13213);
or U15601 (N_15601,N_13318,N_12615);
nor U15602 (N_15602,N_13351,N_13762);
and U15603 (N_15603,N_13177,N_12254);
nand U15604 (N_15604,N_12196,N_13988);
and U15605 (N_15605,N_12895,N_13501);
nand U15606 (N_15606,N_12702,N_12202);
xnor U15607 (N_15607,N_13662,N_13777);
nor U15608 (N_15608,N_13290,N_13272);
nor U15609 (N_15609,N_12454,N_12079);
xnor U15610 (N_15610,N_12605,N_13620);
and U15611 (N_15611,N_13815,N_12692);
and U15612 (N_15612,N_12262,N_13807);
or U15613 (N_15613,N_12004,N_13241);
or U15614 (N_15614,N_13052,N_13891);
nor U15615 (N_15615,N_13337,N_12253);
and U15616 (N_15616,N_13666,N_13820);
xnor U15617 (N_15617,N_12871,N_12355);
or U15618 (N_15618,N_12745,N_12969);
and U15619 (N_15619,N_13465,N_12377);
nand U15620 (N_15620,N_13035,N_13515);
or U15621 (N_15621,N_12540,N_13707);
nand U15622 (N_15622,N_13072,N_12859);
nor U15623 (N_15623,N_13615,N_13208);
nor U15624 (N_15624,N_13799,N_12743);
or U15625 (N_15625,N_13744,N_13690);
xnor U15626 (N_15626,N_12700,N_13083);
nor U15627 (N_15627,N_13348,N_12138);
nand U15628 (N_15628,N_13621,N_13235);
nor U15629 (N_15629,N_12846,N_12415);
or U15630 (N_15630,N_13772,N_12776);
or U15631 (N_15631,N_12228,N_12494);
nor U15632 (N_15632,N_12805,N_13589);
nand U15633 (N_15633,N_13965,N_12194);
nor U15634 (N_15634,N_13537,N_12277);
and U15635 (N_15635,N_12040,N_12574);
and U15636 (N_15636,N_13423,N_13092);
nand U15637 (N_15637,N_13159,N_13888);
nand U15638 (N_15638,N_12943,N_13528);
nor U15639 (N_15639,N_13493,N_12336);
nor U15640 (N_15640,N_12911,N_13274);
nor U15641 (N_15641,N_13476,N_12671);
or U15642 (N_15642,N_12701,N_12720);
and U15643 (N_15643,N_13124,N_12330);
xor U15644 (N_15644,N_13190,N_12960);
xnor U15645 (N_15645,N_13803,N_13825);
or U15646 (N_15646,N_12077,N_13846);
nand U15647 (N_15647,N_12308,N_12904);
xnor U15648 (N_15648,N_12987,N_12268);
nor U15649 (N_15649,N_12275,N_12922);
nor U15650 (N_15650,N_12976,N_13728);
nand U15651 (N_15651,N_13025,N_13069);
nand U15652 (N_15652,N_12272,N_12932);
and U15653 (N_15653,N_12249,N_13204);
nand U15654 (N_15654,N_12295,N_13137);
xnor U15655 (N_15655,N_12879,N_12009);
xor U15656 (N_15656,N_12477,N_12306);
xor U15657 (N_15657,N_13498,N_13839);
or U15658 (N_15658,N_13708,N_13353);
and U15659 (N_15659,N_12271,N_12412);
and U15660 (N_15660,N_13314,N_13970);
or U15661 (N_15661,N_13992,N_13527);
and U15662 (N_15662,N_12248,N_12377);
xnor U15663 (N_15663,N_12267,N_13573);
or U15664 (N_15664,N_13961,N_13774);
nor U15665 (N_15665,N_12863,N_13167);
and U15666 (N_15666,N_12849,N_13378);
nor U15667 (N_15667,N_12944,N_12369);
xnor U15668 (N_15668,N_13784,N_12419);
xor U15669 (N_15669,N_13688,N_13736);
nand U15670 (N_15670,N_13773,N_12261);
or U15671 (N_15671,N_13903,N_12728);
or U15672 (N_15672,N_12249,N_13556);
and U15673 (N_15673,N_12285,N_13698);
xnor U15674 (N_15674,N_12015,N_13208);
nand U15675 (N_15675,N_12257,N_13788);
nand U15676 (N_15676,N_13073,N_13304);
and U15677 (N_15677,N_13707,N_12920);
and U15678 (N_15678,N_12565,N_12654);
nor U15679 (N_15679,N_12046,N_12029);
xnor U15680 (N_15680,N_13829,N_13503);
nand U15681 (N_15681,N_12416,N_12577);
nand U15682 (N_15682,N_13829,N_12751);
nand U15683 (N_15683,N_12587,N_12729);
and U15684 (N_15684,N_12690,N_12450);
and U15685 (N_15685,N_13649,N_12083);
or U15686 (N_15686,N_13752,N_12249);
or U15687 (N_15687,N_12971,N_13398);
or U15688 (N_15688,N_13074,N_13637);
nor U15689 (N_15689,N_12332,N_13827);
xnor U15690 (N_15690,N_12255,N_12908);
nor U15691 (N_15691,N_13391,N_13344);
or U15692 (N_15692,N_12039,N_12106);
nor U15693 (N_15693,N_13689,N_12035);
or U15694 (N_15694,N_12361,N_13712);
or U15695 (N_15695,N_12058,N_12996);
nand U15696 (N_15696,N_12371,N_13267);
nor U15697 (N_15697,N_13932,N_12479);
nand U15698 (N_15698,N_13815,N_12103);
and U15699 (N_15699,N_13167,N_13124);
nand U15700 (N_15700,N_12427,N_12654);
and U15701 (N_15701,N_13655,N_13976);
and U15702 (N_15702,N_12281,N_12243);
or U15703 (N_15703,N_13587,N_13554);
xnor U15704 (N_15704,N_13648,N_13666);
nand U15705 (N_15705,N_13066,N_12604);
and U15706 (N_15706,N_12862,N_13421);
xor U15707 (N_15707,N_13190,N_13364);
or U15708 (N_15708,N_13255,N_12968);
and U15709 (N_15709,N_12431,N_12129);
xor U15710 (N_15710,N_13622,N_12389);
nand U15711 (N_15711,N_13164,N_13210);
and U15712 (N_15712,N_13682,N_13864);
and U15713 (N_15713,N_12992,N_12607);
and U15714 (N_15714,N_12453,N_13785);
and U15715 (N_15715,N_12184,N_13021);
nor U15716 (N_15716,N_13754,N_12963);
nand U15717 (N_15717,N_13237,N_12656);
and U15718 (N_15718,N_12448,N_13239);
and U15719 (N_15719,N_13718,N_12302);
nor U15720 (N_15720,N_12480,N_12700);
xnor U15721 (N_15721,N_12996,N_13967);
nand U15722 (N_15722,N_12257,N_13879);
and U15723 (N_15723,N_13286,N_13841);
nand U15724 (N_15724,N_13953,N_12574);
nand U15725 (N_15725,N_12698,N_12801);
xnor U15726 (N_15726,N_12431,N_12754);
or U15727 (N_15727,N_12062,N_12743);
nand U15728 (N_15728,N_12549,N_13731);
nand U15729 (N_15729,N_13770,N_12321);
xor U15730 (N_15730,N_13126,N_12467);
nor U15731 (N_15731,N_12178,N_13132);
and U15732 (N_15732,N_12613,N_12377);
xnor U15733 (N_15733,N_12912,N_12759);
or U15734 (N_15734,N_12053,N_13708);
or U15735 (N_15735,N_13107,N_13773);
and U15736 (N_15736,N_13783,N_13743);
and U15737 (N_15737,N_13583,N_13245);
nand U15738 (N_15738,N_12235,N_13352);
or U15739 (N_15739,N_13860,N_12054);
nor U15740 (N_15740,N_13863,N_12587);
xnor U15741 (N_15741,N_13475,N_13793);
nor U15742 (N_15742,N_12386,N_12893);
nand U15743 (N_15743,N_13670,N_13258);
xor U15744 (N_15744,N_13366,N_12988);
or U15745 (N_15745,N_13072,N_13244);
or U15746 (N_15746,N_12330,N_13755);
or U15747 (N_15747,N_12252,N_13579);
nor U15748 (N_15748,N_12598,N_12456);
nor U15749 (N_15749,N_13362,N_12931);
or U15750 (N_15750,N_13470,N_12856);
nand U15751 (N_15751,N_13538,N_13707);
nor U15752 (N_15752,N_12740,N_12158);
or U15753 (N_15753,N_12561,N_12184);
and U15754 (N_15754,N_13598,N_12616);
xnor U15755 (N_15755,N_12731,N_13677);
nand U15756 (N_15756,N_13232,N_12659);
nor U15757 (N_15757,N_12854,N_13782);
and U15758 (N_15758,N_13288,N_13992);
and U15759 (N_15759,N_13236,N_12546);
nand U15760 (N_15760,N_12993,N_12639);
and U15761 (N_15761,N_13713,N_13993);
nand U15762 (N_15762,N_13039,N_12059);
and U15763 (N_15763,N_12035,N_12465);
or U15764 (N_15764,N_12488,N_12089);
and U15765 (N_15765,N_12862,N_13510);
nor U15766 (N_15766,N_12279,N_12684);
and U15767 (N_15767,N_13851,N_12313);
and U15768 (N_15768,N_12245,N_12916);
xnor U15769 (N_15769,N_13141,N_13820);
nand U15770 (N_15770,N_13901,N_13326);
and U15771 (N_15771,N_13890,N_12159);
nand U15772 (N_15772,N_13889,N_13655);
nor U15773 (N_15773,N_12406,N_12587);
or U15774 (N_15774,N_13680,N_13263);
and U15775 (N_15775,N_13783,N_13810);
nand U15776 (N_15776,N_12372,N_13464);
and U15777 (N_15777,N_13299,N_12943);
nor U15778 (N_15778,N_12172,N_13538);
nand U15779 (N_15779,N_12989,N_12354);
nand U15780 (N_15780,N_12138,N_13779);
nand U15781 (N_15781,N_12768,N_12757);
or U15782 (N_15782,N_13660,N_12244);
nand U15783 (N_15783,N_13026,N_12670);
xor U15784 (N_15784,N_12548,N_12579);
nor U15785 (N_15785,N_12351,N_13488);
or U15786 (N_15786,N_12526,N_12470);
nor U15787 (N_15787,N_12947,N_13594);
xor U15788 (N_15788,N_13714,N_12439);
xnor U15789 (N_15789,N_12513,N_12746);
or U15790 (N_15790,N_12242,N_13636);
nor U15791 (N_15791,N_13781,N_13315);
or U15792 (N_15792,N_13785,N_12708);
xnor U15793 (N_15793,N_13502,N_12886);
or U15794 (N_15794,N_12905,N_12354);
xor U15795 (N_15795,N_13562,N_13483);
nor U15796 (N_15796,N_12294,N_13015);
nand U15797 (N_15797,N_13060,N_13427);
xnor U15798 (N_15798,N_12484,N_12047);
nand U15799 (N_15799,N_13782,N_13322);
xnor U15800 (N_15800,N_13407,N_13468);
nand U15801 (N_15801,N_12062,N_12936);
xnor U15802 (N_15802,N_13164,N_13285);
xor U15803 (N_15803,N_12731,N_13997);
nor U15804 (N_15804,N_13699,N_12105);
nand U15805 (N_15805,N_12696,N_13880);
xor U15806 (N_15806,N_13388,N_13328);
or U15807 (N_15807,N_12517,N_13353);
and U15808 (N_15808,N_12299,N_13563);
or U15809 (N_15809,N_13580,N_13708);
nand U15810 (N_15810,N_13320,N_12352);
nor U15811 (N_15811,N_12429,N_12610);
nor U15812 (N_15812,N_13660,N_13805);
or U15813 (N_15813,N_13186,N_13436);
nor U15814 (N_15814,N_12934,N_12043);
or U15815 (N_15815,N_13564,N_12086);
nor U15816 (N_15816,N_13519,N_13104);
or U15817 (N_15817,N_13524,N_13079);
nand U15818 (N_15818,N_13057,N_12509);
xor U15819 (N_15819,N_12010,N_12661);
xor U15820 (N_15820,N_13976,N_12033);
nor U15821 (N_15821,N_12261,N_13808);
xnor U15822 (N_15822,N_13620,N_12129);
or U15823 (N_15823,N_13852,N_13460);
xnor U15824 (N_15824,N_12610,N_13885);
xnor U15825 (N_15825,N_13983,N_12055);
nand U15826 (N_15826,N_12439,N_13370);
xnor U15827 (N_15827,N_12903,N_13538);
and U15828 (N_15828,N_13561,N_12271);
nor U15829 (N_15829,N_13984,N_13531);
and U15830 (N_15830,N_12105,N_13243);
or U15831 (N_15831,N_12300,N_12474);
nor U15832 (N_15832,N_13119,N_12094);
nor U15833 (N_15833,N_13873,N_12994);
nand U15834 (N_15834,N_13538,N_13850);
or U15835 (N_15835,N_12925,N_12313);
and U15836 (N_15836,N_13522,N_13392);
xor U15837 (N_15837,N_12515,N_13175);
or U15838 (N_15838,N_12153,N_13417);
or U15839 (N_15839,N_13585,N_12403);
nand U15840 (N_15840,N_12190,N_12002);
nor U15841 (N_15841,N_12584,N_12653);
or U15842 (N_15842,N_12305,N_12294);
xor U15843 (N_15843,N_12909,N_12256);
nor U15844 (N_15844,N_13828,N_13300);
or U15845 (N_15845,N_13370,N_13142);
nor U15846 (N_15846,N_13189,N_12341);
nand U15847 (N_15847,N_13334,N_12171);
nand U15848 (N_15848,N_12512,N_12234);
and U15849 (N_15849,N_12891,N_13669);
xnor U15850 (N_15850,N_12345,N_12839);
nor U15851 (N_15851,N_13259,N_13768);
nand U15852 (N_15852,N_12870,N_13218);
nand U15853 (N_15853,N_12041,N_12298);
nor U15854 (N_15854,N_13487,N_12091);
nor U15855 (N_15855,N_13462,N_12127);
or U15856 (N_15856,N_13946,N_12131);
xnor U15857 (N_15857,N_13630,N_13075);
or U15858 (N_15858,N_13054,N_12884);
or U15859 (N_15859,N_12896,N_13870);
xnor U15860 (N_15860,N_12510,N_12838);
and U15861 (N_15861,N_12123,N_13451);
nor U15862 (N_15862,N_13058,N_12158);
xnor U15863 (N_15863,N_12754,N_12245);
or U15864 (N_15864,N_12029,N_13364);
xor U15865 (N_15865,N_13612,N_13092);
nor U15866 (N_15866,N_12022,N_12335);
or U15867 (N_15867,N_12012,N_13028);
nor U15868 (N_15868,N_12165,N_13406);
and U15869 (N_15869,N_12473,N_13777);
xnor U15870 (N_15870,N_13464,N_12479);
nand U15871 (N_15871,N_12884,N_12810);
or U15872 (N_15872,N_12178,N_13972);
or U15873 (N_15873,N_12351,N_12055);
or U15874 (N_15874,N_12299,N_13320);
and U15875 (N_15875,N_13391,N_13743);
or U15876 (N_15876,N_12368,N_13779);
xnor U15877 (N_15877,N_12652,N_12559);
nor U15878 (N_15878,N_13828,N_13284);
and U15879 (N_15879,N_12650,N_13757);
nand U15880 (N_15880,N_12919,N_13893);
nand U15881 (N_15881,N_13648,N_12922);
or U15882 (N_15882,N_12214,N_13083);
or U15883 (N_15883,N_13838,N_13171);
nor U15884 (N_15884,N_13249,N_13911);
or U15885 (N_15885,N_13499,N_12569);
nor U15886 (N_15886,N_12837,N_13995);
xnor U15887 (N_15887,N_12511,N_13547);
xor U15888 (N_15888,N_12494,N_12790);
nand U15889 (N_15889,N_12417,N_13933);
or U15890 (N_15890,N_12237,N_13611);
xnor U15891 (N_15891,N_12451,N_12941);
or U15892 (N_15892,N_12043,N_12029);
nand U15893 (N_15893,N_13100,N_13482);
nand U15894 (N_15894,N_12360,N_13178);
or U15895 (N_15895,N_13206,N_13234);
or U15896 (N_15896,N_12823,N_13758);
nand U15897 (N_15897,N_12415,N_12618);
xor U15898 (N_15898,N_13889,N_13139);
nor U15899 (N_15899,N_12406,N_13633);
and U15900 (N_15900,N_13668,N_13617);
and U15901 (N_15901,N_13126,N_13328);
nor U15902 (N_15902,N_12893,N_13051);
nor U15903 (N_15903,N_12992,N_12761);
and U15904 (N_15904,N_13240,N_12667);
nand U15905 (N_15905,N_13362,N_12605);
nand U15906 (N_15906,N_13678,N_13172);
nand U15907 (N_15907,N_12210,N_12544);
nand U15908 (N_15908,N_13136,N_13209);
or U15909 (N_15909,N_13495,N_12083);
xor U15910 (N_15910,N_12616,N_13257);
or U15911 (N_15911,N_12841,N_13914);
nand U15912 (N_15912,N_12469,N_13693);
and U15913 (N_15913,N_12896,N_12616);
or U15914 (N_15914,N_12321,N_13678);
nand U15915 (N_15915,N_12103,N_12058);
and U15916 (N_15916,N_12426,N_12661);
nor U15917 (N_15917,N_13679,N_13031);
or U15918 (N_15918,N_12190,N_13481);
or U15919 (N_15919,N_12243,N_13773);
nand U15920 (N_15920,N_13196,N_12314);
or U15921 (N_15921,N_12741,N_12298);
xor U15922 (N_15922,N_12516,N_13828);
and U15923 (N_15923,N_12349,N_12219);
and U15924 (N_15924,N_13106,N_12938);
nor U15925 (N_15925,N_13603,N_12334);
and U15926 (N_15926,N_12253,N_12061);
or U15927 (N_15927,N_12614,N_13728);
nor U15928 (N_15928,N_13874,N_13572);
or U15929 (N_15929,N_13858,N_12856);
nor U15930 (N_15930,N_12327,N_12545);
and U15931 (N_15931,N_13767,N_12621);
xnor U15932 (N_15932,N_13425,N_12949);
nand U15933 (N_15933,N_13385,N_13651);
nand U15934 (N_15934,N_12253,N_12071);
or U15935 (N_15935,N_12128,N_12648);
nor U15936 (N_15936,N_12941,N_13372);
and U15937 (N_15937,N_13783,N_12059);
xor U15938 (N_15938,N_13392,N_12814);
nand U15939 (N_15939,N_13854,N_12491);
or U15940 (N_15940,N_13393,N_13863);
and U15941 (N_15941,N_12810,N_12527);
and U15942 (N_15942,N_12291,N_12825);
nor U15943 (N_15943,N_12170,N_12999);
xnor U15944 (N_15944,N_13075,N_12452);
nor U15945 (N_15945,N_12636,N_12311);
nor U15946 (N_15946,N_12603,N_13336);
nand U15947 (N_15947,N_12866,N_12610);
xnor U15948 (N_15948,N_13275,N_13570);
xnor U15949 (N_15949,N_13755,N_13674);
nand U15950 (N_15950,N_13863,N_13573);
nand U15951 (N_15951,N_12678,N_13940);
nor U15952 (N_15952,N_13534,N_13715);
nor U15953 (N_15953,N_12277,N_13005);
and U15954 (N_15954,N_12077,N_12598);
nor U15955 (N_15955,N_13296,N_12041);
xnor U15956 (N_15956,N_13322,N_13763);
xnor U15957 (N_15957,N_13603,N_12370);
xor U15958 (N_15958,N_12301,N_12736);
xnor U15959 (N_15959,N_12323,N_13940);
and U15960 (N_15960,N_13375,N_12637);
nor U15961 (N_15961,N_12024,N_12903);
and U15962 (N_15962,N_13388,N_12478);
xor U15963 (N_15963,N_12514,N_12218);
nor U15964 (N_15964,N_13372,N_13368);
nor U15965 (N_15965,N_13262,N_13571);
and U15966 (N_15966,N_13788,N_12972);
or U15967 (N_15967,N_12110,N_12453);
and U15968 (N_15968,N_13429,N_13015);
or U15969 (N_15969,N_13109,N_13263);
nor U15970 (N_15970,N_13185,N_13481);
or U15971 (N_15971,N_13160,N_12037);
nor U15972 (N_15972,N_13819,N_12141);
or U15973 (N_15973,N_13195,N_13928);
and U15974 (N_15974,N_12444,N_12784);
xnor U15975 (N_15975,N_13353,N_13358);
xnor U15976 (N_15976,N_13705,N_13668);
and U15977 (N_15977,N_12260,N_12693);
nand U15978 (N_15978,N_13081,N_12835);
or U15979 (N_15979,N_12252,N_12292);
xor U15980 (N_15980,N_12077,N_13509);
xor U15981 (N_15981,N_12191,N_13685);
or U15982 (N_15982,N_12605,N_13060);
or U15983 (N_15983,N_12248,N_13753);
nand U15984 (N_15984,N_13711,N_13077);
and U15985 (N_15985,N_13728,N_12601);
xnor U15986 (N_15986,N_12217,N_12848);
nand U15987 (N_15987,N_13730,N_12247);
nor U15988 (N_15988,N_12184,N_12587);
nor U15989 (N_15989,N_13510,N_13804);
nand U15990 (N_15990,N_12537,N_13863);
xnor U15991 (N_15991,N_12097,N_13081);
or U15992 (N_15992,N_13586,N_12969);
nand U15993 (N_15993,N_12133,N_13547);
nand U15994 (N_15994,N_12187,N_13473);
xnor U15995 (N_15995,N_13733,N_13608);
xnor U15996 (N_15996,N_13684,N_12703);
nand U15997 (N_15997,N_12982,N_12581);
or U15998 (N_15998,N_13986,N_12522);
or U15999 (N_15999,N_12921,N_13220);
xor U16000 (N_16000,N_14808,N_14400);
and U16001 (N_16001,N_14435,N_14510);
and U16002 (N_16002,N_15482,N_14950);
and U16003 (N_16003,N_15293,N_14816);
nand U16004 (N_16004,N_14080,N_14234);
nor U16005 (N_16005,N_14429,N_14191);
nand U16006 (N_16006,N_14927,N_15302);
xnor U16007 (N_16007,N_14056,N_14701);
nand U16008 (N_16008,N_14509,N_14875);
or U16009 (N_16009,N_14320,N_15474);
nand U16010 (N_16010,N_14856,N_14733);
or U16011 (N_16011,N_15696,N_15841);
or U16012 (N_16012,N_14795,N_15211);
and U16013 (N_16013,N_14087,N_15421);
nand U16014 (N_16014,N_14477,N_14712);
xor U16015 (N_16015,N_14592,N_14200);
xor U16016 (N_16016,N_14884,N_15689);
nor U16017 (N_16017,N_15511,N_14189);
and U16018 (N_16018,N_15990,N_15709);
and U16019 (N_16019,N_15833,N_15669);
xnor U16020 (N_16020,N_14730,N_14158);
or U16021 (N_16021,N_14077,N_15250);
nand U16022 (N_16022,N_15783,N_14467);
xor U16023 (N_16023,N_14354,N_15395);
xor U16024 (N_16024,N_14912,N_15255);
or U16025 (N_16025,N_15745,N_14182);
nand U16026 (N_16026,N_14292,N_14492);
and U16027 (N_16027,N_14232,N_14880);
and U16028 (N_16028,N_15595,N_15240);
or U16029 (N_16029,N_14934,N_15080);
nand U16030 (N_16030,N_15367,N_14811);
xnor U16031 (N_16031,N_14657,N_14564);
xnor U16032 (N_16032,N_14129,N_15777);
xor U16033 (N_16033,N_14997,N_14122);
xnor U16034 (N_16034,N_15468,N_15277);
xnor U16035 (N_16035,N_14538,N_14800);
xor U16036 (N_16036,N_14228,N_15016);
nor U16037 (N_16037,N_14041,N_14965);
or U16038 (N_16038,N_15519,N_15134);
xor U16039 (N_16039,N_14656,N_15963);
xnor U16040 (N_16040,N_15611,N_14897);
nor U16041 (N_16041,N_15038,N_15345);
nand U16042 (N_16042,N_14604,N_15284);
nor U16043 (N_16043,N_15007,N_15744);
nor U16044 (N_16044,N_15937,N_14665);
xnor U16045 (N_16045,N_15388,N_15641);
nand U16046 (N_16046,N_15713,N_15300);
or U16047 (N_16047,N_15800,N_14854);
nor U16048 (N_16048,N_14088,N_14379);
nand U16049 (N_16049,N_15181,N_15525);
or U16050 (N_16050,N_14583,N_14031);
or U16051 (N_16051,N_15440,N_14172);
nand U16052 (N_16052,N_15898,N_15050);
nor U16053 (N_16053,N_14209,N_15993);
nand U16054 (N_16054,N_14611,N_15287);
or U16055 (N_16055,N_14334,N_14100);
or U16056 (N_16056,N_15735,N_14150);
xnor U16057 (N_16057,N_14210,N_15798);
nor U16058 (N_16058,N_15625,N_14735);
xor U16059 (N_16059,N_15122,N_15037);
xnor U16060 (N_16060,N_14242,N_15591);
nor U16061 (N_16061,N_15148,N_15527);
xnor U16062 (N_16062,N_14837,N_15810);
and U16063 (N_16063,N_15672,N_14801);
and U16064 (N_16064,N_15149,N_14416);
xnor U16065 (N_16065,N_14393,N_15711);
xnor U16066 (N_16066,N_15093,N_15597);
nor U16067 (N_16067,N_15695,N_15258);
or U16068 (N_16068,N_15054,N_15479);
xnor U16069 (N_16069,N_15423,N_14859);
xor U16070 (N_16070,N_14574,N_15045);
nand U16071 (N_16071,N_15478,N_15807);
xor U16072 (N_16072,N_15512,N_15867);
xor U16073 (N_16073,N_14799,N_14165);
and U16074 (N_16074,N_15307,N_15021);
or U16075 (N_16075,N_14957,N_15852);
or U16076 (N_16076,N_15580,N_14109);
and U16077 (N_16077,N_15064,N_14307);
xnor U16078 (N_16078,N_14970,N_15473);
xnor U16079 (N_16079,N_15958,N_15766);
and U16080 (N_16080,N_14024,N_14969);
xnor U16081 (N_16081,N_14407,N_15815);
nand U16082 (N_16082,N_15506,N_15418);
or U16083 (N_16083,N_14546,N_14527);
nor U16084 (N_16084,N_14148,N_14296);
and U16085 (N_16085,N_14152,N_15427);
or U16086 (N_16086,N_14272,N_15630);
or U16087 (N_16087,N_15504,N_15118);
nand U16088 (N_16088,N_14915,N_15325);
xor U16089 (N_16089,N_14177,N_14882);
and U16090 (N_16090,N_15521,N_15509);
or U16091 (N_16091,N_14782,N_15005);
and U16092 (N_16092,N_14474,N_15551);
and U16093 (N_16093,N_15820,N_14520);
nand U16094 (N_16094,N_14459,N_14271);
or U16095 (N_16095,N_14147,N_14605);
xor U16096 (N_16096,N_15688,N_15916);
nand U16097 (N_16097,N_15896,N_14411);
nor U16098 (N_16098,N_15376,N_15762);
nand U16099 (N_16099,N_14131,N_15004);
and U16100 (N_16100,N_14620,N_15901);
nand U16101 (N_16101,N_14914,N_14140);
nor U16102 (N_16102,N_15319,N_15951);
and U16103 (N_16103,N_14976,N_15053);
and U16104 (N_16104,N_15674,N_14352);
xnor U16105 (N_16105,N_14174,N_14116);
xor U16106 (N_16106,N_15646,N_15985);
xnor U16107 (N_16107,N_14486,N_15905);
nor U16108 (N_16108,N_15095,N_15515);
and U16109 (N_16109,N_14787,N_15514);
and U16110 (N_16110,N_14984,N_15448);
nand U16111 (N_16111,N_14101,N_15880);
xor U16112 (N_16112,N_14476,N_14562);
nand U16113 (N_16113,N_14221,N_14500);
nor U16114 (N_16114,N_14096,N_15529);
nand U16115 (N_16115,N_14702,N_15466);
xnor U16116 (N_16116,N_15772,N_15444);
nand U16117 (N_16117,N_14589,N_14578);
nor U16118 (N_16118,N_15326,N_14504);
nand U16119 (N_16119,N_14081,N_14834);
nor U16120 (N_16120,N_15330,N_15247);
xor U16121 (N_16121,N_14619,N_14185);
and U16122 (N_16122,N_14236,N_14855);
and U16123 (N_16123,N_14378,N_15677);
and U16124 (N_16124,N_15913,N_14905);
and U16125 (N_16125,N_15650,N_14333);
or U16126 (N_16126,N_14532,N_14765);
nor U16127 (N_16127,N_15806,N_15861);
or U16128 (N_16128,N_15865,N_15670);
xor U16129 (N_16129,N_15019,N_14365);
xor U16130 (N_16130,N_14805,N_15671);
or U16131 (N_16131,N_15727,N_15855);
and U16132 (N_16132,N_14732,N_14641);
nand U16133 (N_16133,N_15169,N_15673);
nor U16134 (N_16134,N_15567,N_15006);
and U16135 (N_16135,N_15930,N_15223);
xnor U16136 (N_16136,N_14327,N_14910);
nand U16137 (N_16137,N_14368,N_14469);
or U16138 (N_16138,N_15792,N_15785);
nor U16139 (N_16139,N_15140,N_15133);
nor U16140 (N_16140,N_14194,N_15485);
or U16141 (N_16141,N_14310,N_15540);
xor U16142 (N_16142,N_14291,N_15201);
nor U16143 (N_16143,N_14597,N_14737);
nand U16144 (N_16144,N_15954,N_14420);
and U16145 (N_16145,N_14227,N_14867);
nand U16146 (N_16146,N_14790,N_14642);
xor U16147 (N_16147,N_15795,N_15419);
xor U16148 (N_16148,N_15971,N_14515);
and U16149 (N_16149,N_15831,N_15948);
nor U16150 (N_16150,N_15142,N_15018);
or U16151 (N_16151,N_14149,N_15805);
nand U16152 (N_16152,N_15257,N_15934);
nand U16153 (N_16153,N_15589,N_15168);
nand U16154 (N_16154,N_14306,N_15096);
xnor U16155 (N_16155,N_14507,N_14167);
nor U16156 (N_16156,N_14916,N_15396);
nand U16157 (N_16157,N_15170,N_14279);
xnor U16158 (N_16158,N_14967,N_14481);
and U16159 (N_16159,N_14524,N_15476);
xnor U16160 (N_16160,N_14423,N_14609);
nor U16161 (N_16161,N_14157,N_15398);
or U16162 (N_16162,N_14485,N_14544);
and U16163 (N_16163,N_14678,N_14117);
and U16164 (N_16164,N_15434,N_14806);
xor U16165 (N_16165,N_15318,N_14632);
nand U16166 (N_16166,N_14445,N_15026);
or U16167 (N_16167,N_15743,N_14274);
nand U16168 (N_16168,N_14089,N_14989);
nor U16169 (N_16169,N_14495,N_14044);
nor U16170 (N_16170,N_15887,N_15245);
nor U16171 (N_16171,N_15023,N_14452);
and U16172 (N_16172,N_15289,N_14958);
xor U16173 (N_16173,N_14561,N_15253);
xor U16174 (N_16174,N_15362,N_15294);
and U16175 (N_16175,N_14268,N_14207);
xnor U16176 (N_16176,N_14421,N_15313);
nand U16177 (N_16177,N_14556,N_14062);
and U16178 (N_16178,N_14391,N_14810);
and U16179 (N_16179,N_15978,N_14181);
nand U16180 (N_16180,N_15193,N_14021);
or U16181 (N_16181,N_15781,N_15259);
and U16182 (N_16182,N_15333,N_14830);
and U16183 (N_16183,N_15879,N_14050);
and U16184 (N_16184,N_15417,N_15344);
or U16185 (N_16185,N_15202,N_14410);
xor U16186 (N_16186,N_14282,N_14256);
nand U16187 (N_16187,N_15759,N_14902);
or U16188 (N_16188,N_14534,N_15374);
or U16189 (N_16189,N_14658,N_14076);
or U16190 (N_16190,N_15818,N_15052);
nand U16191 (N_16191,N_14460,N_14253);
or U16192 (N_16192,N_14994,N_15703);
nor U16193 (N_16193,N_14758,N_14093);
nor U16194 (N_16194,N_14612,N_14710);
nor U16195 (N_16195,N_14900,N_14858);
nor U16196 (N_16196,N_14511,N_14223);
xnor U16197 (N_16197,N_15206,N_14708);
xnor U16198 (N_16198,N_14240,N_14362);
nand U16199 (N_16199,N_15203,N_14644);
xor U16200 (N_16200,N_15977,N_14748);
nor U16201 (N_16201,N_15938,N_14224);
xnor U16202 (N_16202,N_15281,N_15182);
nor U16203 (N_16203,N_15178,N_14337);
nor U16204 (N_16204,N_15826,N_14442);
nor U16205 (N_16205,N_15352,N_15477);
nand U16206 (N_16206,N_14304,N_14783);
or U16207 (N_16207,N_14355,N_15288);
nor U16208 (N_16208,N_15651,N_15465);
or U16209 (N_16209,N_15553,N_15129);
and U16210 (N_16210,N_15154,N_15615);
or U16211 (N_16211,N_14968,N_14457);
xnor U16212 (N_16212,N_14462,N_14103);
or U16213 (N_16213,N_14895,N_14012);
xnor U16214 (N_16214,N_15659,N_15397);
nor U16215 (N_16215,N_14284,N_15126);
or U16216 (N_16216,N_14594,N_15059);
xor U16217 (N_16217,N_14659,N_15654);
or U16218 (N_16218,N_15564,N_15997);
xor U16219 (N_16219,N_15243,N_15174);
and U16220 (N_16220,N_14454,N_15234);
or U16221 (N_16221,N_14107,N_15681);
xnor U16222 (N_16222,N_14639,N_14300);
and U16223 (N_16223,N_14071,N_14514);
nor U16224 (N_16224,N_15497,N_15123);
or U16225 (N_16225,N_15014,N_15207);
and U16226 (N_16226,N_14422,N_14051);
xor U16227 (N_16227,N_15882,N_15303);
and U16228 (N_16228,N_15991,N_14332);
nand U16229 (N_16229,N_14105,N_15408);
or U16230 (N_16230,N_15048,N_14536);
and U16231 (N_16231,N_15493,N_15917);
xnor U16232 (N_16232,N_14907,N_15751);
nand U16233 (N_16233,N_14401,N_14666);
nor U16234 (N_16234,N_15623,N_14954);
and U16235 (N_16235,N_14318,N_15124);
and U16236 (N_16236,N_14375,N_15268);
nor U16237 (N_16237,N_15171,N_15046);
nor U16238 (N_16238,N_14052,N_14285);
xor U16239 (N_16239,N_15862,N_14394);
nor U16240 (N_16240,N_14048,N_14829);
nor U16241 (N_16241,N_14246,N_14543);
and U16242 (N_16242,N_15350,N_14086);
xnor U16243 (N_16243,N_14311,N_14010);
nand U16244 (N_16244,N_14668,N_15461);
nand U16245 (N_16245,N_15780,N_15618);
nand U16246 (N_16246,N_15212,N_15543);
or U16247 (N_16247,N_14111,N_14736);
or U16248 (N_16248,N_14697,N_15449);
or U16249 (N_16249,N_14370,N_14962);
and U16250 (N_16250,N_15254,N_14315);
nor U16251 (N_16251,N_15099,N_15020);
nor U16252 (N_16252,N_14894,N_15445);
xor U16253 (N_16253,N_15837,N_14919);
nor U16254 (N_16254,N_15061,N_15517);
and U16255 (N_16255,N_15402,N_14286);
nor U16256 (N_16256,N_15159,N_15378);
xor U16257 (N_16257,N_14385,N_15586);
nor U16258 (N_16258,N_15070,N_14558);
nand U16259 (N_16259,N_14649,N_14535);
nor U16260 (N_16260,N_15803,N_14302);
nor U16261 (N_16261,N_15501,N_15541);
and U16262 (N_16262,N_15370,N_14464);
nor U16263 (N_16263,N_15256,N_14001);
xnor U16264 (N_16264,N_14852,N_15085);
and U16265 (N_16265,N_15507,N_14501);
or U16266 (N_16266,N_15660,N_14453);
xnor U16267 (N_16267,N_14667,N_14933);
xor U16268 (N_16268,N_15731,N_15599);
xor U16269 (N_16269,N_15156,N_14019);
xnor U16270 (N_16270,N_14084,N_15163);
nor U16271 (N_16271,N_15932,N_15283);
xnor U16272 (N_16272,N_14684,N_14386);
and U16273 (N_16273,N_15489,N_15127);
nand U16274 (N_16274,N_15382,N_15612);
or U16275 (N_16275,N_15295,N_15363);
or U16276 (N_16276,N_15875,N_14576);
nand U16277 (N_16277,N_14463,N_15049);
xnor U16278 (N_16278,N_15185,N_15431);
nor U16279 (N_16279,N_15337,N_14653);
xnor U16280 (N_16280,N_15315,N_15779);
nor U16281 (N_16281,N_14142,N_15221);
xnor U16282 (N_16282,N_14709,N_15261);
nand U16283 (N_16283,N_15296,N_15136);
nor U16284 (N_16284,N_15568,N_14254);
and U16285 (N_16285,N_15068,N_15165);
nor U16286 (N_16286,N_14110,N_15964);
and U16287 (N_16287,N_14848,N_14640);
and U16288 (N_16288,N_14049,N_14153);
xnor U16289 (N_16289,N_14565,N_14216);
and U16290 (N_16290,N_14615,N_14714);
xnor U16291 (N_16291,N_15442,N_15897);
or U16292 (N_16292,N_14547,N_15424);
nand U16293 (N_16293,N_14904,N_14408);
and U16294 (N_16294,N_14472,N_14398);
or U16295 (N_16295,N_15106,N_15757);
nor U16296 (N_16296,N_15545,N_15684);
nor U16297 (N_16297,N_15263,N_14582);
or U16298 (N_16298,N_14849,N_15503);
nor U16299 (N_16299,N_15675,N_15317);
and U16300 (N_16300,N_14212,N_14126);
nand U16301 (N_16301,N_14797,N_15384);
xnor U16302 (N_16302,N_14802,N_15336);
nor U16303 (N_16303,N_15983,N_15736);
or U16304 (N_16304,N_15925,N_14804);
or U16305 (N_16305,N_15577,N_15166);
and U16306 (N_16306,N_15225,N_15918);
or U16307 (N_16307,N_14631,N_15531);
or U16308 (N_16308,N_15870,N_15035);
nand U16309 (N_16309,N_15164,N_15583);
xor U16310 (N_16310,N_15919,N_14404);
or U16311 (N_16311,N_15847,N_15566);
nand U16312 (N_16312,N_15789,N_14838);
nand U16313 (N_16313,N_15626,N_14468);
and U16314 (N_16314,N_15393,N_14636);
nor U16315 (N_16315,N_14756,N_14239);
or U16316 (N_16316,N_14045,N_14270);
nor U16317 (N_16317,N_14180,N_15765);
or U16318 (N_16318,N_15112,N_14144);
xor U16319 (N_16319,N_15486,N_14577);
and U16320 (N_16320,N_15346,N_14937);
nor U16321 (N_16321,N_15944,N_14168);
nand U16322 (N_16322,N_14030,N_14193);
nand U16323 (N_16323,N_14585,N_14662);
nand U16324 (N_16324,N_15570,N_15945);
nor U16325 (N_16325,N_14682,N_14186);
nor U16326 (N_16326,N_15399,N_14845);
nor U16327 (N_16327,N_14763,N_15332);
nand U16328 (N_16328,N_15851,N_14889);
nand U16329 (N_16329,N_14357,N_15513);
nor U16330 (N_16330,N_14226,N_15109);
and U16331 (N_16331,N_14343,N_14992);
nor U16332 (N_16332,N_15678,N_15084);
xnor U16333 (N_16333,N_15172,N_14614);
and U16334 (N_16334,N_15455,N_15194);
or U16335 (N_16335,N_14350,N_14528);
and U16336 (N_16336,N_15730,N_15368);
nor U16337 (N_16337,N_15224,N_15377);
or U16338 (N_16338,N_15856,N_14868);
xnor U16339 (N_16339,N_14014,N_14963);
nor U16340 (N_16340,N_15024,N_15372);
or U16341 (N_16341,N_15195,N_14717);
xnor U16342 (N_16342,N_15668,N_14949);
xor U16343 (N_16343,N_14655,N_14687);
nor U16344 (N_16344,N_14784,N_15987);
and U16345 (N_16345,N_14850,N_14006);
nand U16346 (N_16346,N_15644,N_15953);
xnor U16347 (N_16347,N_14586,N_15013);
or U16348 (N_16348,N_14675,N_15797);
nor U16349 (N_16349,N_14057,N_14647);
nor U16350 (N_16350,N_15373,N_15100);
and U16351 (N_16351,N_14112,N_14945);
and U16352 (N_16352,N_15233,N_15547);
nand U16353 (N_16353,N_14898,N_14078);
or U16354 (N_16354,N_14650,N_14027);
xnor U16355 (N_16355,N_14361,N_15305);
nor U16356 (N_16356,N_14190,N_14711);
xor U16357 (N_16357,N_15232,N_15649);
xnor U16358 (N_16358,N_15606,N_14326);
nand U16359 (N_16359,N_14704,N_15146);
nand U16360 (N_16360,N_15082,N_14135);
and U16361 (N_16361,N_15968,N_15537);
xnor U16362 (N_16362,N_15057,N_15770);
xor U16363 (N_16363,N_15416,N_14290);
nor U16364 (N_16364,N_15866,N_15620);
or U16365 (N_16365,N_15998,N_14716);
and U16366 (N_16366,N_15360,N_14940);
and U16367 (N_16367,N_15341,N_14178);
and U16368 (N_16368,N_15188,N_15412);
xor U16369 (N_16369,N_15187,N_14042);
and U16370 (N_16370,N_14262,N_14363);
nand U16371 (N_16371,N_15598,N_15721);
and U16372 (N_16372,N_14584,N_15328);
nand U16373 (N_16373,N_14183,N_14028);
xnor U16374 (N_16374,N_14133,N_14773);
xor U16375 (N_16375,N_14138,N_15450);
nor U16376 (N_16376,N_15927,N_14275);
and U16377 (N_16377,N_14091,N_15957);
and U16378 (N_16378,N_14380,N_15863);
nor U16379 (N_16379,N_15216,N_15697);
nand U16380 (N_16380,N_14247,N_14525);
and U16381 (N_16381,N_15643,N_15602);
and U16382 (N_16382,N_15824,N_15220);
xnor U16383 (N_16383,N_15974,N_14387);
or U16384 (N_16384,N_14599,N_14402);
nand U16385 (N_16385,N_14002,N_14079);
nor U16386 (N_16386,N_15885,N_15839);
xnor U16387 (N_16387,N_15034,N_15874);
or U16388 (N_16388,N_15787,N_14497);
xor U16389 (N_16389,N_14846,N_14690);
or U16390 (N_16390,N_15535,N_15369);
nand U16391 (N_16391,N_15415,N_14860);
or U16392 (N_16392,N_15687,N_14774);
and U16393 (N_16393,N_14269,N_14930);
xor U16394 (N_16394,N_15180,N_15406);
and U16395 (N_16395,N_14513,N_15219);
and U16396 (N_16396,N_15348,N_14211);
xnor U16397 (N_16397,N_15196,N_15558);
or U16398 (N_16398,N_15264,N_15030);
nand U16399 (N_16399,N_14374,N_15158);
nand U16400 (N_16400,N_15522,N_15179);
nor U16401 (N_16401,N_15125,N_15857);
nor U16402 (N_16402,N_14593,N_15949);
or U16403 (N_16403,N_14277,N_14141);
xnor U16404 (N_16404,N_15285,N_15460);
and U16405 (N_16405,N_15813,N_15624);
and U16406 (N_16406,N_14741,N_15446);
or U16407 (N_16407,N_14399,N_15520);
or U16408 (N_16408,N_14499,N_15962);
xor U16409 (N_16409,N_15130,N_14287);
xnor U16410 (N_16410,N_14263,N_15267);
or U16411 (N_16411,N_14616,N_15274);
nand U16412 (N_16412,N_14693,N_14760);
nor U16413 (N_16413,N_15217,N_15055);
nor U16414 (N_16414,N_14466,N_14431);
or U16415 (N_16415,N_14196,N_14099);
and U16416 (N_16416,N_15590,N_15632);
or U16417 (N_16417,N_15955,N_14069);
or U16418 (N_16418,N_15298,N_15989);
nand U16419 (N_16419,N_14624,N_14643);
nand U16420 (N_16420,N_15768,N_14498);
nand U16421 (N_16421,N_14960,N_15593);
xnor U16422 (N_16422,N_14648,N_14156);
nor U16423 (N_16423,N_15510,N_15628);
nand U16424 (N_16424,N_15500,N_14244);
xor U16425 (N_16425,N_14448,N_15720);
nand U16426 (N_16426,N_15011,N_14654);
nor U16427 (N_16427,N_14409,N_15829);
nand U16428 (N_16428,N_15516,N_15808);
nand U16429 (N_16429,N_15755,N_14720);
nor U16430 (N_16430,N_15502,N_15550);
and U16431 (N_16431,N_15942,N_15594);
nand U16432 (N_16432,N_15108,N_15138);
or U16433 (N_16433,N_15043,N_15686);
and U16434 (N_16434,N_14067,N_14841);
xor U16435 (N_16435,N_15992,N_15722);
nand U16436 (N_16436,N_14922,N_14887);
xnor U16437 (N_16437,N_14119,N_14878);
and U16438 (N_16438,N_15959,N_14941);
or U16439 (N_16439,N_14264,N_15028);
and U16440 (N_16440,N_15631,N_15756);
and U16441 (N_16441,N_14389,N_15301);
xnor U16442 (N_16442,N_15761,N_14025);
or U16443 (N_16443,N_15270,N_14202);
nand U16444 (N_16444,N_14696,N_14866);
and U16445 (N_16445,N_15769,N_15290);
or U16446 (N_16446,N_14591,N_15822);
xnor U16447 (N_16447,N_14345,N_15734);
nand U16448 (N_16448,N_15655,N_15680);
and U16449 (N_16449,N_15579,N_15941);
nor U16450 (N_16450,N_14317,N_14455);
nor U16451 (N_16451,N_14348,N_15002);
or U16452 (N_16452,N_14301,N_14392);
nor U16453 (N_16453,N_14935,N_15349);
nor U16454 (N_16454,N_14637,N_15242);
xnor U16455 (N_16455,N_15556,N_14159);
nor U16456 (N_16456,N_15619,N_15157);
or U16457 (N_16457,N_15392,N_14068);
or U16458 (N_16458,N_15036,N_14686);
or U16459 (N_16459,N_15047,N_14596);
and U16460 (N_16460,N_14628,N_15152);
xnor U16461 (N_16461,N_14661,N_14517);
xnor U16462 (N_16462,N_14982,N_14214);
nor U16463 (N_16463,N_15920,N_14746);
xor U16464 (N_16464,N_15717,N_14946);
xor U16465 (N_16465,N_14835,N_14313);
nor U16466 (N_16466,N_15544,N_14503);
or U16467 (N_16467,N_15304,N_15859);
and U16468 (N_16468,N_15884,N_14778);
xor U16469 (N_16469,N_15608,N_15904);
xor U16470 (N_16470,N_14208,N_14447);
nor U16471 (N_16471,N_14891,N_15359);
and U16472 (N_16472,N_15572,N_15139);
xnor U16473 (N_16473,N_15724,N_15058);
or U16474 (N_16474,N_15314,N_14267);
and U16475 (N_16475,N_14231,N_14351);
xnor U16476 (N_16476,N_15389,N_15060);
nand U16477 (N_16477,N_15197,N_15235);
and U16478 (N_16478,N_14502,N_14952);
nor U16479 (N_16479,N_15056,N_14863);
xnor U16480 (N_16480,N_15401,N_14040);
and U16481 (N_16481,N_14925,N_15111);
xor U16482 (N_16482,N_14939,N_15292);
and U16483 (N_16483,N_14098,N_14776);
or U16484 (N_16484,N_14679,N_14324);
nand U16485 (N_16485,N_15355,N_15835);
and U16486 (N_16486,N_15088,N_15471);
nor U16487 (N_16487,N_15524,N_14309);
or U16488 (N_16488,N_15574,N_15252);
or U16489 (N_16489,N_14090,N_15147);
or U16490 (N_16490,N_15864,N_15439);
xnor U16491 (N_16491,N_15872,N_15409);
and U16492 (N_16492,N_15015,N_14102);
or U16493 (N_16493,N_15827,N_15447);
nand U16494 (N_16494,N_14627,N_14998);
and U16495 (N_16495,N_15582,N_14230);
nand U16496 (N_16496,N_15530,N_14871);
nand U16497 (N_16497,N_15533,N_15456);
nand U16498 (N_16498,N_15238,N_14248);
or U16499 (N_16499,N_14623,N_15748);
or U16500 (N_16500,N_15667,N_14066);
nor U16501 (N_16501,N_14171,N_15926);
xnor U16502 (N_16502,N_14794,N_15585);
and U16503 (N_16503,N_15114,N_14166);
or U16504 (N_16504,N_14545,N_14607);
nand U16505 (N_16505,N_15782,N_15708);
xor U16506 (N_16506,N_14229,N_15994);
nor U16507 (N_16507,N_15849,N_14388);
and U16508 (N_16508,N_14413,N_15534);
xnor U16509 (N_16509,N_14222,N_15251);
or U16510 (N_16510,N_14929,N_15413);
nor U16511 (N_16511,N_14289,N_14483);
and U16512 (N_16512,N_15153,N_14322);
and U16513 (N_16513,N_14942,N_15403);
nand U16514 (N_16514,N_14197,N_15210);
or U16515 (N_16515,N_15135,N_15811);
nand U16516 (N_16516,N_15834,N_15183);
and U16517 (N_16517,N_15131,N_15160);
xnor U16518 (N_16518,N_14176,N_14999);
and U16519 (N_16519,N_14983,N_14560);
and U16520 (N_16520,N_14095,N_15546);
nor U16521 (N_16521,N_14831,N_14981);
nand U16522 (N_16522,N_15850,N_14406);
or U16523 (N_16523,N_14698,N_14092);
nor U16524 (N_16524,N_14121,N_15379);
nand U16525 (N_16525,N_14815,N_14053);
and U16526 (N_16526,N_14991,N_15893);
or U16527 (N_16527,N_14673,N_15227);
xor U16528 (N_16528,N_15642,N_14753);
nor U16529 (N_16529,N_15400,N_14974);
nand U16530 (N_16530,N_14874,N_14449);
or U16531 (N_16531,N_14484,N_15454);
or U16532 (N_16532,N_15988,N_15899);
or U16533 (N_16533,N_14956,N_15410);
nor U16534 (N_16534,N_14635,N_14713);
nand U16535 (N_16535,N_15244,N_15331);
xnor U16536 (N_16536,N_15205,N_15262);
and U16537 (N_16537,N_15323,N_14928);
and U16538 (N_16538,N_14634,N_15065);
nand U16539 (N_16539,N_14770,N_14146);
and U16540 (N_16540,N_15664,N_14204);
and U16541 (N_16541,N_14843,N_15895);
nor U16542 (N_16542,N_15032,N_15694);
nand U16543 (N_16543,N_14814,N_15120);
or U16544 (N_16544,N_15639,N_14539);
and U16545 (N_16545,N_15578,N_15812);
nand U16546 (N_16546,N_15072,N_15040);
xnor U16547 (N_16547,N_14670,N_14924);
or U16548 (N_16548,N_14853,N_14729);
xnor U16549 (N_16549,N_15312,N_14134);
and U16550 (N_16550,N_14625,N_15712);
nor U16551 (N_16551,N_15102,N_14793);
xnor U16552 (N_16552,N_14626,N_15796);
nor U16553 (N_16553,N_14781,N_14434);
nor U16554 (N_16554,N_14266,N_14046);
xor U16555 (N_16555,N_15236,N_14015);
and U16556 (N_16556,N_14132,N_15200);
xor U16557 (N_16557,N_14995,N_14836);
or U16558 (N_16558,N_15976,N_15484);
nor U16559 (N_16559,N_14184,N_15749);
nor U16560 (N_16560,N_15707,N_14694);
and U16561 (N_16561,N_14537,N_15799);
xnor U16562 (N_16562,N_14839,N_15973);
nor U16563 (N_16563,N_14683,N_15029);
and U16564 (N_16564,N_14744,N_14342);
and U16565 (N_16565,N_14487,N_15706);
or U16566 (N_16566,N_14518,N_14303);
xnor U16567 (N_16567,N_15890,N_15266);
and U16568 (N_16568,N_15752,N_15764);
xor U16569 (N_16569,N_15433,N_14115);
and U16570 (N_16570,N_15150,N_14340);
and U16571 (N_16571,N_15758,N_14707);
nand U16572 (N_16572,N_15704,N_14825);
nand U16573 (N_16573,N_14424,N_14443);
nand U16574 (N_16574,N_14451,N_15143);
or U16575 (N_16575,N_15271,N_15860);
xor U16576 (N_16576,N_15900,N_14060);
nand U16577 (N_16577,N_14552,N_15386);
or U16578 (N_16578,N_15155,N_14792);
xnor U16579 (N_16579,N_14979,N_15788);
xor U16580 (N_16580,N_14405,N_14260);
nand U16581 (N_16581,N_15074,N_15009);
nor U16582 (N_16582,N_15380,N_15339);
xnor U16583 (N_16583,N_14961,N_15881);
and U16584 (N_16584,N_15871,N_15821);
xnor U16585 (N_16585,N_14299,N_15428);
nand U16586 (N_16586,N_15617,N_15922);
nand U16587 (N_16587,N_15338,N_15740);
nand U16588 (N_16588,N_14938,N_14280);
nor U16589 (N_16589,N_14926,N_15947);
or U16590 (N_16590,N_15414,N_15946);
xnor U16591 (N_16591,N_14570,N_15487);
or U16592 (N_16592,N_14767,N_14890);
nand U16593 (N_16593,N_15498,N_15596);
xor U16594 (N_16594,N_15830,N_15548);
and U16595 (N_16595,N_15366,N_15104);
nor U16596 (N_16596,N_15361,N_14377);
xor U16597 (N_16597,N_15666,N_15483);
xnor U16598 (N_16598,N_14344,N_14948);
nand U16599 (N_16599,N_15719,N_15387);
nand U16600 (N_16600,N_14516,N_15076);
or U16601 (N_16601,N_15033,N_14195);
or U16602 (N_16602,N_14494,N_15260);
xnor U16603 (N_16603,N_14353,N_14947);
xor U16604 (N_16604,N_14298,N_15747);
or U16605 (N_16605,N_14857,N_14251);
and U16606 (N_16606,N_14575,N_14695);
or U16607 (N_16607,N_14726,N_15429);
nand U16608 (N_16608,N_14074,N_14569);
nand U16609 (N_16609,N_15658,N_14143);
or U16610 (N_16610,N_15470,N_15967);
nor U16611 (N_16611,N_14883,N_15679);
nand U16612 (N_16612,N_15723,N_14369);
nor U16613 (N_16613,N_15816,N_15175);
nor U16614 (N_16614,N_15908,N_15275);
or U16615 (N_16615,N_14638,N_14073);
xnor U16616 (N_16616,N_15222,N_14664);
or U16617 (N_16617,N_14734,N_15981);
nand U16618 (N_16618,N_14598,N_14573);
nand U16619 (N_16619,N_15995,N_15031);
xnor U16620 (N_16620,N_14977,N_14550);
nor U16621 (N_16621,N_15552,N_14906);
xor U16622 (N_16622,N_14450,N_14470);
xnor U16623 (N_16623,N_15265,N_15432);
nor U16624 (N_16624,N_15549,N_14376);
nand U16625 (N_16625,N_15280,N_14996);
and U16626 (N_16626,N_14482,N_14540);
xor U16627 (N_16627,N_14331,N_14750);
xor U16628 (N_16628,N_14820,N_15097);
nor U16629 (N_16629,N_14651,N_14441);
nor U16630 (N_16630,N_15802,N_14964);
nand U16631 (N_16631,N_14359,N_14283);
and U16632 (N_16632,N_15451,N_15563);
and U16633 (N_16633,N_15067,N_15001);
nor U16634 (N_16634,N_14786,N_14827);
nor U16635 (N_16635,N_14054,N_15935);
xnor U16636 (N_16636,N_15786,N_14731);
and U16637 (N_16637,N_15610,N_15584);
nor U16638 (N_16638,N_14743,N_15229);
and U16639 (N_16639,N_15273,N_14566);
nand U16640 (N_16640,N_15042,N_14372);
nor U16641 (N_16641,N_15984,N_14440);
and U16642 (N_16642,N_15017,N_15565);
xor U16643 (N_16643,N_15960,N_15132);
xor U16644 (N_16644,N_15066,N_15741);
and U16645 (N_16645,N_15248,N_14061);
and U16646 (N_16646,N_14791,N_15854);
nand U16647 (N_16647,N_14297,N_14745);
and U16648 (N_16648,N_14821,N_15299);
nand U16649 (N_16649,N_14125,N_15508);
nor U16650 (N_16650,N_15891,N_14747);
or U16651 (N_16651,N_14490,N_14003);
and U16652 (N_16652,N_15763,N_14700);
and U16653 (N_16653,N_14308,N_14330);
nand U16654 (N_16654,N_14295,N_14425);
nor U16655 (N_16655,N_15327,N_15966);
and U16656 (N_16656,N_15488,N_15041);
xor U16657 (N_16657,N_14491,N_14779);
xnor U16658 (N_16658,N_14621,N_15750);
xnor U16659 (N_16659,N_15297,N_14718);
and U16660 (N_16660,N_15089,N_15481);
or U16661 (N_16661,N_15701,N_14676);
and U16662 (N_16662,N_14978,N_14798);
and U16663 (N_16663,N_14419,N_14192);
nor U16664 (N_16664,N_14294,N_14873);
nand U16665 (N_16665,N_15121,N_14249);
nand U16666 (N_16666,N_14785,N_15101);
xnor U16667 (N_16667,N_14130,N_15228);
xnor U16668 (N_16668,N_15622,N_14000);
nand U16669 (N_16669,N_14512,N_14601);
or U16670 (N_16670,N_15422,N_14980);
and U16671 (N_16671,N_14329,N_15141);
and U16672 (N_16672,N_14909,N_14699);
and U16673 (N_16673,N_15645,N_15702);
xnor U16674 (N_16674,N_15878,N_15407);
nand U16675 (N_16675,N_15435,N_14590);
nor U16676 (N_16676,N_14618,N_14671);
and U16677 (N_16677,N_14721,N_14465);
xnor U16678 (N_16678,N_14551,N_14738);
nand U16679 (N_16679,N_14258,N_15173);
xor U16680 (N_16680,N_14943,N_15144);
nand U16681 (N_16681,N_15176,N_14473);
nor U16682 (N_16682,N_15956,N_14755);
and U16683 (N_16683,N_15633,N_14522);
nand U16684 (N_16684,N_14766,N_15603);
nand U16685 (N_16685,N_14862,N_15648);
and U16686 (N_16686,N_14986,N_15151);
xnor U16687 (N_16687,N_14217,N_15699);
nand U16688 (N_16688,N_15334,N_14206);
and U16689 (N_16689,N_15969,N_14261);
nand U16690 (N_16690,N_15375,N_14162);
nand U16691 (N_16691,N_15819,N_15554);
nand U16692 (N_16692,N_15716,N_14383);
nor U16693 (N_16693,N_15732,N_14688);
or U16694 (N_16694,N_15354,N_14819);
and U16695 (N_16695,N_14338,N_14011);
nand U16696 (N_16696,N_14439,N_15523);
nand U16697 (N_16697,N_15771,N_14381);
and U16698 (N_16698,N_14706,N_14822);
nor U16699 (N_16699,N_15562,N_14335);
nor U16700 (N_16700,N_15876,N_15576);
and U16701 (N_16701,N_14944,N_15873);
nor U16702 (N_16702,N_15335,N_15801);
nor U16703 (N_16703,N_14506,N_14430);
or U16704 (N_16704,N_14526,N_15430);
or U16705 (N_16705,N_15817,N_15828);
nand U16706 (N_16706,N_14356,N_14505);
nand U16707 (N_16707,N_14321,N_14471);
nand U16708 (N_16708,N_15638,N_15425);
and U16709 (N_16709,N_14951,N_14009);
and U16710 (N_16710,N_15729,N_14273);
nand U16711 (N_16711,N_15943,N_14478);
nand U16712 (N_16712,N_15000,N_15128);
nand U16713 (N_16713,N_15311,N_15613);
or U16714 (N_16714,N_14557,N_15167);
xor U16715 (N_16715,N_14691,N_14059);
nor U16716 (N_16716,N_15685,N_14496);
nor U16717 (N_16717,N_15365,N_14764);
and U16718 (N_16718,N_15437,N_15077);
nand U16719 (N_16719,N_14325,N_15464);
or U16720 (N_16720,N_15776,N_14118);
and U16721 (N_16721,N_14777,N_15737);
xor U16722 (N_16722,N_14579,N_15532);
or U16723 (N_16723,N_15996,N_14237);
nand U16724 (N_16724,N_15105,N_14257);
nand U16725 (N_16725,N_14175,N_15840);
nor U16726 (N_16726,N_14415,N_15869);
nand U16727 (N_16727,N_15342,N_15698);
nand U16728 (N_16728,N_14529,N_14346);
and U16729 (N_16729,N_15980,N_14395);
or U16730 (N_16730,N_14139,N_14971);
or U16731 (N_16731,N_14097,N_15404);
xor U16732 (N_16732,N_14241,N_14931);
or U16733 (N_16733,N_15652,N_14554);
or U16734 (N_16734,N_15069,N_14293);
xnor U16735 (N_16735,N_14201,N_15291);
nand U16736 (N_16736,N_15700,N_15928);
nor U16737 (N_16737,N_14382,N_15117);
nor U16738 (N_16738,N_15090,N_14807);
or U16739 (N_16739,N_14094,N_14493);
xnor U16740 (N_16740,N_14164,N_14187);
xnor U16741 (N_16741,N_14893,N_15356);
nand U16742 (N_16742,N_14692,N_14728);
or U16743 (N_16743,N_14523,N_15888);
nand U16744 (N_16744,N_15086,N_14828);
nor U16745 (N_16745,N_15073,N_15231);
and U16746 (N_16746,N_15555,N_14761);
xnor U16747 (N_16747,N_15078,N_14312);
nor U16748 (N_16748,N_15760,N_15276);
or U16749 (N_16749,N_15791,N_15682);
nand U16750 (N_16750,N_14225,N_15347);
nand U16751 (N_16751,N_15561,N_14771);
xnor U16752 (N_16752,N_15528,N_14757);
or U16753 (N_16753,N_14170,N_15443);
nor U16754 (N_16754,N_15843,N_14123);
and U16755 (N_16755,N_14908,N_15592);
or U16756 (N_16756,N_14879,N_15676);
xnor U16757 (N_16757,N_14173,N_15601);
or U16758 (N_16758,N_15774,N_14358);
and U16759 (N_16759,N_15239,N_14113);
nor U16760 (N_16760,N_15573,N_14276);
xnor U16761 (N_16761,N_15518,N_14740);
nor U16762 (N_16762,N_15634,N_15939);
xor U16763 (N_16763,N_14163,N_14803);
nand U16764 (N_16764,N_14990,N_14371);
nor U16765 (N_16765,N_14036,N_14988);
and U16766 (N_16766,N_14903,N_15814);
or U16767 (N_16767,N_15892,N_14674);
nand U16768 (N_16768,N_14633,N_14339);
and U16769 (N_16769,N_14032,N_15637);
and U16770 (N_16770,N_14703,N_14826);
nand U16771 (N_16771,N_14705,N_14124);
xor U16772 (N_16772,N_14005,N_15950);
nor U16773 (N_16773,N_14437,N_14727);
or U16774 (N_16774,N_14775,N_14681);
or U16775 (N_16775,N_15272,N_15738);
or U16776 (N_16776,N_14058,N_15394);
nor U16777 (N_16777,N_15661,N_15657);
or U16778 (N_16778,N_14219,N_15191);
nor U16779 (N_16779,N_15972,N_15279);
nand U16780 (N_16780,N_15746,N_15538);
nand U16781 (N_16781,N_15640,N_15773);
xor U16782 (N_16782,N_15629,N_15209);
or U16783 (N_16783,N_15308,N_14769);
or U16784 (N_16784,N_15214,N_15003);
and U16785 (N_16785,N_15542,N_14043);
nor U16786 (N_16786,N_15907,N_15975);
nand U16787 (N_16787,N_14151,N_14155);
nand U16788 (N_16788,N_15616,N_14985);
and U16789 (N_16789,N_14923,N_14869);
nor U16790 (N_16790,N_14456,N_14617);
and U16791 (N_16791,N_14932,N_14029);
xor U16792 (N_16792,N_15371,N_14417);
nor U16793 (N_16793,N_15492,N_14328);
and U16794 (N_16794,N_14255,N_15230);
xor U16795 (N_16795,N_14588,N_14595);
nand U16796 (N_16796,N_14022,N_15162);
or U16797 (N_16797,N_14663,N_15912);
and U16798 (N_16798,N_15842,N_14120);
or U16799 (N_16799,N_15911,N_15607);
xnor U16800 (N_16800,N_14959,N_15778);
and U16801 (N_16801,N_15933,N_14911);
and U16802 (N_16802,N_15278,N_15329);
nor U16803 (N_16803,N_14768,N_15062);
and U16804 (N_16804,N_15604,N_15436);
nor U16805 (N_16805,N_15213,N_14652);
nor U16806 (N_16806,N_15071,N_15775);
or U16807 (N_16807,N_15790,N_15081);
or U16808 (N_16808,N_15215,N_14083);
nand U16809 (N_16809,N_15931,N_14955);
nand U16810 (N_16810,N_14812,N_14531);
xnor U16811 (N_16811,N_15636,N_15390);
or U16812 (N_16812,N_15249,N_14064);
and U16813 (N_16813,N_15883,N_14987);
nand U16814 (N_16814,N_14085,N_14877);
nand U16815 (N_16815,N_15915,N_14017);
nand U16816 (N_16816,N_14865,N_14885);
and U16817 (N_16817,N_14136,N_15192);
or U16818 (N_16818,N_14233,N_14851);
or U16819 (N_16819,N_14677,N_15961);
nor U16820 (N_16820,N_14722,N_14480);
and U16821 (N_16821,N_14047,N_14070);
nand U16822 (N_16822,N_15903,N_14613);
nor U16823 (N_16823,N_14600,N_15767);
and U16824 (N_16824,N_14966,N_15526);
or U16825 (N_16825,N_14259,N_14629);
and U16826 (N_16826,N_15838,N_14128);
nand U16827 (N_16827,N_14918,N_14220);
or U16828 (N_16828,N_14809,N_14796);
xor U16829 (N_16829,N_14571,N_14725);
or U16830 (N_16830,N_15846,N_14265);
or U16831 (N_16831,N_14016,N_15909);
or U16832 (N_16832,N_15853,N_14390);
xnor U16833 (N_16833,N_15725,N_15458);
xnor U16834 (N_16834,N_15107,N_15825);
and U16835 (N_16835,N_15539,N_15999);
nor U16836 (N_16836,N_14106,N_14218);
and U16837 (N_16837,N_14892,N_15237);
nand U16838 (N_16838,N_14719,N_15491);
and U16839 (N_16839,N_15010,N_15848);
or U16840 (N_16840,N_14881,N_15965);
nand U16841 (N_16841,N_14788,N_14319);
nand U16842 (N_16842,N_15190,N_14023);
nor U16843 (N_16843,N_15910,N_14739);
nor U16844 (N_16844,N_15340,N_14305);
or U16845 (N_16845,N_15286,N_15198);
and U16846 (N_16846,N_15609,N_14397);
xor U16847 (N_16847,N_14789,N_15269);
xnor U16848 (N_16848,N_14724,N_14314);
nor U16849 (N_16849,N_15683,N_14281);
or U16850 (N_16850,N_15653,N_14444);
nand U16851 (N_16851,N_14993,N_15627);
nor U16852 (N_16852,N_14832,N_15600);
and U16853 (N_16853,N_15426,N_14038);
nand U16854 (N_16854,N_14161,N_14063);
nand U16855 (N_16855,N_15110,N_15587);
xnor U16856 (N_16856,N_15496,N_14913);
and U16857 (N_16857,N_15559,N_14824);
nand U16858 (N_16858,N_15733,N_15189);
and U16859 (N_16859,N_14288,N_14243);
or U16860 (N_16860,N_14082,N_15063);
xnor U16861 (N_16861,N_14818,N_14316);
and U16862 (N_16862,N_15605,N_15690);
nor U16863 (N_16863,N_15438,N_15115);
and U16864 (N_16864,N_15381,N_15457);
xor U16865 (N_16865,N_15309,N_15902);
nor U16866 (N_16866,N_15083,N_15161);
nor U16867 (N_16867,N_15754,N_15351);
nand U16868 (N_16868,N_14567,N_14341);
nor U16869 (N_16869,N_14018,N_15804);
xnor U16870 (N_16870,N_14840,N_15310);
or U16871 (N_16871,N_14414,N_14660);
nor U16872 (N_16872,N_15823,N_15868);
nand U16873 (N_16873,N_15494,N_15343);
nor U16874 (N_16874,N_15621,N_14896);
xnor U16875 (N_16875,N_15635,N_15103);
xor U16876 (N_16876,N_14198,N_14833);
and U16877 (N_16877,N_14366,N_14823);
nand U16878 (N_16878,N_14252,N_14412);
nand U16879 (N_16879,N_14542,N_14917);
nor U16880 (N_16880,N_14323,N_14205);
nor U16881 (N_16881,N_14199,N_15581);
nand U16882 (N_16882,N_15832,N_15588);
nor U16883 (N_16883,N_14075,N_14065);
and U16884 (N_16884,N_15742,N_14160);
nand U16885 (N_16885,N_14817,N_15536);
xnor U16886 (N_16886,N_14035,N_15441);
nor U16887 (N_16887,N_14602,N_14013);
or U16888 (N_16888,N_14780,N_15459);
xnor U16889 (N_16889,N_14973,N_14936);
and U16890 (N_16890,N_14548,N_14521);
nand U16891 (N_16891,N_15012,N_15385);
nand U16892 (N_16892,N_14568,N_14034);
nand U16893 (N_16893,N_14336,N_15647);
and U16894 (N_16894,N_15475,N_14373);
xnor U16895 (N_16895,N_15184,N_14861);
xor U16896 (N_16896,N_14039,N_14572);
nand U16897 (N_16897,N_14672,N_14844);
and U16898 (N_16898,N_15467,N_15358);
nand U16899 (N_16899,N_15116,N_15199);
nor U16900 (N_16900,N_14920,N_15008);
nand U16901 (N_16901,N_14541,N_14519);
or U16902 (N_16902,N_15282,N_14245);
or U16903 (N_16903,N_15411,N_14975);
and U16904 (N_16904,N_14396,N_14426);
or U16905 (N_16905,N_14972,N_14215);
nor U16906 (N_16906,N_14114,N_15614);
xnor U16907 (N_16907,N_15480,N_15145);
nand U16908 (N_16908,N_15079,N_15914);
or U16909 (N_16909,N_15886,N_15499);
and U16910 (N_16910,N_14563,N_14723);
nand U16911 (N_16911,N_14349,N_14347);
and U16912 (N_16912,N_14418,N_15420);
xnor U16913 (N_16913,N_15246,N_15979);
or U16914 (N_16914,N_14367,N_15663);
nor U16915 (N_16915,N_15091,N_15316);
nor U16916 (N_16916,N_14715,N_15982);
nand U16917 (N_16917,N_15656,N_15889);
or U16918 (N_16918,N_14533,N_15952);
and U16919 (N_16919,N_15218,N_14250);
nand U16920 (N_16920,N_14689,N_15324);
nand U16921 (N_16921,N_15691,N_15986);
nor U16922 (N_16922,N_15044,N_15490);
or U16923 (N_16923,N_14458,N_15241);
and U16924 (N_16924,N_15923,N_15662);
nand U16925 (N_16925,N_14622,N_14751);
and U16926 (N_16926,N_15353,N_14680);
or U16927 (N_16927,N_14475,N_15728);
or U16928 (N_16928,N_14438,N_14580);
nor U16929 (N_16929,N_14759,N_14847);
xnor U16930 (N_16930,N_15858,N_15208);
xor U16931 (N_16931,N_15784,N_14581);
nand U16932 (N_16932,N_15844,N_14772);
or U16933 (N_16933,N_14685,N_15845);
and U16934 (N_16934,N_14384,N_14169);
nand U16935 (N_16935,N_15383,N_14553);
and U16936 (N_16936,N_15557,N_14104);
nand U16937 (N_16937,N_14203,N_15094);
xnor U16938 (N_16938,N_14432,N_15472);
xnor U16939 (N_16939,N_14749,N_14630);
xor U16940 (N_16940,N_15794,N_14188);
nand U16941 (N_16941,N_15025,N_14427);
nor U16942 (N_16942,N_14213,N_14145);
xor U16943 (N_16943,N_14108,N_14762);
and U16944 (N_16944,N_14238,N_15320);
xor U16945 (N_16945,N_15113,N_14364);
nand U16946 (N_16946,N_14646,N_14555);
nand U16947 (N_16947,N_14072,N_15894);
or U16948 (N_16948,N_15739,N_14549);
or U16949 (N_16949,N_15715,N_14899);
nor U16950 (N_16950,N_15906,N_14754);
nor U16951 (N_16951,N_14603,N_15921);
nor U16952 (N_16952,N_15571,N_14479);
nand U16953 (N_16953,N_15204,N_14278);
nand U16954 (N_16954,N_14008,N_15039);
nor U16955 (N_16955,N_14886,N_14921);
and U16956 (N_16956,N_14901,N_14559);
xor U16957 (N_16957,N_15929,N_14608);
or U16958 (N_16958,N_14020,N_15718);
xor U16959 (N_16959,N_15186,N_14645);
or U16960 (N_16960,N_15098,N_14752);
and U16961 (N_16961,N_15665,N_14888);
xor U16962 (N_16962,N_14235,N_15575);
and U16963 (N_16963,N_15051,N_14433);
nor U16964 (N_16964,N_14606,N_15924);
xor U16965 (N_16965,N_14842,N_15569);
or U16966 (N_16966,N_14179,N_14669);
nor U16967 (N_16967,N_15793,N_14742);
or U16968 (N_16968,N_14508,N_15692);
xnor U16969 (N_16969,N_14813,N_15087);
xnor U16970 (N_16970,N_15940,N_14428);
and U16971 (N_16971,N_15560,N_15877);
nand U16972 (N_16972,N_15321,N_15469);
nor U16973 (N_16973,N_14360,N_14530);
and U16974 (N_16974,N_15452,N_14033);
or U16975 (N_16975,N_15405,N_14154);
nor U16976 (N_16976,N_15710,N_15836);
or U16977 (N_16977,N_14870,N_14055);
or U16978 (N_16978,N_15322,N_15462);
xnor U16979 (N_16979,N_15970,N_15453);
nor U16980 (N_16980,N_14864,N_15505);
nor U16981 (N_16981,N_15705,N_15119);
xnor U16982 (N_16982,N_15306,N_15726);
xor U16983 (N_16983,N_14610,N_14489);
xnor U16984 (N_16984,N_14461,N_15495);
xor U16985 (N_16985,N_15027,N_15463);
or U16986 (N_16986,N_15357,N_14587);
nand U16987 (N_16987,N_14004,N_15226);
nor U16988 (N_16988,N_15075,N_14037);
and U16989 (N_16989,N_15809,N_15137);
nand U16990 (N_16990,N_15714,N_14953);
and U16991 (N_16991,N_15693,N_14876);
nor U16992 (N_16992,N_14488,N_14007);
nor U16993 (N_16993,N_14446,N_14872);
nand U16994 (N_16994,N_15364,N_15092);
or U16995 (N_16995,N_14403,N_15022);
xnor U16996 (N_16996,N_15936,N_15177);
xnor U16997 (N_16997,N_14137,N_14127);
and U16998 (N_16998,N_15391,N_15753);
or U16999 (N_16999,N_14026,N_14436);
and U17000 (N_17000,N_14818,N_15421);
or U17001 (N_17001,N_15776,N_14934);
nor U17002 (N_17002,N_15264,N_15108);
xnor U17003 (N_17003,N_14141,N_14571);
or U17004 (N_17004,N_14294,N_15049);
nor U17005 (N_17005,N_15961,N_15826);
xor U17006 (N_17006,N_15166,N_14933);
nor U17007 (N_17007,N_14613,N_14798);
nand U17008 (N_17008,N_15404,N_14747);
and U17009 (N_17009,N_15377,N_15782);
nor U17010 (N_17010,N_15552,N_14374);
and U17011 (N_17011,N_14031,N_14727);
xnor U17012 (N_17012,N_14048,N_15032);
nor U17013 (N_17013,N_14823,N_15248);
nand U17014 (N_17014,N_14094,N_15286);
nor U17015 (N_17015,N_15482,N_14344);
nor U17016 (N_17016,N_15785,N_15705);
nand U17017 (N_17017,N_14569,N_14084);
nor U17018 (N_17018,N_15036,N_14394);
xor U17019 (N_17019,N_15949,N_15922);
and U17020 (N_17020,N_14759,N_14641);
nor U17021 (N_17021,N_14755,N_15662);
nand U17022 (N_17022,N_15367,N_15306);
nor U17023 (N_17023,N_14701,N_15315);
xnor U17024 (N_17024,N_15706,N_14922);
or U17025 (N_17025,N_15375,N_15087);
nand U17026 (N_17026,N_14571,N_15885);
or U17027 (N_17027,N_15045,N_14555);
nor U17028 (N_17028,N_15724,N_15118);
nor U17029 (N_17029,N_14238,N_14121);
or U17030 (N_17030,N_15176,N_14145);
nor U17031 (N_17031,N_14007,N_15501);
nand U17032 (N_17032,N_14784,N_15454);
nor U17033 (N_17033,N_14166,N_14664);
nand U17034 (N_17034,N_14035,N_14823);
or U17035 (N_17035,N_15692,N_14863);
nand U17036 (N_17036,N_14243,N_14123);
nand U17037 (N_17037,N_15723,N_14018);
or U17038 (N_17038,N_14604,N_15030);
nand U17039 (N_17039,N_14314,N_15376);
nand U17040 (N_17040,N_14136,N_14355);
nand U17041 (N_17041,N_15598,N_14686);
nand U17042 (N_17042,N_15157,N_15738);
nor U17043 (N_17043,N_15597,N_15327);
xnor U17044 (N_17044,N_14544,N_15340);
nor U17045 (N_17045,N_15583,N_15882);
nor U17046 (N_17046,N_14900,N_14117);
nand U17047 (N_17047,N_15826,N_14639);
xor U17048 (N_17048,N_15593,N_15028);
xor U17049 (N_17049,N_15665,N_15313);
nor U17050 (N_17050,N_15110,N_14521);
nand U17051 (N_17051,N_15817,N_15678);
or U17052 (N_17052,N_14100,N_15736);
and U17053 (N_17053,N_14475,N_14650);
nand U17054 (N_17054,N_14152,N_15291);
xnor U17055 (N_17055,N_14127,N_14536);
nand U17056 (N_17056,N_14748,N_14626);
xnor U17057 (N_17057,N_15996,N_14649);
and U17058 (N_17058,N_15903,N_15518);
and U17059 (N_17059,N_15933,N_14709);
xnor U17060 (N_17060,N_14719,N_15936);
nand U17061 (N_17061,N_14759,N_14429);
nand U17062 (N_17062,N_14843,N_14402);
and U17063 (N_17063,N_14873,N_14936);
nor U17064 (N_17064,N_15357,N_14798);
xnor U17065 (N_17065,N_14751,N_15838);
and U17066 (N_17066,N_14584,N_14452);
nor U17067 (N_17067,N_14947,N_14906);
xnor U17068 (N_17068,N_15568,N_15018);
nor U17069 (N_17069,N_15269,N_14890);
and U17070 (N_17070,N_15756,N_14268);
nand U17071 (N_17071,N_15050,N_14573);
and U17072 (N_17072,N_14668,N_15531);
or U17073 (N_17073,N_14582,N_15132);
nand U17074 (N_17074,N_14227,N_15732);
and U17075 (N_17075,N_15597,N_15585);
and U17076 (N_17076,N_14095,N_14293);
nand U17077 (N_17077,N_15118,N_15824);
or U17078 (N_17078,N_15674,N_14169);
nor U17079 (N_17079,N_14848,N_14192);
or U17080 (N_17080,N_15052,N_14581);
and U17081 (N_17081,N_15355,N_14615);
and U17082 (N_17082,N_14003,N_14795);
nand U17083 (N_17083,N_14471,N_14284);
nor U17084 (N_17084,N_14285,N_14482);
and U17085 (N_17085,N_15790,N_14736);
and U17086 (N_17086,N_14610,N_14199);
nand U17087 (N_17087,N_14174,N_15410);
and U17088 (N_17088,N_15660,N_15624);
or U17089 (N_17089,N_15083,N_14992);
or U17090 (N_17090,N_15331,N_14147);
or U17091 (N_17091,N_15757,N_14397);
xor U17092 (N_17092,N_15111,N_14594);
nand U17093 (N_17093,N_15543,N_14260);
xor U17094 (N_17094,N_15623,N_14878);
and U17095 (N_17095,N_14350,N_15402);
nor U17096 (N_17096,N_15289,N_14592);
and U17097 (N_17097,N_14628,N_14498);
nor U17098 (N_17098,N_14248,N_15839);
xor U17099 (N_17099,N_14274,N_14471);
and U17100 (N_17100,N_14304,N_15392);
or U17101 (N_17101,N_15119,N_14560);
nor U17102 (N_17102,N_15475,N_14406);
nor U17103 (N_17103,N_15182,N_14136);
nand U17104 (N_17104,N_14115,N_15214);
xor U17105 (N_17105,N_15250,N_14889);
nor U17106 (N_17106,N_14322,N_15038);
and U17107 (N_17107,N_14726,N_15102);
and U17108 (N_17108,N_15659,N_15857);
nor U17109 (N_17109,N_15039,N_14839);
xor U17110 (N_17110,N_14612,N_14894);
nor U17111 (N_17111,N_15760,N_14064);
and U17112 (N_17112,N_15967,N_14523);
nor U17113 (N_17113,N_14861,N_15125);
and U17114 (N_17114,N_15814,N_14179);
and U17115 (N_17115,N_15972,N_14395);
and U17116 (N_17116,N_15023,N_14771);
or U17117 (N_17117,N_14024,N_15800);
nand U17118 (N_17118,N_14756,N_15521);
nand U17119 (N_17119,N_15819,N_14886);
xor U17120 (N_17120,N_15762,N_14472);
nand U17121 (N_17121,N_14071,N_15021);
or U17122 (N_17122,N_15679,N_14634);
or U17123 (N_17123,N_15988,N_15968);
and U17124 (N_17124,N_14525,N_15952);
nand U17125 (N_17125,N_15598,N_15890);
nor U17126 (N_17126,N_15664,N_14759);
or U17127 (N_17127,N_15951,N_14915);
and U17128 (N_17128,N_15102,N_15147);
or U17129 (N_17129,N_14868,N_15683);
xor U17130 (N_17130,N_14327,N_15723);
xor U17131 (N_17131,N_15566,N_15664);
and U17132 (N_17132,N_15709,N_15550);
or U17133 (N_17133,N_15094,N_14024);
nor U17134 (N_17134,N_15884,N_14740);
xor U17135 (N_17135,N_15877,N_15323);
and U17136 (N_17136,N_15729,N_15724);
or U17137 (N_17137,N_14396,N_14827);
and U17138 (N_17138,N_15921,N_14412);
and U17139 (N_17139,N_15156,N_14230);
xnor U17140 (N_17140,N_14491,N_14169);
xnor U17141 (N_17141,N_14601,N_15606);
or U17142 (N_17142,N_15381,N_15725);
nor U17143 (N_17143,N_15644,N_15584);
and U17144 (N_17144,N_14896,N_15025);
or U17145 (N_17145,N_14231,N_14184);
xor U17146 (N_17146,N_14497,N_15718);
nand U17147 (N_17147,N_15936,N_15527);
or U17148 (N_17148,N_14270,N_15465);
or U17149 (N_17149,N_14120,N_15186);
nor U17150 (N_17150,N_15100,N_15899);
and U17151 (N_17151,N_14269,N_15476);
and U17152 (N_17152,N_15567,N_14098);
nand U17153 (N_17153,N_15302,N_14887);
or U17154 (N_17154,N_15375,N_15920);
xor U17155 (N_17155,N_15716,N_15257);
nor U17156 (N_17156,N_14415,N_14484);
xnor U17157 (N_17157,N_14909,N_15797);
or U17158 (N_17158,N_14194,N_15804);
nand U17159 (N_17159,N_14620,N_15196);
and U17160 (N_17160,N_14574,N_15090);
nor U17161 (N_17161,N_15827,N_14203);
and U17162 (N_17162,N_14891,N_14187);
or U17163 (N_17163,N_14832,N_15536);
nand U17164 (N_17164,N_14140,N_14000);
and U17165 (N_17165,N_15595,N_14193);
nor U17166 (N_17166,N_14305,N_14711);
nand U17167 (N_17167,N_14556,N_15916);
nor U17168 (N_17168,N_15728,N_14596);
xor U17169 (N_17169,N_15203,N_15599);
nand U17170 (N_17170,N_14244,N_15710);
and U17171 (N_17171,N_14428,N_15168);
nor U17172 (N_17172,N_14210,N_15354);
and U17173 (N_17173,N_15183,N_15042);
or U17174 (N_17174,N_15828,N_14424);
and U17175 (N_17175,N_15843,N_15195);
nor U17176 (N_17176,N_14798,N_15245);
and U17177 (N_17177,N_14759,N_15656);
nand U17178 (N_17178,N_15324,N_14578);
nand U17179 (N_17179,N_14829,N_15783);
or U17180 (N_17180,N_15544,N_15659);
and U17181 (N_17181,N_15502,N_15528);
xor U17182 (N_17182,N_14820,N_14924);
and U17183 (N_17183,N_14284,N_14320);
or U17184 (N_17184,N_14465,N_15437);
nor U17185 (N_17185,N_14217,N_15238);
nor U17186 (N_17186,N_14161,N_15836);
nand U17187 (N_17187,N_15330,N_15646);
and U17188 (N_17188,N_14351,N_15556);
nand U17189 (N_17189,N_15684,N_14113);
nand U17190 (N_17190,N_15619,N_14189);
and U17191 (N_17191,N_14365,N_15079);
nor U17192 (N_17192,N_14849,N_14680);
nand U17193 (N_17193,N_14300,N_15112);
nand U17194 (N_17194,N_15050,N_14747);
and U17195 (N_17195,N_15357,N_14550);
xnor U17196 (N_17196,N_14000,N_15990);
and U17197 (N_17197,N_14673,N_14018);
nor U17198 (N_17198,N_14472,N_14671);
or U17199 (N_17199,N_15776,N_15716);
nor U17200 (N_17200,N_14738,N_14216);
nand U17201 (N_17201,N_14536,N_14783);
nor U17202 (N_17202,N_15633,N_15389);
and U17203 (N_17203,N_14569,N_15372);
nand U17204 (N_17204,N_15280,N_14999);
nor U17205 (N_17205,N_14274,N_15089);
nor U17206 (N_17206,N_15063,N_14726);
xnor U17207 (N_17207,N_14503,N_15751);
nor U17208 (N_17208,N_14443,N_15369);
xnor U17209 (N_17209,N_15816,N_15562);
and U17210 (N_17210,N_15825,N_15957);
nor U17211 (N_17211,N_14488,N_15115);
nor U17212 (N_17212,N_14618,N_14822);
or U17213 (N_17213,N_15160,N_15972);
xnor U17214 (N_17214,N_14979,N_14287);
nor U17215 (N_17215,N_15526,N_15082);
nand U17216 (N_17216,N_15068,N_15314);
xor U17217 (N_17217,N_15474,N_14228);
nor U17218 (N_17218,N_15364,N_15206);
and U17219 (N_17219,N_15917,N_15339);
xnor U17220 (N_17220,N_14648,N_14978);
or U17221 (N_17221,N_14895,N_14382);
nand U17222 (N_17222,N_15296,N_14205);
xor U17223 (N_17223,N_14667,N_14670);
nor U17224 (N_17224,N_14357,N_15791);
nand U17225 (N_17225,N_15224,N_14695);
nand U17226 (N_17226,N_14851,N_14271);
or U17227 (N_17227,N_14126,N_14671);
xnor U17228 (N_17228,N_15982,N_14742);
xor U17229 (N_17229,N_15040,N_15958);
nor U17230 (N_17230,N_14233,N_15689);
and U17231 (N_17231,N_15666,N_14768);
xnor U17232 (N_17232,N_14094,N_14144);
and U17233 (N_17233,N_14886,N_15895);
nor U17234 (N_17234,N_15060,N_14658);
nand U17235 (N_17235,N_15467,N_15651);
nor U17236 (N_17236,N_15237,N_14354);
xor U17237 (N_17237,N_15921,N_14065);
or U17238 (N_17238,N_14550,N_14292);
and U17239 (N_17239,N_14137,N_14109);
or U17240 (N_17240,N_15852,N_14092);
nand U17241 (N_17241,N_15692,N_15582);
nand U17242 (N_17242,N_15231,N_15474);
nor U17243 (N_17243,N_15016,N_15027);
nor U17244 (N_17244,N_15181,N_15974);
or U17245 (N_17245,N_14808,N_15220);
xnor U17246 (N_17246,N_14740,N_14117);
nor U17247 (N_17247,N_14132,N_15705);
or U17248 (N_17248,N_15818,N_15062);
or U17249 (N_17249,N_15423,N_14123);
nand U17250 (N_17250,N_14406,N_15822);
nor U17251 (N_17251,N_14201,N_15428);
and U17252 (N_17252,N_15857,N_14219);
and U17253 (N_17253,N_15469,N_14157);
nor U17254 (N_17254,N_14083,N_15469);
nor U17255 (N_17255,N_14615,N_15803);
and U17256 (N_17256,N_14743,N_14994);
nor U17257 (N_17257,N_14531,N_14367);
or U17258 (N_17258,N_14994,N_15896);
or U17259 (N_17259,N_15097,N_15618);
xnor U17260 (N_17260,N_14007,N_14820);
nand U17261 (N_17261,N_14345,N_14470);
or U17262 (N_17262,N_15584,N_14029);
and U17263 (N_17263,N_14597,N_14586);
xor U17264 (N_17264,N_14159,N_14331);
nor U17265 (N_17265,N_15281,N_14885);
nor U17266 (N_17266,N_15058,N_14214);
nor U17267 (N_17267,N_14641,N_15168);
xor U17268 (N_17268,N_14283,N_15330);
nand U17269 (N_17269,N_14685,N_15093);
and U17270 (N_17270,N_14013,N_15838);
or U17271 (N_17271,N_14302,N_15712);
xnor U17272 (N_17272,N_15282,N_15804);
nand U17273 (N_17273,N_15350,N_14437);
nor U17274 (N_17274,N_14491,N_14462);
and U17275 (N_17275,N_14205,N_14734);
and U17276 (N_17276,N_14939,N_15724);
and U17277 (N_17277,N_14470,N_15125);
or U17278 (N_17278,N_14950,N_14365);
xor U17279 (N_17279,N_15250,N_14043);
or U17280 (N_17280,N_14392,N_15647);
nand U17281 (N_17281,N_15408,N_14881);
nand U17282 (N_17282,N_15332,N_14243);
xnor U17283 (N_17283,N_14642,N_14931);
and U17284 (N_17284,N_14187,N_15865);
nor U17285 (N_17285,N_14639,N_15334);
nand U17286 (N_17286,N_14722,N_15159);
nor U17287 (N_17287,N_15560,N_14231);
nand U17288 (N_17288,N_14360,N_14232);
and U17289 (N_17289,N_14517,N_14189);
xor U17290 (N_17290,N_14845,N_15559);
and U17291 (N_17291,N_15683,N_15949);
or U17292 (N_17292,N_15807,N_15081);
or U17293 (N_17293,N_14444,N_15607);
nor U17294 (N_17294,N_15716,N_15050);
or U17295 (N_17295,N_14170,N_15967);
xnor U17296 (N_17296,N_14958,N_14782);
xnor U17297 (N_17297,N_14837,N_14982);
xnor U17298 (N_17298,N_15996,N_14044);
or U17299 (N_17299,N_15869,N_15901);
nor U17300 (N_17300,N_15376,N_14855);
or U17301 (N_17301,N_14952,N_15384);
xor U17302 (N_17302,N_14294,N_14809);
xor U17303 (N_17303,N_14636,N_14394);
and U17304 (N_17304,N_14952,N_14893);
or U17305 (N_17305,N_15250,N_15263);
and U17306 (N_17306,N_15645,N_14973);
nand U17307 (N_17307,N_14143,N_14651);
or U17308 (N_17308,N_15251,N_14701);
nor U17309 (N_17309,N_15662,N_15107);
nor U17310 (N_17310,N_14742,N_14370);
and U17311 (N_17311,N_14517,N_15906);
or U17312 (N_17312,N_14386,N_14887);
xor U17313 (N_17313,N_14784,N_14988);
nor U17314 (N_17314,N_14429,N_14257);
nand U17315 (N_17315,N_15457,N_15547);
and U17316 (N_17316,N_15824,N_15677);
nand U17317 (N_17317,N_14596,N_14815);
nor U17318 (N_17318,N_15082,N_15478);
nor U17319 (N_17319,N_14600,N_15952);
nand U17320 (N_17320,N_14551,N_14122);
or U17321 (N_17321,N_15418,N_15270);
and U17322 (N_17322,N_15609,N_14086);
xor U17323 (N_17323,N_15617,N_15210);
and U17324 (N_17324,N_14920,N_15033);
or U17325 (N_17325,N_15372,N_14861);
xnor U17326 (N_17326,N_14139,N_14996);
xor U17327 (N_17327,N_14423,N_15538);
and U17328 (N_17328,N_15099,N_15619);
or U17329 (N_17329,N_14711,N_15994);
nor U17330 (N_17330,N_15656,N_14707);
nor U17331 (N_17331,N_15578,N_15087);
and U17332 (N_17332,N_14978,N_15492);
nor U17333 (N_17333,N_14813,N_15513);
nor U17334 (N_17334,N_14147,N_14365);
xor U17335 (N_17335,N_15187,N_14351);
and U17336 (N_17336,N_14392,N_14425);
and U17337 (N_17337,N_15122,N_15698);
nand U17338 (N_17338,N_14632,N_15133);
or U17339 (N_17339,N_14370,N_14569);
xnor U17340 (N_17340,N_14757,N_14248);
xor U17341 (N_17341,N_15470,N_15999);
nor U17342 (N_17342,N_14013,N_14454);
xnor U17343 (N_17343,N_14850,N_14494);
xor U17344 (N_17344,N_15156,N_15673);
xnor U17345 (N_17345,N_14213,N_14343);
and U17346 (N_17346,N_14031,N_14652);
or U17347 (N_17347,N_15293,N_15525);
and U17348 (N_17348,N_15478,N_15165);
and U17349 (N_17349,N_15948,N_15052);
nand U17350 (N_17350,N_15074,N_15407);
nor U17351 (N_17351,N_14161,N_15696);
xnor U17352 (N_17352,N_15966,N_14968);
xnor U17353 (N_17353,N_15854,N_15160);
or U17354 (N_17354,N_15999,N_15900);
or U17355 (N_17355,N_15494,N_14189);
or U17356 (N_17356,N_14992,N_14852);
or U17357 (N_17357,N_15182,N_15788);
nor U17358 (N_17358,N_15586,N_14143);
nor U17359 (N_17359,N_15468,N_15341);
nor U17360 (N_17360,N_15234,N_15494);
nor U17361 (N_17361,N_15030,N_14686);
or U17362 (N_17362,N_14559,N_14854);
xor U17363 (N_17363,N_14719,N_15030);
and U17364 (N_17364,N_14135,N_14049);
or U17365 (N_17365,N_15192,N_14360);
or U17366 (N_17366,N_15478,N_14331);
or U17367 (N_17367,N_14988,N_15396);
and U17368 (N_17368,N_14656,N_15167);
xnor U17369 (N_17369,N_14747,N_14441);
nand U17370 (N_17370,N_15500,N_14214);
or U17371 (N_17371,N_15657,N_14724);
and U17372 (N_17372,N_15226,N_14663);
or U17373 (N_17373,N_15894,N_15634);
or U17374 (N_17374,N_14373,N_14542);
nand U17375 (N_17375,N_15690,N_14533);
or U17376 (N_17376,N_14331,N_15404);
and U17377 (N_17377,N_15157,N_14383);
xor U17378 (N_17378,N_15164,N_15037);
and U17379 (N_17379,N_14024,N_15296);
nand U17380 (N_17380,N_14763,N_15296);
nor U17381 (N_17381,N_14910,N_15575);
and U17382 (N_17382,N_15790,N_14275);
nand U17383 (N_17383,N_14483,N_15820);
nor U17384 (N_17384,N_15744,N_14848);
nor U17385 (N_17385,N_14397,N_15093);
nand U17386 (N_17386,N_14957,N_14567);
nor U17387 (N_17387,N_15038,N_14710);
or U17388 (N_17388,N_14260,N_14192);
xor U17389 (N_17389,N_15115,N_14536);
xnor U17390 (N_17390,N_14091,N_14289);
nand U17391 (N_17391,N_15453,N_15101);
or U17392 (N_17392,N_15615,N_14551);
or U17393 (N_17393,N_15642,N_14951);
nand U17394 (N_17394,N_14976,N_14944);
nor U17395 (N_17395,N_14831,N_15367);
nor U17396 (N_17396,N_15883,N_14083);
nand U17397 (N_17397,N_15738,N_14288);
and U17398 (N_17398,N_14424,N_15126);
nor U17399 (N_17399,N_15560,N_14421);
nor U17400 (N_17400,N_14879,N_15731);
nand U17401 (N_17401,N_15570,N_14410);
nand U17402 (N_17402,N_14311,N_14907);
or U17403 (N_17403,N_14807,N_15894);
xor U17404 (N_17404,N_15019,N_14649);
and U17405 (N_17405,N_14218,N_14016);
nor U17406 (N_17406,N_14670,N_14871);
or U17407 (N_17407,N_15067,N_14982);
nand U17408 (N_17408,N_15578,N_15774);
and U17409 (N_17409,N_14106,N_15520);
nand U17410 (N_17410,N_15327,N_14171);
xnor U17411 (N_17411,N_14743,N_14023);
and U17412 (N_17412,N_14888,N_15530);
nand U17413 (N_17413,N_14491,N_15853);
xnor U17414 (N_17414,N_15735,N_15643);
and U17415 (N_17415,N_15067,N_15480);
nand U17416 (N_17416,N_14697,N_14042);
or U17417 (N_17417,N_15676,N_14083);
nor U17418 (N_17418,N_15298,N_15106);
nand U17419 (N_17419,N_14544,N_14752);
and U17420 (N_17420,N_15932,N_15244);
xor U17421 (N_17421,N_14785,N_15797);
and U17422 (N_17422,N_15066,N_14817);
nor U17423 (N_17423,N_15254,N_14520);
nor U17424 (N_17424,N_14904,N_14335);
nand U17425 (N_17425,N_15743,N_15691);
nand U17426 (N_17426,N_14609,N_15795);
or U17427 (N_17427,N_15822,N_14822);
nor U17428 (N_17428,N_15788,N_15975);
nor U17429 (N_17429,N_14168,N_14878);
nand U17430 (N_17430,N_14211,N_14816);
nand U17431 (N_17431,N_15742,N_14169);
xor U17432 (N_17432,N_15541,N_14965);
nor U17433 (N_17433,N_15690,N_14626);
nor U17434 (N_17434,N_15258,N_14581);
and U17435 (N_17435,N_15849,N_14896);
xor U17436 (N_17436,N_15228,N_15055);
and U17437 (N_17437,N_15192,N_14730);
or U17438 (N_17438,N_15828,N_15525);
nand U17439 (N_17439,N_15098,N_15769);
xnor U17440 (N_17440,N_15751,N_15155);
and U17441 (N_17441,N_15387,N_15768);
nand U17442 (N_17442,N_15705,N_15732);
nor U17443 (N_17443,N_14068,N_14626);
and U17444 (N_17444,N_15239,N_14970);
nand U17445 (N_17445,N_15209,N_14693);
xnor U17446 (N_17446,N_14016,N_14335);
nand U17447 (N_17447,N_15555,N_14624);
nand U17448 (N_17448,N_14517,N_15981);
nor U17449 (N_17449,N_14182,N_15617);
nand U17450 (N_17450,N_14357,N_15717);
and U17451 (N_17451,N_15699,N_14577);
or U17452 (N_17452,N_14563,N_14333);
xor U17453 (N_17453,N_15374,N_15105);
nor U17454 (N_17454,N_15013,N_15322);
nand U17455 (N_17455,N_14353,N_15580);
or U17456 (N_17456,N_14746,N_14882);
nor U17457 (N_17457,N_15327,N_15737);
nand U17458 (N_17458,N_14852,N_14667);
nor U17459 (N_17459,N_14751,N_15680);
and U17460 (N_17460,N_15572,N_15680);
nand U17461 (N_17461,N_15983,N_15826);
and U17462 (N_17462,N_15211,N_14246);
xnor U17463 (N_17463,N_15293,N_14395);
xnor U17464 (N_17464,N_14707,N_15427);
or U17465 (N_17465,N_15693,N_14979);
nor U17466 (N_17466,N_15715,N_14413);
nand U17467 (N_17467,N_15326,N_15969);
and U17468 (N_17468,N_14481,N_14735);
and U17469 (N_17469,N_14865,N_15007);
nor U17470 (N_17470,N_15463,N_15184);
nor U17471 (N_17471,N_14175,N_14209);
or U17472 (N_17472,N_14803,N_14497);
or U17473 (N_17473,N_15274,N_15377);
xnor U17474 (N_17474,N_15193,N_15354);
nand U17475 (N_17475,N_15026,N_14089);
or U17476 (N_17476,N_14035,N_14462);
xnor U17477 (N_17477,N_15312,N_15731);
nand U17478 (N_17478,N_15065,N_14575);
or U17479 (N_17479,N_15001,N_15902);
or U17480 (N_17480,N_15855,N_14494);
nor U17481 (N_17481,N_14959,N_15501);
xor U17482 (N_17482,N_15713,N_15440);
xnor U17483 (N_17483,N_14271,N_14809);
nand U17484 (N_17484,N_14837,N_15415);
nand U17485 (N_17485,N_14246,N_14484);
or U17486 (N_17486,N_14308,N_14388);
nand U17487 (N_17487,N_14301,N_14916);
nand U17488 (N_17488,N_14792,N_14746);
nand U17489 (N_17489,N_15219,N_14271);
nor U17490 (N_17490,N_15931,N_14807);
and U17491 (N_17491,N_14245,N_14629);
xor U17492 (N_17492,N_14909,N_14509);
nor U17493 (N_17493,N_15786,N_14749);
nor U17494 (N_17494,N_14082,N_14709);
nor U17495 (N_17495,N_15506,N_15523);
and U17496 (N_17496,N_14948,N_15950);
xor U17497 (N_17497,N_14409,N_14312);
nor U17498 (N_17498,N_15995,N_14636);
and U17499 (N_17499,N_14656,N_15804);
xor U17500 (N_17500,N_15145,N_14686);
nand U17501 (N_17501,N_15339,N_15963);
xnor U17502 (N_17502,N_15531,N_15649);
nor U17503 (N_17503,N_14340,N_15554);
or U17504 (N_17504,N_15067,N_15815);
nor U17505 (N_17505,N_14181,N_14719);
xnor U17506 (N_17506,N_15849,N_14133);
and U17507 (N_17507,N_15469,N_14051);
or U17508 (N_17508,N_15666,N_14157);
or U17509 (N_17509,N_15005,N_15127);
nand U17510 (N_17510,N_14808,N_14832);
or U17511 (N_17511,N_14123,N_15794);
and U17512 (N_17512,N_15608,N_15957);
xnor U17513 (N_17513,N_14951,N_15919);
nand U17514 (N_17514,N_14993,N_14511);
xor U17515 (N_17515,N_14680,N_14429);
nand U17516 (N_17516,N_14577,N_14441);
and U17517 (N_17517,N_14894,N_15787);
nand U17518 (N_17518,N_15289,N_14928);
nand U17519 (N_17519,N_15792,N_14005);
nor U17520 (N_17520,N_15338,N_15972);
nor U17521 (N_17521,N_14396,N_14740);
nor U17522 (N_17522,N_15043,N_15648);
nand U17523 (N_17523,N_14790,N_14462);
nor U17524 (N_17524,N_14232,N_15317);
nor U17525 (N_17525,N_15890,N_14163);
and U17526 (N_17526,N_14710,N_15018);
and U17527 (N_17527,N_14709,N_15528);
nand U17528 (N_17528,N_15504,N_14959);
and U17529 (N_17529,N_14106,N_15955);
nand U17530 (N_17530,N_14619,N_15794);
xnor U17531 (N_17531,N_14030,N_15094);
nand U17532 (N_17532,N_15882,N_14749);
nor U17533 (N_17533,N_15099,N_14689);
and U17534 (N_17534,N_15981,N_15554);
and U17535 (N_17535,N_15342,N_15002);
and U17536 (N_17536,N_14378,N_14470);
and U17537 (N_17537,N_15918,N_15067);
xor U17538 (N_17538,N_15965,N_15692);
xnor U17539 (N_17539,N_15642,N_14146);
nand U17540 (N_17540,N_15569,N_14712);
and U17541 (N_17541,N_15746,N_14482);
or U17542 (N_17542,N_15770,N_15064);
nor U17543 (N_17543,N_15552,N_15786);
xor U17544 (N_17544,N_14266,N_14005);
nor U17545 (N_17545,N_15519,N_15052);
xor U17546 (N_17546,N_14661,N_14437);
nand U17547 (N_17547,N_15359,N_15446);
nor U17548 (N_17548,N_14649,N_14739);
or U17549 (N_17549,N_14241,N_15297);
or U17550 (N_17550,N_14916,N_14023);
and U17551 (N_17551,N_15148,N_14221);
or U17552 (N_17552,N_14943,N_14123);
and U17553 (N_17553,N_15769,N_15978);
or U17554 (N_17554,N_15469,N_14161);
nand U17555 (N_17555,N_15680,N_14390);
and U17556 (N_17556,N_14623,N_15323);
nand U17557 (N_17557,N_15732,N_15216);
nand U17558 (N_17558,N_14915,N_14105);
nor U17559 (N_17559,N_15954,N_14556);
nor U17560 (N_17560,N_14200,N_14312);
nor U17561 (N_17561,N_14998,N_15265);
nand U17562 (N_17562,N_15475,N_14226);
xor U17563 (N_17563,N_14657,N_14552);
xor U17564 (N_17564,N_15687,N_14080);
nand U17565 (N_17565,N_14187,N_14223);
xor U17566 (N_17566,N_14175,N_15233);
nand U17567 (N_17567,N_14566,N_15583);
and U17568 (N_17568,N_15173,N_15149);
xor U17569 (N_17569,N_15154,N_14246);
or U17570 (N_17570,N_14161,N_15120);
or U17571 (N_17571,N_14432,N_15973);
nand U17572 (N_17572,N_14670,N_14270);
or U17573 (N_17573,N_14221,N_14575);
or U17574 (N_17574,N_14127,N_14163);
nor U17575 (N_17575,N_15509,N_15273);
xnor U17576 (N_17576,N_14800,N_14273);
xnor U17577 (N_17577,N_14779,N_15644);
or U17578 (N_17578,N_15170,N_14024);
nand U17579 (N_17579,N_14101,N_14095);
or U17580 (N_17580,N_14885,N_14351);
nand U17581 (N_17581,N_15442,N_14670);
nor U17582 (N_17582,N_15551,N_14750);
or U17583 (N_17583,N_15449,N_14084);
xor U17584 (N_17584,N_15360,N_14619);
and U17585 (N_17585,N_14468,N_14011);
xor U17586 (N_17586,N_15682,N_14815);
xnor U17587 (N_17587,N_14079,N_15650);
or U17588 (N_17588,N_15705,N_14169);
xor U17589 (N_17589,N_14433,N_15766);
or U17590 (N_17590,N_14903,N_15309);
nand U17591 (N_17591,N_15049,N_15972);
xnor U17592 (N_17592,N_15335,N_14069);
nor U17593 (N_17593,N_14277,N_14902);
nor U17594 (N_17594,N_14901,N_15561);
xor U17595 (N_17595,N_14064,N_14574);
xor U17596 (N_17596,N_14493,N_15088);
and U17597 (N_17597,N_15410,N_14372);
xor U17598 (N_17598,N_14158,N_14530);
nor U17599 (N_17599,N_15793,N_14129);
nor U17600 (N_17600,N_14262,N_14565);
xnor U17601 (N_17601,N_15350,N_14226);
xnor U17602 (N_17602,N_15029,N_14496);
nand U17603 (N_17603,N_15729,N_14368);
and U17604 (N_17604,N_15277,N_14680);
or U17605 (N_17605,N_15190,N_15750);
or U17606 (N_17606,N_14794,N_14748);
xor U17607 (N_17607,N_14783,N_14122);
nand U17608 (N_17608,N_14661,N_14405);
nor U17609 (N_17609,N_15498,N_15909);
or U17610 (N_17610,N_14654,N_15362);
xnor U17611 (N_17611,N_14769,N_14631);
nand U17612 (N_17612,N_14277,N_14065);
xnor U17613 (N_17613,N_15538,N_14528);
nand U17614 (N_17614,N_14328,N_14259);
and U17615 (N_17615,N_14457,N_15905);
and U17616 (N_17616,N_14629,N_15839);
or U17617 (N_17617,N_14440,N_15131);
xnor U17618 (N_17618,N_15671,N_14899);
or U17619 (N_17619,N_14826,N_15323);
xor U17620 (N_17620,N_14478,N_15563);
nor U17621 (N_17621,N_15803,N_15931);
or U17622 (N_17622,N_14283,N_14609);
nor U17623 (N_17623,N_14226,N_15224);
and U17624 (N_17624,N_15608,N_15889);
or U17625 (N_17625,N_15852,N_14116);
nor U17626 (N_17626,N_14977,N_14615);
and U17627 (N_17627,N_15632,N_15328);
nor U17628 (N_17628,N_15854,N_14942);
nand U17629 (N_17629,N_14754,N_15704);
xor U17630 (N_17630,N_14178,N_15406);
and U17631 (N_17631,N_15401,N_14367);
or U17632 (N_17632,N_15481,N_14396);
and U17633 (N_17633,N_15842,N_15887);
nand U17634 (N_17634,N_15348,N_15249);
and U17635 (N_17635,N_14550,N_14258);
nor U17636 (N_17636,N_15909,N_14734);
nand U17637 (N_17637,N_14422,N_15005);
nand U17638 (N_17638,N_14232,N_14554);
nand U17639 (N_17639,N_14060,N_15448);
or U17640 (N_17640,N_15818,N_14865);
or U17641 (N_17641,N_14208,N_15803);
nand U17642 (N_17642,N_15535,N_15874);
nand U17643 (N_17643,N_14733,N_14836);
nand U17644 (N_17644,N_15643,N_15332);
xor U17645 (N_17645,N_15131,N_15426);
or U17646 (N_17646,N_15463,N_15477);
or U17647 (N_17647,N_14249,N_15249);
xor U17648 (N_17648,N_15174,N_14293);
or U17649 (N_17649,N_15683,N_14207);
xor U17650 (N_17650,N_15918,N_14057);
or U17651 (N_17651,N_15841,N_15895);
or U17652 (N_17652,N_15452,N_14830);
or U17653 (N_17653,N_15591,N_15943);
or U17654 (N_17654,N_15436,N_14781);
nand U17655 (N_17655,N_14922,N_15560);
xor U17656 (N_17656,N_15115,N_15979);
nand U17657 (N_17657,N_14167,N_14723);
and U17658 (N_17658,N_15923,N_14210);
nand U17659 (N_17659,N_14829,N_14874);
nor U17660 (N_17660,N_14469,N_15632);
nand U17661 (N_17661,N_15761,N_15530);
and U17662 (N_17662,N_14702,N_14581);
nand U17663 (N_17663,N_15492,N_15401);
xor U17664 (N_17664,N_14478,N_14162);
or U17665 (N_17665,N_15825,N_14515);
nand U17666 (N_17666,N_15314,N_15836);
xor U17667 (N_17667,N_14244,N_15791);
nand U17668 (N_17668,N_14138,N_15939);
or U17669 (N_17669,N_15479,N_15965);
or U17670 (N_17670,N_14098,N_14168);
nor U17671 (N_17671,N_15170,N_14518);
or U17672 (N_17672,N_14881,N_15585);
and U17673 (N_17673,N_14999,N_14504);
and U17674 (N_17674,N_15385,N_15651);
xor U17675 (N_17675,N_14383,N_14251);
and U17676 (N_17676,N_15575,N_15811);
and U17677 (N_17677,N_15516,N_14024);
or U17678 (N_17678,N_15686,N_14544);
xor U17679 (N_17679,N_14204,N_15903);
and U17680 (N_17680,N_14400,N_14399);
xor U17681 (N_17681,N_15483,N_14874);
xor U17682 (N_17682,N_15000,N_15493);
and U17683 (N_17683,N_15799,N_15945);
nand U17684 (N_17684,N_15609,N_14291);
xor U17685 (N_17685,N_14457,N_15602);
xor U17686 (N_17686,N_15102,N_15353);
xnor U17687 (N_17687,N_15319,N_14034);
nor U17688 (N_17688,N_15821,N_15722);
or U17689 (N_17689,N_15470,N_15771);
and U17690 (N_17690,N_15023,N_14545);
xor U17691 (N_17691,N_14343,N_14025);
nor U17692 (N_17692,N_14429,N_14248);
nor U17693 (N_17693,N_15588,N_14780);
nor U17694 (N_17694,N_15672,N_15860);
and U17695 (N_17695,N_14889,N_14940);
or U17696 (N_17696,N_15684,N_14535);
or U17697 (N_17697,N_15182,N_15188);
nand U17698 (N_17698,N_15719,N_15458);
and U17699 (N_17699,N_15707,N_15204);
xor U17700 (N_17700,N_15921,N_15075);
nor U17701 (N_17701,N_15278,N_14620);
or U17702 (N_17702,N_15131,N_14002);
and U17703 (N_17703,N_15131,N_14525);
xor U17704 (N_17704,N_15825,N_15623);
xnor U17705 (N_17705,N_15793,N_15140);
and U17706 (N_17706,N_14984,N_15646);
nand U17707 (N_17707,N_15862,N_15681);
nand U17708 (N_17708,N_15724,N_15977);
or U17709 (N_17709,N_15429,N_14304);
nand U17710 (N_17710,N_15591,N_15411);
and U17711 (N_17711,N_14316,N_14453);
nor U17712 (N_17712,N_15644,N_14225);
nand U17713 (N_17713,N_15616,N_15640);
and U17714 (N_17714,N_15692,N_14616);
xnor U17715 (N_17715,N_14291,N_14428);
nand U17716 (N_17716,N_14326,N_15397);
or U17717 (N_17717,N_15273,N_14558);
nor U17718 (N_17718,N_15362,N_14880);
or U17719 (N_17719,N_14286,N_15252);
or U17720 (N_17720,N_15823,N_15561);
nand U17721 (N_17721,N_14082,N_15275);
and U17722 (N_17722,N_15252,N_14109);
nor U17723 (N_17723,N_15879,N_14518);
xnor U17724 (N_17724,N_15906,N_15944);
nor U17725 (N_17725,N_14940,N_14270);
nand U17726 (N_17726,N_14333,N_14702);
nand U17727 (N_17727,N_14508,N_15513);
nand U17728 (N_17728,N_14704,N_14159);
or U17729 (N_17729,N_15530,N_15576);
nand U17730 (N_17730,N_15866,N_15138);
and U17731 (N_17731,N_15819,N_14303);
nor U17732 (N_17732,N_15763,N_14922);
and U17733 (N_17733,N_15194,N_15276);
nand U17734 (N_17734,N_15014,N_14146);
and U17735 (N_17735,N_14821,N_14210);
nand U17736 (N_17736,N_14351,N_14270);
nor U17737 (N_17737,N_15586,N_15395);
nor U17738 (N_17738,N_14846,N_14694);
nor U17739 (N_17739,N_14177,N_15112);
nand U17740 (N_17740,N_14580,N_14996);
or U17741 (N_17741,N_14952,N_14237);
nand U17742 (N_17742,N_14109,N_14970);
and U17743 (N_17743,N_14537,N_14061);
and U17744 (N_17744,N_15460,N_15911);
nand U17745 (N_17745,N_14888,N_15472);
or U17746 (N_17746,N_15008,N_14470);
and U17747 (N_17747,N_14165,N_15577);
and U17748 (N_17748,N_15814,N_14217);
or U17749 (N_17749,N_15108,N_15670);
nand U17750 (N_17750,N_14376,N_14959);
nor U17751 (N_17751,N_14725,N_15889);
xor U17752 (N_17752,N_14048,N_14450);
or U17753 (N_17753,N_14785,N_14232);
nor U17754 (N_17754,N_15507,N_15141);
or U17755 (N_17755,N_14727,N_14594);
nand U17756 (N_17756,N_14519,N_14662);
or U17757 (N_17757,N_15048,N_14684);
nand U17758 (N_17758,N_15770,N_14652);
nand U17759 (N_17759,N_14429,N_15796);
and U17760 (N_17760,N_14911,N_15752);
and U17761 (N_17761,N_14887,N_14513);
xor U17762 (N_17762,N_15888,N_14327);
or U17763 (N_17763,N_15940,N_14210);
or U17764 (N_17764,N_15501,N_14488);
nor U17765 (N_17765,N_14493,N_14613);
or U17766 (N_17766,N_15833,N_14258);
nand U17767 (N_17767,N_15057,N_14219);
xnor U17768 (N_17768,N_15692,N_15293);
nor U17769 (N_17769,N_14916,N_15295);
nand U17770 (N_17770,N_15457,N_15835);
or U17771 (N_17771,N_15149,N_15103);
nor U17772 (N_17772,N_15046,N_14253);
or U17773 (N_17773,N_15616,N_14432);
nor U17774 (N_17774,N_14267,N_14338);
xnor U17775 (N_17775,N_14151,N_15520);
or U17776 (N_17776,N_14013,N_14669);
nand U17777 (N_17777,N_15535,N_14614);
nor U17778 (N_17778,N_14302,N_15912);
or U17779 (N_17779,N_14559,N_14206);
and U17780 (N_17780,N_14643,N_14562);
xor U17781 (N_17781,N_14078,N_15507);
and U17782 (N_17782,N_14995,N_15256);
and U17783 (N_17783,N_15489,N_15668);
or U17784 (N_17784,N_15846,N_14162);
nor U17785 (N_17785,N_14515,N_14762);
nand U17786 (N_17786,N_15225,N_15159);
nand U17787 (N_17787,N_14021,N_15433);
nor U17788 (N_17788,N_15018,N_15534);
or U17789 (N_17789,N_15260,N_14752);
nor U17790 (N_17790,N_14889,N_15689);
or U17791 (N_17791,N_15480,N_14385);
nand U17792 (N_17792,N_15027,N_14619);
or U17793 (N_17793,N_15001,N_15986);
nor U17794 (N_17794,N_14428,N_14943);
and U17795 (N_17795,N_15080,N_14070);
and U17796 (N_17796,N_14805,N_15131);
nand U17797 (N_17797,N_14604,N_14159);
xor U17798 (N_17798,N_15552,N_15877);
nand U17799 (N_17799,N_15288,N_15009);
and U17800 (N_17800,N_14353,N_14440);
and U17801 (N_17801,N_15308,N_14449);
nand U17802 (N_17802,N_14542,N_15133);
xnor U17803 (N_17803,N_15030,N_15654);
xnor U17804 (N_17804,N_14647,N_15861);
nand U17805 (N_17805,N_15787,N_15512);
nor U17806 (N_17806,N_15376,N_14657);
and U17807 (N_17807,N_14524,N_15711);
and U17808 (N_17808,N_15586,N_15455);
nor U17809 (N_17809,N_14862,N_15182);
xnor U17810 (N_17810,N_14293,N_15310);
nand U17811 (N_17811,N_15452,N_15885);
nand U17812 (N_17812,N_15144,N_15437);
nor U17813 (N_17813,N_14302,N_15515);
or U17814 (N_17814,N_15472,N_14970);
nand U17815 (N_17815,N_15216,N_14558);
nand U17816 (N_17816,N_14189,N_15733);
nor U17817 (N_17817,N_14271,N_15260);
nor U17818 (N_17818,N_15350,N_15401);
nand U17819 (N_17819,N_15165,N_15786);
and U17820 (N_17820,N_15368,N_14856);
or U17821 (N_17821,N_15970,N_15066);
nand U17822 (N_17822,N_14852,N_14391);
nand U17823 (N_17823,N_14078,N_14180);
nor U17824 (N_17824,N_14457,N_14882);
and U17825 (N_17825,N_14878,N_14974);
and U17826 (N_17826,N_14169,N_15734);
and U17827 (N_17827,N_14502,N_14285);
xor U17828 (N_17828,N_14487,N_14917);
nand U17829 (N_17829,N_15915,N_14764);
or U17830 (N_17830,N_14535,N_14039);
or U17831 (N_17831,N_14623,N_15979);
or U17832 (N_17832,N_14063,N_14793);
nand U17833 (N_17833,N_14578,N_15915);
nand U17834 (N_17834,N_14085,N_14348);
or U17835 (N_17835,N_14637,N_14505);
and U17836 (N_17836,N_14729,N_14613);
nand U17837 (N_17837,N_14995,N_15670);
nand U17838 (N_17838,N_14479,N_15265);
xor U17839 (N_17839,N_14446,N_14984);
and U17840 (N_17840,N_14473,N_14621);
nor U17841 (N_17841,N_14656,N_14268);
or U17842 (N_17842,N_15402,N_14274);
nor U17843 (N_17843,N_15670,N_15663);
and U17844 (N_17844,N_14505,N_15075);
xor U17845 (N_17845,N_15462,N_14643);
nor U17846 (N_17846,N_14621,N_14753);
nor U17847 (N_17847,N_14649,N_14471);
xor U17848 (N_17848,N_15038,N_15723);
and U17849 (N_17849,N_15967,N_15743);
and U17850 (N_17850,N_14084,N_14446);
nor U17851 (N_17851,N_14734,N_15719);
nor U17852 (N_17852,N_14973,N_15227);
and U17853 (N_17853,N_14833,N_14694);
and U17854 (N_17854,N_15994,N_15095);
nand U17855 (N_17855,N_15815,N_14820);
nand U17856 (N_17856,N_15878,N_14140);
nor U17857 (N_17857,N_14057,N_14359);
or U17858 (N_17858,N_14216,N_15318);
nand U17859 (N_17859,N_14442,N_15519);
nand U17860 (N_17860,N_14694,N_14484);
and U17861 (N_17861,N_14004,N_15648);
xor U17862 (N_17862,N_15579,N_15424);
xnor U17863 (N_17863,N_14905,N_15843);
nor U17864 (N_17864,N_14599,N_14789);
or U17865 (N_17865,N_15923,N_15831);
nor U17866 (N_17866,N_14638,N_15739);
or U17867 (N_17867,N_15433,N_15984);
or U17868 (N_17868,N_15024,N_15353);
xor U17869 (N_17869,N_15441,N_15034);
nor U17870 (N_17870,N_15737,N_14287);
nand U17871 (N_17871,N_14089,N_14148);
nor U17872 (N_17872,N_15844,N_15267);
nor U17873 (N_17873,N_15736,N_15484);
xor U17874 (N_17874,N_14504,N_14209);
nor U17875 (N_17875,N_14108,N_15886);
or U17876 (N_17876,N_15783,N_15028);
xnor U17877 (N_17877,N_15862,N_14436);
or U17878 (N_17878,N_15504,N_14683);
or U17879 (N_17879,N_14657,N_14082);
or U17880 (N_17880,N_14835,N_15199);
or U17881 (N_17881,N_14848,N_15048);
or U17882 (N_17882,N_14013,N_15933);
or U17883 (N_17883,N_14842,N_14927);
xnor U17884 (N_17884,N_14497,N_15281);
xnor U17885 (N_17885,N_14716,N_14695);
nor U17886 (N_17886,N_14630,N_14133);
and U17887 (N_17887,N_15376,N_15976);
xor U17888 (N_17888,N_14008,N_14570);
and U17889 (N_17889,N_15090,N_14321);
nor U17890 (N_17890,N_14388,N_15954);
xor U17891 (N_17891,N_15694,N_15266);
or U17892 (N_17892,N_14060,N_14632);
or U17893 (N_17893,N_14520,N_15472);
nand U17894 (N_17894,N_15602,N_15530);
xnor U17895 (N_17895,N_15294,N_15906);
or U17896 (N_17896,N_15897,N_14890);
nor U17897 (N_17897,N_14416,N_14806);
nor U17898 (N_17898,N_14750,N_14459);
nand U17899 (N_17899,N_14959,N_14720);
and U17900 (N_17900,N_14823,N_15027);
or U17901 (N_17901,N_15486,N_15315);
nor U17902 (N_17902,N_15578,N_14443);
nor U17903 (N_17903,N_14965,N_15967);
or U17904 (N_17904,N_15832,N_15938);
nor U17905 (N_17905,N_14071,N_15139);
and U17906 (N_17906,N_15247,N_14986);
nand U17907 (N_17907,N_15208,N_15284);
and U17908 (N_17908,N_15302,N_15338);
xor U17909 (N_17909,N_14993,N_15070);
xnor U17910 (N_17910,N_15776,N_14970);
nor U17911 (N_17911,N_14801,N_14915);
xor U17912 (N_17912,N_15430,N_15353);
or U17913 (N_17913,N_14109,N_15511);
or U17914 (N_17914,N_15758,N_15455);
nand U17915 (N_17915,N_14645,N_14882);
nand U17916 (N_17916,N_15188,N_14929);
or U17917 (N_17917,N_14633,N_15696);
or U17918 (N_17918,N_15648,N_14790);
and U17919 (N_17919,N_15742,N_15620);
nor U17920 (N_17920,N_14907,N_14658);
xnor U17921 (N_17921,N_15387,N_15017);
xnor U17922 (N_17922,N_15172,N_14457);
xnor U17923 (N_17923,N_14827,N_15983);
and U17924 (N_17924,N_14217,N_14049);
or U17925 (N_17925,N_14594,N_15236);
or U17926 (N_17926,N_14502,N_15512);
or U17927 (N_17927,N_14578,N_15101);
or U17928 (N_17928,N_15212,N_15856);
xnor U17929 (N_17929,N_15267,N_14743);
xnor U17930 (N_17930,N_14443,N_14327);
xnor U17931 (N_17931,N_14490,N_15893);
xor U17932 (N_17932,N_15712,N_14784);
nor U17933 (N_17933,N_14554,N_14974);
nand U17934 (N_17934,N_14800,N_15072);
nor U17935 (N_17935,N_15346,N_14744);
xor U17936 (N_17936,N_14054,N_14431);
or U17937 (N_17937,N_14864,N_14202);
nor U17938 (N_17938,N_14352,N_15698);
nor U17939 (N_17939,N_14564,N_14963);
nand U17940 (N_17940,N_14856,N_15144);
or U17941 (N_17941,N_14105,N_15127);
xnor U17942 (N_17942,N_15063,N_15645);
nand U17943 (N_17943,N_15493,N_14565);
and U17944 (N_17944,N_14623,N_15868);
nand U17945 (N_17945,N_14563,N_15761);
nor U17946 (N_17946,N_15313,N_14154);
xor U17947 (N_17947,N_14406,N_14293);
nor U17948 (N_17948,N_14309,N_15985);
nand U17949 (N_17949,N_14850,N_14503);
and U17950 (N_17950,N_14708,N_14729);
and U17951 (N_17951,N_15984,N_14129);
nor U17952 (N_17952,N_15039,N_15286);
nor U17953 (N_17953,N_14464,N_15572);
or U17954 (N_17954,N_14077,N_15254);
and U17955 (N_17955,N_14567,N_14742);
xnor U17956 (N_17956,N_14452,N_15252);
or U17957 (N_17957,N_15273,N_14244);
and U17958 (N_17958,N_15582,N_14689);
nand U17959 (N_17959,N_15810,N_15712);
nand U17960 (N_17960,N_14972,N_14270);
and U17961 (N_17961,N_14401,N_14515);
xnor U17962 (N_17962,N_14552,N_15606);
nand U17963 (N_17963,N_15023,N_15326);
nor U17964 (N_17964,N_14883,N_14975);
nand U17965 (N_17965,N_14503,N_15521);
nand U17966 (N_17966,N_14295,N_15278);
and U17967 (N_17967,N_14168,N_15904);
nor U17968 (N_17968,N_15470,N_14747);
nor U17969 (N_17969,N_15563,N_14822);
or U17970 (N_17970,N_14667,N_15503);
or U17971 (N_17971,N_15443,N_15581);
xnor U17972 (N_17972,N_15021,N_14953);
or U17973 (N_17973,N_14608,N_14544);
or U17974 (N_17974,N_15560,N_15930);
or U17975 (N_17975,N_14996,N_14455);
and U17976 (N_17976,N_14283,N_15952);
or U17977 (N_17977,N_14514,N_14304);
and U17978 (N_17978,N_15827,N_14427);
and U17979 (N_17979,N_15208,N_15171);
xnor U17980 (N_17980,N_14802,N_15792);
or U17981 (N_17981,N_14247,N_14794);
or U17982 (N_17982,N_15161,N_15765);
nand U17983 (N_17983,N_15733,N_15331);
nand U17984 (N_17984,N_14305,N_14934);
nor U17985 (N_17985,N_15560,N_15445);
and U17986 (N_17986,N_15416,N_14544);
and U17987 (N_17987,N_15506,N_15171);
nand U17988 (N_17988,N_15834,N_14358);
nand U17989 (N_17989,N_15297,N_14661);
nor U17990 (N_17990,N_14071,N_14420);
nor U17991 (N_17991,N_14934,N_15915);
nand U17992 (N_17992,N_15406,N_14801);
nor U17993 (N_17993,N_14908,N_14003);
nor U17994 (N_17994,N_14866,N_15286);
and U17995 (N_17995,N_14049,N_14271);
and U17996 (N_17996,N_14053,N_15892);
nor U17997 (N_17997,N_15087,N_15912);
and U17998 (N_17998,N_15311,N_15715);
nand U17999 (N_17999,N_15791,N_14763);
xnor U18000 (N_18000,N_17897,N_17640);
and U18001 (N_18001,N_16271,N_17941);
nand U18002 (N_18002,N_16182,N_16969);
nand U18003 (N_18003,N_17929,N_16562);
nand U18004 (N_18004,N_16061,N_17704);
or U18005 (N_18005,N_16167,N_17826);
nor U18006 (N_18006,N_16783,N_17931);
and U18007 (N_18007,N_17273,N_16942);
or U18008 (N_18008,N_16581,N_17377);
nand U18009 (N_18009,N_16899,N_16183);
and U18010 (N_18010,N_16914,N_17946);
nor U18011 (N_18011,N_16999,N_16707);
and U18012 (N_18012,N_16029,N_17658);
or U18013 (N_18013,N_17587,N_16095);
nand U18014 (N_18014,N_16115,N_17042);
nand U18015 (N_18015,N_16127,N_16666);
and U18016 (N_18016,N_16349,N_16203);
nand U18017 (N_18017,N_17951,N_16146);
nand U18018 (N_18018,N_16096,N_16794);
nor U18019 (N_18019,N_17454,N_16173);
nand U18020 (N_18020,N_17609,N_16134);
nand U18021 (N_18021,N_17348,N_17051);
and U18022 (N_18022,N_16943,N_16032);
xnor U18023 (N_18023,N_16194,N_16690);
xor U18024 (N_18024,N_17800,N_17473);
and U18025 (N_18025,N_17821,N_17438);
nand U18026 (N_18026,N_17763,N_16576);
xnor U18027 (N_18027,N_16499,N_17794);
xnor U18028 (N_18028,N_16864,N_16121);
nand U18029 (N_18029,N_16320,N_17329);
xnor U18030 (N_18030,N_17870,N_16423);
nand U18031 (N_18031,N_16250,N_16429);
and U18032 (N_18032,N_16900,N_17391);
nor U18033 (N_18033,N_17521,N_16829);
nand U18034 (N_18034,N_17030,N_16521);
and U18035 (N_18035,N_17410,N_17109);
xnor U18036 (N_18036,N_16972,N_16290);
and U18037 (N_18037,N_17338,N_16059);
and U18038 (N_18038,N_16445,N_16491);
nor U18039 (N_18039,N_16923,N_16520);
nor U18040 (N_18040,N_16856,N_16820);
nor U18041 (N_18041,N_16910,N_16426);
or U18042 (N_18042,N_17633,N_17207);
nor U18043 (N_18043,N_17044,N_17328);
nand U18044 (N_18044,N_16515,N_17599);
nor U18045 (N_18045,N_16201,N_16650);
and U18046 (N_18046,N_16225,N_17049);
and U18047 (N_18047,N_17557,N_16800);
xor U18048 (N_18048,N_16327,N_17646);
nor U18049 (N_18049,N_16427,N_16138);
nand U18050 (N_18050,N_16075,N_16967);
xnor U18051 (N_18051,N_16083,N_16477);
nor U18052 (N_18052,N_17776,N_17107);
nand U18053 (N_18053,N_17515,N_16307);
nor U18054 (N_18054,N_16441,N_17425);
xnor U18055 (N_18055,N_17114,N_16585);
nor U18056 (N_18056,N_17606,N_17072);
or U18057 (N_18057,N_17604,N_17039);
nor U18058 (N_18058,N_17225,N_17289);
or U18059 (N_18059,N_17229,N_16689);
xnor U18060 (N_18060,N_16510,N_17472);
nor U18061 (N_18061,N_16443,N_16681);
and U18062 (N_18062,N_16781,N_17086);
and U18063 (N_18063,N_16645,N_16362);
xnor U18064 (N_18064,N_16335,N_17743);
nand U18065 (N_18065,N_17091,N_17517);
or U18066 (N_18066,N_16748,N_16459);
nor U18067 (N_18067,N_17055,N_16212);
nand U18068 (N_18068,N_16231,N_17943);
nand U18069 (N_18069,N_16209,N_16816);
or U18070 (N_18070,N_16079,N_17475);
nor U18071 (N_18071,N_16357,N_16547);
nand U18072 (N_18072,N_16657,N_17519);
nor U18073 (N_18073,N_16740,N_17296);
and U18074 (N_18074,N_16574,N_16922);
and U18075 (N_18075,N_17585,N_16436);
and U18076 (N_18076,N_16980,N_16221);
or U18077 (N_18077,N_16934,N_16081);
nor U18078 (N_18078,N_17257,N_16695);
or U18079 (N_18079,N_16044,N_17742);
and U18080 (N_18080,N_17195,N_16260);
or U18081 (N_18081,N_16698,N_17550);
or U18082 (N_18082,N_17902,N_17128);
and U18083 (N_18083,N_17908,N_16070);
nor U18084 (N_18084,N_17638,N_17026);
and U18085 (N_18085,N_17809,N_17436);
xor U18086 (N_18086,N_16808,N_17428);
and U18087 (N_18087,N_17570,N_17427);
nand U18088 (N_18088,N_16544,N_17932);
xor U18089 (N_18089,N_16987,N_16045);
nor U18090 (N_18090,N_16950,N_16964);
and U18091 (N_18091,N_16446,N_16289);
or U18092 (N_18092,N_17735,N_17863);
xnor U18093 (N_18093,N_17234,N_16570);
nand U18094 (N_18094,N_17379,N_16909);
and U18095 (N_18095,N_16177,N_16315);
nand U18096 (N_18096,N_17967,N_16814);
and U18097 (N_18097,N_16502,N_17505);
xnor U18098 (N_18098,N_16028,N_17452);
nor U18099 (N_18099,N_16749,N_16918);
nor U18100 (N_18100,N_16546,N_16019);
and U18101 (N_18101,N_16085,N_17303);
or U18102 (N_18102,N_17240,N_17381);
nor U18103 (N_18103,N_16541,N_17441);
and U18104 (N_18104,N_17202,N_17823);
or U18105 (N_18105,N_17656,N_16911);
xnor U18106 (N_18106,N_17966,N_17621);
xor U18107 (N_18107,N_17484,N_16148);
nor U18108 (N_18108,N_16118,N_17117);
nand U18109 (N_18109,N_16669,N_16283);
xnor U18110 (N_18110,N_16471,N_16355);
nor U18111 (N_18111,N_17260,N_16697);
nand U18112 (N_18112,N_17092,N_17615);
xor U18113 (N_18113,N_17050,N_17074);
and U18114 (N_18114,N_17261,N_17188);
xnor U18115 (N_18115,N_16052,N_17817);
and U18116 (N_18116,N_16543,N_17486);
or U18117 (N_18117,N_17525,N_16421);
or U18118 (N_18118,N_17998,N_16601);
nor U18119 (N_18119,N_17458,N_17488);
or U18120 (N_18120,N_17703,N_17903);
xor U18121 (N_18121,N_16178,N_17835);
or U18122 (N_18122,N_17770,N_16878);
or U18123 (N_18123,N_16094,N_17362);
nor U18124 (N_18124,N_16065,N_16852);
nand U18125 (N_18125,N_16640,N_17474);
xnor U18126 (N_18126,N_17737,N_16586);
xnor U18127 (N_18127,N_16353,N_17035);
nand U18128 (N_18128,N_17579,N_16824);
xor U18129 (N_18129,N_16568,N_17244);
nand U18130 (N_18130,N_17022,N_17663);
or U18131 (N_18131,N_16876,N_17090);
and U18132 (N_18132,N_17674,N_16853);
or U18133 (N_18133,N_16235,N_16265);
nor U18134 (N_18134,N_17311,N_16336);
and U18135 (N_18135,N_16627,N_16005);
nor U18136 (N_18136,N_17204,N_17695);
nand U18137 (N_18137,N_17740,N_17848);
nor U18138 (N_18138,N_16830,N_16886);
nand U18139 (N_18139,N_17802,N_17773);
nor U18140 (N_18140,N_17463,N_16993);
and U18141 (N_18141,N_16747,N_17088);
and U18142 (N_18142,N_17972,N_16855);
and U18143 (N_18143,N_16912,N_17720);
nand U18144 (N_18144,N_17561,N_16036);
nand U18145 (N_18145,N_16930,N_17336);
or U18146 (N_18146,N_17219,N_17275);
xor U18147 (N_18147,N_17968,N_17673);
or U18148 (N_18148,N_17567,N_16385);
and U18149 (N_18149,N_16461,N_16483);
xnor U18150 (N_18150,N_16533,N_17723);
nand U18151 (N_18151,N_17098,N_16742);
and U18152 (N_18152,N_17408,N_16206);
and U18153 (N_18153,N_17143,N_16060);
nor U18154 (N_18154,N_16835,N_17918);
or U18155 (N_18155,N_17272,N_17324);
nor U18156 (N_18156,N_16920,N_17165);
nor U18157 (N_18157,N_16957,N_17891);
and U18158 (N_18158,N_16826,N_17559);
xnor U18159 (N_18159,N_17100,N_17191);
and U18160 (N_18160,N_17359,N_17795);
nand U18161 (N_18161,N_17464,N_17502);
or U18162 (N_18162,N_16647,N_16646);
xor U18163 (N_18163,N_17971,N_16376);
or U18164 (N_18164,N_16442,N_17641);
or U18165 (N_18165,N_17015,N_17584);
nand U18166 (N_18166,N_17357,N_17767);
nand U18167 (N_18167,N_17335,N_17712);
nor U18168 (N_18168,N_17524,N_16129);
xnor U18169 (N_18169,N_16809,N_16303);
xor U18170 (N_18170,N_17290,N_17440);
nor U18171 (N_18171,N_17651,N_17546);
nor U18172 (N_18172,N_16846,N_17622);
and U18173 (N_18173,N_17262,N_16825);
nor U18174 (N_18174,N_17144,N_17649);
xor U18175 (N_18175,N_17888,N_17268);
or U18176 (N_18176,N_17554,N_17672);
xor U18177 (N_18177,N_16220,N_16174);
xnor U18178 (N_18178,N_17819,N_16370);
and U18179 (N_18179,N_16453,N_16166);
and U18180 (N_18180,N_16435,N_16014);
and U18181 (N_18181,N_16602,N_16885);
and U18182 (N_18182,N_16831,N_16259);
and U18183 (N_18183,N_17744,N_17405);
xor U18184 (N_18184,N_16401,N_17980);
and U18185 (N_18185,N_16078,N_16311);
or U18186 (N_18186,N_16251,N_17875);
nand U18187 (N_18187,N_16149,N_17116);
xnor U18188 (N_18188,N_16895,N_17416);
xnor U18189 (N_18189,N_16838,N_16295);
xor U18190 (N_18190,N_17921,N_17157);
xnor U18191 (N_18191,N_17243,N_16088);
nand U18192 (N_18192,N_17062,N_16536);
nor U18193 (N_18193,N_16190,N_17730);
nand U18194 (N_18194,N_17677,N_17361);
xnor U18195 (N_18195,N_16230,N_16733);
nand U18196 (N_18196,N_16551,N_16268);
or U18197 (N_18197,N_16252,N_16264);
xor U18198 (N_18198,N_16122,N_16237);
xor U18199 (N_18199,N_17294,N_17893);
nand U18200 (N_18200,N_17302,N_16055);
nor U18201 (N_18201,N_17246,N_16263);
nand U18202 (N_18202,N_17644,N_17779);
nand U18203 (N_18203,N_17937,N_16609);
nor U18204 (N_18204,N_16978,N_16765);
nor U18205 (N_18205,N_16434,N_16309);
nand U18206 (N_18206,N_16915,N_16764);
and U18207 (N_18207,N_17104,N_17686);
or U18208 (N_18208,N_17571,N_16539);
xor U18209 (N_18209,N_17685,N_17129);
or U18210 (N_18210,N_16891,N_16185);
nor U18211 (N_18211,N_16953,N_16973);
nand U18212 (N_18212,N_16236,N_16484);
xor U18213 (N_18213,N_17755,N_17215);
nand U18214 (N_18214,N_17564,N_16365);
nor U18215 (N_18215,N_16960,N_17386);
nor U18216 (N_18216,N_16628,N_17661);
or U18217 (N_18217,N_17719,N_16926);
nand U18218 (N_18218,N_16956,N_17748);
and U18219 (N_18219,N_16242,N_16804);
nand U18220 (N_18220,N_16058,N_16106);
xor U18221 (N_18221,N_16929,N_17083);
or U18222 (N_18222,N_17426,N_16001);
and U18223 (N_18223,N_16590,N_16273);
nand U18224 (N_18224,N_17269,N_17200);
or U18225 (N_18225,N_17983,N_17601);
xnor U18226 (N_18226,N_16992,N_17317);
nand U18227 (N_18227,N_16247,N_17699);
and U18228 (N_18228,N_17807,N_17176);
nor U18229 (N_18229,N_17565,N_17993);
or U18230 (N_18230,N_17510,N_17043);
xnor U18231 (N_18231,N_17694,N_16187);
nor U18232 (N_18232,N_16888,N_16111);
and U18233 (N_18233,N_16965,N_16821);
xnor U18234 (N_18234,N_16977,N_17683);
nor U18235 (N_18235,N_16879,N_16540);
xor U18236 (N_18236,N_17407,N_17247);
nand U18237 (N_18237,N_16812,N_16479);
nand U18238 (N_18238,N_17803,N_17006);
xor U18239 (N_18239,N_17276,N_16974);
nand U18240 (N_18240,N_16644,N_17864);
xor U18241 (N_18241,N_17801,N_16866);
or U18242 (N_18242,N_17681,N_17716);
or U18243 (N_18243,N_17616,N_16205);
xor U18244 (N_18244,N_17798,N_16680);
nor U18245 (N_18245,N_16976,N_17608);
nand U18246 (N_18246,N_17171,N_17047);
or U18247 (N_18247,N_17470,N_17852);
xnor U18248 (N_18248,N_16352,N_16700);
xnor U18249 (N_18249,N_17053,N_16715);
nor U18250 (N_18250,N_17105,N_16169);
or U18251 (N_18251,N_17960,N_17825);
xor U18252 (N_18252,N_17024,N_17182);
and U18253 (N_18253,N_17232,N_17374);
and U18254 (N_18254,N_17534,N_16908);
or U18255 (N_18255,N_16347,N_17871);
nand U18256 (N_18256,N_16392,N_17836);
nand U18257 (N_18257,N_17064,N_16388);
xor U18258 (N_18258,N_16391,N_17493);
nor U18259 (N_18259,N_17827,N_16306);
and U18260 (N_18260,N_16898,N_17617);
nand U18261 (N_18261,N_17573,N_17040);
xnor U18262 (N_18262,N_17990,N_17366);
nor U18263 (N_18263,N_16282,N_17877);
and U18264 (N_18264,N_16982,N_16020);
and U18265 (N_18265,N_17248,N_17859);
nand U18266 (N_18266,N_16501,N_16009);
or U18267 (N_18267,N_16329,N_17976);
and U18268 (N_18268,N_16319,N_17081);
nand U18269 (N_18269,N_16189,N_17293);
nor U18270 (N_18270,N_16763,N_16266);
and U18271 (N_18271,N_17745,N_16648);
xnor U18272 (N_18272,N_16418,N_17793);
nand U18273 (N_18273,N_16463,N_17805);
and U18274 (N_18274,N_17696,N_17964);
and U18275 (N_18275,N_16858,N_17206);
nand U18276 (N_18276,N_16193,N_16507);
or U18277 (N_18277,N_16041,N_17485);
nor U18278 (N_18278,N_16373,N_17291);
xor U18279 (N_18279,N_16968,N_17873);
or U18280 (N_18280,N_17751,N_16276);
nor U18281 (N_18281,N_17340,N_17715);
nand U18282 (N_18282,N_16017,N_17370);
and U18283 (N_18283,N_17368,N_16727);
nand U18284 (N_18284,N_17907,N_16023);
or U18285 (N_18285,N_16344,N_16007);
and U18286 (N_18286,N_17659,N_17156);
and U18287 (N_18287,N_17757,N_17079);
nand U18288 (N_18288,N_17533,N_17230);
nand U18289 (N_18289,N_16619,N_16678);
nand U18290 (N_18290,N_16513,N_16057);
or U18291 (N_18291,N_17245,N_16525);
nand U18292 (N_18292,N_16971,N_16608);
or U18293 (N_18293,N_17196,N_16916);
nor U18294 (N_18294,N_16589,N_16795);
nor U18295 (N_18295,N_16424,N_17738);
nor U18296 (N_18296,N_17791,N_16120);
xor U18297 (N_18297,N_17433,N_17691);
or U18298 (N_18298,N_16863,N_17216);
and U18299 (N_18299,N_16313,N_17319);
nor U18300 (N_18300,N_16304,N_16519);
and U18301 (N_18301,N_17347,N_17162);
nor U18302 (N_18302,N_17306,N_17523);
xor U18303 (N_18303,N_16232,N_16840);
nor U18304 (N_18304,N_16072,N_16557);
nand U18305 (N_18305,N_16626,N_16258);
nor U18306 (N_18306,N_16766,N_17160);
or U18307 (N_18307,N_16383,N_17503);
nor U18308 (N_18308,N_17724,N_17400);
or U18309 (N_18309,N_17671,N_16667);
or U18310 (N_18310,N_16517,N_16124);
xor U18311 (N_18311,N_16696,N_16701);
or U18312 (N_18312,N_17434,N_16013);
and U18313 (N_18313,N_16197,N_17896);
and U18314 (N_18314,N_17457,N_16762);
and U18315 (N_18315,N_17001,N_17278);
nor U18316 (N_18316,N_16310,N_17045);
nand U18317 (N_18317,N_16786,N_16208);
nand U18318 (N_18318,N_16719,N_17477);
or U18319 (N_18319,N_17986,N_16726);
or U18320 (N_18320,N_16716,N_17167);
and U18321 (N_18321,N_16538,N_17183);
xnor U18322 (N_18322,N_17483,N_17149);
and U18323 (N_18323,N_17313,N_17890);
or U18324 (N_18324,N_17298,N_16687);
xnor U18325 (N_18325,N_16822,N_16234);
xnor U18326 (N_18326,N_17342,N_16567);
xnor U18327 (N_18327,N_16255,N_17654);
or U18328 (N_18328,N_17238,N_16529);
or U18329 (N_18329,N_17163,N_16569);
and U18330 (N_18330,N_17529,N_17297);
nor U18331 (N_18331,N_16508,N_16101);
nor U18332 (N_18332,N_16112,N_16358);
xor U18333 (N_18333,N_16622,N_17526);
or U18334 (N_18334,N_16610,N_17038);
and U18335 (N_18335,N_17004,N_16163);
xor U18336 (N_18336,N_17623,N_16312);
nor U18337 (N_18337,N_16287,N_17729);
xor U18338 (N_18338,N_16556,N_17938);
nor U18339 (N_18339,N_16334,N_17936);
or U18340 (N_18340,N_16818,N_16071);
and U18341 (N_18341,N_17127,N_17012);
and U18342 (N_18342,N_16805,N_17912);
or U18343 (N_18343,N_17664,N_17372);
and U18344 (N_18344,N_17507,N_17125);
and U18345 (N_18345,N_16518,N_17613);
and U18346 (N_18346,N_17097,N_16431);
xor U18347 (N_18347,N_17762,N_16559);
nor U18348 (N_18348,N_17070,N_17684);
nand U18349 (N_18349,N_17249,N_17520);
and U18350 (N_18350,N_16555,N_17713);
xnor U18351 (N_18351,N_16514,N_16743);
or U18352 (N_18352,N_17145,N_17430);
nor U18353 (N_18353,N_16847,N_16571);
or U18354 (N_18354,N_16995,N_16654);
xnor U18355 (N_18355,N_17048,N_16870);
xnor U18356 (N_18356,N_16191,N_17333);
nor U18357 (N_18357,N_17179,N_16985);
xnor U18358 (N_18358,N_16789,N_17996);
xor U18359 (N_18359,N_17708,N_17089);
or U18360 (N_18360,N_16988,N_17997);
nand U18361 (N_18361,N_16278,N_17446);
nand U18362 (N_18362,N_16343,N_16175);
xnor U18363 (N_18363,N_17023,N_17810);
nand U18364 (N_18364,N_16940,N_16170);
and U18365 (N_18365,N_17978,N_17420);
xnor U18366 (N_18366,N_16298,N_16371);
and U18367 (N_18367,N_17192,N_17542);
and U18368 (N_18368,N_17197,N_16296);
or U18369 (N_18369,N_17634,N_16474);
xnor U18370 (N_18370,N_17963,N_16238);
nand U18371 (N_18371,N_17292,N_16649);
and U18372 (N_18372,N_17989,N_17108);
or U18373 (N_18373,N_17789,N_16450);
or U18374 (N_18374,N_16425,N_16389);
nor U18375 (N_18375,N_17242,N_17185);
or U18376 (N_18376,N_16767,N_17718);
xnor U18377 (N_18377,N_17412,N_17222);
or U18378 (N_18378,N_17282,N_16399);
or U18379 (N_18379,N_16475,N_17679);
or U18380 (N_18380,N_16887,N_17749);
nor U18381 (N_18381,N_17414,N_17847);
xnor U18382 (N_18382,N_17203,N_17669);
nor U18383 (N_18383,N_17544,N_16535);
and U18384 (N_18384,N_17843,N_17205);
nor U18385 (N_18385,N_17828,N_16369);
nand U18386 (N_18386,N_16164,N_16758);
nand U18387 (N_18387,N_16277,N_16500);
nor U18388 (N_18388,N_17168,N_16051);
nor U18389 (N_18389,N_16098,N_17259);
nor U18390 (N_18390,N_16668,N_17665);
nor U18391 (N_18391,N_16958,N_17027);
nor U18392 (N_18392,N_17581,N_17769);
nand U18393 (N_18393,N_16933,N_17594);
nand U18394 (N_18394,N_16472,N_17459);
nor U18395 (N_18395,N_17310,N_17949);
or U18396 (N_18396,N_17194,N_16834);
nor U18397 (N_18397,N_17625,N_17865);
nand U18398 (N_18398,N_17563,N_17849);
nand U18399 (N_18399,N_17031,N_17432);
xnor U18400 (N_18400,N_16410,N_16093);
nor U18401 (N_18401,N_17214,N_16262);
and U18402 (N_18402,N_16851,N_16875);
nor U18403 (N_18403,N_17142,N_16400);
xor U18404 (N_18404,N_16738,N_16492);
and U18405 (N_18405,N_16975,N_16125);
and U18406 (N_18406,N_17676,N_16135);
or U18407 (N_18407,N_16759,N_16854);
nand U18408 (N_18408,N_17487,N_16359);
nor U18409 (N_18409,N_16222,N_17159);
nand U18410 (N_18410,N_16086,N_16302);
nor U18411 (N_18411,N_16114,N_16186);
and U18412 (N_18412,N_17326,N_17538);
and U18413 (N_18413,N_17878,N_17256);
and U18414 (N_18414,N_17288,N_17147);
and U18415 (N_18415,N_17841,N_17566);
nand U18416 (N_18416,N_16248,N_16677);
xor U18417 (N_18417,N_16021,N_16843);
or U18418 (N_18418,N_16490,N_16606);
xor U18419 (N_18419,N_17330,N_17726);
xnor U18420 (N_18420,N_17777,N_16880);
nand U18421 (N_18421,N_17648,N_17151);
nand U18422 (N_18422,N_17753,N_16054);
nor U18423 (N_18423,N_16006,N_16997);
xor U18424 (N_18424,N_17845,N_17768);
xnor U18425 (N_18425,N_16375,N_17632);
nor U18426 (N_18426,N_16324,N_16671);
or U18427 (N_18427,N_16643,N_16092);
xnor U18428 (N_18428,N_17279,N_16048);
nor U18429 (N_18429,N_16300,N_16670);
xnor U18430 (N_18430,N_16746,N_16550);
xor U18431 (N_18431,N_16133,N_17066);
and U18432 (N_18432,N_16367,N_17922);
and U18433 (N_18433,N_16025,N_17385);
xor U18434 (N_18434,N_17332,N_16600);
nor U18435 (N_18435,N_17073,N_16548);
nor U18436 (N_18436,N_17401,N_16254);
and U18437 (N_18437,N_17255,N_16464);
xor U18438 (N_18438,N_16105,N_16188);
nand U18439 (N_18439,N_17346,N_16040);
and U18440 (N_18440,N_17857,N_17384);
and U18441 (N_18441,N_17509,N_16614);
xnor U18442 (N_18442,N_16892,N_17312);
nor U18443 (N_18443,N_17363,N_17591);
xor U18444 (N_18444,N_17955,N_16480);
nand U18445 (N_18445,N_17115,N_17036);
or U18446 (N_18446,N_16323,N_16952);
nand U18447 (N_18447,N_17861,N_16346);
xor U18448 (N_18448,N_16214,N_17508);
xor U18449 (N_18449,N_17620,N_17842);
or U18450 (N_18450,N_16503,N_16223);
nor U18451 (N_18451,N_17500,N_17927);
or U18452 (N_18452,N_17668,N_16396);
or U18453 (N_18453,N_16598,N_16793);
or U18454 (N_18454,N_17781,N_17834);
or U18455 (N_18455,N_16489,N_16485);
or U18456 (N_18456,N_16176,N_16274);
or U18457 (N_18457,N_17547,N_17506);
and U18458 (N_18458,N_17187,N_16928);
xnor U18459 (N_18459,N_17226,N_17513);
or U18460 (N_18460,N_16414,N_17266);
nor U18461 (N_18461,N_17380,N_17135);
nand U18462 (N_18462,N_16945,N_16713);
or U18463 (N_18463,N_17899,N_17975);
and U18464 (N_18464,N_17184,N_16631);
nor U18465 (N_18465,N_16356,N_17812);
or U18466 (N_18466,N_17924,N_16416);
or U18467 (N_18467,N_16473,N_16239);
nor U18468 (N_18468,N_16000,N_17132);
and U18469 (N_18469,N_16184,N_17840);
nor U18470 (N_18470,N_17909,N_16635);
nand U18471 (N_18471,N_16228,N_16970);
nand U18472 (N_18472,N_17406,N_16168);
and U18473 (N_18473,N_16338,N_16419);
or U18474 (N_18474,N_16452,N_17928);
nand U18475 (N_18475,N_16049,N_16145);
xor U18476 (N_18476,N_16596,N_16718);
or U18477 (N_18477,N_17422,N_16382);
and U18478 (N_18478,N_16267,N_17046);
or U18479 (N_18479,N_16582,N_16703);
nor U18480 (N_18480,N_17754,N_17450);
and U18481 (N_18481,N_17121,N_17732);
or U18482 (N_18482,N_16150,N_16785);
and U18483 (N_18483,N_16224,N_16617);
or U18484 (N_18484,N_16159,N_16776);
and U18485 (N_18485,N_17356,N_16314);
xnor U18486 (N_18486,N_16043,N_16871);
xor U18487 (N_18487,N_16679,N_17830);
xor U18488 (N_18488,N_17378,N_17939);
nor U18489 (N_18489,N_16011,N_17619);
nor U18490 (N_18490,N_16552,N_17592);
nand U18491 (N_18491,N_16566,N_17228);
and U18492 (N_18492,N_17233,N_17037);
nand U18493 (N_18493,N_17977,N_16417);
xnor U18494 (N_18494,N_17596,N_17783);
and U18495 (N_18495,N_17501,N_16637);
and U18496 (N_18496,N_17876,N_16415);
or U18497 (N_18497,N_17467,N_16074);
xor U18498 (N_18498,N_17448,N_17131);
nand U18499 (N_18499,N_16069,N_16272);
nor U18500 (N_18500,N_16849,N_16279);
or U18501 (N_18501,N_17979,N_16097);
nor U18502 (N_18502,N_17423,N_17411);
xnor U18503 (N_18503,N_17627,N_17637);
and U18504 (N_18504,N_16398,N_16522);
or U18505 (N_18505,N_16994,N_17702);
nand U18506 (N_18506,N_17688,N_17479);
xor U18507 (N_18507,N_17575,N_17223);
and U18508 (N_18508,N_17041,N_17920);
xor U18509 (N_18509,N_17879,N_17869);
nor U18510 (N_18510,N_17321,N_16760);
nor U18511 (N_18511,N_16516,N_17058);
nand U18512 (N_18512,N_16297,N_17439);
xor U18513 (N_18513,N_17148,N_17667);
and U18514 (N_18514,N_17007,N_16592);
nor U18515 (N_18515,N_17421,N_16883);
and U18516 (N_18516,N_17786,N_17140);
xnor U18517 (N_18517,N_17172,N_17021);
nor U18518 (N_18518,N_16653,N_17431);
nor U18519 (N_18519,N_16126,N_16673);
and U18520 (N_18520,N_16877,N_17253);
and U18521 (N_18521,N_17019,N_16665);
nor U18522 (N_18522,N_16844,N_16575);
xnor U18523 (N_18523,N_16599,N_17065);
nand U18524 (N_18524,N_16745,N_16664);
nor U18525 (N_18525,N_17945,N_17522);
xor U18526 (N_18526,N_16087,N_17782);
nor U18527 (N_18527,N_16691,N_17258);
nand U18528 (N_18528,N_16868,N_17898);
or U18529 (N_18529,N_17052,N_16064);
xnor U18530 (N_18530,N_16076,N_16583);
nand U18531 (N_18531,N_17806,N_16845);
nand U18532 (N_18532,N_17605,N_17154);
nor U18533 (N_18533,N_16813,N_17106);
and U18534 (N_18534,N_16090,N_16882);
nand U18535 (N_18535,N_17492,N_16534);
nand U18536 (N_18536,N_17352,N_16153);
or U18537 (N_18537,N_16636,N_17224);
and U18538 (N_18538,N_17833,N_17059);
nand U18539 (N_18539,N_17752,N_16941);
nand U18540 (N_18540,N_17209,N_16113);
or U18541 (N_18541,N_17299,N_16100);
and U18542 (N_18542,N_17598,N_16996);
and U18543 (N_18543,N_16739,N_16066);
or U18544 (N_18544,N_16406,N_16806);
nand U18545 (N_18545,N_16591,N_17137);
xnor U18546 (N_18546,N_17150,N_17080);
nand U18547 (N_18547,N_16428,N_17078);
xnor U18548 (N_18548,N_17111,N_17120);
nand U18549 (N_18549,N_16872,N_16897);
and U18550 (N_18550,N_17170,N_16741);
and U18551 (N_18551,N_17787,N_17974);
nor U18552 (N_18552,N_16595,N_16867);
and U18553 (N_18553,N_16067,N_16004);
xor U18554 (N_18554,N_17771,N_17103);
nor U18555 (N_18555,N_17905,N_17655);
nand U18556 (N_18556,N_17014,N_17543);
and U18557 (N_18557,N_16366,N_17250);
xnor U18558 (N_18558,N_16339,N_17495);
or U18559 (N_18559,N_17901,N_17445);
nand U18560 (N_18560,N_16778,N_16938);
xnor U18561 (N_18561,N_16345,N_16889);
xnor U18562 (N_18562,N_17466,N_17832);
and U18563 (N_18563,N_16661,N_16931);
or U18564 (N_18564,N_17327,N_17884);
nor U18565 (N_18565,N_17758,N_16299);
nand U18566 (N_18566,N_17076,N_17540);
xor U18567 (N_18567,N_17295,N_16815);
and U18568 (N_18568,N_17476,N_16913);
and U18569 (N_18569,N_16142,N_17271);
nor U18570 (N_18570,N_16374,N_17856);
nand U18571 (N_18571,N_16465,N_16954);
and U18572 (N_18572,N_17588,N_16672);
nand U18573 (N_18573,N_16629,N_17610);
or U18574 (N_18574,N_16245,N_17734);
xor U18575 (N_18575,N_17532,N_16951);
nor U18576 (N_18576,N_16839,N_16213);
or U18577 (N_18577,N_17639,N_16607);
nor U18578 (N_18578,N_17101,N_16102);
nand U18579 (N_18579,N_16476,N_17186);
and U18580 (N_18580,N_17175,N_17280);
nand U18581 (N_18581,N_16340,N_17947);
and U18582 (N_18582,N_16444,N_16448);
nand U18583 (N_18583,N_17071,N_17398);
or U18584 (N_18584,N_17322,N_17496);
and U18585 (N_18585,N_17136,N_16342);
or U18586 (N_18586,N_17988,N_17636);
nor U18587 (N_18587,N_16998,N_17491);
nand U18588 (N_18588,N_17697,N_17213);
nand U18589 (N_18589,N_17320,N_16243);
xor U18590 (N_18590,N_17872,N_16896);
nand U18591 (N_18591,N_16348,N_17429);
nor U18592 (N_18592,N_16147,N_16862);
xor U18593 (N_18593,N_17662,N_16010);
xnor U18594 (N_18594,N_16906,N_17831);
nand U18595 (N_18595,N_17722,N_16561);
or U18596 (N_18596,N_16901,N_17536);
and U18597 (N_18597,N_17747,N_16615);
and U18598 (N_18598,N_16732,N_17814);
nor U18599 (N_18599,N_16432,N_17887);
or U18600 (N_18600,N_16210,N_17531);
and U18601 (N_18601,N_16381,N_16317);
nand U18602 (N_18602,N_16724,N_16046);
or U18603 (N_18603,N_16409,N_17548);
xor U18604 (N_18604,N_16717,N_16683);
and U18605 (N_18605,N_16038,N_16939);
nand U18606 (N_18606,N_16439,N_17714);
and U18607 (N_18607,N_17480,N_16171);
nand U18608 (N_18608,N_17308,N_17285);
or U18609 (N_18609,N_16154,N_17323);
nor U18610 (N_18610,N_16621,N_17054);
xnor U18611 (N_18611,N_17460,N_16162);
nand U18612 (N_18612,N_16755,N_17958);
nand U18613 (N_18613,N_17389,N_16705);
nand U18614 (N_18614,N_16368,N_17300);
nor U18615 (N_18615,N_17895,N_16777);
nor U18616 (N_18616,N_16280,N_17528);
and U18617 (N_18617,N_17415,N_16291);
xor U18618 (N_18618,N_16156,N_16630);
and U18619 (N_18619,N_16903,N_17647);
and U18620 (N_18620,N_17815,N_16116);
xnor U18621 (N_18621,N_17837,N_16597);
nand U18622 (N_18622,N_16620,N_16305);
or U18623 (N_18623,N_17717,N_17766);
or U18624 (N_18624,N_16729,N_16641);
or U18625 (N_18625,N_16402,N_16395);
and U18626 (N_18626,N_17451,N_17611);
or U18627 (N_18627,N_17727,N_17478);
nor U18628 (N_18628,N_16685,N_16241);
nand U18629 (N_18629,N_16848,N_17822);
or U18630 (N_18630,N_17701,N_16658);
nor U18631 (N_18631,N_16580,N_16377);
xor U18632 (N_18632,N_17449,N_16350);
or U18633 (N_18633,N_16486,N_17930);
or U18634 (N_18634,N_16157,N_17537);
and U18635 (N_18635,N_17553,N_17444);
nor U18636 (N_18636,N_17545,N_17095);
nand U18637 (N_18637,N_16321,N_17874);
nor U18638 (N_18638,N_17746,N_17995);
and U18639 (N_18639,N_16857,N_17469);
or U18640 (N_18640,N_17511,N_17482);
xnor U18641 (N_18641,N_16511,N_16161);
nand U18642 (N_18642,N_16530,N_16686);
nand U18643 (N_18643,N_16728,N_17489);
nor U18644 (N_18644,N_17804,N_17241);
nand U18645 (N_18645,N_16137,N_16393);
xor U18646 (N_18646,N_17630,N_16770);
nor U18647 (N_18647,N_17177,N_17318);
or U18648 (N_18648,N_16565,N_17858);
and U18649 (N_18649,N_16799,N_17353);
nor U18650 (N_18650,N_17367,N_17239);
nand U18651 (N_18651,N_16947,N_16827);
nor U18652 (N_18652,N_16198,N_17504);
or U18653 (N_18653,N_17387,N_16498);
nand U18654 (N_18654,N_17403,N_16158);
or U18655 (N_18655,N_17032,N_16332);
xor U18656 (N_18656,N_16326,N_17251);
xor U18657 (N_18657,N_17028,N_16656);
or U18658 (N_18658,N_17355,N_17334);
and U18659 (N_18659,N_16721,N_17916);
nor U18660 (N_18660,N_17628,N_16788);
or U18661 (N_18661,N_17643,N_17413);
xnor U18662 (N_18662,N_16924,N_16379);
or U18663 (N_18663,N_17354,N_16195);
xor U18664 (N_18664,N_17917,N_17954);
xor U18665 (N_18665,N_16497,N_17792);
xnor U18666 (N_18666,N_16378,N_16364);
or U18667 (N_18667,N_16811,N_17158);
and U18668 (N_18668,N_16790,N_16506);
and U18669 (N_18669,N_16616,N_17210);
nand U18670 (N_18670,N_17307,N_17778);
nand U18671 (N_18671,N_17113,N_17539);
or U18672 (N_18672,N_16593,N_17707);
and U18673 (N_18673,N_16281,N_17867);
or U18674 (N_18674,N_17818,N_16735);
xnor U18675 (N_18675,N_16979,N_16042);
and U18676 (N_18676,N_17382,N_16285);
xnor U18677 (N_18677,N_16932,N_17711);
xnor U18678 (N_18678,N_16625,N_17364);
or U18679 (N_18679,N_16798,N_16505);
and U18680 (N_18680,N_17252,N_16438);
nand U18681 (N_18681,N_17277,N_17494);
or U18682 (N_18682,N_16318,N_17155);
xor U18683 (N_18683,N_17016,N_16524);
xor U18684 (N_18684,N_17018,N_17267);
xnor U18685 (N_18685,N_16179,N_17146);
and U18686 (N_18686,N_16128,N_17093);
and U18687 (N_18687,N_17390,N_17670);
or U18688 (N_18688,N_16963,N_17087);
nor U18689 (N_18689,N_17981,N_16674);
and U18690 (N_18690,N_16604,N_17784);
nor U18691 (N_18691,N_17854,N_17820);
or U18692 (N_18692,N_16068,N_16761);
nand U18693 (N_18693,N_17126,N_16605);
xnor U18694 (N_18694,N_17236,N_17844);
and U18695 (N_18695,N_16652,N_16440);
or U18696 (N_18696,N_16487,N_16962);
xnor U18697 (N_18697,N_17603,N_17760);
nor U18698 (N_18698,N_16246,N_17393);
or U18699 (N_18699,N_16744,N_16012);
and U18700 (N_18700,N_16611,N_16293);
xnor U18701 (N_18701,N_17813,N_16466);
or U18702 (N_18702,N_16151,N_17593);
nand U18703 (N_18703,N_16710,N_17061);
nor U18704 (N_18704,N_16624,N_17265);
and U18705 (N_18705,N_17761,N_16833);
nand U18706 (N_18706,N_17394,N_17190);
nor U18707 (N_18707,N_16308,N_17130);
or U18708 (N_18708,N_17959,N_17577);
nor U18709 (N_18709,N_17556,N_17913);
or U18710 (N_18710,N_16603,N_16482);
nand U18711 (N_18711,N_17582,N_16807);
nand U18712 (N_18712,N_16709,N_16165);
and U18713 (N_18713,N_16578,N_16828);
nand U18714 (N_18714,N_16202,N_16563);
and U18715 (N_18715,N_16284,N_17110);
nor U18716 (N_18716,N_17287,N_16050);
nor U18717 (N_18717,N_17350,N_17211);
and U18718 (N_18718,N_16422,N_17631);
or U18719 (N_18719,N_16140,N_17750);
or U18720 (N_18720,N_17349,N_16117);
and U18721 (N_18721,N_16527,N_17741);
nand U18722 (N_18722,N_17882,N_16774);
and U18723 (N_18723,N_17274,N_17360);
and U18724 (N_18724,N_17029,N_16782);
nor U18725 (N_18725,N_17264,N_17178);
nor U18726 (N_18726,N_16412,N_17011);
xnor U18727 (N_18727,N_16553,N_16084);
and U18728 (N_18728,N_16874,N_16136);
and U18729 (N_18729,N_16144,N_17600);
nand U18730 (N_18730,N_16351,N_17796);
xor U18731 (N_18731,N_17721,N_17642);
nand U18732 (N_18732,N_16706,N_17057);
xor U18733 (N_18733,N_17982,N_17138);
xor U18734 (N_18734,N_17923,N_17635);
xor U18735 (N_18735,N_16244,N_17953);
xnor U18736 (N_18736,N_17010,N_16033);
and U18737 (N_18737,N_17994,N_16413);
or U18738 (N_18738,N_16651,N_16172);
xor U18739 (N_18739,N_16966,N_16256);
nor U18740 (N_18740,N_17085,N_16457);
xnor U18741 (N_18741,N_16233,N_16859);
nand U18742 (N_18742,N_17069,N_16451);
and U18743 (N_18743,N_16372,N_17284);
or U18744 (N_18744,N_17369,N_17574);
nor U18745 (N_18745,N_17700,N_17325);
or U18746 (N_18746,N_17868,N_17910);
and U18747 (N_18747,N_17911,N_16662);
nand U18748 (N_18748,N_16458,N_17660);
or U18749 (N_18749,N_16775,N_17851);
nand U18750 (N_18750,N_17853,N_16131);
or U18751 (N_18751,N_17124,N_16753);
nand U18752 (N_18752,N_17698,N_16080);
nor U18753 (N_18753,N_17569,N_17880);
and U18754 (N_18754,N_16380,N_16768);
nand U18755 (N_18755,N_17133,N_16509);
nor U18756 (N_18756,N_17666,N_17220);
nor U18757 (N_18757,N_16493,N_17008);
nor U18758 (N_18758,N_16832,N_16694);
or U18759 (N_18759,N_16199,N_17442);
and U18760 (N_18760,N_16865,N_16039);
and U18761 (N_18761,N_17653,N_17315);
xnor U18762 (N_18762,N_17985,N_16861);
and U18763 (N_18763,N_17481,N_17435);
or U18764 (N_18764,N_16301,N_17607);
nand U18765 (N_18765,N_16584,N_16949);
xnor U18766 (N_18766,N_16542,N_17404);
nor U18767 (N_18767,N_17134,N_17309);
xnor U18768 (N_18768,N_17925,N_17437);
and U18769 (N_18769,N_16227,N_16160);
nand U18770 (N_18770,N_16523,N_17950);
nand U18771 (N_18771,N_17341,N_16462);
or U18772 (N_18772,N_17855,N_17084);
or U18773 (N_18773,N_16723,N_17935);
xnor U18774 (N_18774,N_17759,N_17235);
nand U18775 (N_18775,N_17552,N_16216);
nor U18776 (N_18776,N_17602,N_16612);
xnor U18777 (N_18777,N_16907,N_17056);
nor U18778 (N_18778,N_17586,N_16269);
nor U18779 (N_18779,N_17399,N_17217);
nand U18780 (N_18780,N_16633,N_17560);
nor U18781 (N_18781,N_16572,N_16333);
and U18782 (N_18782,N_16104,N_16469);
nand U18783 (N_18783,N_16328,N_16130);
nor U18784 (N_18784,N_17396,N_17952);
nor U18785 (N_18785,N_17201,N_16784);
and U18786 (N_18786,N_17578,N_16026);
nand U18787 (N_18787,N_17973,N_16073);
nor U18788 (N_18788,N_17612,N_16089);
nor U18789 (N_18789,N_17645,N_16354);
xor U18790 (N_18790,N_17301,N_16750);
or U18791 (N_18791,N_16736,N_16873);
or U18792 (N_18792,N_17005,N_16618);
xnor U18793 (N_18793,N_16082,N_16261);
and U18794 (N_18794,N_17772,N_16034);
nor U18795 (N_18795,N_17468,N_16196);
xor U18796 (N_18796,N_16817,N_17096);
nand U18797 (N_18797,N_16403,N_17498);
nand U18798 (N_18798,N_17551,N_16881);
nand U18799 (N_18799,N_16008,N_16063);
or U18800 (N_18800,N_17499,N_17675);
nor U18801 (N_18801,N_16655,N_17892);
or U18802 (N_18802,N_17337,N_16682);
nand U18803 (N_18803,N_17915,N_16869);
and U18804 (N_18804,N_16594,N_16779);
or U18805 (N_18805,N_17208,N_16587);
or U18806 (N_18806,N_17518,N_17692);
nand U18807 (N_18807,N_16659,N_16823);
nand U18808 (N_18808,N_17231,N_16558);
xor U18809 (N_18809,N_17991,N_17811);
or U18810 (N_18810,N_17141,N_16325);
nor U18811 (N_18811,N_16015,N_16361);
and U18812 (N_18812,N_17956,N_17376);
xnor U18813 (N_18813,N_17453,N_17705);
or U18814 (N_18814,N_16890,N_16027);
nand U18815 (N_18815,N_16917,N_17112);
xnor U18816 (N_18816,N_17314,N_17497);
nand U18817 (N_18817,N_17424,N_16512);
xnor U18818 (N_18818,N_17583,N_16642);
nand U18819 (N_18819,N_16455,N_16316);
nor U18820 (N_18820,N_16437,N_16810);
xor U18821 (N_18821,N_17680,N_16836);
nor U18822 (N_18822,N_16257,N_17009);
or U18823 (N_18823,N_16545,N_16180);
nor U18824 (N_18824,N_16986,N_17970);
or U18825 (N_18825,N_16240,N_17339);
nor U18826 (N_18826,N_16207,N_16712);
nor U18827 (N_18827,N_16488,N_16948);
nand U18828 (N_18828,N_17756,N_16454);
and U18829 (N_18829,N_17736,N_16564);
or U18830 (N_18830,N_16737,N_17462);
xnor U18831 (N_18831,N_16860,N_16387);
or U18832 (N_18832,N_17198,N_17465);
nor U18833 (N_18833,N_17629,N_16035);
or U18834 (N_18834,N_17780,N_16787);
xor U18835 (N_18835,N_17940,N_17281);
nand U18836 (N_18836,N_16711,N_17094);
nand U18837 (N_18837,N_17580,N_17885);
or U18838 (N_18838,N_17516,N_17189);
and U18839 (N_18839,N_17799,N_17790);
or U18840 (N_18840,N_16003,N_17020);
and U18841 (N_18841,N_16771,N_17512);
nor U18842 (N_18842,N_16959,N_16341);
nor U18843 (N_18843,N_16468,N_16322);
nor U18844 (N_18844,N_16211,N_16363);
nor U18845 (N_18845,N_17862,N_17733);
nand U18846 (N_18846,N_16181,N_17471);
or U18847 (N_18847,N_16053,N_16016);
nand U18848 (N_18848,N_16560,N_16588);
or U18849 (N_18849,N_17838,N_16386);
nand U18850 (N_18850,N_16123,N_17212);
and U18851 (N_18851,N_17344,N_16030);
xnor U18852 (N_18852,N_16819,N_17099);
nor U18853 (N_18853,N_16989,N_17987);
xor U18854 (N_18854,N_17118,N_16676);
nor U18855 (N_18855,N_17304,N_16109);
or U18856 (N_18856,N_16634,N_16720);
and U18857 (N_18857,N_17597,N_17535);
or U18858 (N_18858,N_17063,N_16850);
nand U18859 (N_18859,N_17689,N_16990);
and U18860 (N_18860,N_16983,N_17881);
nor U18861 (N_18861,N_17077,N_17693);
nor U18862 (N_18862,N_16780,N_16791);
or U18863 (N_18863,N_17227,N_17690);
or U18864 (N_18864,N_16331,N_16936);
nor U18865 (N_18865,N_16935,N_16919);
nor U18866 (N_18866,N_17173,N_17808);
and U18867 (N_18867,N_16018,N_16731);
nor U18868 (N_18868,N_16037,N_16430);
nor U18869 (N_18869,N_17000,N_16496);
and U18870 (N_18870,N_17164,N_16639);
xnor U18871 (N_18871,N_17933,N_16722);
nor U18872 (N_18872,N_17254,N_17490);
xor U18873 (N_18873,N_16433,N_17739);
and U18874 (N_18874,N_16360,N_16099);
or U18875 (N_18875,N_17123,N_16408);
nor U18876 (N_18876,N_17934,N_17549);
nor U18877 (N_18877,N_17984,N_17263);
nor U18878 (N_18878,N_17906,N_17846);
xnor U18879 (N_18879,N_17797,N_16420);
xor U18880 (N_18880,N_17161,N_16893);
and U18881 (N_18881,N_17402,N_17237);
and U18882 (N_18882,N_17181,N_16955);
nor U18883 (N_18883,N_16613,N_16684);
and U18884 (N_18884,N_17270,N_16894);
xnor U18885 (N_18885,N_16229,N_16143);
and U18886 (N_18886,N_17725,N_16103);
nand U18887 (N_18887,N_16330,N_16961);
xor U18888 (N_18888,N_17919,N_16062);
xnor U18889 (N_18889,N_16119,N_16218);
xnor U18890 (N_18890,N_16460,N_17961);
or U18891 (N_18891,N_17624,N_16660);
and U18892 (N_18892,N_16532,N_17568);
and U18893 (N_18893,N_16215,N_17166);
xnor U18894 (N_18894,N_17626,N_17678);
nor U18895 (N_18895,N_17025,N_17765);
nor U18896 (N_18896,N_16470,N_16091);
xor U18897 (N_18897,N_16981,N_17002);
nor U18898 (N_18898,N_16405,N_17371);
nand U18899 (N_18899,N_16494,N_16772);
nor U18900 (N_18900,N_16554,N_16754);
nor U18901 (N_18901,N_17942,N_16110);
or U18902 (N_18902,N_16802,N_17358);
xor U18903 (N_18903,N_16725,N_16200);
xnor U18904 (N_18904,N_16397,N_17900);
and U18905 (N_18905,N_17948,N_16047);
or U18906 (N_18906,N_16447,N_16390);
xor U18907 (N_18907,N_17455,N_17785);
nor U18908 (N_18908,N_16921,N_16467);
nand U18909 (N_18909,N_17652,N_16253);
and U18910 (N_18910,N_17764,N_16884);
or U18911 (N_18911,N_16504,N_16132);
and U18912 (N_18912,N_17443,N_17530);
xnor U18913 (N_18913,N_16773,N_16292);
nand U18914 (N_18914,N_17383,N_17119);
or U18915 (N_18915,N_16577,N_17169);
nand U18916 (N_18916,N_17017,N_17590);
and U18917 (N_18917,N_17965,N_17706);
nand U18918 (N_18918,N_17419,N_17886);
or U18919 (N_18919,N_17944,N_16002);
nor U18920 (N_18920,N_17687,N_17562);
xor U18921 (N_18921,N_17409,N_16623);
nand U18922 (N_18922,N_16249,N_16937);
nor U18923 (N_18923,N_16638,N_16286);
xor U18924 (N_18924,N_17576,N_17850);
and U18925 (N_18925,N_16751,N_17286);
or U18926 (N_18926,N_17316,N_17174);
nand U18927 (N_18927,N_16024,N_16688);
or U18928 (N_18928,N_16275,N_17199);
xor U18929 (N_18929,N_17618,N_16756);
and U18930 (N_18930,N_16632,N_16139);
or U18931 (N_18931,N_17003,N_16803);
and U18932 (N_18932,N_16663,N_16693);
nor U18933 (N_18933,N_17033,N_16714);
nor U18934 (N_18934,N_16155,N_17682);
nor U18935 (N_18935,N_16531,N_17775);
nand U18936 (N_18936,N_16384,N_16842);
xor U18937 (N_18937,N_16495,N_16730);
or U18938 (N_18938,N_17331,N_17068);
or U18939 (N_18939,N_16411,N_17388);
nand U18940 (N_18940,N_17889,N_17351);
nor U18941 (N_18941,N_16481,N_16675);
xnor U18942 (N_18942,N_16704,N_16946);
or U18943 (N_18943,N_16927,N_16537);
or U18944 (N_18944,N_17527,N_17709);
nand U18945 (N_18945,N_16692,N_17999);
or U18946 (N_18946,N_16394,N_16905);
nand U18947 (N_18947,N_17883,N_17829);
or U18948 (N_18948,N_16708,N_16022);
and U18949 (N_18949,N_17788,N_16944);
xor U18950 (N_18950,N_17839,N_16792);
nor U18951 (N_18951,N_16449,N_16141);
nand U18952 (N_18952,N_17397,N_16192);
or U18953 (N_18953,N_17122,N_16841);
nand U18954 (N_18954,N_16204,N_16337);
nand U18955 (N_18955,N_16152,N_16796);
nor U18956 (N_18956,N_17373,N_16902);
xor U18957 (N_18957,N_16769,N_17962);
nor U18958 (N_18958,N_16056,N_17710);
or U18959 (N_18959,N_16217,N_16734);
or U18960 (N_18960,N_17731,N_16404);
and U18961 (N_18961,N_16270,N_17418);
and U18962 (N_18962,N_17365,N_16031);
xor U18963 (N_18963,N_17555,N_16573);
or U18964 (N_18964,N_17067,N_17013);
nor U18965 (N_18965,N_16219,N_17102);
nand U18966 (N_18966,N_16526,N_17969);
or U18967 (N_18967,N_16107,N_17957);
nand U18968 (N_18968,N_17657,N_16837);
and U18969 (N_18969,N_17075,N_17595);
nand U18970 (N_18970,N_17461,N_17034);
xnor U18971 (N_18971,N_17395,N_17824);
nor U18972 (N_18972,N_17894,N_16579);
nand U18973 (N_18973,N_16108,N_16984);
and U18974 (N_18974,N_17774,N_17456);
nor U18975 (N_18975,N_17283,N_16294);
nand U18976 (N_18976,N_16702,N_17193);
nor U18977 (N_18977,N_17914,N_17860);
xnor U18978 (N_18978,N_17614,N_16528);
xnor U18979 (N_18979,N_17392,N_17082);
or U18980 (N_18980,N_16991,N_17728);
xor U18981 (N_18981,N_16925,N_17180);
or U18982 (N_18982,N_16699,N_17572);
and U18983 (N_18983,N_17305,N_17926);
and U18984 (N_18984,N_17060,N_16904);
or U18985 (N_18985,N_17866,N_17992);
or U18986 (N_18986,N_17139,N_17447);
and U18987 (N_18987,N_17221,N_16752);
xnor U18988 (N_18988,N_17218,N_17816);
xnor U18989 (N_18989,N_16801,N_17417);
or U18990 (N_18990,N_16226,N_17153);
and U18991 (N_18991,N_17558,N_17514);
xor U18992 (N_18992,N_17152,N_16549);
nor U18993 (N_18993,N_17589,N_16797);
nor U18994 (N_18994,N_16757,N_16456);
nand U18995 (N_18995,N_17904,N_17345);
xor U18996 (N_18996,N_17343,N_16077);
and U18997 (N_18997,N_16478,N_17541);
or U18998 (N_18998,N_16288,N_17650);
and U18999 (N_18999,N_16407,N_17375);
nor U19000 (N_19000,N_17776,N_17687);
nand U19001 (N_19001,N_16848,N_16856);
nand U19002 (N_19002,N_16541,N_17556);
nor U19003 (N_19003,N_16555,N_17153);
nand U19004 (N_19004,N_17438,N_16383);
nor U19005 (N_19005,N_17431,N_16912);
or U19006 (N_19006,N_16694,N_16110);
or U19007 (N_19007,N_17530,N_16224);
xnor U19008 (N_19008,N_17367,N_17730);
xor U19009 (N_19009,N_17292,N_16254);
nand U19010 (N_19010,N_17027,N_17267);
xor U19011 (N_19011,N_16442,N_16768);
xnor U19012 (N_19012,N_16819,N_17388);
or U19013 (N_19013,N_17490,N_17460);
nand U19014 (N_19014,N_16487,N_16853);
nand U19015 (N_19015,N_17701,N_17721);
and U19016 (N_19016,N_16820,N_16175);
or U19017 (N_19017,N_17187,N_16481);
nand U19018 (N_19018,N_17350,N_17694);
xor U19019 (N_19019,N_17061,N_17870);
and U19020 (N_19020,N_16652,N_16706);
and U19021 (N_19021,N_16927,N_16163);
nand U19022 (N_19022,N_16740,N_17149);
and U19023 (N_19023,N_17759,N_17432);
and U19024 (N_19024,N_17254,N_17589);
xor U19025 (N_19025,N_16187,N_17182);
or U19026 (N_19026,N_17073,N_17476);
nand U19027 (N_19027,N_17843,N_16654);
nand U19028 (N_19028,N_16945,N_17012);
and U19029 (N_19029,N_16010,N_17043);
nand U19030 (N_19030,N_17393,N_17564);
nand U19031 (N_19031,N_16279,N_16896);
and U19032 (N_19032,N_17165,N_16667);
and U19033 (N_19033,N_17252,N_17838);
nand U19034 (N_19034,N_17353,N_16525);
nand U19035 (N_19035,N_16566,N_16430);
nand U19036 (N_19036,N_17558,N_16699);
nand U19037 (N_19037,N_17853,N_17085);
and U19038 (N_19038,N_17988,N_17904);
and U19039 (N_19039,N_16464,N_17375);
and U19040 (N_19040,N_17622,N_17172);
nor U19041 (N_19041,N_17403,N_16497);
xnor U19042 (N_19042,N_16805,N_17778);
xnor U19043 (N_19043,N_16246,N_16244);
nand U19044 (N_19044,N_17064,N_17111);
nor U19045 (N_19045,N_16114,N_17595);
nor U19046 (N_19046,N_17910,N_17860);
nand U19047 (N_19047,N_16400,N_16271);
and U19048 (N_19048,N_16199,N_17042);
and U19049 (N_19049,N_17713,N_17870);
and U19050 (N_19050,N_17386,N_16260);
xnor U19051 (N_19051,N_17430,N_17060);
nor U19052 (N_19052,N_17885,N_17585);
or U19053 (N_19053,N_17640,N_16631);
nand U19054 (N_19054,N_17402,N_17839);
xnor U19055 (N_19055,N_17608,N_16874);
nor U19056 (N_19056,N_16441,N_17299);
nand U19057 (N_19057,N_16544,N_16117);
xnor U19058 (N_19058,N_16967,N_17564);
nand U19059 (N_19059,N_17806,N_16125);
nor U19060 (N_19060,N_16294,N_16180);
or U19061 (N_19061,N_17148,N_16869);
nand U19062 (N_19062,N_17218,N_17446);
nor U19063 (N_19063,N_17008,N_17424);
xor U19064 (N_19064,N_16898,N_16331);
nor U19065 (N_19065,N_16727,N_16747);
nor U19066 (N_19066,N_17699,N_17270);
xor U19067 (N_19067,N_16939,N_16393);
nor U19068 (N_19068,N_17726,N_17843);
xnor U19069 (N_19069,N_16513,N_16827);
and U19070 (N_19070,N_17563,N_17112);
nor U19071 (N_19071,N_16212,N_16975);
and U19072 (N_19072,N_17596,N_17380);
nor U19073 (N_19073,N_17315,N_17133);
nand U19074 (N_19074,N_16434,N_17390);
or U19075 (N_19075,N_16424,N_17764);
or U19076 (N_19076,N_17546,N_16750);
xor U19077 (N_19077,N_17057,N_16100);
nor U19078 (N_19078,N_16624,N_17152);
xnor U19079 (N_19079,N_17931,N_17190);
or U19080 (N_19080,N_16242,N_17881);
xnor U19081 (N_19081,N_16529,N_17884);
and U19082 (N_19082,N_17284,N_16816);
xor U19083 (N_19083,N_17026,N_17171);
xnor U19084 (N_19084,N_17500,N_16668);
xnor U19085 (N_19085,N_17287,N_16033);
nor U19086 (N_19086,N_16700,N_16151);
and U19087 (N_19087,N_17197,N_17360);
xnor U19088 (N_19088,N_17584,N_17591);
nand U19089 (N_19089,N_16829,N_17078);
or U19090 (N_19090,N_16351,N_16170);
xnor U19091 (N_19091,N_17939,N_17125);
nand U19092 (N_19092,N_16490,N_17485);
and U19093 (N_19093,N_17002,N_16050);
xnor U19094 (N_19094,N_16668,N_16382);
xor U19095 (N_19095,N_16575,N_17153);
nor U19096 (N_19096,N_16385,N_16527);
nand U19097 (N_19097,N_17197,N_16691);
and U19098 (N_19098,N_16292,N_17877);
and U19099 (N_19099,N_17824,N_16029);
or U19100 (N_19100,N_16716,N_16614);
nor U19101 (N_19101,N_16111,N_16514);
xnor U19102 (N_19102,N_16183,N_17030);
nand U19103 (N_19103,N_16264,N_17200);
xnor U19104 (N_19104,N_17453,N_17249);
xor U19105 (N_19105,N_17685,N_16463);
nand U19106 (N_19106,N_16067,N_17600);
nor U19107 (N_19107,N_16645,N_17877);
nor U19108 (N_19108,N_16440,N_17626);
or U19109 (N_19109,N_17753,N_16881);
nand U19110 (N_19110,N_16470,N_16818);
or U19111 (N_19111,N_17760,N_16303);
nor U19112 (N_19112,N_16800,N_16353);
or U19113 (N_19113,N_17429,N_17209);
xnor U19114 (N_19114,N_17251,N_17013);
or U19115 (N_19115,N_16258,N_17144);
xnor U19116 (N_19116,N_17673,N_16668);
or U19117 (N_19117,N_17802,N_16947);
and U19118 (N_19118,N_16865,N_17506);
nand U19119 (N_19119,N_16206,N_17775);
xnor U19120 (N_19120,N_17754,N_17009);
xor U19121 (N_19121,N_17115,N_17959);
and U19122 (N_19122,N_16993,N_17322);
nand U19123 (N_19123,N_17913,N_16908);
nor U19124 (N_19124,N_17390,N_17010);
and U19125 (N_19125,N_17772,N_17291);
nor U19126 (N_19126,N_16794,N_16036);
and U19127 (N_19127,N_17490,N_16468);
xnor U19128 (N_19128,N_16306,N_17901);
and U19129 (N_19129,N_17363,N_17967);
nand U19130 (N_19130,N_16708,N_17124);
or U19131 (N_19131,N_17682,N_17825);
or U19132 (N_19132,N_16566,N_16967);
nand U19133 (N_19133,N_16168,N_16616);
nand U19134 (N_19134,N_16877,N_17144);
or U19135 (N_19135,N_17585,N_17129);
or U19136 (N_19136,N_16734,N_17243);
or U19137 (N_19137,N_16178,N_17182);
nand U19138 (N_19138,N_16973,N_16227);
nand U19139 (N_19139,N_16703,N_17818);
xor U19140 (N_19140,N_16103,N_16325);
nor U19141 (N_19141,N_16912,N_16511);
and U19142 (N_19142,N_16453,N_16054);
and U19143 (N_19143,N_17014,N_17198);
nor U19144 (N_19144,N_16444,N_16808);
xnor U19145 (N_19145,N_16098,N_16973);
or U19146 (N_19146,N_16693,N_16444);
nand U19147 (N_19147,N_17974,N_17600);
or U19148 (N_19148,N_16766,N_16126);
or U19149 (N_19149,N_17437,N_16963);
and U19150 (N_19150,N_17148,N_16517);
nor U19151 (N_19151,N_16228,N_16877);
and U19152 (N_19152,N_17816,N_16444);
and U19153 (N_19153,N_16637,N_16311);
and U19154 (N_19154,N_16633,N_16940);
xnor U19155 (N_19155,N_17096,N_16233);
and U19156 (N_19156,N_16563,N_17137);
and U19157 (N_19157,N_16405,N_17940);
nand U19158 (N_19158,N_16395,N_16179);
xor U19159 (N_19159,N_16020,N_16183);
xor U19160 (N_19160,N_16731,N_16899);
xnor U19161 (N_19161,N_17839,N_16217);
or U19162 (N_19162,N_16669,N_17906);
nor U19163 (N_19163,N_16132,N_17793);
nand U19164 (N_19164,N_17687,N_17683);
or U19165 (N_19165,N_16282,N_17492);
xor U19166 (N_19166,N_17321,N_16013);
nand U19167 (N_19167,N_16617,N_16785);
or U19168 (N_19168,N_16171,N_17830);
or U19169 (N_19169,N_16889,N_16456);
and U19170 (N_19170,N_17827,N_16828);
xor U19171 (N_19171,N_17165,N_17737);
or U19172 (N_19172,N_17962,N_16110);
xnor U19173 (N_19173,N_17320,N_17666);
and U19174 (N_19174,N_17741,N_17740);
xnor U19175 (N_19175,N_16044,N_16464);
nor U19176 (N_19176,N_17083,N_17493);
nand U19177 (N_19177,N_16487,N_16191);
nor U19178 (N_19178,N_16847,N_17251);
nand U19179 (N_19179,N_17426,N_17699);
or U19180 (N_19180,N_17025,N_17707);
nor U19181 (N_19181,N_17082,N_17977);
xnor U19182 (N_19182,N_17650,N_16443);
nand U19183 (N_19183,N_16940,N_17603);
xor U19184 (N_19184,N_17322,N_17525);
and U19185 (N_19185,N_17754,N_16309);
or U19186 (N_19186,N_17281,N_16984);
nor U19187 (N_19187,N_17479,N_17199);
xor U19188 (N_19188,N_16921,N_17403);
nand U19189 (N_19189,N_17551,N_16432);
or U19190 (N_19190,N_17323,N_16172);
nor U19191 (N_19191,N_16294,N_17696);
nor U19192 (N_19192,N_17215,N_17575);
nor U19193 (N_19193,N_16235,N_17423);
xor U19194 (N_19194,N_16068,N_16339);
and U19195 (N_19195,N_17186,N_17123);
and U19196 (N_19196,N_16335,N_17607);
nor U19197 (N_19197,N_17503,N_17219);
and U19198 (N_19198,N_16279,N_16487);
and U19199 (N_19199,N_16777,N_17792);
xnor U19200 (N_19200,N_17627,N_16871);
nand U19201 (N_19201,N_17155,N_16079);
xnor U19202 (N_19202,N_17451,N_17956);
nor U19203 (N_19203,N_17750,N_16800);
nor U19204 (N_19204,N_16398,N_17394);
nor U19205 (N_19205,N_16479,N_17117);
xnor U19206 (N_19206,N_17500,N_17922);
nand U19207 (N_19207,N_16436,N_17504);
xor U19208 (N_19208,N_16641,N_16260);
and U19209 (N_19209,N_17537,N_16968);
xnor U19210 (N_19210,N_16989,N_17778);
and U19211 (N_19211,N_17672,N_16796);
or U19212 (N_19212,N_16814,N_16591);
nor U19213 (N_19213,N_17089,N_17219);
or U19214 (N_19214,N_16395,N_17374);
and U19215 (N_19215,N_17979,N_16274);
xnor U19216 (N_19216,N_17468,N_17219);
and U19217 (N_19217,N_16634,N_16887);
xor U19218 (N_19218,N_17014,N_17731);
nand U19219 (N_19219,N_17945,N_16882);
nor U19220 (N_19220,N_16623,N_16091);
and U19221 (N_19221,N_16515,N_16026);
and U19222 (N_19222,N_16324,N_17811);
or U19223 (N_19223,N_17241,N_17767);
xor U19224 (N_19224,N_17690,N_16519);
and U19225 (N_19225,N_17674,N_17290);
or U19226 (N_19226,N_17205,N_17806);
and U19227 (N_19227,N_16322,N_17806);
nand U19228 (N_19228,N_16427,N_16676);
nand U19229 (N_19229,N_17798,N_17951);
xor U19230 (N_19230,N_17360,N_17437);
and U19231 (N_19231,N_16118,N_16472);
and U19232 (N_19232,N_16370,N_16456);
nor U19233 (N_19233,N_17423,N_16454);
and U19234 (N_19234,N_16898,N_16120);
nor U19235 (N_19235,N_16112,N_16483);
xnor U19236 (N_19236,N_17563,N_17071);
nand U19237 (N_19237,N_17870,N_17521);
or U19238 (N_19238,N_17416,N_16439);
or U19239 (N_19239,N_16680,N_17123);
xor U19240 (N_19240,N_16791,N_16896);
or U19241 (N_19241,N_17395,N_17972);
nand U19242 (N_19242,N_16316,N_17207);
xor U19243 (N_19243,N_16054,N_16123);
and U19244 (N_19244,N_17340,N_16513);
and U19245 (N_19245,N_16934,N_17315);
and U19246 (N_19246,N_16891,N_16143);
nor U19247 (N_19247,N_17865,N_17781);
or U19248 (N_19248,N_17931,N_16939);
nor U19249 (N_19249,N_16352,N_17591);
xor U19250 (N_19250,N_16428,N_16983);
or U19251 (N_19251,N_17094,N_17714);
nor U19252 (N_19252,N_17200,N_17125);
nor U19253 (N_19253,N_16888,N_17359);
nand U19254 (N_19254,N_17991,N_17292);
and U19255 (N_19255,N_17633,N_17293);
or U19256 (N_19256,N_16887,N_17610);
or U19257 (N_19257,N_16006,N_17293);
or U19258 (N_19258,N_16764,N_16058);
nor U19259 (N_19259,N_17410,N_16812);
nor U19260 (N_19260,N_17069,N_17983);
and U19261 (N_19261,N_17614,N_17380);
xor U19262 (N_19262,N_17141,N_16083);
xor U19263 (N_19263,N_17101,N_17361);
xor U19264 (N_19264,N_16904,N_16329);
nand U19265 (N_19265,N_17997,N_17556);
nor U19266 (N_19266,N_16180,N_16781);
nand U19267 (N_19267,N_16524,N_16586);
nand U19268 (N_19268,N_17189,N_16645);
or U19269 (N_19269,N_16670,N_16997);
nor U19270 (N_19270,N_17495,N_17436);
xor U19271 (N_19271,N_16910,N_17098);
xnor U19272 (N_19272,N_17547,N_17151);
xor U19273 (N_19273,N_16749,N_16731);
xor U19274 (N_19274,N_17780,N_16251);
and U19275 (N_19275,N_16010,N_16961);
and U19276 (N_19276,N_16513,N_16642);
or U19277 (N_19277,N_17268,N_16336);
nand U19278 (N_19278,N_17793,N_16229);
or U19279 (N_19279,N_16145,N_16424);
and U19280 (N_19280,N_17445,N_17394);
or U19281 (N_19281,N_16942,N_16497);
xor U19282 (N_19282,N_16733,N_17633);
nor U19283 (N_19283,N_17075,N_17731);
xor U19284 (N_19284,N_16248,N_17160);
and U19285 (N_19285,N_17849,N_16557);
or U19286 (N_19286,N_16253,N_17130);
nand U19287 (N_19287,N_17178,N_16117);
nand U19288 (N_19288,N_16840,N_16810);
nor U19289 (N_19289,N_17084,N_17367);
nand U19290 (N_19290,N_17161,N_17578);
xnor U19291 (N_19291,N_16137,N_16473);
or U19292 (N_19292,N_17385,N_17988);
nor U19293 (N_19293,N_16866,N_16076);
xor U19294 (N_19294,N_17939,N_16322);
or U19295 (N_19295,N_17697,N_16402);
xor U19296 (N_19296,N_17939,N_16985);
nand U19297 (N_19297,N_17043,N_16238);
nor U19298 (N_19298,N_17825,N_17800);
or U19299 (N_19299,N_17764,N_17507);
and U19300 (N_19300,N_17449,N_17286);
or U19301 (N_19301,N_16738,N_17617);
and U19302 (N_19302,N_17971,N_17362);
or U19303 (N_19303,N_17336,N_16624);
xnor U19304 (N_19304,N_16699,N_16994);
or U19305 (N_19305,N_16189,N_17148);
or U19306 (N_19306,N_16232,N_17443);
nor U19307 (N_19307,N_17371,N_17470);
xnor U19308 (N_19308,N_17048,N_16100);
and U19309 (N_19309,N_17302,N_16554);
and U19310 (N_19310,N_17019,N_16838);
xor U19311 (N_19311,N_17864,N_17173);
or U19312 (N_19312,N_17270,N_16845);
and U19313 (N_19313,N_17512,N_16566);
or U19314 (N_19314,N_17347,N_17266);
nand U19315 (N_19315,N_16307,N_17579);
or U19316 (N_19316,N_17786,N_17522);
nand U19317 (N_19317,N_17662,N_17861);
and U19318 (N_19318,N_16742,N_17425);
nor U19319 (N_19319,N_17854,N_16761);
or U19320 (N_19320,N_17220,N_16684);
nand U19321 (N_19321,N_17249,N_16234);
or U19322 (N_19322,N_17511,N_16544);
or U19323 (N_19323,N_16732,N_16338);
nand U19324 (N_19324,N_17979,N_16008);
and U19325 (N_19325,N_17476,N_16818);
xor U19326 (N_19326,N_16781,N_17558);
xnor U19327 (N_19327,N_17282,N_16091);
nand U19328 (N_19328,N_16955,N_17492);
or U19329 (N_19329,N_17555,N_16151);
or U19330 (N_19330,N_16524,N_16667);
xor U19331 (N_19331,N_17318,N_17330);
nand U19332 (N_19332,N_16644,N_17723);
xor U19333 (N_19333,N_16758,N_17860);
or U19334 (N_19334,N_17971,N_17805);
nor U19335 (N_19335,N_16025,N_17912);
and U19336 (N_19336,N_17104,N_17578);
nor U19337 (N_19337,N_16486,N_17595);
nor U19338 (N_19338,N_17463,N_16431);
xor U19339 (N_19339,N_17685,N_16247);
xor U19340 (N_19340,N_17728,N_17149);
or U19341 (N_19341,N_16497,N_16376);
and U19342 (N_19342,N_17963,N_16979);
nor U19343 (N_19343,N_17437,N_16949);
xnor U19344 (N_19344,N_16750,N_17432);
nor U19345 (N_19345,N_17504,N_16254);
or U19346 (N_19346,N_17123,N_16451);
nand U19347 (N_19347,N_17461,N_16185);
and U19348 (N_19348,N_16735,N_17095);
nand U19349 (N_19349,N_17431,N_16358);
and U19350 (N_19350,N_16780,N_17278);
or U19351 (N_19351,N_16448,N_16601);
or U19352 (N_19352,N_17803,N_16009);
or U19353 (N_19353,N_16010,N_16573);
or U19354 (N_19354,N_16340,N_16535);
and U19355 (N_19355,N_17001,N_17159);
or U19356 (N_19356,N_17157,N_16591);
and U19357 (N_19357,N_16894,N_17978);
and U19358 (N_19358,N_17959,N_17113);
and U19359 (N_19359,N_17897,N_17579);
xor U19360 (N_19360,N_17416,N_16479);
nand U19361 (N_19361,N_17993,N_16452);
nand U19362 (N_19362,N_16534,N_16049);
and U19363 (N_19363,N_16205,N_17152);
and U19364 (N_19364,N_17192,N_16851);
xor U19365 (N_19365,N_17411,N_16397);
nand U19366 (N_19366,N_16752,N_17403);
nor U19367 (N_19367,N_16228,N_16656);
nor U19368 (N_19368,N_16624,N_17143);
nor U19369 (N_19369,N_17122,N_16114);
xor U19370 (N_19370,N_16062,N_17838);
nand U19371 (N_19371,N_16276,N_16464);
nor U19372 (N_19372,N_16976,N_16954);
nand U19373 (N_19373,N_16875,N_16937);
and U19374 (N_19374,N_17614,N_16612);
nand U19375 (N_19375,N_16478,N_17156);
nand U19376 (N_19376,N_17251,N_17540);
nor U19377 (N_19377,N_16794,N_17558);
and U19378 (N_19378,N_16780,N_16913);
or U19379 (N_19379,N_16896,N_16056);
nor U19380 (N_19380,N_17921,N_17903);
nor U19381 (N_19381,N_16817,N_16079);
nand U19382 (N_19382,N_17472,N_16833);
or U19383 (N_19383,N_16475,N_17879);
nor U19384 (N_19384,N_17092,N_17185);
and U19385 (N_19385,N_17745,N_17974);
and U19386 (N_19386,N_17798,N_16893);
nor U19387 (N_19387,N_17091,N_17821);
xor U19388 (N_19388,N_17634,N_17175);
nor U19389 (N_19389,N_17038,N_16487);
or U19390 (N_19390,N_16492,N_17865);
xor U19391 (N_19391,N_16676,N_17680);
and U19392 (N_19392,N_16084,N_16334);
xor U19393 (N_19393,N_16931,N_16385);
and U19394 (N_19394,N_17338,N_16658);
nand U19395 (N_19395,N_17581,N_16359);
or U19396 (N_19396,N_16425,N_17335);
xnor U19397 (N_19397,N_17379,N_17589);
nand U19398 (N_19398,N_16533,N_16919);
nand U19399 (N_19399,N_16653,N_17462);
xor U19400 (N_19400,N_16519,N_17941);
nor U19401 (N_19401,N_17404,N_17325);
nor U19402 (N_19402,N_17197,N_16374);
nand U19403 (N_19403,N_16392,N_17793);
and U19404 (N_19404,N_17947,N_16748);
nor U19405 (N_19405,N_17695,N_16851);
nand U19406 (N_19406,N_16363,N_16827);
nor U19407 (N_19407,N_16516,N_17418);
nand U19408 (N_19408,N_17653,N_16700);
nand U19409 (N_19409,N_17976,N_16433);
and U19410 (N_19410,N_17821,N_17774);
nor U19411 (N_19411,N_17712,N_17113);
and U19412 (N_19412,N_17490,N_17400);
or U19413 (N_19413,N_16680,N_16356);
xnor U19414 (N_19414,N_16492,N_17997);
and U19415 (N_19415,N_16117,N_17960);
and U19416 (N_19416,N_17076,N_17770);
xor U19417 (N_19417,N_16588,N_17762);
and U19418 (N_19418,N_17223,N_16566);
or U19419 (N_19419,N_16192,N_17156);
nor U19420 (N_19420,N_16795,N_17416);
xor U19421 (N_19421,N_17804,N_17772);
nor U19422 (N_19422,N_16460,N_16249);
and U19423 (N_19423,N_17436,N_17157);
nor U19424 (N_19424,N_17406,N_17775);
or U19425 (N_19425,N_16523,N_17991);
and U19426 (N_19426,N_17516,N_16518);
nand U19427 (N_19427,N_17493,N_17551);
nand U19428 (N_19428,N_16671,N_17425);
xor U19429 (N_19429,N_16256,N_16329);
xor U19430 (N_19430,N_17004,N_17931);
or U19431 (N_19431,N_17547,N_17491);
or U19432 (N_19432,N_16590,N_16759);
nor U19433 (N_19433,N_17357,N_17205);
nor U19434 (N_19434,N_17857,N_16431);
nand U19435 (N_19435,N_16364,N_17332);
nand U19436 (N_19436,N_16418,N_17130);
nand U19437 (N_19437,N_16664,N_16141);
or U19438 (N_19438,N_16827,N_17397);
or U19439 (N_19439,N_17642,N_17887);
nand U19440 (N_19440,N_17857,N_16559);
nor U19441 (N_19441,N_16221,N_17841);
or U19442 (N_19442,N_17359,N_16495);
xnor U19443 (N_19443,N_17929,N_17405);
xnor U19444 (N_19444,N_17934,N_16703);
and U19445 (N_19445,N_16964,N_17815);
nand U19446 (N_19446,N_17382,N_17361);
nand U19447 (N_19447,N_16532,N_17692);
nand U19448 (N_19448,N_16212,N_17445);
nand U19449 (N_19449,N_16255,N_17046);
and U19450 (N_19450,N_17216,N_16763);
nand U19451 (N_19451,N_16445,N_16509);
nor U19452 (N_19452,N_17377,N_17976);
or U19453 (N_19453,N_16636,N_17462);
nand U19454 (N_19454,N_17110,N_17958);
or U19455 (N_19455,N_16991,N_16945);
xor U19456 (N_19456,N_16506,N_16419);
xnor U19457 (N_19457,N_16551,N_16113);
and U19458 (N_19458,N_17275,N_17533);
nor U19459 (N_19459,N_17396,N_16622);
and U19460 (N_19460,N_17847,N_17482);
nor U19461 (N_19461,N_16053,N_16972);
and U19462 (N_19462,N_16929,N_16894);
nand U19463 (N_19463,N_17698,N_16619);
or U19464 (N_19464,N_16031,N_17464);
xnor U19465 (N_19465,N_17356,N_17169);
nand U19466 (N_19466,N_17482,N_17911);
nor U19467 (N_19467,N_17336,N_17889);
xor U19468 (N_19468,N_17134,N_17328);
or U19469 (N_19469,N_16720,N_17329);
nand U19470 (N_19470,N_17043,N_16612);
and U19471 (N_19471,N_17873,N_16124);
and U19472 (N_19472,N_17826,N_17992);
and U19473 (N_19473,N_16959,N_17907);
and U19474 (N_19474,N_17907,N_17312);
xor U19475 (N_19475,N_16706,N_17234);
or U19476 (N_19476,N_16223,N_16625);
nor U19477 (N_19477,N_17667,N_16547);
xnor U19478 (N_19478,N_17519,N_17325);
or U19479 (N_19479,N_16554,N_16041);
xor U19480 (N_19480,N_16014,N_17308);
or U19481 (N_19481,N_17229,N_17790);
and U19482 (N_19482,N_16753,N_17063);
and U19483 (N_19483,N_16864,N_17823);
nor U19484 (N_19484,N_16506,N_17587);
nor U19485 (N_19485,N_17896,N_16701);
nand U19486 (N_19486,N_16000,N_17196);
or U19487 (N_19487,N_16358,N_16305);
nor U19488 (N_19488,N_17772,N_16085);
or U19489 (N_19489,N_17411,N_16602);
nor U19490 (N_19490,N_16890,N_16181);
nor U19491 (N_19491,N_16909,N_16565);
and U19492 (N_19492,N_17270,N_17702);
or U19493 (N_19493,N_17489,N_17973);
or U19494 (N_19494,N_16634,N_17008);
and U19495 (N_19495,N_17693,N_16836);
nor U19496 (N_19496,N_16226,N_17501);
nand U19497 (N_19497,N_16721,N_17306);
or U19498 (N_19498,N_16440,N_16893);
nor U19499 (N_19499,N_17135,N_17255);
xor U19500 (N_19500,N_16018,N_16576);
or U19501 (N_19501,N_17235,N_16659);
nand U19502 (N_19502,N_17481,N_17298);
and U19503 (N_19503,N_16037,N_16330);
nand U19504 (N_19504,N_17882,N_17284);
nand U19505 (N_19505,N_16087,N_17903);
nor U19506 (N_19506,N_17624,N_17359);
or U19507 (N_19507,N_17019,N_16781);
and U19508 (N_19508,N_16912,N_17072);
or U19509 (N_19509,N_17014,N_17195);
nand U19510 (N_19510,N_16106,N_17837);
or U19511 (N_19511,N_17887,N_16931);
or U19512 (N_19512,N_17664,N_16045);
nand U19513 (N_19513,N_17118,N_16903);
nor U19514 (N_19514,N_17820,N_17699);
nor U19515 (N_19515,N_17686,N_16413);
nor U19516 (N_19516,N_16537,N_16395);
xnor U19517 (N_19517,N_16260,N_16068);
nor U19518 (N_19518,N_16512,N_17301);
nand U19519 (N_19519,N_16416,N_16243);
xor U19520 (N_19520,N_17292,N_17962);
and U19521 (N_19521,N_16939,N_16545);
or U19522 (N_19522,N_17348,N_17739);
nor U19523 (N_19523,N_16865,N_16758);
and U19524 (N_19524,N_16000,N_16886);
nor U19525 (N_19525,N_16918,N_17483);
nor U19526 (N_19526,N_17065,N_16768);
nor U19527 (N_19527,N_17222,N_17570);
and U19528 (N_19528,N_17070,N_17811);
nand U19529 (N_19529,N_16500,N_16625);
and U19530 (N_19530,N_17058,N_17696);
nand U19531 (N_19531,N_17096,N_17182);
or U19532 (N_19532,N_16746,N_16044);
xor U19533 (N_19533,N_16295,N_17774);
and U19534 (N_19534,N_16912,N_16992);
and U19535 (N_19535,N_17473,N_17383);
nor U19536 (N_19536,N_16771,N_17563);
nor U19537 (N_19537,N_16115,N_16548);
nand U19538 (N_19538,N_16672,N_17341);
xnor U19539 (N_19539,N_16443,N_17478);
nand U19540 (N_19540,N_17311,N_16534);
xnor U19541 (N_19541,N_17294,N_16398);
xor U19542 (N_19542,N_16785,N_16993);
nor U19543 (N_19543,N_17082,N_17294);
xnor U19544 (N_19544,N_17923,N_16613);
nand U19545 (N_19545,N_16979,N_16615);
and U19546 (N_19546,N_17172,N_17958);
nor U19547 (N_19547,N_17902,N_17736);
xor U19548 (N_19548,N_16976,N_17764);
and U19549 (N_19549,N_17479,N_16860);
nor U19550 (N_19550,N_17160,N_17886);
xor U19551 (N_19551,N_16079,N_16698);
xor U19552 (N_19552,N_16768,N_16736);
nor U19553 (N_19553,N_17881,N_16473);
nand U19554 (N_19554,N_16198,N_17000);
and U19555 (N_19555,N_17133,N_17741);
xor U19556 (N_19556,N_17188,N_17420);
xnor U19557 (N_19557,N_16586,N_17862);
nand U19558 (N_19558,N_16015,N_17994);
xnor U19559 (N_19559,N_17392,N_16897);
or U19560 (N_19560,N_16044,N_16783);
nor U19561 (N_19561,N_16713,N_16955);
xnor U19562 (N_19562,N_17147,N_16945);
xnor U19563 (N_19563,N_16917,N_17370);
and U19564 (N_19564,N_16558,N_16408);
nand U19565 (N_19565,N_16657,N_16411);
and U19566 (N_19566,N_17819,N_17945);
xor U19567 (N_19567,N_16165,N_17539);
nor U19568 (N_19568,N_17908,N_16943);
and U19569 (N_19569,N_17638,N_16999);
nand U19570 (N_19570,N_16017,N_17713);
nand U19571 (N_19571,N_16121,N_16404);
xnor U19572 (N_19572,N_16443,N_17177);
nand U19573 (N_19573,N_17708,N_16186);
nor U19574 (N_19574,N_16163,N_16067);
and U19575 (N_19575,N_17232,N_17665);
or U19576 (N_19576,N_16595,N_16263);
or U19577 (N_19577,N_16835,N_16028);
nand U19578 (N_19578,N_17090,N_17131);
or U19579 (N_19579,N_17651,N_17194);
or U19580 (N_19580,N_17494,N_16332);
xnor U19581 (N_19581,N_16746,N_16353);
xor U19582 (N_19582,N_17876,N_16150);
xnor U19583 (N_19583,N_17978,N_16691);
and U19584 (N_19584,N_16244,N_17649);
xor U19585 (N_19585,N_17118,N_17488);
xor U19586 (N_19586,N_16148,N_17948);
nand U19587 (N_19587,N_17895,N_17792);
nor U19588 (N_19588,N_16942,N_16964);
or U19589 (N_19589,N_16112,N_17248);
xor U19590 (N_19590,N_17391,N_16190);
nor U19591 (N_19591,N_17129,N_16440);
xnor U19592 (N_19592,N_17929,N_17581);
nand U19593 (N_19593,N_17764,N_16388);
nand U19594 (N_19594,N_16368,N_17725);
nor U19595 (N_19595,N_17155,N_17211);
and U19596 (N_19596,N_17980,N_17313);
or U19597 (N_19597,N_16311,N_17392);
nor U19598 (N_19598,N_16898,N_16359);
xor U19599 (N_19599,N_17790,N_17476);
or U19600 (N_19600,N_17219,N_17742);
and U19601 (N_19601,N_17613,N_17974);
nor U19602 (N_19602,N_17557,N_16405);
and U19603 (N_19603,N_17082,N_17174);
nor U19604 (N_19604,N_17464,N_16202);
and U19605 (N_19605,N_16940,N_17072);
or U19606 (N_19606,N_17027,N_17560);
nand U19607 (N_19607,N_16931,N_16749);
nor U19608 (N_19608,N_17555,N_17256);
nand U19609 (N_19609,N_17330,N_16920);
or U19610 (N_19610,N_16292,N_17512);
xor U19611 (N_19611,N_16344,N_17746);
xor U19612 (N_19612,N_17003,N_17627);
nor U19613 (N_19613,N_17796,N_16661);
or U19614 (N_19614,N_17621,N_16758);
xor U19615 (N_19615,N_16508,N_17052);
xor U19616 (N_19616,N_16978,N_16930);
nand U19617 (N_19617,N_17821,N_16669);
nor U19618 (N_19618,N_16720,N_17761);
nand U19619 (N_19619,N_17481,N_17923);
or U19620 (N_19620,N_16338,N_17056);
nor U19621 (N_19621,N_17422,N_16701);
nor U19622 (N_19622,N_16645,N_17946);
xor U19623 (N_19623,N_16593,N_17410);
and U19624 (N_19624,N_16978,N_17961);
nor U19625 (N_19625,N_17318,N_16641);
xor U19626 (N_19626,N_16157,N_17498);
nand U19627 (N_19627,N_16371,N_17551);
or U19628 (N_19628,N_16315,N_16841);
nand U19629 (N_19629,N_17437,N_16692);
xor U19630 (N_19630,N_16988,N_16366);
xor U19631 (N_19631,N_17193,N_17372);
or U19632 (N_19632,N_16643,N_17818);
and U19633 (N_19633,N_16528,N_16322);
nor U19634 (N_19634,N_17151,N_16359);
nor U19635 (N_19635,N_17660,N_16331);
xor U19636 (N_19636,N_17261,N_17135);
nor U19637 (N_19637,N_16304,N_17997);
xor U19638 (N_19638,N_16673,N_17499);
nand U19639 (N_19639,N_16056,N_17862);
xor U19640 (N_19640,N_16504,N_16584);
nand U19641 (N_19641,N_17182,N_16202);
and U19642 (N_19642,N_17726,N_17697);
nand U19643 (N_19643,N_16504,N_16483);
and U19644 (N_19644,N_17431,N_16682);
or U19645 (N_19645,N_16519,N_16977);
or U19646 (N_19646,N_17193,N_16650);
xor U19647 (N_19647,N_16628,N_16994);
nor U19648 (N_19648,N_16875,N_16599);
and U19649 (N_19649,N_16463,N_16026);
and U19650 (N_19650,N_17928,N_16481);
or U19651 (N_19651,N_16752,N_16148);
or U19652 (N_19652,N_17367,N_17811);
or U19653 (N_19653,N_16736,N_16504);
and U19654 (N_19654,N_16000,N_16189);
xor U19655 (N_19655,N_16470,N_17328);
nand U19656 (N_19656,N_16499,N_16524);
and U19657 (N_19657,N_17005,N_16057);
or U19658 (N_19658,N_16091,N_17351);
nor U19659 (N_19659,N_17443,N_16112);
nand U19660 (N_19660,N_17296,N_16621);
xnor U19661 (N_19661,N_17966,N_17702);
nand U19662 (N_19662,N_16798,N_17354);
and U19663 (N_19663,N_17958,N_17589);
and U19664 (N_19664,N_17850,N_17641);
nand U19665 (N_19665,N_16229,N_17767);
xor U19666 (N_19666,N_17732,N_16424);
and U19667 (N_19667,N_17623,N_16974);
and U19668 (N_19668,N_16276,N_16571);
xnor U19669 (N_19669,N_17561,N_17244);
nand U19670 (N_19670,N_17878,N_17774);
nand U19671 (N_19671,N_16521,N_16245);
nand U19672 (N_19672,N_16471,N_17759);
or U19673 (N_19673,N_17875,N_17758);
nor U19674 (N_19674,N_17212,N_17018);
nand U19675 (N_19675,N_16777,N_16576);
xor U19676 (N_19676,N_17373,N_17854);
or U19677 (N_19677,N_16663,N_16196);
nor U19678 (N_19678,N_17850,N_17104);
and U19679 (N_19679,N_16059,N_16020);
and U19680 (N_19680,N_17452,N_17512);
nand U19681 (N_19681,N_16005,N_16553);
xor U19682 (N_19682,N_16182,N_16569);
nand U19683 (N_19683,N_16315,N_16379);
nor U19684 (N_19684,N_16606,N_16430);
or U19685 (N_19685,N_16337,N_16520);
nand U19686 (N_19686,N_16661,N_16328);
xor U19687 (N_19687,N_17046,N_17444);
or U19688 (N_19688,N_16611,N_16033);
xnor U19689 (N_19689,N_17490,N_17452);
and U19690 (N_19690,N_17445,N_16203);
or U19691 (N_19691,N_16807,N_17431);
nand U19692 (N_19692,N_16857,N_16899);
or U19693 (N_19693,N_16682,N_17626);
or U19694 (N_19694,N_17123,N_16868);
or U19695 (N_19695,N_17459,N_17807);
or U19696 (N_19696,N_16400,N_17717);
or U19697 (N_19697,N_17808,N_17072);
or U19698 (N_19698,N_17184,N_16547);
and U19699 (N_19699,N_17310,N_16695);
nor U19700 (N_19700,N_16046,N_17318);
or U19701 (N_19701,N_17257,N_16064);
nand U19702 (N_19702,N_16939,N_17422);
nand U19703 (N_19703,N_17043,N_16202);
and U19704 (N_19704,N_16025,N_17796);
and U19705 (N_19705,N_17998,N_17613);
and U19706 (N_19706,N_16654,N_17736);
xor U19707 (N_19707,N_16951,N_17263);
nand U19708 (N_19708,N_16270,N_16088);
or U19709 (N_19709,N_17518,N_17781);
xor U19710 (N_19710,N_16669,N_16503);
nand U19711 (N_19711,N_17388,N_16747);
or U19712 (N_19712,N_17591,N_17314);
or U19713 (N_19713,N_16296,N_17142);
nand U19714 (N_19714,N_16774,N_16898);
nor U19715 (N_19715,N_16829,N_17392);
xor U19716 (N_19716,N_17839,N_16962);
nand U19717 (N_19717,N_16521,N_16414);
nand U19718 (N_19718,N_16809,N_17894);
and U19719 (N_19719,N_17466,N_17508);
nand U19720 (N_19720,N_16508,N_17087);
nor U19721 (N_19721,N_17717,N_17006);
nand U19722 (N_19722,N_17372,N_17346);
and U19723 (N_19723,N_16677,N_17314);
and U19724 (N_19724,N_16725,N_17859);
nand U19725 (N_19725,N_17638,N_17969);
nor U19726 (N_19726,N_17859,N_16855);
xor U19727 (N_19727,N_16795,N_16432);
xor U19728 (N_19728,N_16208,N_17295);
nand U19729 (N_19729,N_17588,N_16477);
nand U19730 (N_19730,N_16792,N_17449);
or U19731 (N_19731,N_16975,N_16873);
xor U19732 (N_19732,N_16947,N_17722);
or U19733 (N_19733,N_17163,N_16311);
or U19734 (N_19734,N_16437,N_16049);
nor U19735 (N_19735,N_16483,N_16546);
nand U19736 (N_19736,N_17895,N_16412);
xnor U19737 (N_19737,N_17253,N_17989);
nor U19738 (N_19738,N_16812,N_16866);
nand U19739 (N_19739,N_16468,N_16155);
or U19740 (N_19740,N_16661,N_17935);
and U19741 (N_19741,N_16353,N_16152);
nand U19742 (N_19742,N_17239,N_16213);
nor U19743 (N_19743,N_16013,N_16084);
nor U19744 (N_19744,N_16969,N_16616);
and U19745 (N_19745,N_17450,N_17111);
or U19746 (N_19746,N_17861,N_16728);
xor U19747 (N_19747,N_17699,N_16809);
xnor U19748 (N_19748,N_17281,N_16330);
and U19749 (N_19749,N_17968,N_17326);
nand U19750 (N_19750,N_17966,N_17261);
nor U19751 (N_19751,N_16062,N_17050);
nand U19752 (N_19752,N_16962,N_17021);
or U19753 (N_19753,N_17179,N_16241);
and U19754 (N_19754,N_16037,N_16811);
or U19755 (N_19755,N_17881,N_16119);
and U19756 (N_19756,N_17054,N_17911);
and U19757 (N_19757,N_16596,N_17589);
or U19758 (N_19758,N_17405,N_17141);
xor U19759 (N_19759,N_17015,N_16276);
nand U19760 (N_19760,N_16031,N_17361);
xor U19761 (N_19761,N_16741,N_17691);
nor U19762 (N_19762,N_17251,N_17174);
nand U19763 (N_19763,N_17598,N_16992);
or U19764 (N_19764,N_16804,N_16755);
nand U19765 (N_19765,N_17511,N_16236);
xor U19766 (N_19766,N_17096,N_16338);
nand U19767 (N_19767,N_16432,N_16632);
or U19768 (N_19768,N_17611,N_16563);
nor U19769 (N_19769,N_17121,N_17924);
xnor U19770 (N_19770,N_16767,N_17439);
nor U19771 (N_19771,N_16543,N_16746);
and U19772 (N_19772,N_16390,N_16994);
nand U19773 (N_19773,N_16225,N_16654);
and U19774 (N_19774,N_17383,N_17553);
or U19775 (N_19775,N_16675,N_17432);
nor U19776 (N_19776,N_17938,N_17201);
or U19777 (N_19777,N_16971,N_17265);
or U19778 (N_19778,N_16899,N_16885);
and U19779 (N_19779,N_16365,N_16934);
or U19780 (N_19780,N_17382,N_17752);
and U19781 (N_19781,N_17246,N_17178);
xnor U19782 (N_19782,N_17264,N_17078);
or U19783 (N_19783,N_16825,N_17751);
xnor U19784 (N_19784,N_16834,N_17799);
nor U19785 (N_19785,N_16418,N_17354);
nand U19786 (N_19786,N_17657,N_16717);
nor U19787 (N_19787,N_17490,N_17868);
nor U19788 (N_19788,N_16934,N_16300);
nand U19789 (N_19789,N_16829,N_17616);
nand U19790 (N_19790,N_17767,N_16019);
and U19791 (N_19791,N_16213,N_16897);
xor U19792 (N_19792,N_16788,N_16398);
or U19793 (N_19793,N_16729,N_16972);
nor U19794 (N_19794,N_17904,N_16294);
nand U19795 (N_19795,N_17015,N_17883);
or U19796 (N_19796,N_16493,N_16537);
nor U19797 (N_19797,N_17648,N_16181);
nor U19798 (N_19798,N_17590,N_16443);
nand U19799 (N_19799,N_16309,N_17971);
xor U19800 (N_19800,N_16603,N_16091);
and U19801 (N_19801,N_17715,N_16821);
nor U19802 (N_19802,N_17040,N_17287);
xor U19803 (N_19803,N_17344,N_17655);
and U19804 (N_19804,N_17933,N_16054);
or U19805 (N_19805,N_17125,N_16833);
nor U19806 (N_19806,N_17371,N_16052);
xnor U19807 (N_19807,N_16135,N_17850);
or U19808 (N_19808,N_16661,N_16215);
nand U19809 (N_19809,N_16714,N_17707);
nor U19810 (N_19810,N_16758,N_16803);
or U19811 (N_19811,N_17947,N_17087);
xor U19812 (N_19812,N_16196,N_17572);
and U19813 (N_19813,N_16605,N_16671);
xor U19814 (N_19814,N_17973,N_17676);
or U19815 (N_19815,N_17915,N_16658);
and U19816 (N_19816,N_17130,N_16316);
nand U19817 (N_19817,N_16192,N_16296);
and U19818 (N_19818,N_17038,N_17740);
nand U19819 (N_19819,N_17091,N_16840);
xor U19820 (N_19820,N_16727,N_17901);
nand U19821 (N_19821,N_17108,N_17352);
xnor U19822 (N_19822,N_17711,N_16979);
xor U19823 (N_19823,N_16087,N_17692);
nor U19824 (N_19824,N_16795,N_17073);
or U19825 (N_19825,N_17856,N_17049);
nor U19826 (N_19826,N_17716,N_17965);
and U19827 (N_19827,N_17679,N_17917);
and U19828 (N_19828,N_16535,N_17406);
or U19829 (N_19829,N_16453,N_17597);
nor U19830 (N_19830,N_16622,N_16367);
and U19831 (N_19831,N_16236,N_17732);
or U19832 (N_19832,N_16905,N_17503);
or U19833 (N_19833,N_16097,N_16261);
xor U19834 (N_19834,N_16741,N_16585);
nor U19835 (N_19835,N_17898,N_17756);
or U19836 (N_19836,N_17026,N_16301);
xnor U19837 (N_19837,N_16229,N_17393);
nand U19838 (N_19838,N_17499,N_16217);
or U19839 (N_19839,N_17776,N_17674);
nand U19840 (N_19840,N_16818,N_17869);
nor U19841 (N_19841,N_16699,N_17328);
xor U19842 (N_19842,N_17016,N_16493);
nor U19843 (N_19843,N_17029,N_16430);
and U19844 (N_19844,N_16236,N_16853);
xor U19845 (N_19845,N_16952,N_17562);
xor U19846 (N_19846,N_17449,N_16338);
xnor U19847 (N_19847,N_16999,N_17978);
nor U19848 (N_19848,N_17242,N_16546);
and U19849 (N_19849,N_17885,N_17026);
and U19850 (N_19850,N_16464,N_16058);
and U19851 (N_19851,N_17423,N_17953);
nand U19852 (N_19852,N_16460,N_16662);
and U19853 (N_19853,N_16809,N_16268);
and U19854 (N_19854,N_16062,N_16329);
or U19855 (N_19855,N_16560,N_16104);
nand U19856 (N_19856,N_17270,N_16671);
nand U19857 (N_19857,N_17126,N_16431);
nand U19858 (N_19858,N_17420,N_16103);
or U19859 (N_19859,N_16490,N_17439);
xor U19860 (N_19860,N_16918,N_16492);
or U19861 (N_19861,N_17355,N_16853);
nor U19862 (N_19862,N_17771,N_16364);
or U19863 (N_19863,N_16566,N_17027);
nand U19864 (N_19864,N_16912,N_16355);
nor U19865 (N_19865,N_17251,N_17524);
or U19866 (N_19866,N_17713,N_16496);
and U19867 (N_19867,N_17873,N_17417);
or U19868 (N_19868,N_17522,N_17973);
xnor U19869 (N_19869,N_16730,N_17670);
nor U19870 (N_19870,N_17711,N_16140);
nand U19871 (N_19871,N_16186,N_16918);
nand U19872 (N_19872,N_17577,N_16416);
nor U19873 (N_19873,N_16751,N_17460);
xnor U19874 (N_19874,N_16464,N_17641);
xnor U19875 (N_19875,N_16311,N_16168);
or U19876 (N_19876,N_17266,N_16965);
and U19877 (N_19877,N_16241,N_17413);
and U19878 (N_19878,N_16669,N_16603);
or U19879 (N_19879,N_17129,N_16957);
nor U19880 (N_19880,N_17190,N_16017);
xnor U19881 (N_19881,N_16806,N_17355);
and U19882 (N_19882,N_17741,N_16924);
xor U19883 (N_19883,N_17950,N_17218);
xor U19884 (N_19884,N_16218,N_17102);
nor U19885 (N_19885,N_16020,N_16234);
nand U19886 (N_19886,N_16115,N_17674);
nand U19887 (N_19887,N_16283,N_16596);
nor U19888 (N_19888,N_17217,N_17617);
nand U19889 (N_19889,N_17098,N_16584);
xor U19890 (N_19890,N_17267,N_16173);
nand U19891 (N_19891,N_16028,N_16733);
and U19892 (N_19892,N_16377,N_17424);
nand U19893 (N_19893,N_17177,N_16614);
nand U19894 (N_19894,N_16479,N_17719);
or U19895 (N_19895,N_16754,N_16169);
and U19896 (N_19896,N_17410,N_16614);
or U19897 (N_19897,N_16667,N_17874);
xnor U19898 (N_19898,N_16258,N_17078);
xnor U19899 (N_19899,N_16488,N_17647);
or U19900 (N_19900,N_17790,N_16941);
nand U19901 (N_19901,N_17380,N_16117);
xnor U19902 (N_19902,N_17135,N_17957);
xor U19903 (N_19903,N_17118,N_17212);
and U19904 (N_19904,N_17221,N_17639);
nor U19905 (N_19905,N_17198,N_17719);
xnor U19906 (N_19906,N_17878,N_17670);
xnor U19907 (N_19907,N_17844,N_16815);
xnor U19908 (N_19908,N_17289,N_16683);
nor U19909 (N_19909,N_17512,N_17207);
nor U19910 (N_19910,N_17467,N_16346);
or U19911 (N_19911,N_16269,N_17646);
xnor U19912 (N_19912,N_16477,N_16313);
nor U19913 (N_19913,N_17659,N_17940);
nand U19914 (N_19914,N_17070,N_16709);
xnor U19915 (N_19915,N_17630,N_17108);
nand U19916 (N_19916,N_17544,N_17194);
nor U19917 (N_19917,N_17060,N_16911);
and U19918 (N_19918,N_16062,N_16737);
xnor U19919 (N_19919,N_17753,N_16365);
and U19920 (N_19920,N_17437,N_16800);
nand U19921 (N_19921,N_16324,N_17740);
and U19922 (N_19922,N_17350,N_16892);
nand U19923 (N_19923,N_17304,N_17174);
nor U19924 (N_19924,N_16282,N_17229);
and U19925 (N_19925,N_17618,N_16290);
xnor U19926 (N_19926,N_16918,N_16175);
nor U19927 (N_19927,N_17257,N_17176);
xnor U19928 (N_19928,N_16262,N_16399);
nand U19929 (N_19929,N_17865,N_17790);
nand U19930 (N_19930,N_17064,N_17076);
nor U19931 (N_19931,N_17481,N_17275);
xor U19932 (N_19932,N_17125,N_16184);
and U19933 (N_19933,N_16074,N_17809);
nor U19934 (N_19934,N_17602,N_17907);
nor U19935 (N_19935,N_17745,N_17242);
or U19936 (N_19936,N_17543,N_17339);
and U19937 (N_19937,N_16731,N_17444);
nand U19938 (N_19938,N_17878,N_17008);
xor U19939 (N_19939,N_16418,N_17176);
xnor U19940 (N_19940,N_16926,N_16380);
nor U19941 (N_19941,N_17894,N_16581);
and U19942 (N_19942,N_16702,N_16542);
or U19943 (N_19943,N_17488,N_17108);
or U19944 (N_19944,N_17510,N_16713);
and U19945 (N_19945,N_17141,N_17396);
nand U19946 (N_19946,N_16517,N_17215);
and U19947 (N_19947,N_16999,N_16386);
nor U19948 (N_19948,N_17591,N_17472);
or U19949 (N_19949,N_16972,N_17806);
nor U19950 (N_19950,N_17315,N_16814);
nor U19951 (N_19951,N_16966,N_16245);
nor U19952 (N_19952,N_17903,N_17690);
or U19953 (N_19953,N_17153,N_16698);
and U19954 (N_19954,N_17180,N_17170);
nor U19955 (N_19955,N_17735,N_16851);
and U19956 (N_19956,N_16870,N_16847);
nand U19957 (N_19957,N_16891,N_16762);
nor U19958 (N_19958,N_17814,N_16338);
or U19959 (N_19959,N_17739,N_17330);
nand U19960 (N_19960,N_17779,N_16706);
nand U19961 (N_19961,N_17022,N_16611);
and U19962 (N_19962,N_16830,N_17160);
or U19963 (N_19963,N_17199,N_17060);
or U19964 (N_19964,N_17390,N_16356);
nor U19965 (N_19965,N_16636,N_17982);
xnor U19966 (N_19966,N_17821,N_17172);
or U19967 (N_19967,N_17445,N_17277);
nand U19968 (N_19968,N_17185,N_17316);
nor U19969 (N_19969,N_16185,N_16817);
nand U19970 (N_19970,N_16907,N_17194);
xor U19971 (N_19971,N_17375,N_16311);
nand U19972 (N_19972,N_17978,N_17988);
nor U19973 (N_19973,N_17573,N_17044);
or U19974 (N_19974,N_17833,N_17248);
or U19975 (N_19975,N_16787,N_16509);
nand U19976 (N_19976,N_17405,N_16083);
or U19977 (N_19977,N_17392,N_16891);
xor U19978 (N_19978,N_16614,N_16678);
nor U19979 (N_19979,N_17520,N_17560);
nand U19980 (N_19980,N_17714,N_16415);
and U19981 (N_19981,N_16126,N_17762);
nor U19982 (N_19982,N_17269,N_17133);
or U19983 (N_19983,N_16101,N_17857);
nand U19984 (N_19984,N_16549,N_17126);
and U19985 (N_19985,N_16988,N_16716);
xnor U19986 (N_19986,N_17490,N_17509);
or U19987 (N_19987,N_16738,N_17044);
or U19988 (N_19988,N_16773,N_16525);
nor U19989 (N_19989,N_17768,N_16597);
or U19990 (N_19990,N_17005,N_17756);
nor U19991 (N_19991,N_17367,N_16399);
xnor U19992 (N_19992,N_16663,N_16031);
and U19993 (N_19993,N_17352,N_16884);
nor U19994 (N_19994,N_16232,N_17306);
xor U19995 (N_19995,N_16885,N_17050);
nor U19996 (N_19996,N_16418,N_16170);
nor U19997 (N_19997,N_16095,N_17578);
nand U19998 (N_19998,N_16722,N_16912);
nand U19999 (N_19999,N_17396,N_16772);
nor U20000 (N_20000,N_18044,N_19999);
and U20001 (N_20001,N_18474,N_19328);
nor U20002 (N_20002,N_19067,N_18369);
xnor U20003 (N_20003,N_18439,N_18705);
and U20004 (N_20004,N_18921,N_18870);
xor U20005 (N_20005,N_18942,N_19831);
xnor U20006 (N_20006,N_18106,N_18946);
or U20007 (N_20007,N_18438,N_18774);
nand U20008 (N_20008,N_18624,N_18547);
nand U20009 (N_20009,N_18877,N_19962);
nor U20010 (N_20010,N_19174,N_18536);
and U20011 (N_20011,N_19112,N_19772);
and U20012 (N_20012,N_19062,N_19269);
xnor U20013 (N_20013,N_19037,N_19776);
or U20014 (N_20014,N_18286,N_18113);
nand U20015 (N_20015,N_19353,N_18288);
nand U20016 (N_20016,N_18268,N_18794);
and U20017 (N_20017,N_19770,N_19581);
and U20018 (N_20018,N_19003,N_19424);
xor U20019 (N_20019,N_19966,N_19885);
xor U20020 (N_20020,N_19171,N_19431);
and U20021 (N_20021,N_19276,N_18267);
and U20022 (N_20022,N_18737,N_18098);
nor U20023 (N_20023,N_18460,N_19050);
xor U20024 (N_20024,N_18445,N_19463);
nand U20025 (N_20025,N_19822,N_19702);
nand U20026 (N_20026,N_19231,N_19645);
xnor U20027 (N_20027,N_18918,N_18147);
or U20028 (N_20028,N_19049,N_19658);
nand U20029 (N_20029,N_18763,N_19586);
or U20030 (N_20030,N_18433,N_19677);
or U20031 (N_20031,N_19434,N_18564);
xnor U20032 (N_20032,N_19198,N_18152);
and U20033 (N_20033,N_18049,N_18718);
xnor U20034 (N_20034,N_18879,N_19116);
xor U20035 (N_20035,N_18404,N_19107);
and U20036 (N_20036,N_18487,N_18990);
nand U20037 (N_20037,N_18695,N_18694);
and U20038 (N_20038,N_19407,N_19460);
or U20039 (N_20039,N_19259,N_18191);
nand U20040 (N_20040,N_18262,N_18137);
nand U20041 (N_20041,N_18804,N_19135);
nor U20042 (N_20042,N_18349,N_19488);
and U20043 (N_20043,N_19388,N_19444);
nand U20044 (N_20044,N_18760,N_19589);
or U20045 (N_20045,N_19871,N_18999);
nor U20046 (N_20046,N_19010,N_19760);
or U20047 (N_20047,N_18724,N_18340);
or U20048 (N_20048,N_18593,N_18220);
xnor U20049 (N_20049,N_19859,N_18630);
or U20050 (N_20050,N_18689,N_19004);
or U20051 (N_20051,N_19188,N_19143);
and U20052 (N_20052,N_19798,N_18135);
nor U20053 (N_20053,N_19949,N_18308);
xor U20054 (N_20054,N_18443,N_18352);
and U20055 (N_20055,N_18755,N_19857);
and U20056 (N_20056,N_18773,N_18463);
xor U20057 (N_20057,N_19638,N_18780);
xnor U20058 (N_20058,N_19138,N_19780);
or U20059 (N_20059,N_19425,N_18577);
nor U20060 (N_20060,N_18754,N_18895);
nand U20061 (N_20061,N_18112,N_18298);
nand U20062 (N_20062,N_18775,N_18448);
and U20063 (N_20063,N_19142,N_19741);
xor U20064 (N_20064,N_19855,N_19311);
and U20065 (N_20065,N_19828,N_19480);
or U20066 (N_20066,N_19244,N_19453);
nor U20067 (N_20067,N_19367,N_19160);
nand U20068 (N_20068,N_18528,N_19342);
or U20069 (N_20069,N_19181,N_19764);
xnor U20070 (N_20070,N_18243,N_18567);
nor U20071 (N_20071,N_19560,N_19291);
or U20072 (N_20072,N_18249,N_18892);
or U20073 (N_20073,N_19043,N_19597);
nand U20074 (N_20074,N_18465,N_18255);
xor U20075 (N_20075,N_19118,N_19787);
nand U20076 (N_20076,N_18066,N_19528);
xnor U20077 (N_20077,N_19700,N_19295);
nor U20078 (N_20078,N_19646,N_19614);
nor U20079 (N_20079,N_18477,N_19921);
and U20080 (N_20080,N_18893,N_18708);
or U20081 (N_20081,N_19662,N_18955);
or U20082 (N_20082,N_18852,N_18886);
and U20083 (N_20083,N_19249,N_18618);
or U20084 (N_20084,N_18123,N_19555);
xor U20085 (N_20085,N_19268,N_18983);
nor U20086 (N_20086,N_18684,N_19066);
or U20087 (N_20087,N_18525,N_18681);
xor U20088 (N_20088,N_19930,N_18508);
nor U20089 (N_20089,N_18746,N_18292);
xor U20090 (N_20090,N_18411,N_18576);
or U20091 (N_20091,N_19364,N_19647);
and U20092 (N_20092,N_18813,N_18102);
xor U20093 (N_20093,N_19209,N_19551);
and U20094 (N_20094,N_18984,N_19925);
and U20095 (N_20095,N_19687,N_18712);
and U20096 (N_20096,N_19515,N_18876);
nor U20097 (N_20097,N_18207,N_19001);
nor U20098 (N_20098,N_19162,N_19907);
or U20099 (N_20099,N_18836,N_19680);
or U20100 (N_20100,N_18166,N_18851);
or U20101 (N_20101,N_18764,N_19455);
nor U20102 (N_20102,N_19296,N_18998);
xnor U20103 (N_20103,N_19409,N_19566);
or U20104 (N_20104,N_18041,N_18076);
xor U20105 (N_20105,N_19771,N_18840);
nor U20106 (N_20106,N_19029,N_19018);
or U20107 (N_20107,N_19876,N_18226);
nand U20108 (N_20108,N_19232,N_18731);
or U20109 (N_20109,N_18488,N_19493);
xor U20110 (N_20110,N_19158,N_19071);
or U20111 (N_20111,N_19681,N_19627);
and U20112 (N_20112,N_18301,N_18874);
xnor U20113 (N_20113,N_18186,N_19334);
xnor U20114 (N_20114,N_18108,N_19304);
or U20115 (N_20115,N_19452,N_18093);
nand U20116 (N_20116,N_18450,N_18252);
or U20117 (N_20117,N_19090,N_18168);
nand U20118 (N_20118,N_19078,N_19571);
xor U20119 (N_20119,N_18165,N_19746);
and U20120 (N_20120,N_19222,N_18073);
nand U20121 (N_20121,N_18502,N_19752);
nand U20122 (N_20122,N_18526,N_19239);
or U20123 (N_20123,N_19149,N_19631);
nand U20124 (N_20124,N_18675,N_18100);
xnor U20125 (N_20125,N_18274,N_19385);
and U20126 (N_20126,N_19192,N_18784);
nand U20127 (N_20127,N_18406,N_19405);
nor U20128 (N_20128,N_18745,N_18189);
nor U20129 (N_20129,N_18659,N_18825);
or U20130 (N_20130,N_18674,N_18619);
and U20131 (N_20131,N_18798,N_19319);
xnor U20132 (N_20132,N_19769,N_19306);
and U20133 (N_20133,N_18492,N_19469);
and U20134 (N_20134,N_19387,N_18936);
nor U20135 (N_20135,N_19114,N_19301);
and U20136 (N_20136,N_18235,N_18322);
and U20137 (N_20137,N_18177,N_19689);
nand U20138 (N_20138,N_19950,N_19877);
nor U20139 (N_20139,N_19710,N_19499);
and U20140 (N_20140,N_19747,N_18699);
nor U20141 (N_20141,N_18449,N_19755);
or U20142 (N_20142,N_18738,N_19056);
and U20143 (N_20143,N_19817,N_18201);
xor U20144 (N_20144,N_18361,N_18461);
xnor U20145 (N_20145,N_19363,N_18723);
nor U20146 (N_20146,N_19185,N_19894);
or U20147 (N_20147,N_19781,N_19314);
xnor U20148 (N_20148,N_18582,N_19691);
nor U20149 (N_20149,N_18812,N_18862);
or U20150 (N_20150,N_18617,N_19603);
or U20151 (N_20151,N_18398,N_18698);
nand U20152 (N_20152,N_19718,N_18493);
xor U20153 (N_20153,N_18640,N_18966);
xnor U20154 (N_20154,N_18861,N_18590);
and U20155 (N_20155,N_18293,N_18822);
nor U20156 (N_20156,N_18156,N_19380);
xnor U20157 (N_20157,N_18560,N_18107);
and U20158 (N_20158,N_18504,N_19795);
xor U20159 (N_20159,N_18848,N_19823);
nor U20160 (N_20160,N_19454,N_19240);
nor U20161 (N_20161,N_19176,N_18383);
xor U20162 (N_20162,N_19500,N_18552);
nor U20163 (N_20163,N_18683,N_19675);
xor U20164 (N_20164,N_19663,N_18482);
nor U20165 (N_20165,N_19038,N_18557);
nand U20166 (N_20166,N_19322,N_18407);
or U20167 (N_20167,N_18602,N_18163);
nand U20168 (N_20168,N_19613,N_19882);
xor U20169 (N_20169,N_18896,N_18522);
or U20170 (N_20170,N_18070,N_18200);
or U20171 (N_20171,N_18103,N_19208);
xor U20172 (N_20172,N_18996,N_18595);
nor U20173 (N_20173,N_19046,N_18769);
xnor U20174 (N_20174,N_19419,N_18062);
nor U20175 (N_20175,N_19835,N_19292);
nand U20176 (N_20176,N_19890,N_19624);
xnor U20177 (N_20177,N_18133,N_18359);
nor U20178 (N_20178,N_19262,N_18647);
nand U20179 (N_20179,N_18673,N_18434);
or U20180 (N_20180,N_19525,N_18136);
xnor U20181 (N_20181,N_18815,N_19811);
xor U20182 (N_20182,N_18722,N_18141);
nand U20183 (N_20183,N_18211,N_18223);
and U20184 (N_20184,N_19006,N_19970);
or U20185 (N_20185,N_19852,N_19895);
nor U20186 (N_20186,N_18266,N_19836);
nor U20187 (N_20187,N_18279,N_19111);
and U20188 (N_20188,N_18923,N_18858);
xnor U20189 (N_20189,N_18244,N_19355);
nor U20190 (N_20190,N_18765,N_18909);
xor U20191 (N_20191,N_19850,N_18258);
nand U20192 (N_20192,N_19507,N_19509);
xnor U20193 (N_20193,N_18097,N_19375);
xnor U20194 (N_20194,N_19720,N_18426);
or U20195 (N_20195,N_18654,N_19540);
nand U20196 (N_20196,N_19829,N_19513);
and U20197 (N_20197,N_19327,N_18700);
xnor U20198 (N_20198,N_18187,N_19651);
nor U20199 (N_20199,N_19124,N_19941);
nand U20200 (N_20200,N_19806,N_18803);
xnor U20201 (N_20201,N_19219,N_18238);
and U20202 (N_20202,N_19341,N_18037);
xor U20203 (N_20203,N_18489,N_18767);
and U20204 (N_20204,N_18117,N_18190);
and U20205 (N_20205,N_19481,N_19803);
nand U20206 (N_20206,N_19931,N_18579);
or U20207 (N_20207,N_19640,N_19261);
and U20208 (N_20208,N_19115,N_19315);
nor U20209 (N_20209,N_18598,N_18132);
and U20210 (N_20210,N_18585,N_19035);
or U20211 (N_20211,N_19072,N_19478);
or U20212 (N_20212,N_19556,N_19552);
nand U20213 (N_20213,N_19081,N_19754);
and U20214 (N_20214,N_19462,N_18328);
xor U20215 (N_20215,N_19329,N_18029);
nand U20216 (N_20216,N_19523,N_18641);
nor U20217 (N_20217,N_18897,N_19674);
or U20218 (N_20218,N_19473,N_18912);
or U20219 (N_20219,N_18545,N_18417);
nor U20220 (N_20220,N_18204,N_19669);
nand U20221 (N_20221,N_19022,N_19553);
nand U20222 (N_20222,N_18360,N_18196);
and U20223 (N_20223,N_18458,N_19324);
or U20224 (N_20224,N_18134,N_18437);
nor U20225 (N_20225,N_19935,N_18973);
nor U20226 (N_20226,N_18748,N_18884);
and U20227 (N_20227,N_18807,N_19830);
or U20228 (N_20228,N_18086,N_18563);
and U20229 (N_20229,N_19492,N_18986);
nor U20230 (N_20230,N_19336,N_18741);
nor U20231 (N_20231,N_19740,N_19709);
xor U20232 (N_20232,N_19542,N_18188);
xnor U20233 (N_20233,N_19800,N_18385);
xnor U20234 (N_20234,N_18727,N_18372);
xor U20235 (N_20235,N_19748,N_19007);
and U20236 (N_20236,N_18074,N_19359);
nor U20237 (N_20237,N_19750,N_18843);
nand U20238 (N_20238,N_19578,N_19153);
or U20239 (N_20239,N_18664,N_19574);
nand U20240 (N_20240,N_19888,N_18703);
xor U20241 (N_20241,N_18922,N_19526);
nor U20242 (N_20242,N_18580,N_18149);
or U20243 (N_20243,N_19957,N_18625);
xnor U20244 (N_20244,N_18900,N_19942);
nand U20245 (N_20245,N_18957,N_19190);
nor U20246 (N_20246,N_19096,N_19456);
and U20247 (N_20247,N_19602,N_19002);
and U20248 (N_20248,N_19634,N_18272);
and U20249 (N_20249,N_18658,N_18033);
and U20250 (N_20250,N_18915,N_18393);
nor U20251 (N_20251,N_19896,N_19486);
xor U20252 (N_20252,N_19694,N_18325);
nand U20253 (N_20253,N_18549,N_18758);
xor U20254 (N_20254,N_19101,N_18820);
nor U20255 (N_20255,N_18729,N_18838);
nand U20256 (N_20256,N_18311,N_18048);
nor U20257 (N_20257,N_19796,N_19713);
nor U20258 (N_20258,N_18985,N_18358);
and U20259 (N_20259,N_19053,N_19382);
xnor U20260 (N_20260,N_19904,N_19177);
nor U20261 (N_20261,N_19719,N_19260);
xnor U20262 (N_20262,N_18863,N_19938);
or U20263 (N_20263,N_18115,N_19994);
nand U20264 (N_20264,N_19576,N_18356);
xnor U20265 (N_20265,N_19333,N_19762);
or U20266 (N_20266,N_19263,N_18339);
nand U20267 (N_20267,N_18122,N_19641);
and U20268 (N_20268,N_19370,N_18092);
nand U20269 (N_20269,N_19287,N_18779);
and U20270 (N_20270,N_19607,N_19502);
xnor U20271 (N_20271,N_19695,N_18534);
and U20272 (N_20272,N_19042,N_19841);
nor U20273 (N_20273,N_19435,N_19496);
xor U20274 (N_20274,N_19622,N_18987);
nor U20275 (N_20275,N_19923,N_19178);
nor U20276 (N_20276,N_18316,N_18941);
xor U20277 (N_20277,N_18656,N_19832);
xor U20278 (N_20278,N_19632,N_19693);
and U20279 (N_20279,N_18786,N_19983);
or U20280 (N_20280,N_19365,N_18629);
xor U20281 (N_20281,N_18355,N_18085);
nand U20282 (N_20282,N_18256,N_19620);
xnor U20283 (N_20283,N_18761,N_19459);
or U20284 (N_20284,N_18424,N_19298);
nor U20285 (N_20285,N_19110,N_19723);
nor U20286 (N_20286,N_18828,N_19784);
nor U20287 (N_20287,N_18982,N_18559);
or U20288 (N_20288,N_19751,N_19237);
xor U20289 (N_20289,N_18883,N_18665);
nor U20290 (N_20290,N_18390,N_19494);
or U20291 (N_20291,N_19963,N_18890);
and U20292 (N_20292,N_18173,N_18759);
nand U20293 (N_20293,N_18846,N_18179);
xnor U20294 (N_20294,N_18975,N_19608);
or U20295 (N_20295,N_19075,N_18792);
nand U20296 (N_20296,N_18533,N_19168);
xor U20297 (N_20297,N_19182,N_18193);
nand U20298 (N_20298,N_19057,N_18739);
and U20299 (N_20299,N_19959,N_19362);
and U20300 (N_20300,N_19320,N_18965);
or U20301 (N_20301,N_19025,N_19792);
nor U20302 (N_20302,N_19973,N_18806);
and U20303 (N_20303,N_18199,N_19449);
and U20304 (N_20304,N_18810,N_18752);
and U20305 (N_20305,N_19349,N_19340);
and U20306 (N_20306,N_19476,N_18198);
nand U20307 (N_20307,N_19849,N_19443);
xor U20308 (N_20308,N_19736,N_18027);
nand U20309 (N_20309,N_19582,N_18735);
xor U20310 (N_20310,N_19284,N_18976);
or U20311 (N_20311,N_19186,N_19428);
nand U20312 (N_20312,N_18725,N_19332);
xnor U20313 (N_20313,N_19898,N_18704);
nand U20314 (N_20314,N_18970,N_19475);
nand U20315 (N_20315,N_19401,N_19753);
nor U20316 (N_20316,N_19863,N_18910);
nand U20317 (N_20317,N_18878,N_18042);
and U20318 (N_20318,N_18370,N_19733);
xnor U20319 (N_20319,N_18081,N_19878);
or U20320 (N_20320,N_18818,N_18904);
nor U20321 (N_20321,N_18180,N_19900);
nand U20322 (N_20322,N_18270,N_19464);
and U20323 (N_20323,N_19778,N_19583);
nand U20324 (N_20324,N_19157,N_18969);
or U20325 (N_20325,N_18264,N_19837);
nor U20326 (N_20326,N_19732,N_18587);
xor U20327 (N_20327,N_18194,N_18344);
and U20328 (N_20328,N_19163,N_18195);
nor U20329 (N_20329,N_19164,N_19381);
nand U20330 (N_20330,N_18206,N_19965);
and U20331 (N_20331,N_19285,N_19908);
and U20332 (N_20332,N_19791,N_18109);
and U20333 (N_20333,N_19442,N_19678);
nor U20334 (N_20334,N_19672,N_18202);
nand U20335 (N_20335,N_19580,N_19212);
nand U20336 (N_20336,N_18906,N_18105);
and U20337 (N_20337,N_19785,N_18523);
and U20338 (N_20338,N_18594,N_19399);
xor U20339 (N_20339,N_18138,N_19313);
nor U20340 (N_20340,N_19846,N_18399);
and U20341 (N_20341,N_19601,N_19977);
nand U20342 (N_20342,N_18480,N_18591);
nand U20343 (N_20343,N_18413,N_18857);
and U20344 (N_20344,N_19708,N_18320);
nor U20345 (N_20345,N_18678,N_19000);
and U20346 (N_20346,N_19703,N_19490);
xnor U20347 (N_20347,N_18979,N_18470);
nor U20348 (N_20348,N_18733,N_19447);
or U20349 (N_20349,N_19044,N_18155);
nand U20350 (N_20350,N_18373,N_19482);
and U20351 (N_20351,N_19549,N_18510);
and U20352 (N_20352,N_19737,N_18351);
xnor U20353 (N_20353,N_18333,N_19570);
xor U20354 (N_20354,N_18079,N_19100);
nor U20355 (N_20355,N_18289,N_19848);
xnor U20356 (N_20356,N_19953,N_19120);
and U20357 (N_20357,N_18422,N_19531);
xnor U20358 (N_20358,N_19166,N_18063);
or U20359 (N_20359,N_18307,N_18467);
or U20360 (N_20360,N_18428,N_19972);
and U20361 (N_20361,N_18677,N_19061);
xnor U20362 (N_20362,N_19400,N_18475);
and U20363 (N_20363,N_18309,N_18484);
nand U20364 (N_20364,N_18254,N_18012);
nor U20365 (N_20365,N_19465,N_18860);
or U20366 (N_20366,N_18844,N_19517);
and U20367 (N_20367,N_19406,N_19416);
xnor U20368 (N_20368,N_19881,N_18964);
or U20369 (N_20369,N_19151,N_19346);
or U20370 (N_20370,N_18817,N_19954);
nand U20371 (N_20371,N_18571,N_19202);
nand U20372 (N_20372,N_19461,N_19532);
nand U20373 (N_20373,N_18521,N_19105);
and U20374 (N_20374,N_18535,N_19193);
nand U20375 (N_20375,N_18651,N_19706);
xor U20376 (N_20376,N_19592,N_19643);
and U20377 (N_20377,N_19901,N_19217);
xnor U20378 (N_20378,N_19246,N_19724);
or U20379 (N_20379,N_19749,N_19548);
nand U20380 (N_20380,N_19595,N_18887);
or U20381 (N_20381,N_18281,N_19477);
or U20382 (N_20382,N_19150,N_18430);
and U20383 (N_20383,N_18781,N_18770);
xor U20384 (N_20384,N_18217,N_19816);
xnor U20385 (N_20385,N_18635,N_19130);
and U20386 (N_20386,N_18575,N_18690);
nor U20387 (N_20387,N_18816,N_18365);
or U20388 (N_20388,N_19253,N_18153);
nor U20389 (N_20389,N_18772,N_18130);
nor U20390 (N_20390,N_19248,N_19758);
or U20391 (N_20391,N_18253,N_19238);
and U20392 (N_20392,N_18544,N_19225);
xor U20393 (N_20393,N_18078,N_18671);
nor U20394 (N_20394,N_18888,N_18701);
nand U20395 (N_20395,N_18558,N_18284);
xor U20396 (N_20396,N_19541,N_19682);
nand U20397 (N_20397,N_19446,N_19169);
nor U20398 (N_20398,N_18621,N_18329);
or U20399 (N_20399,N_19412,N_18553);
xor U20400 (N_20400,N_19893,N_19373);
or U20401 (N_20401,N_18150,N_18080);
and U20402 (N_20402,N_19676,N_19300);
nand U20403 (N_20403,N_18962,N_19489);
xnor U20404 (N_20404,N_18231,N_18929);
xor U20405 (N_20405,N_18084,N_19255);
and U20406 (N_20406,N_18000,N_19550);
xnor U20407 (N_20407,N_18511,N_19670);
nand U20408 (N_20408,N_18176,N_19666);
nand U20409 (N_20409,N_18148,N_18315);
nand U20410 (N_20410,N_18436,N_19922);
xnor U20411 (N_20411,N_19199,N_18916);
nor U20412 (N_20412,N_19985,N_19191);
xnor U20413 (N_20413,N_18788,N_18364);
or U20414 (N_20414,N_18007,N_18660);
xnor U20415 (N_20415,N_18043,N_19064);
xor U20416 (N_20416,N_19247,N_18959);
and U20417 (N_20417,N_19865,N_19854);
and U20418 (N_20418,N_18599,N_18911);
and U20419 (N_20419,N_18841,N_18757);
nor U20420 (N_20420,N_18403,N_18686);
or U20421 (N_20421,N_19099,N_19673);
and U20422 (N_20422,N_18299,N_18350);
nand U20423 (N_20423,N_18010,N_18503);
nor U20424 (N_20424,N_19369,N_18055);
and U20425 (N_20425,N_19827,N_18958);
nand U20426 (N_20426,N_18023,N_19390);
nand U20427 (N_20427,N_19014,N_19266);
nand U20428 (N_20428,N_18913,N_19082);
xnor U20429 (N_20429,N_19273,N_18490);
or U20430 (N_20430,N_18127,N_19979);
nand U20431 (N_20431,N_18090,N_18456);
and U20432 (N_20432,N_18072,N_18732);
nor U20433 (N_20433,N_19448,N_19964);
xor U20434 (N_20434,N_19402,N_19630);
or U20435 (N_20435,N_19080,N_18405);
xnor U20436 (N_20436,N_18357,N_18494);
and U20437 (N_20437,N_19794,N_18295);
and U20438 (N_20438,N_19906,N_18145);
and U20439 (N_20439,N_19783,N_18795);
xor U20440 (N_20440,N_18291,N_18920);
nor U20441 (N_20441,N_19372,N_19122);
nor U20442 (N_20442,N_18940,N_18605);
or U20443 (N_20443,N_19184,N_19495);
xnor U20444 (N_20444,N_19577,N_19487);
nor U20445 (N_20445,N_18688,N_19361);
or U20446 (N_20446,N_19197,N_19337);
nand U20447 (N_20447,N_18110,N_18622);
nand U20448 (N_20448,N_18290,N_19913);
xnor U20449 (N_20449,N_19637,N_18069);
nand U20450 (N_20450,N_18319,N_19230);
nor U20451 (N_20451,N_19521,N_18766);
nor U20452 (N_20452,N_18856,N_18230);
and U20453 (N_20453,N_19512,N_18551);
and U20454 (N_20454,N_18294,N_18971);
nor U20455 (N_20455,N_19290,N_18991);
xor U20456 (N_20456,N_18014,N_18586);
xnor U20457 (N_20457,N_18431,N_19330);
and U20458 (N_20458,N_19861,N_18019);
or U20459 (N_20459,N_18039,N_19012);
nand U20460 (N_20460,N_18937,N_19216);
nor U20461 (N_20461,N_18919,N_19221);
or U20462 (N_20462,N_19429,N_19123);
or U20463 (N_20463,N_19383,N_18989);
nand U20464 (N_20464,N_18992,N_19413);
nor U20465 (N_20465,N_18516,N_19927);
nand U20466 (N_20466,N_19339,N_19030);
xor U20467 (N_20467,N_18185,N_19782);
nand U20468 (N_20468,N_18444,N_19939);
nor U20469 (N_20469,N_19524,N_18047);
nand U20470 (N_20470,N_19505,N_19932);
and U20471 (N_20471,N_18974,N_19699);
or U20472 (N_20472,N_18378,N_18050);
nand U20473 (N_20473,N_19376,N_18866);
nand U20474 (N_20474,N_19839,N_19704);
or U20475 (N_20475,N_18901,N_18696);
and U20476 (N_20476,N_18347,N_18616);
or U20477 (N_20477,N_18057,N_18053);
and U20478 (N_20478,N_18539,N_18184);
or U20479 (N_20479,N_18607,N_18570);
xor U20480 (N_20480,N_19267,N_19205);
nor U20481 (N_20481,N_19036,N_18823);
xnor U20482 (N_20482,N_18692,N_18046);
xnor U20483 (N_20483,N_19104,N_19611);
or U20484 (N_20484,N_18853,N_18013);
nand U20485 (N_20485,N_18022,N_18239);
xor U20486 (N_20486,N_19229,N_18330);
nand U20487 (N_20487,N_18945,N_19154);
and U20488 (N_20488,N_18483,N_19201);
and U20489 (N_20489,N_19529,N_19270);
xnor U20490 (N_20490,N_19251,N_18143);
nand U20491 (N_20491,N_19305,N_18652);
nor U20492 (N_20492,N_19996,N_19048);
nand U20493 (N_20493,N_18608,N_18719);
nand U20494 (N_20494,N_19590,N_18248);
and U20495 (N_20495,N_18847,N_19874);
nor U20496 (N_20496,N_18960,N_19498);
nor U20497 (N_20497,N_19520,N_19879);
xnor U20498 (N_20498,N_18953,N_18233);
nor U20499 (N_20499,N_18697,N_18620);
nand U20500 (N_20500,N_19224,N_18026);
nor U20501 (N_20501,N_18574,N_18905);
or U20502 (N_20502,N_18814,N_19392);
nor U20503 (N_20503,N_18596,N_18229);
or U20504 (N_20504,N_19833,N_18051);
nand U20505 (N_20505,N_19605,N_18059);
or U20506 (N_20506,N_19812,N_19858);
xor U20507 (N_20507,N_18855,N_18031);
and U20508 (N_20508,N_19968,N_18353);
xor U20509 (N_20509,N_19639,N_19288);
xnor U20510 (N_20510,N_19427,N_18395);
xor U20511 (N_20511,N_18245,N_18182);
xor U20512 (N_20512,N_19289,N_18015);
nand U20513 (N_20513,N_19310,N_18710);
xor U20514 (N_20514,N_18386,N_19420);
nand U20515 (N_20515,N_19335,N_19196);
xnor U20516 (N_20516,N_18834,N_19187);
and U20517 (N_20517,N_19137,N_19027);
nor U20518 (N_20518,N_19819,N_19623);
and U20519 (N_20519,N_19629,N_18583);
nand U20520 (N_20520,N_18627,N_19148);
nor U20521 (N_20521,N_18902,N_19739);
or U20522 (N_20522,N_19068,N_18777);
xnor U20523 (N_20523,N_19374,N_19766);
nor U20524 (N_20524,N_18327,N_18715);
or U20525 (N_20525,N_18342,N_18091);
nor U20526 (N_20526,N_18400,N_18396);
or U20527 (N_20527,N_19411,N_18016);
nand U20528 (N_20528,N_19960,N_19033);
xor U20529 (N_20529,N_19585,N_19325);
or U20530 (N_20530,N_18332,N_19562);
nor U20531 (N_20531,N_18183,N_19656);
nand U20532 (N_20532,N_18939,N_19474);
nand U20533 (N_20533,N_18529,N_19019);
or U20534 (N_20534,N_18845,N_19307);
or U20535 (N_20535,N_18837,N_19272);
or U20536 (N_20536,N_18935,N_18131);
nor U20537 (N_20537,N_18273,N_18161);
or U20538 (N_20538,N_19089,N_19910);
nor U20539 (N_20539,N_19810,N_18011);
nand U20540 (N_20540,N_19055,N_19648);
or U20541 (N_20541,N_19527,N_19323);
xnor U20542 (N_20542,N_19936,N_19023);
or U20543 (N_20543,N_18337,N_19626);
xnor U20544 (N_20544,N_19534,N_18144);
nand U20545 (N_20545,N_18832,N_19093);
nor U20546 (N_20546,N_18121,N_19357);
nand U20547 (N_20547,N_19257,N_18214);
and U20548 (N_20548,N_18657,N_19696);
nand U20549 (N_20549,N_19020,N_19155);
and U20550 (N_20550,N_19617,N_19086);
nand U20551 (N_20551,N_18821,N_19711);
nor U20552 (N_20552,N_18572,N_19206);
and U20553 (N_20553,N_19351,N_18280);
nand U20554 (N_20554,N_19873,N_18943);
nand U20555 (N_20555,N_18499,N_19657);
nor U20556 (N_20556,N_19554,N_19133);
nand U20557 (N_20557,N_19379,N_19993);
nand U20558 (N_20558,N_18082,N_19085);
or U20559 (N_20559,N_19073,N_18213);
nor U20560 (N_20560,N_19914,N_18303);
and U20561 (N_20561,N_19514,N_19271);
nand U20562 (N_20562,N_18800,N_19956);
nand U20563 (N_20563,N_18776,N_19141);
xnor U20564 (N_20564,N_18172,N_19604);
xor U20565 (N_20565,N_19466,N_19761);
nor U20566 (N_20566,N_18568,N_18783);
nand U20567 (N_20567,N_19200,N_19485);
xor U20568 (N_20568,N_19911,N_19790);
and U20569 (N_20569,N_19126,N_18524);
nor U20570 (N_20570,N_18067,N_18116);
nand U20571 (N_20571,N_18471,N_19242);
nand U20572 (N_20572,N_19536,N_19843);
nand U20573 (N_20573,N_18676,N_19293);
xnor U20574 (N_20574,N_18614,N_18285);
nor U20575 (N_20575,N_19978,N_19113);
or U20576 (N_20576,N_18881,N_19660);
or U20577 (N_20577,N_19692,N_18397);
nand U20578 (N_20578,N_18197,N_18453);
xnor U20579 (N_20579,N_18415,N_19279);
nor U20580 (N_20580,N_19805,N_18030);
xor U20581 (N_20581,N_19432,N_18334);
nor U20582 (N_20582,N_19844,N_18561);
or U20583 (N_20583,N_18251,N_18867);
nand U20584 (N_20584,N_18429,N_18466);
xnor U20585 (N_20585,N_19880,N_19450);
and U20586 (N_20586,N_18446,N_18017);
or U20587 (N_20587,N_18476,N_19032);
nand U20588 (N_20588,N_18653,N_18597);
nand U20589 (N_20589,N_18392,N_18645);
xor U20590 (N_20590,N_18721,N_18025);
and U20591 (N_20591,N_18859,N_19228);
and U20592 (N_20592,N_19483,N_19779);
nand U20593 (N_20593,N_18178,N_19568);
nor U20594 (N_20594,N_19902,N_18882);
xor U20595 (N_20595,N_19087,N_19134);
nor U20596 (N_20596,N_18125,N_18164);
or U20597 (N_20597,N_19884,N_18237);
nor U20598 (N_20598,N_18793,N_18040);
and U20599 (N_20599,N_18662,N_19912);
nand U20600 (N_20600,N_18457,N_19653);
nand U20601 (N_20601,N_18667,N_18124);
nor U20602 (N_20602,N_19569,N_18993);
xor U20603 (N_20603,N_19918,N_18451);
and U20604 (N_20604,N_18687,N_19088);
or U20605 (N_20605,N_19159,N_19744);
nand U20606 (N_20606,N_18782,N_19802);
or U20607 (N_20607,N_18633,N_19840);
nor U20608 (N_20608,N_19807,N_18032);
nor U20609 (N_20609,N_19804,N_18672);
nand U20610 (N_20610,N_19788,N_18242);
and U20611 (N_20611,N_19650,N_18368);
xor U20612 (N_20612,N_18799,N_18297);
nand U20613 (N_20613,N_18509,N_19017);
or U20614 (N_20614,N_18421,N_19933);
and U20615 (N_20615,N_18928,N_19929);
or U20616 (N_20616,N_18427,N_18060);
xnor U20617 (N_20617,N_19981,N_19765);
and U20618 (N_20618,N_19417,N_18872);
or U20619 (N_20619,N_19423,N_19258);
and U20620 (N_20620,N_19354,N_19097);
xnor U20621 (N_20621,N_19070,N_19725);
and U20622 (N_20622,N_19140,N_18903);
or U20623 (N_20623,N_19106,N_18265);
xnor U20624 (N_20624,N_19326,N_19945);
nand U20625 (N_20625,N_19920,N_19866);
nor U20626 (N_20626,N_18506,N_19047);
nor U20627 (N_20627,N_19971,N_18495);
and U20628 (N_20628,N_18871,N_18412);
or U20629 (N_20629,N_18338,N_18604);
nand U20630 (N_20630,N_18498,N_19275);
nor U20631 (N_20631,N_18612,N_18980);
xnor U20632 (N_20632,N_19842,N_19610);
or U20633 (N_20633,N_18008,N_18452);
or U20634 (N_20634,N_19815,N_19280);
or U20635 (N_20635,N_19661,N_19059);
or U20636 (N_20636,N_18868,N_19045);
xnor U20637 (N_20637,N_19491,N_19976);
nor U20638 (N_20638,N_18306,N_19961);
nor U20639 (N_20639,N_19726,N_18538);
or U20640 (N_20640,N_18829,N_19108);
xnor U20641 (N_20641,N_18791,N_18158);
and U20642 (N_20642,N_18346,N_18247);
or U20643 (N_20643,N_18743,N_19683);
or U20644 (N_20644,N_19479,N_19243);
and U20645 (N_20645,N_19299,N_18321);
xor U20646 (N_20646,N_19664,N_18512);
nand U20647 (N_20647,N_19995,N_19926);
nand U20648 (N_20648,N_19937,N_18707);
or U20649 (N_20649,N_18496,N_18240);
nand U20650 (N_20650,N_19179,N_18740);
nor U20651 (N_20651,N_18418,N_18442);
nand U20652 (N_20652,N_18382,N_18899);
and U20653 (N_20653,N_19628,N_19659);
nand U20654 (N_20654,N_19026,N_19868);
xnor U20655 (N_20655,N_19102,N_19294);
xnor U20656 (N_20656,N_19074,N_19697);
nand U20657 (N_20657,N_18628,N_18260);
and U20658 (N_20658,N_18215,N_19421);
nor U20659 (N_20659,N_18668,N_19410);
or U20660 (N_20660,N_18685,N_18514);
nand U20661 (N_20661,N_18278,N_19109);
xor U20662 (N_20662,N_18151,N_18753);
nor U20663 (N_20663,N_18842,N_18331);
nor U20664 (N_20664,N_19083,N_19619);
and U20665 (N_20665,N_18850,N_18796);
nor U20666 (N_20666,N_19204,N_19774);
nand U20667 (N_20667,N_19125,N_18550);
nand U20668 (N_20668,N_18566,N_18835);
nor U20669 (N_20669,N_18626,N_18925);
nor U20670 (N_20670,N_18801,N_18827);
nor U20671 (N_20671,N_18104,N_18811);
or U20672 (N_20672,N_18569,N_19144);
nand U20673 (N_20673,N_19853,N_18018);
xnor U20674 (N_20674,N_18556,N_18259);
and U20675 (N_20675,N_19808,N_18680);
and U20676 (N_20676,N_18304,N_19593);
and U20677 (N_20677,N_19173,N_18345);
or U20678 (N_20678,N_19358,N_19845);
nand U20679 (N_20679,N_19203,N_19547);
xnor U20680 (N_20680,N_18035,N_19439);
and U20681 (N_20681,N_18520,N_19430);
or U20682 (N_20682,N_18648,N_19282);
or U20683 (N_20683,N_19127,N_19321);
and U20684 (N_20684,N_19872,N_19655);
nor U20685 (N_20685,N_19445,N_19987);
or U20686 (N_20686,N_18894,N_19944);
and U20687 (N_20687,N_18169,N_19226);
nand U20688 (N_20688,N_19404,N_18714);
xor U20689 (N_20689,N_19303,N_18824);
and U20690 (N_20690,N_19690,N_19063);
and U20691 (N_20691,N_18638,N_18805);
nor U20692 (N_20692,N_18111,N_18730);
or U20693 (N_20693,N_18435,N_19975);
nand U20694 (N_20694,N_18236,N_19860);
nand U20695 (N_20695,N_19175,N_18720);
or U20696 (N_20696,N_19457,N_19990);
nor U20697 (N_20697,N_18414,N_18377);
nor U20698 (N_20698,N_18632,N_18146);
xnor U20699 (N_20699,N_18058,N_19518);
or U20700 (N_20700,N_19398,N_18726);
and U20701 (N_20701,N_19360,N_19742);
nor U20702 (N_20702,N_18313,N_19767);
xnor U20703 (N_20703,N_18314,N_19701);
nor U20704 (N_20704,N_19714,N_19538);
and U20705 (N_20705,N_19565,N_18934);
nand U20706 (N_20706,N_18831,N_19715);
or U20707 (N_20707,N_18374,N_18241);
or U20708 (N_20708,N_19437,N_19573);
nand U20709 (N_20709,N_19584,N_18907);
nor U20710 (N_20710,N_18898,N_19283);
or U20711 (N_20711,N_18589,N_19543);
nand U20712 (N_20712,N_18513,N_18228);
xnor U20713 (N_20713,N_19039,N_19211);
nand U20714 (N_20714,N_19947,N_18409);
nand U20715 (N_20715,N_18056,N_18606);
nand U20716 (N_20716,N_19722,N_18343);
and U20717 (N_20717,N_18140,N_19516);
xnor U20718 (N_20718,N_19403,N_18978);
and U20719 (N_20719,N_18854,N_18216);
nor U20720 (N_20720,N_18120,N_19522);
or U20721 (N_20721,N_18028,N_19621);
nand U20722 (N_20722,N_18530,N_19743);
and U20723 (N_20723,N_19183,N_18642);
and U20724 (N_20724,N_19052,N_19905);
nor U20725 (N_20725,N_18388,N_19265);
or U20726 (N_20726,N_18603,N_18317);
xnor U20727 (N_20727,N_18275,N_19559);
nor U20728 (N_20728,N_19564,N_19095);
and U20729 (N_20729,N_19756,N_19396);
xor U20730 (N_20730,N_19152,N_19069);
nand U20731 (N_20731,N_19533,N_19727);
nand U20732 (N_20732,N_19992,N_18643);
xor U20733 (N_20733,N_19546,N_19233);
or U20734 (N_20734,N_19915,N_19503);
nor U20735 (N_20735,N_19934,N_18263);
nand U20736 (N_20736,N_19426,N_19318);
xor U20737 (N_20737,N_19982,N_19236);
nand U20738 (N_20738,N_18300,N_18554);
and U20739 (N_20739,N_18501,N_18785);
nor U20740 (N_20740,N_19834,N_18750);
or U20741 (N_20741,N_18192,N_19838);
nor U20742 (N_20742,N_18952,N_18543);
xor U20743 (N_20743,N_19484,N_19129);
nor U20744 (N_20744,N_19356,N_19951);
or U20745 (N_20745,N_18650,N_19825);
xor U20746 (N_20746,N_19472,N_19234);
or U20747 (N_20747,N_18376,N_18972);
xor U20748 (N_20748,N_18988,N_18305);
and U20749 (N_20749,N_19441,N_19241);
or U20750 (N_20750,N_19316,N_19286);
or U20751 (N_20751,N_19958,N_19277);
and U20752 (N_20752,N_19967,N_19009);
nand U20753 (N_20753,N_18402,N_18408);
or U20754 (N_20754,N_18478,N_18669);
or U20755 (N_20755,N_19599,N_19887);
or U20756 (N_20756,N_18954,N_18283);
nor U20757 (N_20757,N_19575,N_18588);
nand U20758 (N_20758,N_18089,N_19389);
nor U20759 (N_20759,N_18366,N_18968);
nor U20760 (N_20760,N_18768,N_19974);
nand U20761 (N_20761,N_19856,N_18717);
nor U20762 (N_20762,N_18174,N_18096);
nand U20763 (N_20763,N_18789,N_19773);
nor U20764 (N_20764,N_18646,N_18491);
xor U20765 (N_20765,N_18849,N_18967);
and U20766 (N_20766,N_18581,N_18038);
nor U20767 (N_20767,N_18302,N_19864);
nand U20768 (N_20768,N_18469,N_18977);
and U20769 (N_20769,N_18875,N_19685);
and U20770 (N_20770,N_19139,N_19587);
and U20771 (N_20771,N_19511,N_18203);
nand U20772 (N_20772,N_19501,N_19909);
nand U20773 (N_20773,N_18778,N_18927);
and U20774 (N_20774,N_18462,N_19705);
nand U20775 (N_20775,N_18702,N_18873);
xnor U20776 (N_20776,N_18497,N_18312);
xor U20777 (N_20777,N_18271,N_19254);
and U20778 (N_20778,N_19092,N_18088);
and U20779 (N_20779,N_19223,N_18003);
and U20780 (N_20780,N_18930,N_18170);
and U20781 (N_20781,N_19309,N_18584);
xor U20782 (N_20782,N_18071,N_19386);
or U20783 (N_20783,N_18797,N_18926);
or U20784 (N_20784,N_19654,N_18734);
and U20785 (N_20785,N_18001,N_19215);
nand U20786 (N_20786,N_19609,N_18809);
nand U20787 (N_20787,N_19686,N_19031);
nor U20788 (N_20788,N_19730,N_19028);
xnor U20789 (N_20789,N_19331,N_19789);
nand U20790 (N_20790,N_18749,N_19058);
nor U20791 (N_20791,N_19079,N_19768);
and U20792 (N_20792,N_19065,N_19098);
nand U20793 (N_20793,N_18615,N_19826);
or U20794 (N_20794,N_18336,N_18375);
nand U20795 (N_20795,N_19763,N_19809);
nand U20796 (N_20796,N_18995,N_18600);
nand U20797 (N_20797,N_18087,N_19615);
nor U20798 (N_20798,N_18277,N_18416);
or U20799 (N_20799,N_19777,N_18505);
and U20800 (N_20800,N_18997,N_19814);
nor U20801 (N_20801,N_19635,N_18441);
nor U20802 (N_20802,N_18679,N_18649);
nand U20803 (N_20803,N_18613,N_19471);
nand U20804 (N_20804,N_18517,N_18819);
and U20805 (N_20805,N_18548,N_18227);
nand U20806 (N_20806,N_18045,N_18956);
or U20807 (N_20807,N_19136,N_19189);
xor U20808 (N_20808,N_19545,N_19530);
nor U20809 (N_20809,N_19899,N_19707);
nor U20810 (N_20810,N_18706,N_19679);
nand U20811 (N_20811,N_18004,N_18542);
xor U20812 (N_20812,N_18869,N_18771);
nand U20813 (N_20813,N_18167,N_19665);
xor U20814 (N_20814,N_19504,N_18736);
and U20815 (N_20815,N_19015,N_19094);
nor U20816 (N_20816,N_19438,N_19813);
nor U20817 (N_20817,N_18639,N_19984);
and U20818 (N_20818,N_19557,N_18885);
nor U20819 (N_20819,N_18234,N_19869);
nand U20820 (N_20820,N_19652,N_18889);
xor U20821 (N_20821,N_18276,N_19008);
nor U20822 (N_20822,N_18068,N_19775);
and U20823 (N_20823,N_18257,N_19235);
and U20824 (N_20824,N_19180,N_19821);
nor U20825 (N_20825,N_19344,N_19649);
nor U20826 (N_20826,N_19506,N_18573);
and U20827 (N_20827,N_19642,N_19579);
nor U20828 (N_20828,N_19537,N_18468);
and U20829 (N_20829,N_19350,N_19470);
nor U20830 (N_20830,N_19948,N_19824);
nand U20831 (N_20831,N_19588,N_19563);
or U20832 (N_20832,N_19227,N_19598);
xor U20833 (N_20833,N_18742,N_18099);
nor U20834 (N_20834,N_18114,N_19117);
and U20835 (N_20835,N_18440,N_19011);
or U20836 (N_20836,N_18693,N_18951);
nand U20837 (N_20837,N_18932,N_19717);
and U20838 (N_20838,N_19745,N_19348);
nor U20839 (N_20839,N_18728,N_18367);
nor U20840 (N_20840,N_19510,N_19060);
and U20841 (N_20841,N_19377,N_19757);
nand U20842 (N_20842,N_19264,N_18447);
xor U20843 (N_20843,N_18611,N_19818);
nor U20844 (N_20844,N_19986,N_18515);
nor U20845 (N_20845,N_19721,N_19734);
or U20846 (N_20846,N_18634,N_18341);
and U20847 (N_20847,N_19759,N_19468);
or U20848 (N_20848,N_18222,N_18938);
nand U20849 (N_20849,N_18389,N_19671);
and U20850 (N_20850,N_18519,N_18083);
and U20851 (N_20851,N_19698,N_18432);
xor U20852 (N_20852,N_18171,N_18540);
or U20853 (N_20853,N_19218,N_19600);
nor U20854 (N_20854,N_19875,N_18094);
nand U20855 (N_20855,N_18808,N_19147);
and U20856 (N_20856,N_18713,N_18479);
xnor U20857 (N_20857,N_19395,N_18655);
and U20858 (N_20858,N_19731,N_19916);
or U20859 (N_20859,N_19040,N_18384);
and U20860 (N_20860,N_19886,N_19969);
nor U20861 (N_20861,N_18209,N_18391);
nor U20862 (N_20862,N_19606,N_19024);
nor U20863 (N_20863,N_18949,N_19195);
nor U20864 (N_20864,N_19005,N_18839);
nor U20865 (N_20865,N_18326,N_18142);
or U20866 (N_20866,N_19572,N_18691);
nand U20867 (N_20867,N_19497,N_18024);
nand U20868 (N_20868,N_18095,N_18420);
or U20869 (N_20869,N_19919,N_19245);
and U20870 (N_20870,N_19667,N_18666);
nor U20871 (N_20871,N_18947,N_18565);
nor U20872 (N_20872,N_19891,N_18065);
and U20873 (N_20873,N_19312,N_18826);
xnor U20874 (N_20874,N_18002,N_18455);
or U20875 (N_20875,N_18610,N_19213);
or U20876 (N_20876,N_18790,N_18129);
and U20877 (N_20877,N_19451,N_19440);
nor U20878 (N_20878,N_19084,N_19352);
nor U20879 (N_20879,N_19343,N_19034);
nand U20880 (N_20880,N_19618,N_19567);
nor U20881 (N_20881,N_19738,N_19594);
nand U20882 (N_20882,N_19146,N_19436);
xnor U20883 (N_20883,N_19414,N_19644);
xnor U20884 (N_20884,N_18518,N_19668);
xnor U20885 (N_20885,N_18379,N_19897);
nand U20886 (N_20886,N_18541,N_19366);
nand U20887 (N_20887,N_18891,N_19422);
and U20888 (N_20888,N_18394,N_18154);
and U20889 (N_20889,N_19596,N_19889);
nor U20890 (N_20890,N_19418,N_18631);
nand U20891 (N_20891,N_18425,N_18401);
xor U20892 (N_20892,N_18380,N_18532);
nand U20893 (N_20893,N_18208,N_18981);
and U20894 (N_20894,N_18219,N_19616);
or U20895 (N_20895,N_18250,N_19021);
nor U20896 (N_20896,N_18537,N_19345);
nand U20897 (N_20897,N_18077,N_19128);
nor U20898 (N_20898,N_18101,N_19274);
xor U20899 (N_20899,N_18410,N_18948);
nand U20900 (N_20900,N_18944,N_18473);
nor U20901 (N_20901,N_18716,N_18933);
xor U20902 (N_20902,N_18126,N_19712);
nand U20903 (N_20903,N_19997,N_18751);
nand U20904 (N_20904,N_19371,N_18128);
nand U20905 (N_20905,N_19544,N_19467);
xor U20906 (N_20906,N_18296,N_19847);
nand U20907 (N_20907,N_18931,N_18052);
or U20908 (N_20908,N_19943,N_19252);
and U20909 (N_20909,N_19338,N_18864);
nand U20910 (N_20910,N_18034,N_19998);
and U20911 (N_20911,N_18246,N_18802);
nand U20912 (N_20912,N_19988,N_19633);
nand U20913 (N_20913,N_18747,N_18354);
xnor U20914 (N_20914,N_19302,N_18323);
nor U20915 (N_20915,N_19728,N_19051);
xor U20916 (N_20916,N_19991,N_18036);
and U20917 (N_20917,N_18961,N_19591);
nand U20918 (N_20918,N_19799,N_19170);
and U20919 (N_20919,N_18261,N_19867);
or U20920 (N_20920,N_18636,N_19539);
xnor U20921 (N_20921,N_19612,N_19347);
nand U20922 (N_20922,N_19131,N_18787);
nor U20923 (N_20923,N_19393,N_18061);
or U20924 (N_20924,N_18924,N_19797);
or U20925 (N_20925,N_18218,N_19210);
nor U20926 (N_20926,N_19207,N_18670);
or U20927 (N_20927,N_18181,N_18711);
nor U20928 (N_20928,N_19132,N_19946);
and U20929 (N_20929,N_18020,N_19214);
xnor U20930 (N_20930,N_19076,N_19793);
nand U20931 (N_20931,N_18009,N_18507);
nor U20932 (N_20932,N_18472,N_19903);
nor U20933 (N_20933,N_18159,N_18221);
or U20934 (N_20934,N_19989,N_18318);
nor U20935 (N_20935,N_18682,N_18064);
xnor U20936 (N_20936,N_18963,N_18756);
xnor U20937 (N_20937,N_19194,N_19684);
nor U20938 (N_20938,N_19016,N_19145);
or U20939 (N_20939,N_19172,N_18205);
and U20940 (N_20940,N_19729,N_18601);
nand U20941 (N_20941,N_19433,N_19561);
and U20942 (N_20942,N_19535,N_19156);
and U20943 (N_20943,N_18865,N_18075);
or U20944 (N_20944,N_18914,N_18663);
or U20945 (N_20945,N_18224,N_18609);
nand U20946 (N_20946,N_18644,N_19013);
or U20947 (N_20947,N_18021,N_18175);
or U20948 (N_20948,N_18637,N_18454);
nor U20949 (N_20949,N_18324,N_18762);
and U20950 (N_20950,N_19892,N_18833);
nand U20951 (N_20951,N_19167,N_19250);
nor U20952 (N_20952,N_19415,N_19917);
and U20953 (N_20953,N_18880,N_19384);
or U20954 (N_20954,N_19636,N_19980);
and U20955 (N_20955,N_18269,N_18348);
xor U20956 (N_20956,N_19688,N_18546);
and U20957 (N_20957,N_19955,N_18210);
xor U20958 (N_20958,N_19054,N_19220);
or U20959 (N_20959,N_19924,N_19862);
nor U20960 (N_20960,N_18160,N_18459);
xnor U20961 (N_20961,N_18335,N_18481);
nand U20962 (N_20962,N_18623,N_18464);
nand U20963 (N_20963,N_18500,N_19308);
nor U20964 (N_20964,N_19077,N_19735);
or U20965 (N_20965,N_18310,N_19851);
nand U20966 (N_20966,N_19928,N_18661);
xnor U20967 (N_20967,N_19378,N_18282);
or U20968 (N_20968,N_18162,N_19458);
or U20969 (N_20969,N_18423,N_19801);
xnor U20970 (N_20970,N_19161,N_18485);
xor U20971 (N_20971,N_19317,N_19952);
nand U20972 (N_20972,N_19558,N_19121);
nand U20973 (N_20973,N_19091,N_18225);
nand U20974 (N_20974,N_19408,N_19041);
xor U20975 (N_20975,N_18419,N_19281);
xnor U20976 (N_20976,N_18054,N_19297);
xnor U20977 (N_20977,N_19870,N_18908);
nor U20978 (N_20978,N_19786,N_18830);
xnor U20979 (N_20979,N_18363,N_18006);
and U20980 (N_20980,N_19391,N_19397);
xnor U20981 (N_20981,N_18157,N_18232);
nor U20982 (N_20982,N_19716,N_19820);
nor U20983 (N_20983,N_19103,N_19519);
nand U20984 (N_20984,N_18139,N_19394);
or U20985 (N_20985,N_18592,N_19256);
nand U20986 (N_20986,N_18555,N_19278);
nand U20987 (N_20987,N_18287,N_19883);
xor U20988 (N_20988,N_18486,N_18994);
nor U20989 (N_20989,N_18950,N_19119);
nand U20990 (N_20990,N_18381,N_18917);
nor U20991 (N_20991,N_18005,N_19368);
or U20992 (N_20992,N_18212,N_18119);
xor U20993 (N_20993,N_19165,N_18562);
or U20994 (N_20994,N_19940,N_18118);
xnor U20995 (N_20995,N_18744,N_19625);
nor U20996 (N_20996,N_19508,N_18371);
and U20997 (N_20997,N_18527,N_18578);
or U20998 (N_20998,N_18387,N_18709);
nand U20999 (N_20999,N_18362,N_18531);
or U21000 (N_21000,N_19996,N_19775);
xor U21001 (N_21001,N_18139,N_19338);
nor U21002 (N_21002,N_18936,N_19545);
or U21003 (N_21003,N_19158,N_18664);
and U21004 (N_21004,N_19476,N_18414);
nand U21005 (N_21005,N_18512,N_19402);
nand U21006 (N_21006,N_18573,N_18556);
nor U21007 (N_21007,N_19810,N_18540);
nor U21008 (N_21008,N_18960,N_18696);
and U21009 (N_21009,N_19242,N_18672);
nor U21010 (N_21010,N_18572,N_18299);
nor U21011 (N_21011,N_18487,N_18322);
nor U21012 (N_21012,N_18495,N_18191);
or U21013 (N_21013,N_19914,N_19095);
nand U21014 (N_21014,N_19254,N_19537);
xnor U21015 (N_21015,N_18890,N_19306);
nor U21016 (N_21016,N_18593,N_19424);
and U21017 (N_21017,N_18961,N_18528);
or U21018 (N_21018,N_18567,N_19287);
nand U21019 (N_21019,N_19047,N_18900);
or U21020 (N_21020,N_19486,N_19293);
and U21021 (N_21021,N_19066,N_19920);
and U21022 (N_21022,N_19430,N_19335);
xor U21023 (N_21023,N_19787,N_19572);
xor U21024 (N_21024,N_18784,N_18606);
and U21025 (N_21025,N_18705,N_19178);
or U21026 (N_21026,N_19964,N_18173);
nand U21027 (N_21027,N_19670,N_18171);
xnor U21028 (N_21028,N_19128,N_19815);
xnor U21029 (N_21029,N_19901,N_19182);
nor U21030 (N_21030,N_19754,N_19865);
xnor U21031 (N_21031,N_18561,N_18396);
or U21032 (N_21032,N_18700,N_19785);
xor U21033 (N_21033,N_19335,N_19096);
nor U21034 (N_21034,N_18362,N_18904);
and U21035 (N_21035,N_18191,N_18133);
nor U21036 (N_21036,N_19892,N_18080);
nand U21037 (N_21037,N_19137,N_19985);
and U21038 (N_21038,N_18917,N_19619);
xnor U21039 (N_21039,N_19030,N_19088);
or U21040 (N_21040,N_19155,N_18544);
or U21041 (N_21041,N_19104,N_18417);
nand U21042 (N_21042,N_18709,N_19736);
nor U21043 (N_21043,N_18435,N_19847);
and U21044 (N_21044,N_19840,N_18649);
and U21045 (N_21045,N_19982,N_18267);
xor U21046 (N_21046,N_18842,N_18235);
nand U21047 (N_21047,N_19182,N_18017);
or U21048 (N_21048,N_19725,N_18443);
xnor U21049 (N_21049,N_18635,N_18636);
or U21050 (N_21050,N_18309,N_19855);
xor U21051 (N_21051,N_18455,N_19282);
nand U21052 (N_21052,N_18203,N_19037);
or U21053 (N_21053,N_19294,N_19236);
xor U21054 (N_21054,N_19300,N_19295);
nor U21055 (N_21055,N_19029,N_19470);
nand U21056 (N_21056,N_19541,N_18830);
and U21057 (N_21057,N_19855,N_18889);
or U21058 (N_21058,N_19148,N_18517);
and U21059 (N_21059,N_18990,N_19594);
or U21060 (N_21060,N_19790,N_19307);
or U21061 (N_21061,N_18988,N_18019);
or U21062 (N_21062,N_19227,N_18358);
and U21063 (N_21063,N_19378,N_19085);
and U21064 (N_21064,N_18895,N_18334);
or U21065 (N_21065,N_18273,N_19321);
nand U21066 (N_21066,N_18163,N_18434);
nor U21067 (N_21067,N_19189,N_19106);
nor U21068 (N_21068,N_18060,N_19552);
nor U21069 (N_21069,N_19152,N_18528);
and U21070 (N_21070,N_19421,N_19711);
and U21071 (N_21071,N_18594,N_18877);
or U21072 (N_21072,N_19052,N_18560);
or U21073 (N_21073,N_19277,N_19144);
xor U21074 (N_21074,N_18715,N_18724);
nand U21075 (N_21075,N_18766,N_19836);
nor U21076 (N_21076,N_18625,N_19166);
xor U21077 (N_21077,N_19617,N_19839);
nor U21078 (N_21078,N_19873,N_19828);
xnor U21079 (N_21079,N_19198,N_18574);
nand U21080 (N_21080,N_19355,N_18030);
or U21081 (N_21081,N_19161,N_19255);
xnor U21082 (N_21082,N_19669,N_19154);
nand U21083 (N_21083,N_19036,N_19481);
nor U21084 (N_21084,N_18785,N_18760);
xnor U21085 (N_21085,N_19730,N_19009);
or U21086 (N_21086,N_19564,N_19635);
and U21087 (N_21087,N_18228,N_19509);
xnor U21088 (N_21088,N_19192,N_19775);
or U21089 (N_21089,N_19170,N_19440);
nor U21090 (N_21090,N_19196,N_18609);
nor U21091 (N_21091,N_19514,N_18296);
or U21092 (N_21092,N_19909,N_18851);
xor U21093 (N_21093,N_18808,N_19969);
nand U21094 (N_21094,N_18661,N_19956);
xnor U21095 (N_21095,N_19836,N_18844);
nand U21096 (N_21096,N_19974,N_19773);
or U21097 (N_21097,N_19274,N_19961);
nor U21098 (N_21098,N_18803,N_19359);
nor U21099 (N_21099,N_18406,N_19356);
or U21100 (N_21100,N_19057,N_19310);
and U21101 (N_21101,N_18580,N_19808);
and U21102 (N_21102,N_19870,N_19236);
or U21103 (N_21103,N_19050,N_18455);
xnor U21104 (N_21104,N_19899,N_18844);
xor U21105 (N_21105,N_18444,N_18021);
nor U21106 (N_21106,N_19356,N_18653);
nor U21107 (N_21107,N_19273,N_18408);
xnor U21108 (N_21108,N_19393,N_19930);
xor U21109 (N_21109,N_18683,N_18276);
nand U21110 (N_21110,N_18960,N_18569);
and U21111 (N_21111,N_18250,N_18370);
xnor U21112 (N_21112,N_18579,N_19103);
and U21113 (N_21113,N_18284,N_18271);
and U21114 (N_21114,N_19343,N_19844);
xor U21115 (N_21115,N_18696,N_19902);
and U21116 (N_21116,N_19417,N_18371);
xnor U21117 (N_21117,N_19453,N_18510);
xor U21118 (N_21118,N_19889,N_19252);
nand U21119 (N_21119,N_18881,N_18213);
xnor U21120 (N_21120,N_19192,N_18645);
nor U21121 (N_21121,N_18996,N_18249);
or U21122 (N_21122,N_18314,N_18578);
and U21123 (N_21123,N_19766,N_19210);
xor U21124 (N_21124,N_19666,N_18089);
or U21125 (N_21125,N_18861,N_19910);
nand U21126 (N_21126,N_18487,N_18256);
nor U21127 (N_21127,N_19424,N_18854);
xnor U21128 (N_21128,N_19543,N_19134);
nand U21129 (N_21129,N_18345,N_18446);
nor U21130 (N_21130,N_18944,N_18765);
xnor U21131 (N_21131,N_19314,N_18558);
nand U21132 (N_21132,N_19377,N_18483);
nor U21133 (N_21133,N_18373,N_18499);
nand U21134 (N_21134,N_19077,N_18804);
xnor U21135 (N_21135,N_18516,N_19154);
or U21136 (N_21136,N_19810,N_19291);
xor U21137 (N_21137,N_19759,N_18936);
and U21138 (N_21138,N_19204,N_19980);
and U21139 (N_21139,N_18758,N_18012);
xnor U21140 (N_21140,N_19481,N_19534);
xnor U21141 (N_21141,N_19394,N_19119);
or U21142 (N_21142,N_18744,N_19323);
and U21143 (N_21143,N_18126,N_19694);
or U21144 (N_21144,N_18338,N_19160);
xnor U21145 (N_21145,N_18999,N_19399);
and U21146 (N_21146,N_19776,N_19597);
xnor U21147 (N_21147,N_18486,N_19988);
nor U21148 (N_21148,N_19480,N_19359);
nand U21149 (N_21149,N_18659,N_18027);
nor U21150 (N_21150,N_18783,N_19137);
and U21151 (N_21151,N_19014,N_19574);
nand U21152 (N_21152,N_18581,N_18998);
and U21153 (N_21153,N_18845,N_18822);
nor U21154 (N_21154,N_19098,N_18303);
nand U21155 (N_21155,N_18379,N_19802);
or U21156 (N_21156,N_18247,N_19921);
nor U21157 (N_21157,N_19825,N_19493);
xnor U21158 (N_21158,N_18466,N_19873);
nor U21159 (N_21159,N_19248,N_18381);
or U21160 (N_21160,N_19028,N_19300);
and U21161 (N_21161,N_19510,N_18568);
or U21162 (N_21162,N_18601,N_18108);
and U21163 (N_21163,N_19159,N_18957);
xor U21164 (N_21164,N_19640,N_18356);
nand U21165 (N_21165,N_19883,N_18327);
and U21166 (N_21166,N_19342,N_19936);
and U21167 (N_21167,N_19718,N_19673);
nand U21168 (N_21168,N_18179,N_18076);
xnor U21169 (N_21169,N_19625,N_19974);
nand U21170 (N_21170,N_19889,N_18408);
and U21171 (N_21171,N_19818,N_19276);
nor U21172 (N_21172,N_19908,N_18700);
nor U21173 (N_21173,N_19618,N_18924);
or U21174 (N_21174,N_18637,N_18963);
or U21175 (N_21175,N_18967,N_18976);
xor U21176 (N_21176,N_18341,N_19836);
or U21177 (N_21177,N_18875,N_18017);
and U21178 (N_21178,N_18900,N_19293);
nand U21179 (N_21179,N_19356,N_18257);
and U21180 (N_21180,N_19351,N_19137);
nor U21181 (N_21181,N_19826,N_19591);
nand U21182 (N_21182,N_19753,N_19446);
nand U21183 (N_21183,N_18023,N_18796);
and U21184 (N_21184,N_18738,N_18612);
nor U21185 (N_21185,N_18610,N_18439);
nand U21186 (N_21186,N_19134,N_18798);
xnor U21187 (N_21187,N_18570,N_19249);
xor U21188 (N_21188,N_19456,N_19252);
or U21189 (N_21189,N_19960,N_19373);
xor U21190 (N_21190,N_19977,N_18570);
nand U21191 (N_21191,N_19977,N_18325);
or U21192 (N_21192,N_19405,N_19153);
xnor U21193 (N_21193,N_18229,N_19849);
nand U21194 (N_21194,N_18181,N_19031);
xor U21195 (N_21195,N_19087,N_19368);
xor U21196 (N_21196,N_18830,N_19878);
nor U21197 (N_21197,N_18152,N_18979);
xnor U21198 (N_21198,N_19652,N_18340);
and U21199 (N_21199,N_19462,N_18157);
nor U21200 (N_21200,N_19700,N_19428);
or U21201 (N_21201,N_18408,N_18621);
or U21202 (N_21202,N_19078,N_19822);
or U21203 (N_21203,N_18772,N_19182);
nand U21204 (N_21204,N_18572,N_19809);
nor U21205 (N_21205,N_18664,N_19186);
and U21206 (N_21206,N_19984,N_19633);
nor U21207 (N_21207,N_19295,N_19459);
and U21208 (N_21208,N_18305,N_19773);
and U21209 (N_21209,N_19972,N_18884);
nand U21210 (N_21210,N_18941,N_18792);
and U21211 (N_21211,N_18316,N_19263);
or U21212 (N_21212,N_18586,N_18968);
or U21213 (N_21213,N_19248,N_18387);
and U21214 (N_21214,N_18746,N_19672);
nor U21215 (N_21215,N_18599,N_19451);
nand U21216 (N_21216,N_18615,N_19772);
or U21217 (N_21217,N_19811,N_19681);
nand U21218 (N_21218,N_18485,N_19508);
nand U21219 (N_21219,N_18421,N_19371);
nand U21220 (N_21220,N_19277,N_19316);
xnor U21221 (N_21221,N_19927,N_19518);
nand U21222 (N_21222,N_18362,N_19178);
nor U21223 (N_21223,N_19432,N_19925);
and U21224 (N_21224,N_19649,N_19758);
and U21225 (N_21225,N_18023,N_18240);
nand U21226 (N_21226,N_18279,N_18035);
or U21227 (N_21227,N_19864,N_19148);
or U21228 (N_21228,N_18328,N_18945);
xnor U21229 (N_21229,N_18644,N_18992);
or U21230 (N_21230,N_19377,N_19937);
nand U21231 (N_21231,N_18364,N_19408);
and U21232 (N_21232,N_19919,N_19758);
nand U21233 (N_21233,N_19860,N_19708);
nor U21234 (N_21234,N_18146,N_18848);
and U21235 (N_21235,N_18112,N_19381);
and U21236 (N_21236,N_19708,N_19218);
nand U21237 (N_21237,N_19865,N_19070);
xor U21238 (N_21238,N_19534,N_19758);
xnor U21239 (N_21239,N_19566,N_18313);
and U21240 (N_21240,N_19961,N_19645);
or U21241 (N_21241,N_19843,N_19303);
nand U21242 (N_21242,N_19545,N_19397);
xnor U21243 (N_21243,N_18692,N_18372);
nor U21244 (N_21244,N_18959,N_19619);
xor U21245 (N_21245,N_19033,N_19250);
xnor U21246 (N_21246,N_19888,N_18314);
xnor U21247 (N_21247,N_18868,N_19081);
xnor U21248 (N_21248,N_18590,N_19234);
or U21249 (N_21249,N_19008,N_19325);
or U21250 (N_21250,N_18297,N_18052);
nor U21251 (N_21251,N_18536,N_19402);
nand U21252 (N_21252,N_18970,N_19924);
and U21253 (N_21253,N_19857,N_18899);
or U21254 (N_21254,N_19474,N_18106);
nand U21255 (N_21255,N_18567,N_18294);
nand U21256 (N_21256,N_18807,N_18806);
nand U21257 (N_21257,N_19971,N_19070);
xor U21258 (N_21258,N_19179,N_19904);
nand U21259 (N_21259,N_19982,N_18202);
xnor U21260 (N_21260,N_18832,N_19013);
and U21261 (N_21261,N_19057,N_19437);
nor U21262 (N_21262,N_18757,N_19432);
and U21263 (N_21263,N_19514,N_19575);
nand U21264 (N_21264,N_19926,N_18748);
nand U21265 (N_21265,N_18306,N_19194);
and U21266 (N_21266,N_19899,N_19936);
nor U21267 (N_21267,N_18143,N_18141);
nand U21268 (N_21268,N_19771,N_18357);
and U21269 (N_21269,N_18460,N_19119);
or U21270 (N_21270,N_19966,N_18635);
xor U21271 (N_21271,N_19941,N_19504);
nand U21272 (N_21272,N_19102,N_18564);
nor U21273 (N_21273,N_18767,N_18098);
nor U21274 (N_21274,N_19882,N_18210);
nand U21275 (N_21275,N_18728,N_19128);
nand U21276 (N_21276,N_19664,N_18454);
nand U21277 (N_21277,N_18364,N_19352);
xnor U21278 (N_21278,N_18971,N_19386);
nand U21279 (N_21279,N_18645,N_19100);
nand U21280 (N_21280,N_19448,N_18628);
nand U21281 (N_21281,N_18208,N_18910);
and U21282 (N_21282,N_18609,N_18517);
xnor U21283 (N_21283,N_19281,N_19929);
nor U21284 (N_21284,N_19526,N_18057);
or U21285 (N_21285,N_19661,N_19738);
nand U21286 (N_21286,N_19887,N_19010);
nor U21287 (N_21287,N_19306,N_18077);
nor U21288 (N_21288,N_19903,N_19100);
nor U21289 (N_21289,N_19716,N_19354);
and U21290 (N_21290,N_19814,N_18809);
or U21291 (N_21291,N_19526,N_19223);
nand U21292 (N_21292,N_18490,N_18371);
and U21293 (N_21293,N_18355,N_18126);
xnor U21294 (N_21294,N_19756,N_19580);
or U21295 (N_21295,N_18571,N_19603);
and U21296 (N_21296,N_18482,N_18323);
xor U21297 (N_21297,N_18383,N_19166);
and U21298 (N_21298,N_18579,N_19035);
and U21299 (N_21299,N_19212,N_18799);
or U21300 (N_21300,N_18933,N_18400);
xor U21301 (N_21301,N_19293,N_19455);
or U21302 (N_21302,N_19428,N_18923);
nor U21303 (N_21303,N_18773,N_19210);
and U21304 (N_21304,N_18136,N_18323);
nor U21305 (N_21305,N_18863,N_19522);
xor U21306 (N_21306,N_18691,N_18440);
and U21307 (N_21307,N_18690,N_19711);
nand U21308 (N_21308,N_18310,N_18077);
nor U21309 (N_21309,N_18710,N_19064);
and U21310 (N_21310,N_19040,N_19696);
or U21311 (N_21311,N_19833,N_18381);
nor U21312 (N_21312,N_18630,N_19990);
or U21313 (N_21313,N_18729,N_19760);
nand U21314 (N_21314,N_18925,N_19790);
nor U21315 (N_21315,N_18033,N_18867);
nor U21316 (N_21316,N_18092,N_19557);
nor U21317 (N_21317,N_18024,N_18881);
nand U21318 (N_21318,N_19115,N_19267);
and U21319 (N_21319,N_19792,N_18783);
or U21320 (N_21320,N_18856,N_18035);
or U21321 (N_21321,N_18563,N_19323);
and U21322 (N_21322,N_19300,N_19630);
or U21323 (N_21323,N_18923,N_19577);
or U21324 (N_21324,N_18301,N_19480);
nand U21325 (N_21325,N_18914,N_18772);
and U21326 (N_21326,N_18790,N_18832);
nor U21327 (N_21327,N_18638,N_19583);
nand U21328 (N_21328,N_19181,N_19214);
nand U21329 (N_21329,N_19734,N_19780);
and U21330 (N_21330,N_19486,N_19085);
nand U21331 (N_21331,N_18599,N_19617);
or U21332 (N_21332,N_18237,N_19618);
xor U21333 (N_21333,N_19474,N_19505);
nor U21334 (N_21334,N_19821,N_18396);
and U21335 (N_21335,N_19543,N_18874);
xor U21336 (N_21336,N_18001,N_19022);
or U21337 (N_21337,N_18574,N_18553);
xor U21338 (N_21338,N_19570,N_18718);
nand U21339 (N_21339,N_18608,N_18698);
nor U21340 (N_21340,N_18058,N_19701);
xor U21341 (N_21341,N_19361,N_18397);
xnor U21342 (N_21342,N_18686,N_19817);
nand U21343 (N_21343,N_19246,N_19558);
xnor U21344 (N_21344,N_19709,N_18966);
nor U21345 (N_21345,N_19386,N_19128);
nor U21346 (N_21346,N_19577,N_18206);
nand U21347 (N_21347,N_19922,N_18247);
or U21348 (N_21348,N_18164,N_19084);
or U21349 (N_21349,N_18784,N_19220);
and U21350 (N_21350,N_18127,N_18714);
nor U21351 (N_21351,N_18335,N_18310);
nor U21352 (N_21352,N_18020,N_18118);
and U21353 (N_21353,N_19278,N_18409);
and U21354 (N_21354,N_19488,N_18056);
nand U21355 (N_21355,N_18702,N_19972);
and U21356 (N_21356,N_18798,N_18912);
xor U21357 (N_21357,N_19953,N_19060);
and U21358 (N_21358,N_18666,N_19148);
xor U21359 (N_21359,N_19211,N_18486);
or U21360 (N_21360,N_18866,N_19491);
and U21361 (N_21361,N_18127,N_19605);
nor U21362 (N_21362,N_19897,N_19314);
nand U21363 (N_21363,N_18486,N_18521);
xor U21364 (N_21364,N_19579,N_19332);
nor U21365 (N_21365,N_19829,N_19401);
or U21366 (N_21366,N_18870,N_18454);
or U21367 (N_21367,N_19363,N_18911);
and U21368 (N_21368,N_19301,N_18395);
or U21369 (N_21369,N_18906,N_18882);
nand U21370 (N_21370,N_18214,N_18110);
and U21371 (N_21371,N_19265,N_18005);
and U21372 (N_21372,N_19923,N_18962);
or U21373 (N_21373,N_18332,N_18381);
nand U21374 (N_21374,N_18208,N_18252);
nor U21375 (N_21375,N_19774,N_18473);
and U21376 (N_21376,N_19914,N_19840);
nor U21377 (N_21377,N_18443,N_18255);
xor U21378 (N_21378,N_19677,N_18994);
nor U21379 (N_21379,N_19750,N_19385);
nor U21380 (N_21380,N_19309,N_18324);
nor U21381 (N_21381,N_18989,N_18473);
nand U21382 (N_21382,N_18621,N_18017);
nand U21383 (N_21383,N_19442,N_19680);
and U21384 (N_21384,N_18994,N_18226);
xor U21385 (N_21385,N_18106,N_18786);
and U21386 (N_21386,N_18427,N_18815);
and U21387 (N_21387,N_18018,N_18868);
nor U21388 (N_21388,N_19471,N_19049);
nor U21389 (N_21389,N_19971,N_18137);
nand U21390 (N_21390,N_19555,N_19947);
and U21391 (N_21391,N_19773,N_19428);
xor U21392 (N_21392,N_18399,N_18879);
and U21393 (N_21393,N_19411,N_18949);
or U21394 (N_21394,N_19102,N_19953);
nand U21395 (N_21395,N_19717,N_18999);
xnor U21396 (N_21396,N_19982,N_18407);
or U21397 (N_21397,N_18384,N_18793);
nand U21398 (N_21398,N_18100,N_18950);
or U21399 (N_21399,N_19974,N_18021);
nand U21400 (N_21400,N_18707,N_18540);
nand U21401 (N_21401,N_18856,N_18026);
and U21402 (N_21402,N_19927,N_18335);
nor U21403 (N_21403,N_19407,N_19081);
or U21404 (N_21404,N_18412,N_19916);
nand U21405 (N_21405,N_19172,N_18076);
xor U21406 (N_21406,N_18767,N_18998);
and U21407 (N_21407,N_19254,N_19314);
and U21408 (N_21408,N_19955,N_18312);
xor U21409 (N_21409,N_19696,N_19535);
and U21410 (N_21410,N_18896,N_18810);
nor U21411 (N_21411,N_19213,N_18425);
and U21412 (N_21412,N_19462,N_19232);
nor U21413 (N_21413,N_18049,N_19106);
or U21414 (N_21414,N_19873,N_18436);
or U21415 (N_21415,N_18753,N_18371);
or U21416 (N_21416,N_19583,N_18005);
or U21417 (N_21417,N_18817,N_18126);
nand U21418 (N_21418,N_18022,N_19111);
and U21419 (N_21419,N_18184,N_18417);
nor U21420 (N_21420,N_19813,N_19968);
xor U21421 (N_21421,N_18424,N_19834);
or U21422 (N_21422,N_18217,N_18365);
nand U21423 (N_21423,N_18230,N_18310);
nand U21424 (N_21424,N_18904,N_18113);
or U21425 (N_21425,N_19883,N_18964);
xor U21426 (N_21426,N_18502,N_19218);
nand U21427 (N_21427,N_19541,N_18238);
nand U21428 (N_21428,N_18687,N_19511);
nand U21429 (N_21429,N_18419,N_19271);
nor U21430 (N_21430,N_19405,N_19056);
xor U21431 (N_21431,N_19051,N_18108);
nand U21432 (N_21432,N_19607,N_19994);
or U21433 (N_21433,N_19347,N_18048);
nand U21434 (N_21434,N_19942,N_18085);
xnor U21435 (N_21435,N_18935,N_18836);
nand U21436 (N_21436,N_19351,N_19933);
nand U21437 (N_21437,N_18531,N_19358);
nor U21438 (N_21438,N_18114,N_18688);
and U21439 (N_21439,N_19210,N_19366);
nor U21440 (N_21440,N_18878,N_19423);
nand U21441 (N_21441,N_19841,N_18392);
nor U21442 (N_21442,N_18964,N_19436);
xnor U21443 (N_21443,N_18480,N_19254);
nand U21444 (N_21444,N_18067,N_18234);
xnor U21445 (N_21445,N_19805,N_18447);
xor U21446 (N_21446,N_18617,N_19700);
or U21447 (N_21447,N_18342,N_18462);
nor U21448 (N_21448,N_19013,N_19765);
xor U21449 (N_21449,N_18061,N_18186);
nand U21450 (N_21450,N_18174,N_18161);
nand U21451 (N_21451,N_18769,N_19045);
and U21452 (N_21452,N_19760,N_19322);
nand U21453 (N_21453,N_19780,N_19944);
nor U21454 (N_21454,N_19495,N_18135);
nand U21455 (N_21455,N_19377,N_19486);
nor U21456 (N_21456,N_18989,N_18104);
nor U21457 (N_21457,N_18191,N_18196);
xor U21458 (N_21458,N_19859,N_18187);
and U21459 (N_21459,N_19787,N_19054);
nand U21460 (N_21460,N_19322,N_18971);
or U21461 (N_21461,N_18183,N_19960);
or U21462 (N_21462,N_19765,N_19301);
nand U21463 (N_21463,N_18392,N_18922);
nor U21464 (N_21464,N_19232,N_19202);
nand U21465 (N_21465,N_19669,N_19490);
nand U21466 (N_21466,N_18905,N_19567);
xor U21467 (N_21467,N_19904,N_18485);
and U21468 (N_21468,N_19774,N_18107);
xnor U21469 (N_21469,N_18548,N_18511);
or U21470 (N_21470,N_19910,N_18507);
nand U21471 (N_21471,N_19893,N_19031);
nand U21472 (N_21472,N_18176,N_18443);
xnor U21473 (N_21473,N_19813,N_19667);
nand U21474 (N_21474,N_19603,N_19639);
nor U21475 (N_21475,N_19280,N_18291);
or U21476 (N_21476,N_18982,N_19449);
nor U21477 (N_21477,N_18117,N_18158);
or U21478 (N_21478,N_18813,N_19118);
xor U21479 (N_21479,N_19915,N_18552);
nand U21480 (N_21480,N_19839,N_18695);
or U21481 (N_21481,N_19940,N_18184);
and U21482 (N_21482,N_18761,N_19444);
and U21483 (N_21483,N_18504,N_19403);
and U21484 (N_21484,N_19622,N_18773);
xor U21485 (N_21485,N_19984,N_18502);
and U21486 (N_21486,N_18857,N_19528);
nand U21487 (N_21487,N_19898,N_18070);
nor U21488 (N_21488,N_18766,N_18649);
or U21489 (N_21489,N_18033,N_19002);
or U21490 (N_21490,N_18400,N_19540);
xnor U21491 (N_21491,N_19165,N_18864);
and U21492 (N_21492,N_19211,N_18127);
nor U21493 (N_21493,N_19384,N_19158);
nand U21494 (N_21494,N_18023,N_18392);
xnor U21495 (N_21495,N_19951,N_18112);
nor U21496 (N_21496,N_19654,N_19541);
nor U21497 (N_21497,N_18760,N_18137);
xor U21498 (N_21498,N_19619,N_18488);
nor U21499 (N_21499,N_19187,N_18156);
and U21500 (N_21500,N_18703,N_19962);
nor U21501 (N_21501,N_18556,N_18300);
nor U21502 (N_21502,N_18815,N_18866);
and U21503 (N_21503,N_19356,N_18615);
and U21504 (N_21504,N_19868,N_18543);
nand U21505 (N_21505,N_18935,N_19693);
xor U21506 (N_21506,N_19948,N_18288);
nor U21507 (N_21507,N_19143,N_19110);
and U21508 (N_21508,N_19820,N_19088);
nand U21509 (N_21509,N_18187,N_18707);
nand U21510 (N_21510,N_18726,N_18395);
nand U21511 (N_21511,N_19779,N_19895);
and U21512 (N_21512,N_19964,N_18476);
nand U21513 (N_21513,N_18526,N_18110);
or U21514 (N_21514,N_19271,N_18713);
or U21515 (N_21515,N_19569,N_19075);
nor U21516 (N_21516,N_18076,N_18921);
or U21517 (N_21517,N_19095,N_18187);
or U21518 (N_21518,N_18534,N_19844);
nor U21519 (N_21519,N_18383,N_18246);
nor U21520 (N_21520,N_18739,N_19094);
nor U21521 (N_21521,N_18662,N_18450);
xnor U21522 (N_21522,N_19647,N_19961);
or U21523 (N_21523,N_18211,N_18120);
nor U21524 (N_21524,N_18544,N_18445);
xor U21525 (N_21525,N_18364,N_18853);
xnor U21526 (N_21526,N_18204,N_18929);
and U21527 (N_21527,N_19721,N_18184);
xor U21528 (N_21528,N_19958,N_18321);
or U21529 (N_21529,N_19849,N_19978);
and U21530 (N_21530,N_19511,N_18121);
or U21531 (N_21531,N_18921,N_18249);
nor U21532 (N_21532,N_18131,N_19011);
and U21533 (N_21533,N_19723,N_18838);
xnor U21534 (N_21534,N_19820,N_18451);
nor U21535 (N_21535,N_18491,N_19270);
nor U21536 (N_21536,N_19194,N_18702);
and U21537 (N_21537,N_19215,N_19978);
nand U21538 (N_21538,N_18266,N_19724);
xor U21539 (N_21539,N_18306,N_19545);
or U21540 (N_21540,N_19737,N_19756);
nor U21541 (N_21541,N_19671,N_18606);
or U21542 (N_21542,N_18659,N_18912);
nor U21543 (N_21543,N_18085,N_19499);
xnor U21544 (N_21544,N_18667,N_19469);
nand U21545 (N_21545,N_18965,N_18203);
nand U21546 (N_21546,N_19161,N_18616);
nor U21547 (N_21547,N_18483,N_18294);
xnor U21548 (N_21548,N_18108,N_19499);
or U21549 (N_21549,N_18162,N_19524);
or U21550 (N_21550,N_19882,N_18868);
nor U21551 (N_21551,N_18750,N_18628);
and U21552 (N_21552,N_18823,N_19998);
nand U21553 (N_21553,N_18167,N_19986);
xnor U21554 (N_21554,N_19011,N_18723);
nand U21555 (N_21555,N_18302,N_18258);
or U21556 (N_21556,N_18088,N_19703);
or U21557 (N_21557,N_18473,N_19538);
and U21558 (N_21558,N_18311,N_19523);
nand U21559 (N_21559,N_19788,N_18301);
xor U21560 (N_21560,N_18279,N_19705);
nor U21561 (N_21561,N_19891,N_18680);
and U21562 (N_21562,N_18142,N_18092);
and U21563 (N_21563,N_19556,N_18217);
nand U21564 (N_21564,N_18820,N_18680);
nand U21565 (N_21565,N_18267,N_19981);
xnor U21566 (N_21566,N_18527,N_18547);
and U21567 (N_21567,N_19856,N_18089);
or U21568 (N_21568,N_19074,N_19037);
or U21569 (N_21569,N_19502,N_18428);
nor U21570 (N_21570,N_18297,N_19344);
nand U21571 (N_21571,N_19756,N_18079);
xor U21572 (N_21572,N_19328,N_19737);
nand U21573 (N_21573,N_19271,N_19650);
nor U21574 (N_21574,N_19629,N_19165);
and U21575 (N_21575,N_18735,N_18142);
and U21576 (N_21576,N_19399,N_18433);
nor U21577 (N_21577,N_19924,N_18453);
or U21578 (N_21578,N_19283,N_19966);
or U21579 (N_21579,N_19478,N_18219);
nor U21580 (N_21580,N_19285,N_19577);
xnor U21581 (N_21581,N_18674,N_19351);
or U21582 (N_21582,N_19029,N_18222);
nor U21583 (N_21583,N_18070,N_18512);
or U21584 (N_21584,N_18466,N_18957);
xnor U21585 (N_21585,N_18199,N_19590);
and U21586 (N_21586,N_19479,N_18984);
nor U21587 (N_21587,N_18032,N_18773);
xor U21588 (N_21588,N_19879,N_18015);
and U21589 (N_21589,N_18894,N_18767);
nor U21590 (N_21590,N_19689,N_18190);
or U21591 (N_21591,N_19734,N_18786);
and U21592 (N_21592,N_19766,N_18925);
xor U21593 (N_21593,N_18807,N_18699);
xor U21594 (N_21594,N_19708,N_19244);
xnor U21595 (N_21595,N_18798,N_19430);
and U21596 (N_21596,N_18842,N_19161);
and U21597 (N_21597,N_19524,N_18060);
nand U21598 (N_21598,N_18452,N_19403);
nor U21599 (N_21599,N_19443,N_19706);
and U21600 (N_21600,N_18890,N_18892);
xnor U21601 (N_21601,N_19237,N_18000);
or U21602 (N_21602,N_18456,N_18015);
and U21603 (N_21603,N_18221,N_18795);
or U21604 (N_21604,N_18499,N_19539);
xor U21605 (N_21605,N_19846,N_18608);
xor U21606 (N_21606,N_18713,N_19524);
nor U21607 (N_21607,N_19819,N_18442);
nand U21608 (N_21608,N_19724,N_19308);
and U21609 (N_21609,N_19518,N_18348);
and U21610 (N_21610,N_19756,N_18596);
and U21611 (N_21611,N_19588,N_19004);
nand U21612 (N_21612,N_19563,N_19692);
or U21613 (N_21613,N_18790,N_18165);
nor U21614 (N_21614,N_19932,N_18649);
or U21615 (N_21615,N_19120,N_19988);
xnor U21616 (N_21616,N_18425,N_19468);
xor U21617 (N_21617,N_19708,N_19760);
or U21618 (N_21618,N_18421,N_18717);
nor U21619 (N_21619,N_19822,N_19153);
xor U21620 (N_21620,N_18652,N_19171);
nand U21621 (N_21621,N_19069,N_18239);
xnor U21622 (N_21622,N_18653,N_18572);
or U21623 (N_21623,N_18002,N_18741);
nand U21624 (N_21624,N_18929,N_18604);
xor U21625 (N_21625,N_19778,N_18763);
xnor U21626 (N_21626,N_18068,N_18055);
nor U21627 (N_21627,N_18502,N_18590);
xnor U21628 (N_21628,N_18077,N_18751);
and U21629 (N_21629,N_18889,N_19215);
nor U21630 (N_21630,N_19547,N_18583);
nor U21631 (N_21631,N_19247,N_19396);
nor U21632 (N_21632,N_18798,N_18165);
nor U21633 (N_21633,N_19364,N_18900);
nand U21634 (N_21634,N_19109,N_18130);
xnor U21635 (N_21635,N_19683,N_19746);
xnor U21636 (N_21636,N_19220,N_18675);
nor U21637 (N_21637,N_18783,N_19217);
nor U21638 (N_21638,N_18462,N_19238);
or U21639 (N_21639,N_19587,N_18312);
or U21640 (N_21640,N_19453,N_18979);
and U21641 (N_21641,N_19750,N_18132);
or U21642 (N_21642,N_18999,N_18350);
nor U21643 (N_21643,N_19603,N_18776);
xnor U21644 (N_21644,N_18117,N_19022);
xor U21645 (N_21645,N_19154,N_19075);
nand U21646 (N_21646,N_18808,N_19585);
or U21647 (N_21647,N_18079,N_19137);
nor U21648 (N_21648,N_19822,N_19218);
or U21649 (N_21649,N_19971,N_19978);
or U21650 (N_21650,N_18821,N_18667);
nor U21651 (N_21651,N_18184,N_19705);
nor U21652 (N_21652,N_19682,N_19236);
xnor U21653 (N_21653,N_19394,N_19866);
or U21654 (N_21654,N_18867,N_18269);
nand U21655 (N_21655,N_18179,N_19809);
nand U21656 (N_21656,N_19497,N_19776);
nand U21657 (N_21657,N_18403,N_19342);
and U21658 (N_21658,N_19850,N_18531);
nor U21659 (N_21659,N_18307,N_19678);
xnor U21660 (N_21660,N_19210,N_18666);
xor U21661 (N_21661,N_18492,N_18041);
nand U21662 (N_21662,N_19040,N_19421);
or U21663 (N_21663,N_19320,N_18366);
nor U21664 (N_21664,N_18585,N_19590);
nand U21665 (N_21665,N_18801,N_18588);
nor U21666 (N_21666,N_19775,N_18550);
and U21667 (N_21667,N_19496,N_18899);
xnor U21668 (N_21668,N_18519,N_19344);
nand U21669 (N_21669,N_19925,N_19464);
or U21670 (N_21670,N_18297,N_19916);
xor U21671 (N_21671,N_18691,N_19568);
nand U21672 (N_21672,N_18554,N_19802);
nand U21673 (N_21673,N_19914,N_19660);
nand U21674 (N_21674,N_19025,N_19513);
nor U21675 (N_21675,N_19735,N_19547);
and U21676 (N_21676,N_18367,N_18188);
nand U21677 (N_21677,N_19314,N_18305);
and U21678 (N_21678,N_18782,N_18246);
or U21679 (N_21679,N_19926,N_19270);
and U21680 (N_21680,N_18127,N_18865);
and U21681 (N_21681,N_19555,N_18866);
or U21682 (N_21682,N_19839,N_19029);
nand U21683 (N_21683,N_18685,N_19459);
nor U21684 (N_21684,N_19954,N_19410);
nand U21685 (N_21685,N_19620,N_19327);
nand U21686 (N_21686,N_18886,N_18069);
nand U21687 (N_21687,N_19479,N_19864);
and U21688 (N_21688,N_19752,N_18693);
nand U21689 (N_21689,N_18752,N_18744);
nand U21690 (N_21690,N_19595,N_18880);
xnor U21691 (N_21691,N_19348,N_19453);
nand U21692 (N_21692,N_19310,N_18800);
xor U21693 (N_21693,N_18375,N_19177);
xor U21694 (N_21694,N_18943,N_19670);
nor U21695 (N_21695,N_18853,N_18005);
xnor U21696 (N_21696,N_18760,N_18586);
and U21697 (N_21697,N_19937,N_19276);
or U21698 (N_21698,N_19393,N_19024);
and U21699 (N_21699,N_18056,N_19877);
nand U21700 (N_21700,N_18626,N_19326);
nor U21701 (N_21701,N_18121,N_18570);
and U21702 (N_21702,N_19306,N_19526);
and U21703 (N_21703,N_18822,N_19549);
or U21704 (N_21704,N_19712,N_18087);
and U21705 (N_21705,N_19484,N_19810);
and U21706 (N_21706,N_19111,N_18921);
nand U21707 (N_21707,N_19883,N_19027);
nand U21708 (N_21708,N_18680,N_18586);
or U21709 (N_21709,N_18805,N_18735);
nor U21710 (N_21710,N_18884,N_18472);
xor U21711 (N_21711,N_19737,N_18889);
and U21712 (N_21712,N_18559,N_18333);
nor U21713 (N_21713,N_19352,N_18738);
and U21714 (N_21714,N_18092,N_19854);
xnor U21715 (N_21715,N_18535,N_19153);
xor U21716 (N_21716,N_19372,N_18696);
nand U21717 (N_21717,N_18760,N_18280);
or U21718 (N_21718,N_18629,N_19852);
xor U21719 (N_21719,N_18135,N_19097);
or U21720 (N_21720,N_18499,N_19303);
or U21721 (N_21721,N_18018,N_19124);
and U21722 (N_21722,N_18510,N_18104);
nor U21723 (N_21723,N_19827,N_19840);
nor U21724 (N_21724,N_19999,N_18711);
and U21725 (N_21725,N_18643,N_18335);
nand U21726 (N_21726,N_18468,N_19658);
xor U21727 (N_21727,N_18374,N_19725);
or U21728 (N_21728,N_18888,N_19219);
nand U21729 (N_21729,N_18945,N_19067);
nor U21730 (N_21730,N_18931,N_19657);
nor U21731 (N_21731,N_18847,N_18092);
or U21732 (N_21732,N_19110,N_18886);
xor U21733 (N_21733,N_19216,N_19616);
nor U21734 (N_21734,N_19095,N_19368);
and U21735 (N_21735,N_19492,N_18814);
nor U21736 (N_21736,N_19955,N_19023);
or U21737 (N_21737,N_19890,N_18141);
or U21738 (N_21738,N_18086,N_18534);
nor U21739 (N_21739,N_18535,N_18886);
or U21740 (N_21740,N_18766,N_18010);
nor U21741 (N_21741,N_18547,N_19628);
nor U21742 (N_21742,N_19502,N_18655);
nand U21743 (N_21743,N_19377,N_19754);
and U21744 (N_21744,N_19486,N_18730);
or U21745 (N_21745,N_19945,N_18114);
nor U21746 (N_21746,N_19730,N_19188);
or U21747 (N_21747,N_19946,N_19899);
nor U21748 (N_21748,N_19276,N_19836);
or U21749 (N_21749,N_19758,N_18521);
and U21750 (N_21750,N_19842,N_18918);
or U21751 (N_21751,N_18178,N_18357);
nand U21752 (N_21752,N_19055,N_19880);
and U21753 (N_21753,N_19631,N_18827);
or U21754 (N_21754,N_19745,N_19402);
and U21755 (N_21755,N_18442,N_19579);
and U21756 (N_21756,N_19569,N_18027);
xor U21757 (N_21757,N_18385,N_18553);
and U21758 (N_21758,N_18479,N_19914);
nand U21759 (N_21759,N_19466,N_19773);
nand U21760 (N_21760,N_19031,N_19962);
xnor U21761 (N_21761,N_18848,N_19849);
nand U21762 (N_21762,N_18372,N_19967);
nand U21763 (N_21763,N_18747,N_19803);
nor U21764 (N_21764,N_18023,N_18895);
or U21765 (N_21765,N_18423,N_18415);
and U21766 (N_21766,N_18232,N_18930);
or U21767 (N_21767,N_18055,N_18706);
nor U21768 (N_21768,N_18711,N_18468);
xor U21769 (N_21769,N_18106,N_18113);
xnor U21770 (N_21770,N_18566,N_19316);
or U21771 (N_21771,N_18112,N_19388);
or U21772 (N_21772,N_19305,N_19324);
and U21773 (N_21773,N_18431,N_19669);
nand U21774 (N_21774,N_18953,N_18593);
or U21775 (N_21775,N_18715,N_18956);
or U21776 (N_21776,N_19905,N_19325);
xnor U21777 (N_21777,N_19338,N_18048);
nand U21778 (N_21778,N_18754,N_19901);
xnor U21779 (N_21779,N_19331,N_18771);
and U21780 (N_21780,N_19141,N_19420);
nand U21781 (N_21781,N_19849,N_18697);
or U21782 (N_21782,N_19840,N_18202);
or U21783 (N_21783,N_18413,N_18751);
nor U21784 (N_21784,N_19241,N_19369);
nor U21785 (N_21785,N_19663,N_19005);
nand U21786 (N_21786,N_18282,N_19897);
nor U21787 (N_21787,N_18920,N_19351);
nor U21788 (N_21788,N_18828,N_18476);
nand U21789 (N_21789,N_18170,N_19660);
or U21790 (N_21790,N_19129,N_19499);
and U21791 (N_21791,N_19436,N_19591);
nand U21792 (N_21792,N_18783,N_18877);
nand U21793 (N_21793,N_18520,N_18125);
or U21794 (N_21794,N_19096,N_19498);
nor U21795 (N_21795,N_18296,N_19313);
nor U21796 (N_21796,N_19428,N_18266);
or U21797 (N_21797,N_19642,N_18846);
xor U21798 (N_21798,N_18733,N_19387);
xnor U21799 (N_21799,N_19468,N_19702);
or U21800 (N_21800,N_19021,N_18648);
nand U21801 (N_21801,N_18826,N_18513);
nand U21802 (N_21802,N_19721,N_18769);
and U21803 (N_21803,N_19712,N_19995);
nand U21804 (N_21804,N_18063,N_18516);
or U21805 (N_21805,N_18423,N_19805);
nor U21806 (N_21806,N_18102,N_18275);
and U21807 (N_21807,N_19104,N_18006);
and U21808 (N_21808,N_18407,N_18573);
nor U21809 (N_21809,N_18279,N_18558);
or U21810 (N_21810,N_18490,N_18775);
or U21811 (N_21811,N_18618,N_19983);
nand U21812 (N_21812,N_19311,N_18782);
xnor U21813 (N_21813,N_18421,N_19247);
nor U21814 (N_21814,N_18981,N_19795);
xor U21815 (N_21815,N_18090,N_18945);
nand U21816 (N_21816,N_18236,N_18099);
nor U21817 (N_21817,N_18790,N_19408);
nor U21818 (N_21818,N_19846,N_19575);
nor U21819 (N_21819,N_19287,N_19098);
xnor U21820 (N_21820,N_18618,N_18483);
nand U21821 (N_21821,N_19396,N_19045);
and U21822 (N_21822,N_18678,N_19907);
and U21823 (N_21823,N_19797,N_18670);
nor U21824 (N_21824,N_18385,N_18701);
xor U21825 (N_21825,N_19201,N_18777);
nor U21826 (N_21826,N_18201,N_19885);
nand U21827 (N_21827,N_18571,N_19657);
and U21828 (N_21828,N_18671,N_18857);
nand U21829 (N_21829,N_19163,N_19291);
nand U21830 (N_21830,N_19258,N_19215);
or U21831 (N_21831,N_19583,N_19924);
or U21832 (N_21832,N_19010,N_18867);
or U21833 (N_21833,N_18114,N_18117);
nand U21834 (N_21834,N_19804,N_18988);
nor U21835 (N_21835,N_18201,N_18988);
or U21836 (N_21836,N_19710,N_18205);
or U21837 (N_21837,N_18761,N_18137);
xor U21838 (N_21838,N_18972,N_19055);
or U21839 (N_21839,N_18742,N_19119);
or U21840 (N_21840,N_18581,N_19511);
nand U21841 (N_21841,N_18388,N_18782);
nand U21842 (N_21842,N_18672,N_19245);
nor U21843 (N_21843,N_19087,N_18132);
or U21844 (N_21844,N_18782,N_19955);
xnor U21845 (N_21845,N_18080,N_18647);
nand U21846 (N_21846,N_18805,N_19259);
and U21847 (N_21847,N_18339,N_18604);
nor U21848 (N_21848,N_19300,N_18639);
nor U21849 (N_21849,N_18771,N_18592);
and U21850 (N_21850,N_18396,N_19506);
xor U21851 (N_21851,N_19952,N_18674);
or U21852 (N_21852,N_19284,N_19827);
or U21853 (N_21853,N_18225,N_18738);
nand U21854 (N_21854,N_18601,N_18491);
nand U21855 (N_21855,N_19059,N_19583);
and U21856 (N_21856,N_18902,N_18102);
nor U21857 (N_21857,N_18482,N_19826);
and U21858 (N_21858,N_19552,N_19821);
nand U21859 (N_21859,N_19196,N_18429);
nor U21860 (N_21860,N_19554,N_19070);
xnor U21861 (N_21861,N_19573,N_19923);
and U21862 (N_21862,N_18578,N_18291);
nand U21863 (N_21863,N_19548,N_19666);
nand U21864 (N_21864,N_18944,N_18735);
xnor U21865 (N_21865,N_19251,N_18703);
or U21866 (N_21866,N_19315,N_18467);
and U21867 (N_21867,N_19363,N_19133);
or U21868 (N_21868,N_18171,N_18134);
xor U21869 (N_21869,N_18368,N_19610);
and U21870 (N_21870,N_19560,N_18095);
xor U21871 (N_21871,N_19945,N_18176);
and U21872 (N_21872,N_19811,N_19369);
nand U21873 (N_21873,N_19720,N_18202);
nand U21874 (N_21874,N_18704,N_18522);
and U21875 (N_21875,N_19894,N_19884);
nor U21876 (N_21876,N_19937,N_18449);
and U21877 (N_21877,N_18188,N_18517);
or U21878 (N_21878,N_18487,N_18995);
xor U21879 (N_21879,N_19091,N_19599);
nor U21880 (N_21880,N_19148,N_19012);
or U21881 (N_21881,N_18952,N_18592);
or U21882 (N_21882,N_19856,N_18312);
xnor U21883 (N_21883,N_19477,N_18936);
or U21884 (N_21884,N_18456,N_18615);
nor U21885 (N_21885,N_19932,N_19411);
nand U21886 (N_21886,N_19140,N_19517);
xor U21887 (N_21887,N_19514,N_18453);
xnor U21888 (N_21888,N_19074,N_19605);
xnor U21889 (N_21889,N_18247,N_18641);
nor U21890 (N_21890,N_19450,N_19486);
nand U21891 (N_21891,N_18600,N_18407);
or U21892 (N_21892,N_19223,N_19850);
and U21893 (N_21893,N_19081,N_18019);
or U21894 (N_21894,N_19395,N_19796);
and U21895 (N_21895,N_18608,N_18629);
nor U21896 (N_21896,N_19974,N_18090);
and U21897 (N_21897,N_19703,N_19296);
and U21898 (N_21898,N_18820,N_18486);
and U21899 (N_21899,N_19914,N_19217);
xnor U21900 (N_21900,N_18812,N_18796);
nor U21901 (N_21901,N_19201,N_19692);
xnor U21902 (N_21902,N_18595,N_19969);
nand U21903 (N_21903,N_19851,N_19601);
nor U21904 (N_21904,N_18014,N_18640);
nand U21905 (N_21905,N_19934,N_18444);
nor U21906 (N_21906,N_19800,N_19165);
nor U21907 (N_21907,N_18612,N_18685);
or U21908 (N_21908,N_18454,N_19300);
nand U21909 (N_21909,N_18301,N_18866);
or U21910 (N_21910,N_19846,N_18962);
nor U21911 (N_21911,N_19345,N_18578);
and U21912 (N_21912,N_18342,N_19721);
and U21913 (N_21913,N_18031,N_18822);
or U21914 (N_21914,N_18737,N_18047);
nor U21915 (N_21915,N_18052,N_19670);
xor U21916 (N_21916,N_18823,N_18125);
nor U21917 (N_21917,N_19267,N_19961);
or U21918 (N_21918,N_18942,N_19656);
nand U21919 (N_21919,N_19867,N_18202);
xnor U21920 (N_21920,N_19377,N_18378);
nand U21921 (N_21921,N_18308,N_18378);
nor U21922 (N_21922,N_19827,N_19388);
nand U21923 (N_21923,N_19011,N_18279);
nand U21924 (N_21924,N_18525,N_19458);
or U21925 (N_21925,N_18862,N_19372);
or U21926 (N_21926,N_18577,N_18222);
nand U21927 (N_21927,N_18492,N_19925);
nand U21928 (N_21928,N_18529,N_18517);
xor U21929 (N_21929,N_19385,N_19725);
xnor U21930 (N_21930,N_19193,N_19652);
nand U21931 (N_21931,N_18009,N_19925);
xor U21932 (N_21932,N_18867,N_19886);
xnor U21933 (N_21933,N_19852,N_18953);
xnor U21934 (N_21934,N_19904,N_19804);
nor U21935 (N_21935,N_19076,N_18245);
and U21936 (N_21936,N_18001,N_18502);
nor U21937 (N_21937,N_18918,N_18899);
nor U21938 (N_21938,N_18291,N_19978);
nand U21939 (N_21939,N_18450,N_18792);
and U21940 (N_21940,N_19333,N_19443);
xnor U21941 (N_21941,N_19897,N_19512);
and U21942 (N_21942,N_18112,N_18724);
nand U21943 (N_21943,N_19822,N_18830);
and U21944 (N_21944,N_18753,N_18992);
xor U21945 (N_21945,N_19736,N_19903);
nor U21946 (N_21946,N_18694,N_19986);
and U21947 (N_21947,N_18907,N_19291);
nor U21948 (N_21948,N_18483,N_19532);
or U21949 (N_21949,N_19022,N_19371);
nor U21950 (N_21950,N_18214,N_18607);
and U21951 (N_21951,N_19023,N_19862);
and U21952 (N_21952,N_18075,N_19974);
nand U21953 (N_21953,N_19966,N_18339);
nand U21954 (N_21954,N_19117,N_19632);
and U21955 (N_21955,N_19885,N_19821);
nand U21956 (N_21956,N_19160,N_19887);
xnor U21957 (N_21957,N_19595,N_19648);
nand U21958 (N_21958,N_19375,N_18054);
or U21959 (N_21959,N_19321,N_19016);
and U21960 (N_21960,N_18293,N_18786);
nand U21961 (N_21961,N_19917,N_18063);
xor U21962 (N_21962,N_18163,N_19754);
or U21963 (N_21963,N_18171,N_19760);
nand U21964 (N_21964,N_19386,N_18640);
or U21965 (N_21965,N_19701,N_18935);
xnor U21966 (N_21966,N_18055,N_19290);
and U21967 (N_21967,N_19189,N_18555);
and U21968 (N_21968,N_18783,N_19466);
and U21969 (N_21969,N_19831,N_19071);
nand U21970 (N_21970,N_18597,N_19661);
nor U21971 (N_21971,N_19364,N_18930);
or U21972 (N_21972,N_19550,N_19806);
xor U21973 (N_21973,N_19423,N_19693);
nand U21974 (N_21974,N_19457,N_18284);
nor U21975 (N_21975,N_18476,N_18493);
nand U21976 (N_21976,N_19537,N_19894);
nand U21977 (N_21977,N_18300,N_18035);
or U21978 (N_21978,N_18482,N_19146);
or U21979 (N_21979,N_18897,N_18033);
nor U21980 (N_21980,N_19551,N_19838);
or U21981 (N_21981,N_18329,N_18744);
nand U21982 (N_21982,N_19902,N_18548);
or U21983 (N_21983,N_18638,N_19704);
nor U21984 (N_21984,N_18917,N_18107);
and U21985 (N_21985,N_19027,N_18036);
nor U21986 (N_21986,N_18841,N_19619);
and U21987 (N_21987,N_18879,N_18814);
nand U21988 (N_21988,N_19049,N_19340);
xnor U21989 (N_21989,N_18904,N_18482);
nand U21990 (N_21990,N_18119,N_19931);
and U21991 (N_21991,N_18705,N_18196);
nand U21992 (N_21992,N_19839,N_19748);
nor U21993 (N_21993,N_18406,N_19403);
nand U21994 (N_21994,N_19461,N_18545);
and U21995 (N_21995,N_18857,N_18888);
or U21996 (N_21996,N_19813,N_19608);
nor U21997 (N_21997,N_19993,N_19992);
and U21998 (N_21998,N_19580,N_19836);
nand U21999 (N_21999,N_19415,N_19717);
and U22000 (N_22000,N_21225,N_21499);
xnor U22001 (N_22001,N_20242,N_21368);
and U22002 (N_22002,N_20299,N_21553);
and U22003 (N_22003,N_21566,N_21985);
or U22004 (N_22004,N_21458,N_20567);
nand U22005 (N_22005,N_20525,N_21496);
xor U22006 (N_22006,N_21949,N_20026);
xor U22007 (N_22007,N_21526,N_20589);
xnor U22008 (N_22008,N_20392,N_20877);
and U22009 (N_22009,N_21835,N_20894);
or U22010 (N_22010,N_21461,N_20427);
xnor U22011 (N_22011,N_20259,N_21495);
xor U22012 (N_22012,N_21989,N_20924);
nor U22013 (N_22013,N_21921,N_20043);
nor U22014 (N_22014,N_21884,N_20393);
nand U22015 (N_22015,N_21044,N_21264);
nor U22016 (N_22016,N_20433,N_20241);
and U22017 (N_22017,N_20276,N_21250);
nor U22018 (N_22018,N_20733,N_21279);
or U22019 (N_22019,N_20926,N_20155);
nand U22020 (N_22020,N_20701,N_21518);
xor U22021 (N_22021,N_21951,N_21386);
and U22022 (N_22022,N_20278,N_20360);
or U22023 (N_22023,N_21986,N_21163);
and U22024 (N_22024,N_21826,N_20157);
or U22025 (N_22025,N_21789,N_20267);
and U22026 (N_22026,N_20871,N_21018);
nand U22027 (N_22027,N_20369,N_21750);
or U22028 (N_22028,N_20725,N_20576);
or U22029 (N_22029,N_21669,N_20014);
or U22030 (N_22030,N_20072,N_20847);
or U22031 (N_22031,N_21093,N_21374);
or U22032 (N_22032,N_21142,N_20657);
nor U22033 (N_22033,N_20776,N_21110);
and U22034 (N_22034,N_21085,N_20321);
xnor U22035 (N_22035,N_21170,N_21497);
xor U22036 (N_22036,N_20874,N_20731);
or U22037 (N_22037,N_21628,N_21603);
nand U22038 (N_22038,N_21684,N_21530);
nand U22039 (N_22039,N_20575,N_20958);
or U22040 (N_22040,N_20688,N_21622);
nand U22041 (N_22041,N_21737,N_20068);
and U22042 (N_22042,N_20250,N_21834);
nand U22043 (N_22043,N_21854,N_21840);
or U22044 (N_22044,N_21412,N_20969);
xnor U22045 (N_22045,N_20451,N_21094);
and U22046 (N_22046,N_21886,N_21008);
nand U22047 (N_22047,N_20206,N_20856);
xor U22048 (N_22048,N_20312,N_21166);
xor U22049 (N_22049,N_21697,N_21156);
nor U22050 (N_22050,N_20448,N_20109);
xnor U22051 (N_22051,N_20234,N_20006);
and U22052 (N_22052,N_21892,N_20611);
nand U22053 (N_22053,N_20236,N_20971);
and U22054 (N_22054,N_20495,N_21539);
nand U22055 (N_22055,N_21514,N_21294);
nor U22056 (N_22056,N_21792,N_21592);
or U22057 (N_22057,N_20459,N_20395);
or U22058 (N_22058,N_21925,N_21708);
or U22059 (N_22059,N_21210,N_21372);
xnor U22060 (N_22060,N_20141,N_21355);
or U22061 (N_22061,N_20474,N_21720);
and U22062 (N_22062,N_21274,N_20097);
nand U22063 (N_22063,N_20981,N_21425);
xor U22064 (N_22064,N_21112,N_20119);
nand U22065 (N_22065,N_21994,N_21842);
nand U22066 (N_22066,N_21390,N_20309);
or U22067 (N_22067,N_20516,N_21931);
xnor U22068 (N_22068,N_20686,N_20216);
nand U22069 (N_22069,N_21626,N_20202);
or U22070 (N_22070,N_21005,N_20770);
or U22071 (N_22071,N_20316,N_21290);
and U22072 (N_22072,N_20844,N_21984);
or U22073 (N_22073,N_20934,N_20983);
nor U22074 (N_22074,N_21728,N_20005);
xor U22075 (N_22075,N_20868,N_21455);
nand U22076 (N_22076,N_20092,N_21379);
nand U22077 (N_22077,N_20801,N_20698);
nand U22078 (N_22078,N_21267,N_20809);
and U22079 (N_22079,N_21158,N_20573);
xor U22080 (N_22080,N_21464,N_21689);
and U22081 (N_22081,N_20941,N_20923);
or U22082 (N_22082,N_20358,N_20619);
and U22083 (N_22083,N_20491,N_21024);
xnor U22084 (N_22084,N_20830,N_20446);
and U22085 (N_22085,N_21117,N_20886);
xor U22086 (N_22086,N_20115,N_21244);
and U22087 (N_22087,N_21492,N_20381);
and U22088 (N_22088,N_20936,N_21908);
or U22089 (N_22089,N_21895,N_20489);
and U22090 (N_22090,N_21661,N_20722);
xnor U22091 (N_22091,N_21215,N_21263);
nand U22092 (N_22092,N_21269,N_21249);
nand U22093 (N_22093,N_21585,N_21467);
and U22094 (N_22094,N_21508,N_20948);
and U22095 (N_22095,N_21993,N_20633);
nor U22096 (N_22096,N_21111,N_21798);
and U22097 (N_22097,N_20728,N_20095);
nor U22098 (N_22098,N_21659,N_21043);
and U22099 (N_22099,N_20838,N_21680);
nand U22100 (N_22100,N_21183,N_20214);
nor U22101 (N_22101,N_21880,N_21990);
nor U22102 (N_22102,N_20270,N_21871);
or U22103 (N_22103,N_20704,N_21296);
xor U22104 (N_22104,N_21820,N_21309);
xor U22105 (N_22105,N_21120,N_20080);
or U22106 (N_22106,N_21890,N_21083);
nand U22107 (N_22107,N_21050,N_21021);
nand U22108 (N_22108,N_21724,N_20246);
xnor U22109 (N_22109,N_21791,N_20028);
and U22110 (N_22110,N_20646,N_20314);
nor U22111 (N_22111,N_20001,N_20930);
nor U22112 (N_22112,N_21786,N_21537);
or U22113 (N_22113,N_21955,N_21741);
xnor U22114 (N_22114,N_21647,N_21541);
and U22115 (N_22115,N_20519,N_20558);
and U22116 (N_22116,N_21169,N_20238);
or U22117 (N_22117,N_21318,N_21181);
nand U22118 (N_22118,N_20617,N_21174);
or U22119 (N_22119,N_20424,N_21284);
or U22120 (N_22120,N_21730,N_21644);
or U22121 (N_22121,N_21221,N_20134);
or U22122 (N_22122,N_21838,N_21608);
and U22123 (N_22123,N_21339,N_21431);
or U22124 (N_22124,N_20213,N_20697);
and U22125 (N_22125,N_21002,N_20747);
or U22126 (N_22126,N_20771,N_20494);
xor U22127 (N_22127,N_21575,N_21056);
xor U22128 (N_22128,N_20088,N_21382);
and U22129 (N_22129,N_21247,N_21565);
xor U22130 (N_22130,N_21062,N_21883);
nand U22131 (N_22131,N_20414,N_21576);
nor U22132 (N_22132,N_20866,N_20881);
nor U22133 (N_22133,N_21941,N_21872);
and U22134 (N_22134,N_20305,N_20665);
nor U22135 (N_22135,N_21591,N_20779);
and U22136 (N_22136,N_21639,N_20922);
or U22137 (N_22137,N_20681,N_21362);
nor U22138 (N_22138,N_21573,N_21594);
xor U22139 (N_22139,N_20857,N_20648);
or U22140 (N_22140,N_20493,N_21630);
xor U22141 (N_22141,N_21175,N_20498);
nor U22142 (N_22142,N_21995,N_20501);
nand U22143 (N_22143,N_21182,N_20811);
or U22144 (N_22144,N_21760,N_21731);
and U22145 (N_22145,N_20029,N_20327);
or U22146 (N_22146,N_21303,N_20711);
nor U22147 (N_22147,N_21747,N_21195);
or U22148 (N_22148,N_21453,N_20613);
xor U22149 (N_22149,N_21223,N_21810);
nor U22150 (N_22150,N_21653,N_21818);
nor U22151 (N_22151,N_21119,N_20663);
xnor U22152 (N_22152,N_20917,N_21057);
or U22153 (N_22153,N_21329,N_21971);
and U22154 (N_22154,N_20705,N_20901);
xnor U22155 (N_22155,N_21700,N_21114);
nor U22156 (N_22156,N_20712,N_21214);
xor U22157 (N_22157,N_21668,N_21969);
and U22158 (N_22158,N_20222,N_21206);
and U22159 (N_22159,N_21462,N_20060);
or U22160 (N_22160,N_21614,N_21781);
nor U22161 (N_22161,N_20790,N_21729);
xnor U22162 (N_22162,N_20815,N_20081);
and U22163 (N_22163,N_21765,N_21635);
nor U22164 (N_22164,N_20674,N_21306);
nor U22165 (N_22165,N_21926,N_21652);
and U22166 (N_22166,N_20470,N_21547);
xnor U22167 (N_22167,N_20330,N_21634);
xor U22168 (N_22168,N_21108,N_21754);
or U22169 (N_22169,N_21470,N_21506);
or U22170 (N_22170,N_20162,N_20891);
or U22171 (N_22171,N_20528,N_20846);
and U22172 (N_22172,N_21270,N_21715);
or U22173 (N_22173,N_20129,N_21444);
nor U22174 (N_22174,N_21580,N_21289);
and U22175 (N_22175,N_21784,N_20375);
or U22176 (N_22176,N_20145,N_20825);
or U22177 (N_22177,N_20376,N_20650);
and U22178 (N_22178,N_20927,N_21437);
or U22179 (N_22179,N_20438,N_20773);
and U22180 (N_22180,N_21367,N_21681);
and U22181 (N_22181,N_21098,N_20428);
nand U22182 (N_22182,N_21824,N_21611);
xnor U22183 (N_22183,N_20535,N_21405);
nand U22184 (N_22184,N_21173,N_21920);
xor U22185 (N_22185,N_21293,N_20780);
and U22186 (N_22186,N_21311,N_20002);
or U22187 (N_22187,N_20911,N_20571);
nand U22188 (N_22188,N_21416,N_21945);
nor U22189 (N_22189,N_21651,N_20925);
nand U22190 (N_22190,N_20099,N_20378);
nand U22191 (N_22191,N_21755,N_20797);
nand U22192 (N_22192,N_21102,N_21642);
xnor U22193 (N_22193,N_20166,N_20082);
and U22194 (N_22194,N_21924,N_20398);
xor U22195 (N_22195,N_20225,N_21371);
or U22196 (N_22196,N_20729,N_20695);
xnor U22197 (N_22197,N_20091,N_21707);
and U22198 (N_22198,N_20070,N_21343);
and U22199 (N_22199,N_20892,N_21740);
and U22200 (N_22200,N_20828,N_21940);
and U22201 (N_22201,N_21189,N_20337);
nor U22202 (N_22202,N_21194,N_20929);
and U22203 (N_22203,N_21888,N_21488);
nand U22204 (N_22204,N_20518,N_20356);
or U22205 (N_22205,N_20384,N_21161);
xnor U22206 (N_22206,N_21099,N_21404);
xor U22207 (N_22207,N_21192,N_21352);
nor U22208 (N_22208,N_21947,N_20123);
or U22209 (N_22209,N_21507,N_20996);
nor U22210 (N_22210,N_20850,N_20713);
xor U22211 (N_22211,N_21257,N_20980);
nor U22212 (N_22212,N_20536,N_21275);
nand U22213 (N_22213,N_20757,N_21906);
or U22214 (N_22214,N_21430,N_20715);
nand U22215 (N_22215,N_20775,N_20986);
nor U22216 (N_22216,N_20034,N_20565);
nand U22217 (N_22217,N_21930,N_20122);
xor U22218 (N_22218,N_20689,N_21153);
nor U22219 (N_22219,N_20207,N_20482);
nor U22220 (N_22220,N_20346,N_20172);
and U22221 (N_22221,N_21191,N_21735);
and U22222 (N_22222,N_20988,N_21570);
or U22223 (N_22223,N_21751,N_20197);
and U22224 (N_22224,N_21678,N_20671);
and U22225 (N_22225,N_20921,N_20906);
xor U22226 (N_22226,N_20635,N_20508);
nand U22227 (N_22227,N_21271,N_20707);
nand U22228 (N_22228,N_20416,N_21889);
nand U22229 (N_22229,N_20914,N_20605);
nand U22230 (N_22230,N_20455,N_21481);
nand U22231 (N_22231,N_21616,N_20198);
nand U22232 (N_22232,N_21604,N_21615);
or U22233 (N_22233,N_20554,N_21956);
xnor U22234 (N_22234,N_21471,N_21081);
nor U22235 (N_22235,N_20945,N_20691);
nand U22236 (N_22236,N_20870,N_21981);
nor U22237 (N_22237,N_20177,N_21353);
and U22238 (N_22238,N_21109,N_20180);
nor U22239 (N_22239,N_20767,N_20763);
nor U22240 (N_22240,N_21685,N_21832);
nand U22241 (N_22241,N_21772,N_20593);
nand U22242 (N_22242,N_21693,N_20545);
nand U22243 (N_22243,N_21665,N_21236);
xnor U22244 (N_22244,N_20199,N_21843);
xnor U22245 (N_22245,N_21233,N_20908);
xnor U22246 (N_22246,N_21934,N_20677);
xnor U22247 (N_22247,N_21836,N_21746);
nor U22248 (N_22248,N_20984,N_21641);
nand U22249 (N_22249,N_20151,N_21314);
xnor U22250 (N_22250,N_20739,N_20524);
nor U22251 (N_22251,N_21793,N_21503);
nor U22252 (N_22252,N_20616,N_21426);
and U22253 (N_22253,N_21076,N_20461);
or U22254 (N_22254,N_21384,N_20897);
nand U22255 (N_22255,N_20916,N_20237);
nand U22256 (N_22256,N_21113,N_20702);
nor U22257 (N_22257,N_20140,N_21691);
and U22258 (N_22258,N_21582,N_21452);
nor U22259 (N_22259,N_21361,N_21330);
nor U22260 (N_22260,N_20253,N_20560);
and U22261 (N_22261,N_20003,N_21702);
or U22262 (N_22262,N_20890,N_21852);
or U22263 (N_22263,N_20420,N_21066);
xnor U22264 (N_22264,N_21317,N_20228);
xor U22265 (N_22265,N_20121,N_20302);
xor U22266 (N_22266,N_20319,N_20456);
nor U22267 (N_22267,N_20765,N_20585);
nor U22268 (N_22268,N_20840,N_21280);
and U22269 (N_22269,N_20506,N_20004);
and U22270 (N_22270,N_21992,N_21897);
nor U22271 (N_22271,N_20740,N_21283);
xnor U22272 (N_22272,N_20561,N_20854);
nor U22273 (N_22273,N_20709,N_21596);
xnor U22274 (N_22274,N_20872,N_21288);
or U22275 (N_22275,N_20876,N_21465);
nand U22276 (N_22276,N_21605,N_20325);
or U22277 (N_22277,N_20730,N_21184);
nor U22278 (N_22278,N_21898,N_21501);
nor U22279 (N_22279,N_21959,N_21468);
xnor U22280 (N_22280,N_20789,N_20193);
and U22281 (N_22281,N_20895,N_21116);
or U22282 (N_22282,N_21562,N_20557);
or U22283 (N_22283,N_21325,N_20819);
and U22284 (N_22284,N_20219,N_21917);
nor U22285 (N_22285,N_20544,N_20035);
and U22286 (N_22286,N_20694,N_20951);
nor U22287 (N_22287,N_21469,N_21082);
xor U22288 (N_22288,N_20053,N_21766);
nor U22289 (N_22289,N_21268,N_21694);
nand U22290 (N_22290,N_21428,N_20549);
xor U22291 (N_22291,N_21858,N_21645);
xor U22292 (N_22292,N_20226,N_20837);
xnor U22293 (N_22293,N_21138,N_20297);
and U22294 (N_22294,N_20653,N_20317);
nand U22295 (N_22295,N_20659,N_21127);
and U22296 (N_22296,N_21004,N_21176);
and U22297 (N_22297,N_20989,N_21996);
xnor U22298 (N_22298,N_21019,N_21509);
or U22299 (N_22299,N_21770,N_20614);
nand U22300 (N_22300,N_20723,N_20902);
and U22301 (N_22301,N_20362,N_20748);
or U22302 (N_22302,N_21429,N_20204);
nor U22303 (N_22303,N_20529,N_21866);
nand U22304 (N_22304,N_20161,N_20443);
nand U22305 (N_22305,N_21851,N_20371);
nand U22306 (N_22306,N_20056,N_20531);
xnor U22307 (N_22307,N_21479,N_20012);
nor U22308 (N_22308,N_21121,N_21736);
nand U22309 (N_22309,N_20301,N_20853);
or U22310 (N_22310,N_21891,N_21086);
nor U22311 (N_22311,N_20964,N_20859);
xor U22312 (N_22312,N_21409,N_20103);
nand U22313 (N_22313,N_21837,N_21391);
or U22314 (N_22314,N_20402,N_21060);
nor U22315 (N_22315,N_21683,N_20133);
and U22316 (N_22316,N_20511,N_21983);
or U22317 (N_22317,N_21473,N_21491);
and U22318 (N_22318,N_21017,N_20793);
or U22319 (N_22319,N_20232,N_21434);
nor U22320 (N_22320,N_21618,N_20435);
nand U22321 (N_22321,N_21126,N_20700);
and U22322 (N_22322,N_20230,N_20823);
nand U22323 (N_22323,N_20192,N_20311);
nor U22324 (N_22324,N_21831,N_21915);
xor U22325 (N_22325,N_20696,N_20548);
nand U22326 (N_22326,N_20794,N_21738);
and U22327 (N_22327,N_21803,N_21145);
and U22328 (N_22328,N_20915,N_21699);
and U22329 (N_22329,N_21532,N_20386);
xnor U22330 (N_22330,N_20212,N_20104);
or U22331 (N_22331,N_21548,N_21540);
or U22332 (N_22332,N_20065,N_20553);
nor U22333 (N_22333,N_21159,N_20432);
nor U22334 (N_22334,N_21744,N_21726);
nor U22335 (N_22335,N_21900,N_20569);
and U22336 (N_22336,N_21037,N_20919);
xnor U22337 (N_22337,N_21240,N_20954);
and U22338 (N_22338,N_20734,N_20298);
nor U22339 (N_22339,N_21551,N_21725);
and U22340 (N_22340,N_20022,N_20750);
xnor U22341 (N_22341,N_21748,N_20799);
and U22342 (N_22342,N_20512,N_21717);
nand U22343 (N_22343,N_20982,N_21821);
nor U22344 (N_22344,N_21403,N_21870);
and U22345 (N_22345,N_20594,N_21305);
xor U22346 (N_22346,N_21273,N_20867);
and U22347 (N_22347,N_20188,N_20599);
xnor U22348 (N_22348,N_20062,N_21448);
or U22349 (N_22349,N_20785,N_21599);
nand U22350 (N_22350,N_21067,N_20306);
xnor U22351 (N_22351,N_20510,N_20946);
nand U22352 (N_22352,N_20810,N_20547);
xor U22353 (N_22353,N_20735,N_21690);
xor U22354 (N_22354,N_21131,N_21672);
and U22355 (N_22355,N_20135,N_21410);
and U22356 (N_22356,N_21734,N_20487);
and U22357 (N_22357,N_20274,N_21130);
nor U22358 (N_22358,N_20261,N_20963);
and U22359 (N_22359,N_21643,N_20751);
or U22360 (N_22360,N_21485,N_21331);
xor U22361 (N_22361,N_20910,N_20596);
or U22362 (N_22362,N_20503,N_20777);
or U22363 (N_22363,N_21047,N_20147);
or U22364 (N_22364,N_20634,N_20168);
xor U22365 (N_22365,N_20873,N_20607);
and U22366 (N_22366,N_21912,N_21122);
and U22367 (N_22367,N_21764,N_20318);
nand U22368 (N_22368,N_20935,N_21077);
xor U22369 (N_22369,N_21795,N_20466);
or U22370 (N_22370,N_21046,N_21529);
or U22371 (N_22371,N_21733,N_21761);
nand U22372 (N_22372,N_20111,N_21459);
nand U22373 (N_22373,N_21790,N_20724);
xor U22374 (N_22374,N_20673,N_20268);
nor U22375 (N_22375,N_20453,N_21922);
or U22376 (N_22376,N_20139,N_21543);
or U22377 (N_22377,N_21199,N_20628);
nor U22378 (N_22378,N_21524,N_20149);
nand U22379 (N_22379,N_20154,N_20505);
and U22380 (N_22380,N_20431,N_20087);
nor U22381 (N_22381,N_21349,N_21100);
nor U22382 (N_22382,N_21177,N_20422);
or U22383 (N_22383,N_20639,N_21711);
nand U22384 (N_22384,N_20079,N_20841);
nor U22385 (N_22385,N_21976,N_20366);
nand U22386 (N_22386,N_20879,N_21029);
xor U22387 (N_22387,N_20184,N_21172);
or U22388 (N_22388,N_20521,N_20025);
nand U22389 (N_22389,N_20559,N_20224);
nor U22390 (N_22390,N_20348,N_20442);
nand U22391 (N_22391,N_20760,N_21943);
or U22392 (N_22392,N_21476,N_21567);
or U22393 (N_22393,N_20608,N_21844);
nor U22394 (N_22394,N_20664,N_21337);
nand U22395 (N_22395,N_20441,N_20181);
xnor U22396 (N_22396,N_21814,N_21493);
or U22397 (N_22397,N_20208,N_21973);
nor U22398 (N_22398,N_21073,N_20820);
nor U22399 (N_22399,N_21395,N_20998);
nor U22400 (N_22400,N_21419,N_21065);
xor U22401 (N_22401,N_20351,N_20651);
nor U22402 (N_22402,N_21010,N_20862);
nand U22403 (N_22403,N_21406,N_21150);
and U22404 (N_22404,N_20174,N_20292);
and U22405 (N_22405,N_21646,N_21638);
xnor U22406 (N_22406,N_20640,N_20164);
and U22407 (N_22407,N_20486,N_20762);
or U22408 (N_22408,N_21967,N_21778);
and U22409 (N_22409,N_20452,N_21327);
or U22410 (N_22410,N_21187,N_21519);
nand U22411 (N_22411,N_20832,N_20128);
or U22412 (N_22412,N_21938,N_20200);
and U22413 (N_22413,N_20500,N_20050);
nor U22414 (N_22414,N_20737,N_20061);
and U22415 (N_22415,N_20514,N_21512);
and U22416 (N_22416,N_20584,N_20738);
nor U22417 (N_22417,N_20315,N_20160);
and U22418 (N_22418,N_20156,N_20552);
nand U22419 (N_22419,N_20173,N_20266);
or U22420 (N_22420,N_21400,N_21020);
or U22421 (N_22421,N_21775,N_20627);
nand U22422 (N_22422,N_21097,N_21165);
xor U22423 (N_22423,N_20235,N_20275);
or U22424 (N_22424,N_20011,N_21282);
and U22425 (N_22425,N_21682,N_21204);
and U22426 (N_22426,N_21217,N_20522);
nor U22427 (N_22427,N_21052,N_20262);
nor U22428 (N_22428,N_21797,N_20293);
or U22429 (N_22429,N_21197,N_21801);
and U22430 (N_22430,N_20687,N_21261);
nor U22431 (N_22431,N_21650,N_20816);
nand U22432 (N_22432,N_20426,N_20804);
nand U22433 (N_22433,N_20716,N_20419);
xnor U22434 (N_22434,N_20397,N_20203);
and U22435 (N_22435,N_20331,N_20974);
or U22436 (N_22436,N_21074,N_21799);
and U22437 (N_22437,N_20622,N_20023);
nand U22438 (N_22438,N_20995,N_21291);
nand U22439 (N_22439,N_21713,N_21961);
and U22440 (N_22440,N_21460,N_20372);
nor U22441 (N_22441,N_21149,N_20499);
or U22442 (N_22442,N_20834,N_21987);
xnor U22443 (N_22443,N_20772,N_21511);
nand U22444 (N_22444,N_20256,N_20753);
and U22445 (N_22445,N_21558,N_20033);
and U22446 (N_22446,N_21045,N_21847);
or U22447 (N_22447,N_21171,N_21230);
and U22448 (N_22448,N_21334,N_20215);
nor U22449 (N_22449,N_21433,N_21220);
nor U22450 (N_22450,N_21151,N_21721);
xor U22451 (N_22451,N_20625,N_21857);
nand U22452 (N_22452,N_20685,N_21709);
nand U22453 (N_22453,N_20105,N_21440);
nor U22454 (N_22454,N_20024,N_20720);
xor U22455 (N_22455,N_21299,N_20630);
nand U22456 (N_22456,N_21103,N_21226);
nor U22457 (N_22457,N_20187,N_21144);
nand U22458 (N_22458,N_20684,N_20822);
nand U22459 (N_22459,N_21723,N_20106);
and U22460 (N_22460,N_21782,N_20165);
xor U22461 (N_22461,N_20296,N_21124);
nor U22462 (N_22462,N_20107,N_21246);
or U22463 (N_22463,N_20336,N_20907);
or U22464 (N_22464,N_20347,N_20690);
nand U22465 (N_22465,N_21904,N_20880);
nor U22466 (N_22466,N_20572,N_20534);
xnor U22467 (N_22467,N_21388,N_20796);
or U22468 (N_22468,N_21397,N_21688);
nand U22469 (N_22469,N_21063,N_20959);
or U22470 (N_22470,N_21028,N_20460);
or U22471 (N_22471,N_20313,N_21783);
and U22472 (N_22472,N_21773,N_21861);
nand U22473 (N_22473,N_20254,N_21032);
nand U22474 (N_22474,N_20117,N_21907);
xnor U22475 (N_22475,N_20600,N_21482);
and U22476 (N_22476,N_21185,N_20836);
xnor U22477 (N_22477,N_20756,N_21160);
and U22478 (N_22478,N_21878,N_20805);
nand U22479 (N_22479,N_20076,N_21439);
and U22480 (N_22480,N_21716,N_20654);
nor U22481 (N_22481,N_20387,N_20132);
and U22482 (N_22482,N_20239,N_21013);
xor U22483 (N_22483,N_21104,N_21960);
or U22484 (N_22484,N_20802,N_20742);
nor U22485 (N_22485,N_21025,N_21001);
xor U22486 (N_22486,N_20581,N_20363);
nor U22487 (N_22487,N_20307,N_20477);
or U22488 (N_22488,N_20365,N_21319);
nand U22489 (N_22489,N_21869,N_20167);
and U22490 (N_22490,N_20171,N_21295);
nor U22491 (N_22491,N_20471,N_20411);
or U22492 (N_22492,N_21344,N_21164);
nor U22493 (N_22493,N_21718,N_21322);
and U22494 (N_22494,N_20736,N_21146);
nor U22495 (N_22495,N_21281,N_20992);
nor U22496 (N_22496,N_20638,N_20434);
xor U22497 (N_22497,N_21968,N_21923);
nor U22498 (N_22498,N_21787,N_21040);
xnor U22499 (N_22499,N_21038,N_21027);
and U22500 (N_22500,N_20719,N_21602);
nor U22501 (N_22501,N_20469,N_20462);
xnor U22502 (N_22502,N_20143,N_20304);
xor U22503 (N_22503,N_20774,N_20579);
and U22504 (N_22504,N_21359,N_21875);
nand U22505 (N_22505,N_20710,N_20112);
or U22506 (N_22506,N_20333,N_20086);
xor U22507 (N_22507,N_21675,N_20643);
and U22508 (N_22508,N_20803,N_20485);
or U22509 (N_22509,N_21964,N_21213);
nand U22510 (N_22510,N_21583,N_21266);
xnor U22511 (N_22511,N_20842,N_20798);
xor U22512 (N_22512,N_21757,N_20764);
nor U22513 (N_22513,N_21954,N_20620);
and U22514 (N_22514,N_20039,N_20990);
xor U22515 (N_22515,N_21023,N_21415);
nand U22516 (N_22516,N_20642,N_20741);
and U22517 (N_22517,N_20978,N_21377);
and U22518 (N_22518,N_20976,N_21483);
and U22519 (N_22519,N_21712,N_20041);
nor U22520 (N_22520,N_20656,N_20813);
and U22521 (N_22521,N_20676,N_20631);
xnor U22522 (N_22522,N_21633,N_20182);
nor U22523 (N_22523,N_20644,N_20288);
and U22524 (N_22524,N_21198,N_20975);
nand U22525 (N_22525,N_20394,N_20812);
or U22526 (N_22526,N_21515,N_21914);
nor U22527 (N_22527,N_20714,N_20067);
or U22528 (N_22528,N_20205,N_21636);
or U22529 (N_22529,N_20932,N_20271);
xor U22530 (N_22530,N_20679,N_20973);
xnor U22531 (N_22531,N_20944,N_21815);
xor U22532 (N_22532,N_20513,N_21649);
and U22533 (N_22533,N_21902,N_20110);
nand U22534 (N_22534,N_21549,N_20036);
and U22535 (N_22535,N_21340,N_21536);
and U22536 (N_22536,N_21527,N_20623);
nor U22537 (N_22537,N_21609,N_20537);
nor U22538 (N_22538,N_21243,N_20413);
xor U22539 (N_22539,N_21078,N_21051);
and U22540 (N_22540,N_21059,N_21796);
xor U22541 (N_22541,N_21375,N_20377);
xor U22542 (N_22542,N_20473,N_20328);
nor U22543 (N_22543,N_21053,N_20985);
nand U22544 (N_22544,N_21180,N_20883);
xnor U22545 (N_22545,N_21360,N_21999);
nor U22546 (N_22546,N_21788,N_20000);
xnor U22547 (N_22547,N_20905,N_21178);
nor U22548 (N_22548,N_20950,N_21357);
nand U22549 (N_22549,N_20179,N_21418);
xnor U22550 (N_22550,N_21061,N_20968);
xor U22551 (N_22551,N_21498,N_20415);
xnor U22552 (N_22552,N_20058,N_21935);
nor U22553 (N_22553,N_21776,N_20017);
and U22554 (N_22554,N_21436,N_21590);
xnor U22555 (N_22555,N_21022,N_21432);
nand U22556 (N_22556,N_20152,N_20090);
xor U22557 (N_22557,N_21560,N_20588);
xnor U22558 (N_22558,N_20444,N_20176);
and U22559 (N_22559,N_20287,N_21107);
nand U22560 (N_22560,N_21664,N_21648);
xor U22561 (N_22561,N_20185,N_20940);
and U22562 (N_22562,N_20610,N_21321);
nand U22563 (N_22563,N_20196,N_21137);
and U22564 (N_22564,N_20410,N_20417);
and U22565 (N_22565,N_21356,N_20609);
nand U22566 (N_22566,N_20884,N_20692);
nand U22567 (N_22567,N_21850,N_21070);
and U22568 (N_22568,N_20009,N_21033);
xnor U22569 (N_22569,N_20354,N_21157);
and U22570 (N_22570,N_20098,N_20124);
nor U22571 (N_22571,N_21779,N_20647);
xor U22572 (N_22572,N_21896,N_21637);
xnor U22573 (N_22573,N_20277,N_20795);
nor U22574 (N_22574,N_21817,N_20766);
nor U22575 (N_22575,N_21903,N_20031);
xnor U22576 (N_22576,N_21401,N_21297);
xnor U22577 (N_22577,N_20146,N_21480);
nor U22578 (N_22578,N_21301,N_20340);
or U22579 (N_22579,N_21188,N_21154);
or U22580 (N_22580,N_21600,N_21420);
and U22581 (N_22581,N_21811,N_21962);
or U22582 (N_22582,N_21253,N_21979);
xnor U22583 (N_22583,N_21545,N_21865);
or U22584 (N_22584,N_21015,N_20279);
nand U22585 (N_22585,N_21011,N_20972);
and U22586 (N_22586,N_20784,N_20515);
nand U22587 (N_22587,N_21115,N_20960);
xor U22588 (N_22588,N_21833,N_20158);
nor U22589 (N_22589,N_21285,N_21978);
xor U22590 (N_22590,N_21186,N_20632);
or U22591 (N_22591,N_20746,N_20057);
xnor U22592 (N_22592,N_20264,N_20852);
nor U22593 (N_22593,N_21394,N_20782);
or U22594 (N_22594,N_20562,N_20855);
nand U22595 (N_22595,N_20808,N_21816);
or U22596 (N_22596,N_20680,N_21679);
and U22597 (N_22597,N_21095,N_21561);
nor U22598 (N_22598,N_21474,N_20223);
xor U22599 (N_22599,N_21451,N_20051);
or U22600 (N_22600,N_20045,N_21655);
xnor U22601 (N_22601,N_20032,N_21490);
or U22602 (N_22602,N_21813,N_20178);
xnor U22603 (N_22603,N_21885,N_21332);
nand U22604 (N_22604,N_20865,N_21676);
nand U22605 (N_22605,N_20074,N_21202);
and U22606 (N_22606,N_20211,N_21933);
nor U22607 (N_22607,N_21862,N_21805);
xnor U22608 (N_22608,N_20400,N_21014);
and U22609 (N_22609,N_20555,N_20273);
nor U22610 (N_22610,N_20851,N_20745);
nand U22611 (N_22611,N_21774,N_21849);
nand U22612 (N_22612,N_21245,N_20483);
nor U22613 (N_22613,N_20191,N_20999);
nand U22614 (N_22614,N_20412,N_21620);
nand U22615 (N_22615,N_21000,N_21864);
or U22616 (N_22616,N_21106,N_21800);
nand U22617 (N_22617,N_21229,N_21342);
or U22618 (N_22618,N_20114,N_21048);
and U22619 (N_22619,N_21581,N_21911);
xnor U22620 (N_22620,N_21564,N_20282);
nor U22621 (N_22621,N_20476,N_20436);
nand U22622 (N_22622,N_20170,N_21392);
and U22623 (N_22623,N_21841,N_21631);
or U22624 (N_22624,N_20675,N_21556);
xor U22625 (N_22625,N_21307,N_20492);
nor U22626 (N_22626,N_20574,N_21312);
nand U22627 (N_22627,N_21196,N_20520);
nand U22628 (N_22628,N_20020,N_21393);
and U22629 (N_22629,N_21132,N_21704);
or U22630 (N_22630,N_21373,N_20563);
and U22631 (N_22631,N_20717,N_21538);
nor U22632 (N_22632,N_20450,N_20882);
and U22633 (N_22633,N_20457,N_20353);
nor U22634 (N_22634,N_21222,N_21147);
xor U22635 (N_22635,N_20153,N_21874);
xnor U22636 (N_22636,N_21597,N_21913);
or U22637 (N_22637,N_20126,N_20368);
xnor U22638 (N_22638,N_21167,N_20094);
nor U22639 (N_22639,N_20332,N_21856);
nor U22640 (N_22640,N_21088,N_21463);
xnor U22641 (N_22641,N_20447,N_21398);
nor U22642 (N_22642,N_21657,N_20931);
and U22643 (N_22643,N_20439,N_20150);
xor U22644 (N_22644,N_21135,N_21087);
nand U22645 (N_22645,N_21877,N_20408);
nand U22646 (N_22646,N_21328,N_21965);
or U22647 (N_22647,N_21698,N_20939);
and U22648 (N_22648,N_21071,N_20845);
and U22649 (N_22649,N_20385,N_20858);
nor U22650 (N_22650,N_20624,N_21258);
and U22651 (N_22651,N_21640,N_21612);
xor U22652 (N_22652,N_20889,N_20083);
or U22653 (N_22653,N_20046,N_20148);
or U22654 (N_22654,N_20370,N_20201);
or U22655 (N_22655,N_21929,N_21068);
and U22656 (N_22656,N_21607,N_21030);
or U22657 (N_22657,N_21619,N_21089);
nor U22658 (N_22658,N_20030,N_20382);
nor U22659 (N_22659,N_20142,N_20626);
nor U22660 (N_22660,N_20860,N_21963);
and U22661 (N_22661,N_21867,N_21621);
and U22662 (N_22662,N_20015,N_21407);
or U22663 (N_22663,N_21887,N_20130);
nor U22664 (N_22664,N_21617,N_20502);
nand U22665 (N_22665,N_20281,N_20357);
nor U22666 (N_22666,N_20344,N_20885);
nand U22667 (N_22667,N_21075,N_20038);
or U22668 (N_22668,N_20590,N_21232);
and U22669 (N_22669,N_21256,N_20551);
xnor U22670 (N_22670,N_20478,N_20418);
xor U22671 (N_22671,N_20229,N_20582);
xor U22672 (N_22672,N_21839,N_21882);
nand U22673 (N_22673,N_21587,N_21513);
or U22674 (N_22674,N_20835,N_21193);
and U22675 (N_22675,N_20550,N_21055);
xnor U22676 (N_22676,N_21414,N_21823);
xor U22677 (N_22677,N_21141,N_21853);
or U22678 (N_22678,N_20993,N_20055);
and U22679 (N_22679,N_20652,N_21829);
nand U22680 (N_22680,N_21695,N_20814);
or U22681 (N_22681,N_20994,N_20504);
or U22682 (N_22682,N_21588,N_20977);
xor U22683 (N_22683,N_21324,N_21016);
or U22684 (N_22684,N_20324,N_21278);
nor U22685 (N_22685,N_20373,N_21466);
nor U22686 (N_22686,N_20645,N_21054);
and U22687 (N_22687,N_21554,N_20027);
xor U22688 (N_22688,N_21228,N_21936);
or U22689 (N_22689,N_20089,N_20364);
or U22690 (N_22690,N_20388,N_20343);
and U22691 (N_22691,N_20096,N_21980);
nor U22692 (N_22692,N_21845,N_20044);
nand U22693 (N_22693,N_20578,N_20021);
xor U22694 (N_22694,N_21502,N_20217);
or U22695 (N_22695,N_21399,N_21606);
xnor U22696 (N_22696,N_21363,N_20818);
xor U22697 (N_22697,N_21510,N_21625);
nand U22698 (N_22698,N_21091,N_21007);
and U22699 (N_22699,N_20898,N_20933);
xor U22700 (N_22700,N_20577,N_20064);
or U22701 (N_22701,N_21486,N_21830);
nand U22702 (N_22702,N_21449,N_20244);
and U22703 (N_22703,N_20943,N_20339);
xor U22704 (N_22704,N_20286,N_20440);
and U22705 (N_22705,N_21710,N_21552);
xnor U22706 (N_22706,N_20116,N_20570);
nor U22707 (N_22707,N_21208,N_20066);
nor U22708 (N_22708,N_20612,N_21096);
nor U22709 (N_22709,N_20792,N_20918);
nand U22710 (N_22710,N_20660,N_21868);
nor U22711 (N_22711,N_20285,N_21218);
and U22712 (N_22712,N_20425,N_20839);
or U22713 (N_22713,N_21494,N_20938);
or U22714 (N_22714,N_20303,N_21739);
and U22715 (N_22715,N_20329,N_21944);
or U22716 (N_22716,N_21860,N_21298);
and U22717 (N_22717,N_21991,N_20290);
nand U22718 (N_22718,N_21366,N_20019);
nor U22719 (N_22719,N_21155,N_20403);
or U22720 (N_22720,N_21686,N_20131);
nand U22721 (N_22721,N_20606,N_21677);
nor U22722 (N_22722,N_21624,N_20190);
xnor U22723 (N_22723,N_21162,N_21732);
nor U22724 (N_22724,N_21517,N_20059);
nand U22725 (N_22725,N_21118,N_21255);
nand U22726 (N_22726,N_20338,N_20769);
nand U22727 (N_22727,N_21881,N_21975);
and U22728 (N_22728,N_20247,N_20120);
xnor U22729 (N_22729,N_20824,N_21316);
nand U22730 (N_22730,N_21205,N_20669);
and U22731 (N_22731,N_20758,N_20849);
and U22732 (N_22732,N_20248,N_20672);
xnor U22733 (N_22733,N_21674,N_20284);
xnor U22734 (N_22734,N_21381,N_20308);
or U22735 (N_22735,N_20291,N_20833);
nor U22736 (N_22736,N_21928,N_20320);
xor U22737 (N_22737,N_20240,N_20546);
nand U22738 (N_22738,N_21338,N_20615);
or U22739 (N_22739,N_20595,N_20069);
nand U22740 (N_22740,N_20040,N_21190);
nand U22741 (N_22741,N_21216,N_20586);
or U22742 (N_22742,N_20875,N_21041);
and U22743 (N_22743,N_21632,N_20183);
nand U22744 (N_22744,N_21489,N_20490);
and U22745 (N_22745,N_20125,N_21952);
nor U22746 (N_22746,N_20962,N_21478);
and U22747 (N_22747,N_20864,N_21424);
nand U22748 (N_22748,N_20396,N_20399);
xnor U22749 (N_22749,N_20054,N_21825);
nor U22750 (N_22750,N_20678,N_20602);
xnor U22751 (N_22751,N_21542,N_20118);
xor U22752 (N_22752,N_21828,N_20300);
nor U22753 (N_22753,N_20821,N_21802);
or U22754 (N_22754,N_21031,N_20806);
or U22755 (N_22755,N_21148,N_20621);
nand U22756 (N_22756,N_21988,N_20334);
nor U22757 (N_22757,N_21345,N_20108);
or U22758 (N_22758,N_21950,N_21819);
nand U22759 (N_22759,N_20953,N_20636);
or U22760 (N_22760,N_20289,N_21893);
and U22761 (N_22761,N_21932,N_20007);
nand U22762 (N_22762,N_20604,N_21336);
and U22763 (N_22763,N_20468,N_20018);
xor U22764 (N_22764,N_20601,N_21251);
or U22765 (N_22765,N_20269,N_21333);
xnor U22766 (N_22766,N_21069,N_21347);
or U22767 (N_22767,N_20791,N_20538);
and U22768 (N_22768,N_20591,N_21629);
or U22769 (N_22769,N_21413,N_21354);
nand U22770 (N_22770,N_20718,N_20942);
nor U22771 (N_22771,N_20540,N_21533);
nand U22772 (N_22772,N_21383,N_20265);
and U22773 (N_22773,N_20662,N_21706);
or U22774 (N_22774,N_20075,N_21876);
or U22775 (N_22775,N_21673,N_20429);
nand U22776 (N_22776,N_21227,N_20255);
nand U22777 (N_22777,N_21528,N_21520);
or U22778 (N_22778,N_20603,N_20817);
nand U22779 (N_22779,N_21762,N_20668);
xor U22780 (N_22780,N_21671,N_21237);
nor U22781 (N_22781,N_21937,N_21039);
nand U22782 (N_22782,N_21313,N_21351);
xor U22783 (N_22783,N_20136,N_20727);
xnor U22784 (N_22784,N_21231,N_21660);
and U22785 (N_22785,N_21894,N_21722);
nor U22786 (N_22786,N_21254,N_20260);
nand U22787 (N_22787,N_20754,N_20404);
nor U22788 (N_22788,N_21557,N_21806);
or U22789 (N_22789,N_20568,N_21447);
nand U22790 (N_22790,N_20580,N_21211);
nand U22791 (N_22791,N_21209,N_21207);
nand U22792 (N_22792,N_21572,N_21417);
or U22793 (N_22793,N_21304,N_20661);
nand U22794 (N_22794,N_21457,N_21358);
xor U22795 (N_22795,N_20220,N_21248);
or U22796 (N_22796,N_20481,N_20682);
or U22797 (N_22797,N_21662,N_21445);
nand U22798 (N_22798,N_21569,N_21438);
nor U22799 (N_22799,N_21079,N_20218);
or U22800 (N_22800,N_21219,N_21504);
and U22801 (N_22801,N_21200,N_20144);
xor U22802 (N_22802,N_21234,N_21435);
nand U22803 (N_22803,N_20699,N_20052);
or U22804 (N_22804,N_21531,N_21942);
nor U22805 (N_22805,N_20869,N_21378);
nand U22806 (N_22806,N_21598,N_20861);
and U22807 (N_22807,N_21859,N_20743);
nand U22808 (N_22808,N_21080,N_21003);
nor U22809 (N_22809,N_21769,N_20761);
or U22810 (N_22810,N_21918,N_20472);
nand U22811 (N_22811,N_20194,N_20484);
nor U22812 (N_22812,N_20159,N_20010);
nand U22813 (N_22813,N_20101,N_21260);
nand U22814 (N_22814,N_20667,N_20991);
or U22815 (N_22815,N_21136,N_21034);
and U22816 (N_22816,N_20749,N_20526);
nor U22817 (N_22817,N_21262,N_21550);
nor U22818 (N_22818,N_20464,N_21302);
nor U22819 (N_22819,N_21364,N_20583);
nor U22820 (N_22820,N_20827,N_21235);
xor U22821 (N_22821,N_21446,N_20138);
nand U22822 (N_22822,N_20463,N_21974);
nand U22823 (N_22823,N_21701,N_20093);
nand U22824 (N_22824,N_21982,N_21212);
and U22825 (N_22825,N_20913,N_21777);
and U22826 (N_22826,N_20666,N_20243);
xnor U22827 (N_22827,N_21756,N_21910);
xnor U22828 (N_22828,N_21012,N_20920);
and U22829 (N_22829,N_21522,N_20113);
nand U22830 (N_22830,N_20788,N_21123);
nor U22831 (N_22831,N_21380,N_20517);
or U22832 (N_22832,N_20359,N_20454);
xnor U22833 (N_22833,N_21092,N_21939);
nand U22834 (N_22834,N_21320,N_20406);
nand U22835 (N_22835,N_21456,N_20530);
nor U22836 (N_22836,N_20532,N_20310);
xor U22837 (N_22837,N_21534,N_21348);
xor U22838 (N_22838,N_21559,N_20496);
or U22839 (N_22839,N_21310,N_21026);
nor U22840 (N_22840,N_20037,N_20263);
nand U22841 (N_22841,N_20016,N_20987);
and U22842 (N_22842,N_20077,N_21326);
nand U22843 (N_22843,N_20421,N_21812);
nand U22844 (N_22844,N_20649,N_21252);
nand U22845 (N_22845,N_20063,N_20084);
and U22846 (N_22846,N_20787,N_21899);
and U22847 (N_22847,N_20670,N_20175);
and U22848 (N_22848,N_21422,N_20071);
nor U22849 (N_22849,N_20342,N_20407);
and U22850 (N_22850,N_21516,N_20744);
or U22851 (N_22851,N_20361,N_20479);
or U22852 (N_22852,N_21442,N_20480);
xnor U22853 (N_22853,N_20937,N_20888);
nor U22854 (N_22854,N_21421,N_20209);
xor U22855 (N_22855,N_20947,N_20597);
and U22856 (N_22856,N_20405,N_20283);
xor U22857 (N_22857,N_20863,N_21105);
or U22858 (N_22858,N_21767,N_21927);
or U22859 (N_22859,N_20195,N_21749);
xnor U22860 (N_22860,N_21703,N_21705);
or U22861 (N_22861,N_20533,N_21571);
and U22862 (N_22862,N_21768,N_21287);
nand U22863 (N_22863,N_20233,N_20800);
nand U22864 (N_22864,N_20961,N_20997);
or U22865 (N_22865,N_20956,N_21958);
nand U22866 (N_22866,N_20843,N_20475);
or U22867 (N_22867,N_21441,N_20900);
and U22868 (N_22868,N_20509,N_20249);
nand U22869 (N_22869,N_21376,N_20783);
or U22870 (N_22870,N_21846,N_20322);
xor U22871 (N_22871,N_20409,N_21759);
and U22872 (N_22872,N_20252,N_20759);
and U22873 (N_22873,N_21696,N_20928);
nand U22874 (N_22874,N_21084,N_20258);
nor U22875 (N_22875,N_21593,N_20085);
or U22876 (N_22876,N_21133,N_21670);
or U22877 (N_22877,N_20896,N_21224);
xnor U22878 (N_22878,N_21544,N_20967);
or U22879 (N_22879,N_21341,N_20658);
and U22880 (N_22880,N_21579,N_21134);
xor U22881 (N_22881,N_21966,N_20383);
nand U22882 (N_22882,N_20379,N_21049);
or U22883 (N_22883,N_21719,N_20904);
and U22884 (N_22884,N_21745,N_20189);
or U22885 (N_22885,N_21408,N_21905);
nand U22886 (N_22886,N_20732,N_20210);
nand U22887 (N_22887,N_20912,N_21785);
and U22888 (N_22888,N_20272,N_21450);
xnor U22889 (N_22889,N_20047,N_20367);
nor U22890 (N_22890,N_20949,N_20323);
and U22891 (N_22891,N_21758,N_21125);
and U22892 (N_22892,N_20708,N_21919);
or U22893 (N_22893,N_21714,N_20350);
and U22894 (N_22894,N_21286,N_21323);
xnor U22895 (N_22895,N_20497,N_21577);
xor U22896 (N_22896,N_21692,N_20227);
nand U22897 (N_22897,N_20355,N_21500);
or U22898 (N_22898,N_20048,N_20465);
xnor U22899 (N_22899,N_20013,N_20541);
nor U22900 (N_22900,N_21595,N_20543);
or U22901 (N_22901,N_21389,N_20629);
nor U22902 (N_22902,N_21035,N_20445);
or U22903 (N_22903,N_21848,N_21946);
xor U22904 (N_22904,N_20231,N_20437);
xnor U22905 (N_22905,N_20127,N_20523);
and U22906 (N_22906,N_21101,N_20169);
nor U22907 (N_22907,N_21346,N_20778);
xnor U22908 (N_22908,N_20979,N_21879);
nand U22909 (N_22909,N_20618,N_20102);
nand U22910 (N_22910,N_21743,N_21239);
xor U22911 (N_22911,N_20280,N_21315);
xor U22912 (N_22912,N_21916,N_21654);
xor U22913 (N_22913,N_21058,N_21687);
nand U22914 (N_22914,N_20389,N_21259);
and U22915 (N_22915,N_20186,N_21613);
or U22916 (N_22916,N_20955,N_21423);
and U22917 (N_22917,N_21292,N_21152);
or U22918 (N_22918,N_20294,N_20137);
and U22919 (N_22919,N_21804,N_20049);
or U22920 (N_22920,N_21036,N_20726);
or U22921 (N_22921,N_20683,N_21742);
xor U22922 (N_22922,N_20752,N_20335);
xor U22923 (N_22923,N_20349,N_21535);
nor U22924 (N_22924,N_21627,N_21272);
and U22925 (N_22925,N_21505,N_20655);
nand U22926 (N_22926,N_20341,N_20899);
or U22927 (N_22927,N_21129,N_20251);
nand U22928 (N_22928,N_21546,N_21335);
nor U22929 (N_22929,N_20957,N_20467);
nor U22930 (N_22930,N_20295,N_21610);
xnor U22931 (N_22931,N_20073,N_21667);
and U22932 (N_22932,N_20693,N_21238);
xnor U22933 (N_22933,N_21998,N_21977);
and U22934 (N_22934,N_21484,N_20326);
or U22935 (N_22935,N_20527,N_20374);
xnor U22936 (N_22936,N_20706,N_21563);
xnor U22937 (N_22937,N_21589,N_21584);
nand U22938 (N_22938,N_21574,N_21179);
xnor U22939 (N_22939,N_20807,N_20831);
or U22940 (N_22940,N_21350,N_21555);
and U22941 (N_22941,N_21477,N_20826);
nor U22942 (N_22942,N_20401,N_21402);
or U22943 (N_22943,N_20952,N_21277);
xnor U22944 (N_22944,N_21568,N_21168);
nor U22945 (N_22945,N_21427,N_21753);
or U22946 (N_22946,N_21300,N_21901);
and U22947 (N_22947,N_20556,N_21064);
or U22948 (N_22948,N_20641,N_20965);
nor U22949 (N_22949,N_20566,N_21807);
or U22950 (N_22950,N_21863,N_20564);
xnor U22951 (N_22951,N_20423,N_20078);
xor U22952 (N_22952,N_21752,N_21265);
or U22953 (N_22953,N_20592,N_20345);
nand U22954 (N_22954,N_21369,N_20352);
or U22955 (N_22955,N_20100,N_21242);
or U22956 (N_22956,N_21727,N_21822);
xnor U22957 (N_22957,N_21953,N_21809);
xor U22958 (N_22958,N_20909,N_20893);
or U22959 (N_22959,N_20768,N_21601);
xor U22960 (N_22960,N_21140,N_21909);
or U22961 (N_22961,N_21525,N_21578);
nor U22962 (N_22962,N_21308,N_21443);
or U22963 (N_22963,N_20703,N_20755);
nor U22964 (N_22964,N_21365,N_21656);
nand U22965 (N_22965,N_21763,N_21948);
xnor U22966 (N_22966,N_20721,N_21387);
xor U22967 (N_22967,N_21139,N_21970);
or U22968 (N_22968,N_21780,N_21957);
or U22969 (N_22969,N_20008,N_21090);
nand U22970 (N_22970,N_21411,N_20878);
nand U22971 (N_22971,N_21006,N_21396);
xor U22972 (N_22972,N_20848,N_21997);
nor U22973 (N_22973,N_21808,N_20966);
xnor U22974 (N_22974,N_20391,N_20637);
or U22975 (N_22975,N_21370,N_21873);
nand U22976 (N_22976,N_21487,N_21203);
and U22977 (N_22977,N_21827,N_20539);
nor U22978 (N_22978,N_21658,N_20257);
or U22979 (N_22979,N_20781,N_21072);
and U22980 (N_22980,N_20542,N_20163);
nand U22981 (N_22981,N_20829,N_21586);
xnor U22982 (N_22982,N_21009,N_21666);
nand U22983 (N_22983,N_20587,N_20903);
or U22984 (N_22984,N_21385,N_21241);
nand U22985 (N_22985,N_21521,N_20390);
and U22986 (N_22986,N_20221,N_20786);
nor U22987 (N_22987,N_21771,N_21623);
xnor U22988 (N_22988,N_20887,N_21042);
nor U22989 (N_22989,N_21454,N_21794);
nor U22990 (N_22990,N_21201,N_21276);
nor U22991 (N_22991,N_21128,N_20380);
nor U22992 (N_22992,N_20598,N_20507);
nand U22993 (N_22993,N_21855,N_21472);
and U22994 (N_22994,N_21972,N_20449);
xnor U22995 (N_22995,N_21663,N_21523);
or U22996 (N_22996,N_20430,N_20042);
nor U22997 (N_22997,N_20970,N_20245);
xnor U22998 (N_22998,N_21475,N_21143);
xor U22999 (N_22999,N_20488,N_20458);
and U23000 (N_23000,N_20095,N_20270);
xnor U23001 (N_23001,N_20605,N_20760);
and U23002 (N_23002,N_20770,N_21687);
nand U23003 (N_23003,N_20374,N_21822);
and U23004 (N_23004,N_21058,N_21509);
or U23005 (N_23005,N_21851,N_21301);
nor U23006 (N_23006,N_20632,N_20438);
and U23007 (N_23007,N_20761,N_21435);
nand U23008 (N_23008,N_21953,N_21900);
or U23009 (N_23009,N_20063,N_20531);
nand U23010 (N_23010,N_21515,N_21832);
and U23011 (N_23011,N_20167,N_20483);
and U23012 (N_23012,N_21050,N_21616);
xnor U23013 (N_23013,N_20899,N_20905);
nor U23014 (N_23014,N_21091,N_20811);
or U23015 (N_23015,N_21839,N_21037);
or U23016 (N_23016,N_20644,N_21430);
xor U23017 (N_23017,N_21575,N_21870);
or U23018 (N_23018,N_21141,N_20828);
nand U23019 (N_23019,N_21266,N_21221);
and U23020 (N_23020,N_21863,N_20633);
nor U23021 (N_23021,N_21348,N_21133);
nor U23022 (N_23022,N_21326,N_20211);
nand U23023 (N_23023,N_20836,N_20766);
nand U23024 (N_23024,N_20537,N_21666);
xnor U23025 (N_23025,N_20977,N_21194);
xnor U23026 (N_23026,N_21097,N_21089);
nand U23027 (N_23027,N_20772,N_21495);
or U23028 (N_23028,N_20253,N_21039);
or U23029 (N_23029,N_20761,N_20656);
or U23030 (N_23030,N_20711,N_21379);
and U23031 (N_23031,N_21906,N_20029);
and U23032 (N_23032,N_20833,N_20237);
or U23033 (N_23033,N_20945,N_21091);
xnor U23034 (N_23034,N_21476,N_21232);
xor U23035 (N_23035,N_20626,N_21498);
or U23036 (N_23036,N_21096,N_21607);
and U23037 (N_23037,N_21261,N_20871);
or U23038 (N_23038,N_21936,N_21824);
nand U23039 (N_23039,N_21343,N_20416);
nor U23040 (N_23040,N_21272,N_21815);
or U23041 (N_23041,N_21155,N_20829);
xor U23042 (N_23042,N_20280,N_20387);
nor U23043 (N_23043,N_21280,N_20746);
xnor U23044 (N_23044,N_21971,N_20579);
nor U23045 (N_23045,N_21765,N_20840);
xor U23046 (N_23046,N_21235,N_21855);
xor U23047 (N_23047,N_20777,N_21148);
nor U23048 (N_23048,N_21451,N_21725);
xnor U23049 (N_23049,N_21553,N_20921);
xnor U23050 (N_23050,N_21839,N_20086);
xnor U23051 (N_23051,N_20323,N_21029);
or U23052 (N_23052,N_20574,N_20867);
nor U23053 (N_23053,N_21050,N_21047);
nand U23054 (N_23054,N_20417,N_21316);
nor U23055 (N_23055,N_20619,N_20300);
nor U23056 (N_23056,N_20726,N_21873);
nor U23057 (N_23057,N_20609,N_20409);
nand U23058 (N_23058,N_20028,N_21804);
and U23059 (N_23059,N_20820,N_20025);
or U23060 (N_23060,N_21234,N_20946);
nand U23061 (N_23061,N_21211,N_21101);
nor U23062 (N_23062,N_20585,N_21309);
nor U23063 (N_23063,N_20591,N_21484);
xor U23064 (N_23064,N_20342,N_21835);
and U23065 (N_23065,N_20286,N_20802);
xnor U23066 (N_23066,N_21965,N_21725);
or U23067 (N_23067,N_21023,N_21802);
or U23068 (N_23068,N_21736,N_20665);
xor U23069 (N_23069,N_20144,N_20523);
nor U23070 (N_23070,N_20382,N_20333);
and U23071 (N_23071,N_21356,N_20867);
nand U23072 (N_23072,N_21570,N_21511);
and U23073 (N_23073,N_20197,N_21441);
or U23074 (N_23074,N_20147,N_20289);
nor U23075 (N_23075,N_21339,N_21262);
nor U23076 (N_23076,N_21299,N_20957);
xor U23077 (N_23077,N_21419,N_21747);
or U23078 (N_23078,N_21068,N_21556);
nand U23079 (N_23079,N_20373,N_20076);
and U23080 (N_23080,N_21044,N_20640);
nand U23081 (N_23081,N_20788,N_20332);
nand U23082 (N_23082,N_21347,N_21601);
and U23083 (N_23083,N_20867,N_20722);
xor U23084 (N_23084,N_20276,N_20295);
or U23085 (N_23085,N_21243,N_21765);
or U23086 (N_23086,N_20200,N_21136);
nor U23087 (N_23087,N_20588,N_20642);
nand U23088 (N_23088,N_20125,N_20071);
nand U23089 (N_23089,N_20761,N_21934);
and U23090 (N_23090,N_21777,N_21940);
nor U23091 (N_23091,N_21639,N_21568);
or U23092 (N_23092,N_20482,N_20128);
nand U23093 (N_23093,N_20582,N_21884);
or U23094 (N_23094,N_21644,N_21194);
xor U23095 (N_23095,N_21708,N_20938);
nor U23096 (N_23096,N_20705,N_21988);
nand U23097 (N_23097,N_20796,N_20251);
nor U23098 (N_23098,N_21579,N_20712);
nor U23099 (N_23099,N_20358,N_21718);
and U23100 (N_23100,N_20679,N_20562);
xor U23101 (N_23101,N_20151,N_20026);
nor U23102 (N_23102,N_20714,N_21355);
nand U23103 (N_23103,N_20593,N_21360);
xnor U23104 (N_23104,N_20655,N_21334);
or U23105 (N_23105,N_21160,N_21041);
nand U23106 (N_23106,N_21559,N_20950);
nor U23107 (N_23107,N_20627,N_20238);
and U23108 (N_23108,N_20539,N_20395);
xor U23109 (N_23109,N_21242,N_21303);
and U23110 (N_23110,N_20424,N_21690);
or U23111 (N_23111,N_20921,N_20187);
and U23112 (N_23112,N_21052,N_20089);
xor U23113 (N_23113,N_20925,N_21189);
xnor U23114 (N_23114,N_21239,N_20432);
or U23115 (N_23115,N_20799,N_21801);
nand U23116 (N_23116,N_21591,N_21177);
nand U23117 (N_23117,N_20705,N_21542);
xnor U23118 (N_23118,N_21691,N_21921);
and U23119 (N_23119,N_21311,N_20694);
or U23120 (N_23120,N_20277,N_20838);
or U23121 (N_23121,N_20614,N_20106);
nand U23122 (N_23122,N_21213,N_20770);
nand U23123 (N_23123,N_21025,N_20704);
nor U23124 (N_23124,N_21097,N_20511);
xnor U23125 (N_23125,N_20041,N_21555);
nand U23126 (N_23126,N_21247,N_20588);
nand U23127 (N_23127,N_20835,N_21373);
or U23128 (N_23128,N_20108,N_21285);
xnor U23129 (N_23129,N_20581,N_21296);
and U23130 (N_23130,N_21804,N_21013);
nor U23131 (N_23131,N_20173,N_21762);
or U23132 (N_23132,N_20835,N_20819);
nor U23133 (N_23133,N_20187,N_20098);
xor U23134 (N_23134,N_20476,N_21923);
nand U23135 (N_23135,N_21469,N_20422);
xor U23136 (N_23136,N_20677,N_20373);
nand U23137 (N_23137,N_20221,N_20693);
nor U23138 (N_23138,N_20855,N_21173);
xnor U23139 (N_23139,N_21435,N_20224);
and U23140 (N_23140,N_20473,N_20500);
and U23141 (N_23141,N_21313,N_20513);
and U23142 (N_23142,N_21871,N_20684);
xor U23143 (N_23143,N_20835,N_21118);
nor U23144 (N_23144,N_20710,N_21294);
nand U23145 (N_23145,N_21471,N_21390);
and U23146 (N_23146,N_21935,N_21728);
xor U23147 (N_23147,N_21230,N_20023);
nor U23148 (N_23148,N_20054,N_21632);
or U23149 (N_23149,N_21243,N_21075);
xor U23150 (N_23150,N_20841,N_20353);
nand U23151 (N_23151,N_20643,N_20826);
nor U23152 (N_23152,N_21514,N_21702);
or U23153 (N_23153,N_21202,N_20244);
or U23154 (N_23154,N_20942,N_20874);
nand U23155 (N_23155,N_20018,N_21354);
xnor U23156 (N_23156,N_20303,N_20418);
xor U23157 (N_23157,N_21132,N_21744);
and U23158 (N_23158,N_20820,N_21599);
nand U23159 (N_23159,N_20516,N_21853);
xnor U23160 (N_23160,N_20468,N_20172);
or U23161 (N_23161,N_20244,N_20446);
xor U23162 (N_23162,N_21035,N_21087);
and U23163 (N_23163,N_21803,N_20729);
nand U23164 (N_23164,N_20388,N_21307);
nand U23165 (N_23165,N_21766,N_21037);
xor U23166 (N_23166,N_21849,N_21920);
xnor U23167 (N_23167,N_21345,N_21171);
xnor U23168 (N_23168,N_20991,N_20239);
or U23169 (N_23169,N_21169,N_20392);
xnor U23170 (N_23170,N_20595,N_20385);
and U23171 (N_23171,N_21354,N_21351);
nor U23172 (N_23172,N_20149,N_20819);
or U23173 (N_23173,N_21237,N_20263);
xnor U23174 (N_23174,N_20494,N_21779);
or U23175 (N_23175,N_21486,N_20074);
nand U23176 (N_23176,N_20220,N_21942);
or U23177 (N_23177,N_21151,N_20030);
nor U23178 (N_23178,N_21220,N_20595);
xor U23179 (N_23179,N_21203,N_21650);
nor U23180 (N_23180,N_20045,N_20619);
and U23181 (N_23181,N_21385,N_20067);
and U23182 (N_23182,N_20991,N_20010);
or U23183 (N_23183,N_21636,N_21712);
nand U23184 (N_23184,N_20041,N_21081);
xnor U23185 (N_23185,N_20094,N_20244);
and U23186 (N_23186,N_21864,N_21040);
xnor U23187 (N_23187,N_21940,N_21736);
or U23188 (N_23188,N_20360,N_20984);
nand U23189 (N_23189,N_20098,N_21542);
nor U23190 (N_23190,N_20375,N_20085);
nand U23191 (N_23191,N_20496,N_20803);
or U23192 (N_23192,N_21177,N_21048);
and U23193 (N_23193,N_21568,N_20735);
and U23194 (N_23194,N_21898,N_20216);
and U23195 (N_23195,N_21191,N_20521);
and U23196 (N_23196,N_21777,N_20379);
and U23197 (N_23197,N_20379,N_20641);
xnor U23198 (N_23198,N_21607,N_20163);
and U23199 (N_23199,N_21632,N_20045);
nor U23200 (N_23200,N_21916,N_20727);
xor U23201 (N_23201,N_21056,N_20851);
or U23202 (N_23202,N_20232,N_20617);
and U23203 (N_23203,N_20660,N_21692);
nand U23204 (N_23204,N_21556,N_21448);
and U23205 (N_23205,N_21885,N_20023);
or U23206 (N_23206,N_21961,N_20744);
nand U23207 (N_23207,N_20870,N_20455);
xnor U23208 (N_23208,N_20806,N_20918);
and U23209 (N_23209,N_20365,N_20634);
and U23210 (N_23210,N_21191,N_20241);
and U23211 (N_23211,N_21639,N_20827);
or U23212 (N_23212,N_21908,N_21277);
and U23213 (N_23213,N_20135,N_20790);
and U23214 (N_23214,N_21064,N_20785);
or U23215 (N_23215,N_21437,N_21947);
xor U23216 (N_23216,N_21210,N_20138);
nand U23217 (N_23217,N_20287,N_20317);
or U23218 (N_23218,N_21434,N_21465);
and U23219 (N_23219,N_21498,N_21635);
or U23220 (N_23220,N_20331,N_21297);
and U23221 (N_23221,N_20077,N_21259);
and U23222 (N_23222,N_20706,N_21735);
nor U23223 (N_23223,N_21674,N_21250);
and U23224 (N_23224,N_21598,N_21244);
and U23225 (N_23225,N_20359,N_21131);
or U23226 (N_23226,N_20531,N_20278);
or U23227 (N_23227,N_21190,N_21515);
or U23228 (N_23228,N_20961,N_21581);
or U23229 (N_23229,N_21719,N_20572);
nor U23230 (N_23230,N_20938,N_20236);
nand U23231 (N_23231,N_20646,N_21920);
nor U23232 (N_23232,N_20691,N_21820);
nor U23233 (N_23233,N_21670,N_20317);
nand U23234 (N_23234,N_20792,N_21842);
and U23235 (N_23235,N_20088,N_21020);
nand U23236 (N_23236,N_21181,N_21865);
nand U23237 (N_23237,N_21414,N_20399);
or U23238 (N_23238,N_20041,N_20424);
or U23239 (N_23239,N_21444,N_21075);
xor U23240 (N_23240,N_20807,N_21338);
or U23241 (N_23241,N_20426,N_20879);
and U23242 (N_23242,N_21292,N_21867);
or U23243 (N_23243,N_21349,N_21719);
xor U23244 (N_23244,N_20573,N_20126);
or U23245 (N_23245,N_20088,N_21101);
xnor U23246 (N_23246,N_20454,N_21856);
nor U23247 (N_23247,N_21272,N_21954);
nor U23248 (N_23248,N_21366,N_20210);
and U23249 (N_23249,N_20566,N_20866);
xor U23250 (N_23250,N_20839,N_20716);
or U23251 (N_23251,N_20073,N_21070);
and U23252 (N_23252,N_21056,N_21256);
nor U23253 (N_23253,N_20008,N_21397);
or U23254 (N_23254,N_20861,N_20405);
xor U23255 (N_23255,N_20193,N_21328);
xor U23256 (N_23256,N_21062,N_21264);
nand U23257 (N_23257,N_20904,N_20820);
nand U23258 (N_23258,N_20972,N_20420);
or U23259 (N_23259,N_20211,N_20602);
and U23260 (N_23260,N_20463,N_21810);
or U23261 (N_23261,N_20223,N_20687);
nor U23262 (N_23262,N_20352,N_21682);
nand U23263 (N_23263,N_21978,N_20291);
and U23264 (N_23264,N_21011,N_21015);
or U23265 (N_23265,N_20236,N_21535);
xor U23266 (N_23266,N_20757,N_20725);
nand U23267 (N_23267,N_21549,N_21476);
or U23268 (N_23268,N_21650,N_20937);
nand U23269 (N_23269,N_20952,N_21712);
nand U23270 (N_23270,N_20792,N_21972);
or U23271 (N_23271,N_21027,N_21101);
xnor U23272 (N_23272,N_20627,N_21918);
and U23273 (N_23273,N_21713,N_21247);
nor U23274 (N_23274,N_21608,N_20776);
nand U23275 (N_23275,N_21305,N_21490);
nor U23276 (N_23276,N_20341,N_20215);
nand U23277 (N_23277,N_21578,N_21821);
or U23278 (N_23278,N_20611,N_20757);
nor U23279 (N_23279,N_20411,N_21228);
nand U23280 (N_23280,N_21613,N_20210);
nor U23281 (N_23281,N_20578,N_20468);
and U23282 (N_23282,N_20159,N_21553);
nand U23283 (N_23283,N_21457,N_20649);
xnor U23284 (N_23284,N_21421,N_21469);
or U23285 (N_23285,N_21940,N_20415);
nand U23286 (N_23286,N_21551,N_21569);
or U23287 (N_23287,N_21279,N_20594);
or U23288 (N_23288,N_20745,N_21905);
or U23289 (N_23289,N_21363,N_21798);
nand U23290 (N_23290,N_20333,N_21277);
or U23291 (N_23291,N_20938,N_21761);
nor U23292 (N_23292,N_21605,N_20116);
xor U23293 (N_23293,N_21908,N_21051);
xnor U23294 (N_23294,N_21953,N_21815);
xor U23295 (N_23295,N_20364,N_20990);
or U23296 (N_23296,N_21826,N_21200);
xnor U23297 (N_23297,N_20757,N_21814);
xnor U23298 (N_23298,N_20129,N_20348);
nor U23299 (N_23299,N_21586,N_21603);
nor U23300 (N_23300,N_21843,N_20567);
xnor U23301 (N_23301,N_20590,N_21059);
and U23302 (N_23302,N_20608,N_21030);
nand U23303 (N_23303,N_21615,N_21550);
or U23304 (N_23304,N_21003,N_21393);
xor U23305 (N_23305,N_20088,N_21665);
or U23306 (N_23306,N_20281,N_20346);
nand U23307 (N_23307,N_21569,N_20798);
and U23308 (N_23308,N_20088,N_20529);
or U23309 (N_23309,N_20022,N_20997);
nor U23310 (N_23310,N_21688,N_21637);
or U23311 (N_23311,N_21137,N_21885);
and U23312 (N_23312,N_21447,N_20322);
nand U23313 (N_23313,N_21661,N_20050);
and U23314 (N_23314,N_20766,N_21368);
or U23315 (N_23315,N_21468,N_20408);
and U23316 (N_23316,N_21493,N_20165);
nor U23317 (N_23317,N_21319,N_21453);
and U23318 (N_23318,N_20103,N_21663);
nand U23319 (N_23319,N_20634,N_20522);
or U23320 (N_23320,N_20657,N_21213);
nand U23321 (N_23321,N_21239,N_20954);
and U23322 (N_23322,N_20518,N_21197);
or U23323 (N_23323,N_20225,N_21140);
nor U23324 (N_23324,N_21247,N_20963);
nand U23325 (N_23325,N_21128,N_21902);
and U23326 (N_23326,N_21741,N_20200);
nand U23327 (N_23327,N_20017,N_20106);
nor U23328 (N_23328,N_21738,N_21382);
nor U23329 (N_23329,N_21174,N_21247);
or U23330 (N_23330,N_20869,N_21320);
nor U23331 (N_23331,N_21825,N_21389);
or U23332 (N_23332,N_21410,N_20564);
or U23333 (N_23333,N_21964,N_20798);
nand U23334 (N_23334,N_21855,N_21625);
or U23335 (N_23335,N_21638,N_21418);
or U23336 (N_23336,N_21625,N_21085);
or U23337 (N_23337,N_21088,N_21709);
nor U23338 (N_23338,N_21324,N_21920);
nand U23339 (N_23339,N_21123,N_20528);
nor U23340 (N_23340,N_20635,N_20502);
or U23341 (N_23341,N_21541,N_20968);
and U23342 (N_23342,N_20119,N_20229);
and U23343 (N_23343,N_21418,N_21874);
xnor U23344 (N_23344,N_20272,N_21537);
and U23345 (N_23345,N_20947,N_21055);
nand U23346 (N_23346,N_20999,N_21311);
nand U23347 (N_23347,N_20384,N_21523);
xor U23348 (N_23348,N_21573,N_21477);
nor U23349 (N_23349,N_20519,N_20479);
nand U23350 (N_23350,N_21759,N_21819);
nor U23351 (N_23351,N_21559,N_20468);
nor U23352 (N_23352,N_20424,N_21770);
or U23353 (N_23353,N_20031,N_21390);
or U23354 (N_23354,N_20784,N_20738);
xnor U23355 (N_23355,N_20437,N_21985);
or U23356 (N_23356,N_20920,N_21811);
and U23357 (N_23357,N_21805,N_20571);
xor U23358 (N_23358,N_20061,N_21068);
xnor U23359 (N_23359,N_20753,N_21878);
xor U23360 (N_23360,N_21966,N_20648);
and U23361 (N_23361,N_21730,N_21508);
nor U23362 (N_23362,N_21579,N_21814);
and U23363 (N_23363,N_20136,N_20599);
nand U23364 (N_23364,N_21147,N_20514);
nor U23365 (N_23365,N_21195,N_21447);
nand U23366 (N_23366,N_20933,N_21084);
or U23367 (N_23367,N_20150,N_20255);
xor U23368 (N_23368,N_21861,N_20539);
nor U23369 (N_23369,N_20553,N_21944);
nor U23370 (N_23370,N_21470,N_20343);
xor U23371 (N_23371,N_21906,N_21023);
xnor U23372 (N_23372,N_21180,N_21766);
xnor U23373 (N_23373,N_20821,N_21135);
or U23374 (N_23374,N_21820,N_20382);
and U23375 (N_23375,N_21468,N_20343);
nor U23376 (N_23376,N_21713,N_20498);
xor U23377 (N_23377,N_20923,N_20409);
and U23378 (N_23378,N_21089,N_20211);
nand U23379 (N_23379,N_21643,N_21456);
nand U23380 (N_23380,N_20214,N_21785);
or U23381 (N_23381,N_21898,N_20650);
nor U23382 (N_23382,N_21090,N_21679);
and U23383 (N_23383,N_21168,N_20552);
xnor U23384 (N_23384,N_21151,N_20145);
and U23385 (N_23385,N_21144,N_20871);
or U23386 (N_23386,N_21474,N_20467);
and U23387 (N_23387,N_21737,N_21390);
nand U23388 (N_23388,N_20127,N_20398);
and U23389 (N_23389,N_20441,N_20074);
nand U23390 (N_23390,N_20422,N_21997);
or U23391 (N_23391,N_21661,N_20998);
xnor U23392 (N_23392,N_21259,N_20907);
or U23393 (N_23393,N_21753,N_20084);
nor U23394 (N_23394,N_21218,N_21035);
nor U23395 (N_23395,N_20201,N_21245);
nor U23396 (N_23396,N_20738,N_21688);
nand U23397 (N_23397,N_21897,N_21675);
or U23398 (N_23398,N_20821,N_21916);
nor U23399 (N_23399,N_21085,N_20962);
nand U23400 (N_23400,N_20401,N_21439);
nor U23401 (N_23401,N_20486,N_21677);
nand U23402 (N_23402,N_20703,N_20196);
or U23403 (N_23403,N_21872,N_20842);
and U23404 (N_23404,N_20875,N_21518);
xor U23405 (N_23405,N_20293,N_21933);
nand U23406 (N_23406,N_20809,N_21085);
nand U23407 (N_23407,N_21617,N_20309);
nor U23408 (N_23408,N_20889,N_20772);
or U23409 (N_23409,N_20512,N_21338);
xor U23410 (N_23410,N_21894,N_20329);
xnor U23411 (N_23411,N_20279,N_21688);
nand U23412 (N_23412,N_21445,N_20324);
and U23413 (N_23413,N_21473,N_20001);
xor U23414 (N_23414,N_21081,N_21328);
nand U23415 (N_23415,N_20303,N_21102);
nor U23416 (N_23416,N_21561,N_21499);
and U23417 (N_23417,N_21812,N_20491);
nor U23418 (N_23418,N_20862,N_21571);
and U23419 (N_23419,N_21846,N_20380);
or U23420 (N_23420,N_20303,N_21140);
and U23421 (N_23421,N_20186,N_21644);
nor U23422 (N_23422,N_20446,N_21817);
nor U23423 (N_23423,N_21266,N_20381);
nor U23424 (N_23424,N_21327,N_21361);
nor U23425 (N_23425,N_21049,N_21627);
xnor U23426 (N_23426,N_21246,N_21525);
or U23427 (N_23427,N_21914,N_20338);
and U23428 (N_23428,N_20551,N_21084);
and U23429 (N_23429,N_21915,N_21399);
and U23430 (N_23430,N_21006,N_21223);
nand U23431 (N_23431,N_21731,N_21911);
and U23432 (N_23432,N_21356,N_20670);
nand U23433 (N_23433,N_21785,N_21136);
nand U23434 (N_23434,N_21972,N_20263);
nor U23435 (N_23435,N_21485,N_21570);
and U23436 (N_23436,N_20923,N_20348);
or U23437 (N_23437,N_21590,N_21612);
xnor U23438 (N_23438,N_21379,N_20947);
or U23439 (N_23439,N_21260,N_20657);
nor U23440 (N_23440,N_20253,N_21283);
nand U23441 (N_23441,N_21628,N_21093);
nand U23442 (N_23442,N_21659,N_20579);
xnor U23443 (N_23443,N_21197,N_21051);
nand U23444 (N_23444,N_21625,N_20256);
or U23445 (N_23445,N_20523,N_20153);
xnor U23446 (N_23446,N_20195,N_21563);
xnor U23447 (N_23447,N_20196,N_21999);
xnor U23448 (N_23448,N_20171,N_21716);
and U23449 (N_23449,N_21230,N_20864);
nor U23450 (N_23450,N_20966,N_21887);
xnor U23451 (N_23451,N_21007,N_20863);
nor U23452 (N_23452,N_21079,N_21897);
xnor U23453 (N_23453,N_21479,N_20368);
xor U23454 (N_23454,N_20691,N_21472);
or U23455 (N_23455,N_21743,N_20789);
nand U23456 (N_23456,N_20017,N_20973);
nor U23457 (N_23457,N_21750,N_20544);
or U23458 (N_23458,N_20239,N_21143);
or U23459 (N_23459,N_21923,N_21915);
nand U23460 (N_23460,N_21062,N_20073);
or U23461 (N_23461,N_20915,N_21559);
or U23462 (N_23462,N_21117,N_21052);
nor U23463 (N_23463,N_21673,N_21352);
and U23464 (N_23464,N_20640,N_21377);
or U23465 (N_23465,N_21242,N_21647);
nor U23466 (N_23466,N_20684,N_21063);
or U23467 (N_23467,N_21319,N_21672);
nand U23468 (N_23468,N_20807,N_21167);
and U23469 (N_23469,N_20533,N_21918);
or U23470 (N_23470,N_21745,N_21425);
and U23471 (N_23471,N_20101,N_20663);
and U23472 (N_23472,N_20738,N_21693);
or U23473 (N_23473,N_21220,N_20229);
nor U23474 (N_23474,N_20978,N_20952);
nor U23475 (N_23475,N_21108,N_20896);
xor U23476 (N_23476,N_20164,N_20957);
and U23477 (N_23477,N_20411,N_21453);
nor U23478 (N_23478,N_21643,N_20640);
nand U23479 (N_23479,N_21413,N_20188);
nand U23480 (N_23480,N_20433,N_20038);
and U23481 (N_23481,N_20399,N_20799);
xor U23482 (N_23482,N_21478,N_21362);
nor U23483 (N_23483,N_20655,N_21527);
xor U23484 (N_23484,N_21277,N_21604);
nand U23485 (N_23485,N_20751,N_21186);
xnor U23486 (N_23486,N_21957,N_21613);
or U23487 (N_23487,N_20424,N_20352);
or U23488 (N_23488,N_21720,N_20234);
nand U23489 (N_23489,N_20185,N_20179);
and U23490 (N_23490,N_21591,N_21160);
and U23491 (N_23491,N_21185,N_21655);
nor U23492 (N_23492,N_21405,N_21575);
and U23493 (N_23493,N_20126,N_20305);
and U23494 (N_23494,N_20638,N_20507);
and U23495 (N_23495,N_20917,N_20566);
nand U23496 (N_23496,N_20007,N_21504);
or U23497 (N_23497,N_20565,N_21079);
or U23498 (N_23498,N_20479,N_20360);
or U23499 (N_23499,N_21920,N_21534);
nand U23500 (N_23500,N_21056,N_20145);
and U23501 (N_23501,N_21619,N_21667);
xor U23502 (N_23502,N_20751,N_20765);
nand U23503 (N_23503,N_20274,N_20343);
or U23504 (N_23504,N_20653,N_21039);
nor U23505 (N_23505,N_21401,N_20964);
nor U23506 (N_23506,N_21774,N_20807);
or U23507 (N_23507,N_21776,N_21742);
and U23508 (N_23508,N_21897,N_21527);
or U23509 (N_23509,N_21130,N_20670);
xor U23510 (N_23510,N_21057,N_21656);
nand U23511 (N_23511,N_21288,N_20372);
nor U23512 (N_23512,N_20712,N_21357);
nor U23513 (N_23513,N_20734,N_20056);
and U23514 (N_23514,N_21041,N_20623);
or U23515 (N_23515,N_20782,N_21973);
nor U23516 (N_23516,N_21000,N_20734);
or U23517 (N_23517,N_21347,N_21748);
nor U23518 (N_23518,N_21934,N_21854);
nand U23519 (N_23519,N_21151,N_20147);
nand U23520 (N_23520,N_20587,N_20985);
nand U23521 (N_23521,N_20485,N_21144);
and U23522 (N_23522,N_21440,N_20562);
nor U23523 (N_23523,N_21620,N_20622);
nor U23524 (N_23524,N_20890,N_21435);
nor U23525 (N_23525,N_21075,N_21858);
nand U23526 (N_23526,N_20489,N_20267);
nand U23527 (N_23527,N_20852,N_21219);
or U23528 (N_23528,N_20958,N_20158);
xor U23529 (N_23529,N_20145,N_21116);
or U23530 (N_23530,N_21097,N_21666);
and U23531 (N_23531,N_21317,N_20635);
xnor U23532 (N_23532,N_21501,N_21810);
xor U23533 (N_23533,N_21549,N_20914);
xor U23534 (N_23534,N_20761,N_21750);
or U23535 (N_23535,N_21332,N_20588);
nand U23536 (N_23536,N_20961,N_20676);
nor U23537 (N_23537,N_20935,N_20968);
nand U23538 (N_23538,N_21957,N_20495);
or U23539 (N_23539,N_21513,N_21859);
xnor U23540 (N_23540,N_21223,N_20283);
nor U23541 (N_23541,N_20107,N_21845);
nor U23542 (N_23542,N_20905,N_21686);
nor U23543 (N_23543,N_21560,N_21338);
nand U23544 (N_23544,N_20795,N_20885);
xnor U23545 (N_23545,N_21534,N_20729);
nor U23546 (N_23546,N_21840,N_21470);
xor U23547 (N_23547,N_21548,N_21724);
xor U23548 (N_23548,N_20958,N_20876);
and U23549 (N_23549,N_20454,N_21129);
or U23550 (N_23550,N_20597,N_21267);
and U23551 (N_23551,N_21918,N_20738);
or U23552 (N_23552,N_20619,N_21242);
nor U23553 (N_23553,N_21290,N_21081);
or U23554 (N_23554,N_20837,N_20345);
or U23555 (N_23555,N_20286,N_20835);
and U23556 (N_23556,N_20052,N_21786);
nor U23557 (N_23557,N_20252,N_20602);
nand U23558 (N_23558,N_21508,N_21386);
nand U23559 (N_23559,N_20377,N_20891);
or U23560 (N_23560,N_21448,N_20958);
or U23561 (N_23561,N_21145,N_21190);
and U23562 (N_23562,N_20338,N_20451);
or U23563 (N_23563,N_20503,N_21292);
nand U23564 (N_23564,N_20260,N_21302);
or U23565 (N_23565,N_20947,N_21784);
nor U23566 (N_23566,N_21458,N_21221);
nand U23567 (N_23567,N_20851,N_21952);
xor U23568 (N_23568,N_21142,N_21754);
xnor U23569 (N_23569,N_21960,N_21281);
nand U23570 (N_23570,N_21412,N_20646);
nor U23571 (N_23571,N_20486,N_21287);
or U23572 (N_23572,N_20922,N_21712);
nand U23573 (N_23573,N_20413,N_21427);
xnor U23574 (N_23574,N_20829,N_20270);
nand U23575 (N_23575,N_20209,N_20917);
nor U23576 (N_23576,N_20269,N_20520);
and U23577 (N_23577,N_20214,N_20376);
nor U23578 (N_23578,N_21044,N_21951);
nand U23579 (N_23579,N_20888,N_21097);
nor U23580 (N_23580,N_20467,N_21287);
or U23581 (N_23581,N_20790,N_20059);
xor U23582 (N_23582,N_21205,N_20122);
nor U23583 (N_23583,N_20555,N_21217);
or U23584 (N_23584,N_20892,N_21693);
xnor U23585 (N_23585,N_21411,N_20022);
and U23586 (N_23586,N_20374,N_21640);
and U23587 (N_23587,N_21983,N_21370);
and U23588 (N_23588,N_20053,N_21388);
nor U23589 (N_23589,N_20780,N_21219);
and U23590 (N_23590,N_21407,N_20224);
or U23591 (N_23591,N_21754,N_20053);
xor U23592 (N_23592,N_21681,N_21626);
nand U23593 (N_23593,N_20200,N_20245);
nor U23594 (N_23594,N_20000,N_20346);
nand U23595 (N_23595,N_21766,N_21357);
xor U23596 (N_23596,N_20208,N_20812);
or U23597 (N_23597,N_20809,N_21452);
or U23598 (N_23598,N_20954,N_20475);
nand U23599 (N_23599,N_20153,N_20537);
xnor U23600 (N_23600,N_21245,N_20804);
or U23601 (N_23601,N_20641,N_21640);
nor U23602 (N_23602,N_20220,N_20017);
nand U23603 (N_23603,N_20154,N_20089);
nand U23604 (N_23604,N_21875,N_20165);
nand U23605 (N_23605,N_20111,N_21528);
nor U23606 (N_23606,N_20429,N_21176);
xnor U23607 (N_23607,N_21911,N_21258);
nor U23608 (N_23608,N_20183,N_21136);
or U23609 (N_23609,N_20413,N_20085);
nand U23610 (N_23610,N_21803,N_20670);
and U23611 (N_23611,N_21684,N_21148);
nand U23612 (N_23612,N_20487,N_20966);
and U23613 (N_23613,N_21796,N_21444);
or U23614 (N_23614,N_21338,N_21760);
nand U23615 (N_23615,N_20904,N_20328);
and U23616 (N_23616,N_21710,N_21506);
and U23617 (N_23617,N_21950,N_20558);
and U23618 (N_23618,N_20721,N_21383);
or U23619 (N_23619,N_20903,N_20139);
nand U23620 (N_23620,N_20220,N_20747);
and U23621 (N_23621,N_20219,N_21073);
or U23622 (N_23622,N_21023,N_20051);
nor U23623 (N_23623,N_20321,N_20594);
and U23624 (N_23624,N_21330,N_20494);
and U23625 (N_23625,N_21598,N_21619);
xnor U23626 (N_23626,N_20875,N_20593);
or U23627 (N_23627,N_21351,N_20420);
or U23628 (N_23628,N_20986,N_21995);
and U23629 (N_23629,N_20051,N_21143);
xor U23630 (N_23630,N_20564,N_20609);
and U23631 (N_23631,N_20689,N_21543);
nor U23632 (N_23632,N_20293,N_21754);
and U23633 (N_23633,N_21730,N_21619);
and U23634 (N_23634,N_21054,N_21720);
xor U23635 (N_23635,N_20828,N_21142);
nand U23636 (N_23636,N_21184,N_20597);
nand U23637 (N_23637,N_20954,N_20458);
xnor U23638 (N_23638,N_20513,N_20354);
nand U23639 (N_23639,N_21673,N_21106);
or U23640 (N_23640,N_20762,N_20837);
nand U23641 (N_23641,N_21559,N_21428);
and U23642 (N_23642,N_20775,N_21494);
xnor U23643 (N_23643,N_21899,N_20641);
and U23644 (N_23644,N_20394,N_21428);
or U23645 (N_23645,N_21523,N_21617);
and U23646 (N_23646,N_20827,N_21664);
xor U23647 (N_23647,N_21593,N_20324);
nor U23648 (N_23648,N_21059,N_20413);
and U23649 (N_23649,N_21439,N_20624);
or U23650 (N_23650,N_20118,N_20978);
nand U23651 (N_23651,N_21790,N_21844);
and U23652 (N_23652,N_20655,N_21542);
nand U23653 (N_23653,N_21529,N_20912);
nor U23654 (N_23654,N_21044,N_20270);
nor U23655 (N_23655,N_21043,N_21505);
and U23656 (N_23656,N_20419,N_20566);
or U23657 (N_23657,N_20408,N_20643);
nor U23658 (N_23658,N_21610,N_20681);
nor U23659 (N_23659,N_20408,N_21582);
and U23660 (N_23660,N_21205,N_20286);
and U23661 (N_23661,N_20083,N_20039);
or U23662 (N_23662,N_20031,N_21602);
nor U23663 (N_23663,N_20624,N_21569);
nand U23664 (N_23664,N_20127,N_21704);
xor U23665 (N_23665,N_21362,N_21228);
nand U23666 (N_23666,N_21051,N_21772);
xor U23667 (N_23667,N_21519,N_21302);
nand U23668 (N_23668,N_21759,N_21350);
or U23669 (N_23669,N_21568,N_20041);
nor U23670 (N_23670,N_20854,N_20261);
and U23671 (N_23671,N_20851,N_21013);
xor U23672 (N_23672,N_20689,N_20523);
nand U23673 (N_23673,N_21560,N_21710);
and U23674 (N_23674,N_21735,N_20118);
and U23675 (N_23675,N_21040,N_20493);
and U23676 (N_23676,N_20081,N_21146);
or U23677 (N_23677,N_21902,N_21186);
and U23678 (N_23678,N_21522,N_21327);
nand U23679 (N_23679,N_21979,N_21982);
nor U23680 (N_23680,N_21144,N_20209);
nor U23681 (N_23681,N_20519,N_20474);
and U23682 (N_23682,N_20466,N_20741);
and U23683 (N_23683,N_21370,N_21905);
nand U23684 (N_23684,N_21978,N_21472);
nor U23685 (N_23685,N_21821,N_20462);
nand U23686 (N_23686,N_20993,N_20277);
xor U23687 (N_23687,N_20075,N_20403);
xnor U23688 (N_23688,N_20316,N_21499);
xor U23689 (N_23689,N_20928,N_20498);
and U23690 (N_23690,N_20680,N_21599);
xnor U23691 (N_23691,N_20687,N_21456);
xnor U23692 (N_23692,N_21867,N_20951);
nor U23693 (N_23693,N_20786,N_20498);
xnor U23694 (N_23694,N_20639,N_20758);
or U23695 (N_23695,N_20132,N_20908);
xnor U23696 (N_23696,N_21058,N_21406);
nor U23697 (N_23697,N_20841,N_21459);
nor U23698 (N_23698,N_20484,N_21698);
and U23699 (N_23699,N_21813,N_21407);
nor U23700 (N_23700,N_20756,N_20053);
xnor U23701 (N_23701,N_21102,N_21803);
xnor U23702 (N_23702,N_20310,N_20164);
xnor U23703 (N_23703,N_21838,N_20958);
nor U23704 (N_23704,N_20963,N_20885);
and U23705 (N_23705,N_21180,N_20713);
or U23706 (N_23706,N_20327,N_21177);
or U23707 (N_23707,N_21848,N_21253);
and U23708 (N_23708,N_21428,N_21195);
xnor U23709 (N_23709,N_21589,N_20337);
xor U23710 (N_23710,N_20144,N_21167);
nor U23711 (N_23711,N_21168,N_20630);
and U23712 (N_23712,N_20792,N_20688);
nor U23713 (N_23713,N_21480,N_21586);
xnor U23714 (N_23714,N_21921,N_21562);
nor U23715 (N_23715,N_20146,N_20887);
nor U23716 (N_23716,N_21287,N_20793);
nand U23717 (N_23717,N_20977,N_21945);
nand U23718 (N_23718,N_21055,N_21460);
nor U23719 (N_23719,N_21990,N_21485);
xor U23720 (N_23720,N_21257,N_21428);
or U23721 (N_23721,N_21157,N_21154);
and U23722 (N_23722,N_20773,N_21711);
and U23723 (N_23723,N_20026,N_21241);
nand U23724 (N_23724,N_20843,N_21540);
xnor U23725 (N_23725,N_21740,N_20958);
nor U23726 (N_23726,N_21145,N_21482);
nor U23727 (N_23727,N_20677,N_21156);
xor U23728 (N_23728,N_20322,N_21220);
and U23729 (N_23729,N_21617,N_21041);
nand U23730 (N_23730,N_21244,N_20496);
and U23731 (N_23731,N_21224,N_20746);
xor U23732 (N_23732,N_20991,N_21081);
nand U23733 (N_23733,N_21194,N_20684);
xnor U23734 (N_23734,N_21402,N_21460);
nand U23735 (N_23735,N_21377,N_21181);
and U23736 (N_23736,N_20322,N_21964);
nand U23737 (N_23737,N_20632,N_20936);
nor U23738 (N_23738,N_20767,N_21836);
or U23739 (N_23739,N_20238,N_20770);
xnor U23740 (N_23740,N_21508,N_21216);
or U23741 (N_23741,N_21842,N_21873);
nor U23742 (N_23742,N_21445,N_21357);
and U23743 (N_23743,N_21981,N_21254);
and U23744 (N_23744,N_21511,N_20537);
and U23745 (N_23745,N_21074,N_20315);
and U23746 (N_23746,N_21925,N_21530);
or U23747 (N_23747,N_21349,N_21488);
nand U23748 (N_23748,N_21900,N_21403);
nand U23749 (N_23749,N_20643,N_21058);
nand U23750 (N_23750,N_20768,N_20853);
xor U23751 (N_23751,N_21206,N_21664);
or U23752 (N_23752,N_21789,N_21199);
nand U23753 (N_23753,N_21950,N_20396);
nand U23754 (N_23754,N_20620,N_20645);
or U23755 (N_23755,N_20666,N_21387);
or U23756 (N_23756,N_21499,N_20390);
nand U23757 (N_23757,N_21832,N_21331);
xnor U23758 (N_23758,N_21661,N_20606);
and U23759 (N_23759,N_21574,N_21398);
and U23760 (N_23760,N_21307,N_21880);
xor U23761 (N_23761,N_21735,N_21929);
or U23762 (N_23762,N_20820,N_20075);
nor U23763 (N_23763,N_20621,N_20488);
xnor U23764 (N_23764,N_21449,N_20868);
xor U23765 (N_23765,N_21961,N_20816);
and U23766 (N_23766,N_20384,N_21551);
or U23767 (N_23767,N_21251,N_20513);
and U23768 (N_23768,N_21252,N_20869);
nor U23769 (N_23769,N_20394,N_21788);
xnor U23770 (N_23770,N_20067,N_20680);
or U23771 (N_23771,N_20415,N_21140);
xnor U23772 (N_23772,N_20102,N_21072);
nor U23773 (N_23773,N_20156,N_21635);
and U23774 (N_23774,N_20514,N_21899);
nor U23775 (N_23775,N_20369,N_20992);
and U23776 (N_23776,N_20734,N_21674);
nor U23777 (N_23777,N_21786,N_21532);
or U23778 (N_23778,N_21885,N_21229);
nor U23779 (N_23779,N_20094,N_21644);
xor U23780 (N_23780,N_21423,N_20799);
xor U23781 (N_23781,N_21611,N_21442);
xnor U23782 (N_23782,N_20565,N_20501);
or U23783 (N_23783,N_21611,N_21095);
and U23784 (N_23784,N_21670,N_21546);
xnor U23785 (N_23785,N_21771,N_20172);
nand U23786 (N_23786,N_21891,N_20725);
nand U23787 (N_23787,N_20006,N_21010);
xnor U23788 (N_23788,N_20263,N_20853);
xor U23789 (N_23789,N_21099,N_20851);
xnor U23790 (N_23790,N_20241,N_20755);
nand U23791 (N_23791,N_20373,N_21021);
and U23792 (N_23792,N_21288,N_21553);
nand U23793 (N_23793,N_21113,N_20280);
nor U23794 (N_23794,N_21287,N_21937);
or U23795 (N_23795,N_21021,N_20201);
nor U23796 (N_23796,N_21997,N_20065);
or U23797 (N_23797,N_21502,N_20143);
or U23798 (N_23798,N_20565,N_21236);
nand U23799 (N_23799,N_20466,N_21822);
xnor U23800 (N_23800,N_20041,N_20309);
and U23801 (N_23801,N_21852,N_20512);
or U23802 (N_23802,N_20227,N_21666);
xnor U23803 (N_23803,N_20919,N_20384);
nand U23804 (N_23804,N_21449,N_21128);
nor U23805 (N_23805,N_21169,N_21072);
and U23806 (N_23806,N_21931,N_21191);
and U23807 (N_23807,N_20716,N_21617);
and U23808 (N_23808,N_21686,N_20172);
xnor U23809 (N_23809,N_21681,N_21114);
and U23810 (N_23810,N_20898,N_20573);
xor U23811 (N_23811,N_20759,N_21069);
or U23812 (N_23812,N_21662,N_21537);
nor U23813 (N_23813,N_21617,N_20807);
and U23814 (N_23814,N_20166,N_20654);
xor U23815 (N_23815,N_20751,N_20841);
or U23816 (N_23816,N_21730,N_20864);
xnor U23817 (N_23817,N_20728,N_21091);
or U23818 (N_23818,N_20521,N_20763);
or U23819 (N_23819,N_20174,N_21613);
nor U23820 (N_23820,N_21315,N_21424);
or U23821 (N_23821,N_20073,N_21479);
or U23822 (N_23822,N_20149,N_21333);
nor U23823 (N_23823,N_21732,N_21680);
nor U23824 (N_23824,N_20785,N_20143);
and U23825 (N_23825,N_20999,N_21057);
or U23826 (N_23826,N_20364,N_21245);
xor U23827 (N_23827,N_21026,N_21994);
nor U23828 (N_23828,N_20338,N_20525);
or U23829 (N_23829,N_21882,N_20966);
nor U23830 (N_23830,N_20882,N_20675);
nor U23831 (N_23831,N_20471,N_21971);
nor U23832 (N_23832,N_21948,N_21448);
and U23833 (N_23833,N_21330,N_21459);
nand U23834 (N_23834,N_20402,N_20054);
xnor U23835 (N_23835,N_20845,N_20645);
or U23836 (N_23836,N_21038,N_20026);
and U23837 (N_23837,N_21419,N_21082);
and U23838 (N_23838,N_21946,N_20625);
or U23839 (N_23839,N_20373,N_20802);
nor U23840 (N_23840,N_21497,N_21590);
nand U23841 (N_23841,N_21924,N_21146);
nand U23842 (N_23842,N_20800,N_21590);
and U23843 (N_23843,N_20421,N_21593);
nor U23844 (N_23844,N_20791,N_20410);
nor U23845 (N_23845,N_20699,N_21341);
nor U23846 (N_23846,N_21288,N_20153);
or U23847 (N_23847,N_21682,N_20023);
xor U23848 (N_23848,N_20898,N_20497);
xor U23849 (N_23849,N_20184,N_20075);
xnor U23850 (N_23850,N_21970,N_20481);
nor U23851 (N_23851,N_20524,N_20068);
nor U23852 (N_23852,N_20187,N_20344);
xnor U23853 (N_23853,N_20056,N_20622);
and U23854 (N_23854,N_21091,N_20447);
xnor U23855 (N_23855,N_21333,N_20123);
nor U23856 (N_23856,N_21988,N_21610);
nand U23857 (N_23857,N_21429,N_21261);
or U23858 (N_23858,N_20147,N_20381);
and U23859 (N_23859,N_21965,N_21817);
nand U23860 (N_23860,N_21478,N_21411);
or U23861 (N_23861,N_20912,N_20397);
nor U23862 (N_23862,N_21699,N_21766);
or U23863 (N_23863,N_20239,N_21478);
and U23864 (N_23864,N_21953,N_21052);
and U23865 (N_23865,N_20672,N_21271);
nand U23866 (N_23866,N_21946,N_20142);
xnor U23867 (N_23867,N_20553,N_20064);
nand U23868 (N_23868,N_21501,N_21847);
and U23869 (N_23869,N_20010,N_21780);
or U23870 (N_23870,N_20339,N_20556);
nor U23871 (N_23871,N_21293,N_21487);
xnor U23872 (N_23872,N_21525,N_21122);
xor U23873 (N_23873,N_20353,N_20466);
nor U23874 (N_23874,N_20047,N_20211);
nor U23875 (N_23875,N_21515,N_20933);
or U23876 (N_23876,N_21650,N_20812);
or U23877 (N_23877,N_21190,N_21573);
xor U23878 (N_23878,N_20984,N_21228);
nor U23879 (N_23879,N_20103,N_20353);
xor U23880 (N_23880,N_20837,N_21435);
or U23881 (N_23881,N_21975,N_20468);
nor U23882 (N_23882,N_20060,N_20840);
xor U23883 (N_23883,N_20439,N_20586);
and U23884 (N_23884,N_20141,N_21421);
xor U23885 (N_23885,N_20234,N_20074);
and U23886 (N_23886,N_21580,N_20685);
nor U23887 (N_23887,N_21867,N_20620);
and U23888 (N_23888,N_20916,N_20569);
or U23889 (N_23889,N_20454,N_20280);
nor U23890 (N_23890,N_21653,N_21186);
nor U23891 (N_23891,N_21151,N_20732);
or U23892 (N_23892,N_20182,N_20372);
nor U23893 (N_23893,N_20125,N_20505);
nand U23894 (N_23894,N_20027,N_21023);
or U23895 (N_23895,N_21785,N_20602);
and U23896 (N_23896,N_20571,N_21196);
nor U23897 (N_23897,N_21299,N_21753);
nor U23898 (N_23898,N_20091,N_20854);
or U23899 (N_23899,N_20740,N_20729);
and U23900 (N_23900,N_20925,N_21604);
nor U23901 (N_23901,N_20976,N_20847);
xnor U23902 (N_23902,N_21769,N_21903);
or U23903 (N_23903,N_21687,N_21541);
and U23904 (N_23904,N_21438,N_21445);
xnor U23905 (N_23905,N_20577,N_20818);
and U23906 (N_23906,N_21689,N_21494);
or U23907 (N_23907,N_21611,N_20902);
nor U23908 (N_23908,N_20712,N_21275);
xnor U23909 (N_23909,N_20008,N_21148);
xor U23910 (N_23910,N_20723,N_21645);
or U23911 (N_23911,N_20014,N_20553);
nand U23912 (N_23912,N_20500,N_20441);
xnor U23913 (N_23913,N_21800,N_20579);
nor U23914 (N_23914,N_20667,N_20327);
xor U23915 (N_23915,N_21509,N_20281);
nand U23916 (N_23916,N_20117,N_20833);
xor U23917 (N_23917,N_21118,N_21012);
nand U23918 (N_23918,N_20554,N_20548);
xnor U23919 (N_23919,N_21711,N_21281);
and U23920 (N_23920,N_21913,N_21093);
and U23921 (N_23921,N_21513,N_21591);
and U23922 (N_23922,N_21580,N_21007);
nand U23923 (N_23923,N_21939,N_21541);
and U23924 (N_23924,N_20946,N_20807);
nor U23925 (N_23925,N_21791,N_21906);
xor U23926 (N_23926,N_20527,N_20193);
xnor U23927 (N_23927,N_20007,N_21464);
xnor U23928 (N_23928,N_20238,N_21275);
and U23929 (N_23929,N_20944,N_21777);
nor U23930 (N_23930,N_21000,N_21892);
or U23931 (N_23931,N_21760,N_21804);
nand U23932 (N_23932,N_20991,N_21626);
nor U23933 (N_23933,N_20178,N_21578);
or U23934 (N_23934,N_20575,N_21900);
nor U23935 (N_23935,N_21931,N_21915);
or U23936 (N_23936,N_20591,N_20551);
nor U23937 (N_23937,N_21315,N_21751);
nand U23938 (N_23938,N_21728,N_21179);
or U23939 (N_23939,N_20827,N_21806);
nand U23940 (N_23940,N_21914,N_21975);
and U23941 (N_23941,N_21199,N_21141);
or U23942 (N_23942,N_21976,N_20881);
or U23943 (N_23943,N_21916,N_20190);
nor U23944 (N_23944,N_20122,N_20916);
nand U23945 (N_23945,N_20153,N_21373);
nor U23946 (N_23946,N_21623,N_20078);
nand U23947 (N_23947,N_21595,N_20954);
nor U23948 (N_23948,N_21766,N_21007);
nand U23949 (N_23949,N_21295,N_21053);
nor U23950 (N_23950,N_20231,N_21528);
nor U23951 (N_23951,N_21935,N_20400);
nand U23952 (N_23952,N_21434,N_21488);
or U23953 (N_23953,N_21721,N_21289);
and U23954 (N_23954,N_20535,N_20349);
xor U23955 (N_23955,N_20057,N_20697);
xnor U23956 (N_23956,N_20153,N_20735);
xor U23957 (N_23957,N_21693,N_21905);
and U23958 (N_23958,N_20811,N_21620);
and U23959 (N_23959,N_20017,N_21861);
and U23960 (N_23960,N_20021,N_20776);
nand U23961 (N_23961,N_20494,N_21198);
xor U23962 (N_23962,N_21799,N_21695);
nor U23963 (N_23963,N_21725,N_21846);
nor U23964 (N_23964,N_20961,N_20832);
or U23965 (N_23965,N_20315,N_21966);
or U23966 (N_23966,N_20670,N_21586);
nor U23967 (N_23967,N_21138,N_21056);
and U23968 (N_23968,N_21150,N_20234);
and U23969 (N_23969,N_20874,N_20614);
xnor U23970 (N_23970,N_21351,N_21500);
xor U23971 (N_23971,N_21113,N_21351);
xnor U23972 (N_23972,N_20173,N_21885);
nand U23973 (N_23973,N_21738,N_21071);
or U23974 (N_23974,N_21265,N_21942);
xor U23975 (N_23975,N_20128,N_21221);
or U23976 (N_23976,N_20886,N_21326);
xnor U23977 (N_23977,N_21857,N_20417);
xor U23978 (N_23978,N_21076,N_20983);
nor U23979 (N_23979,N_20718,N_21054);
nor U23980 (N_23980,N_20363,N_21874);
xnor U23981 (N_23981,N_21145,N_21558);
nor U23982 (N_23982,N_21633,N_20775);
or U23983 (N_23983,N_21456,N_21071);
or U23984 (N_23984,N_20659,N_20011);
and U23985 (N_23985,N_20082,N_20948);
xnor U23986 (N_23986,N_20951,N_20524);
or U23987 (N_23987,N_20937,N_21816);
xnor U23988 (N_23988,N_21990,N_21259);
nor U23989 (N_23989,N_20376,N_20338);
xor U23990 (N_23990,N_20237,N_21994);
or U23991 (N_23991,N_21092,N_20167);
and U23992 (N_23992,N_20750,N_20450);
nor U23993 (N_23993,N_21325,N_21903);
nand U23994 (N_23994,N_21327,N_20048);
xor U23995 (N_23995,N_20806,N_21749);
or U23996 (N_23996,N_21743,N_21110);
or U23997 (N_23997,N_21328,N_20935);
or U23998 (N_23998,N_20639,N_20149);
xor U23999 (N_23999,N_21117,N_21985);
nand U24000 (N_24000,N_22480,N_23837);
nand U24001 (N_24001,N_22798,N_23111);
xnor U24002 (N_24002,N_23532,N_22255);
nand U24003 (N_24003,N_23106,N_22324);
xnor U24004 (N_24004,N_23434,N_22010);
xnor U24005 (N_24005,N_23988,N_22006);
xnor U24006 (N_24006,N_22829,N_22364);
nand U24007 (N_24007,N_22081,N_23744);
nor U24008 (N_24008,N_23573,N_23139);
and U24009 (N_24009,N_22143,N_22688);
or U24010 (N_24010,N_22115,N_22648);
or U24011 (N_24011,N_22151,N_23323);
or U24012 (N_24012,N_23456,N_22557);
or U24013 (N_24013,N_22745,N_23529);
or U24014 (N_24014,N_22504,N_22879);
nor U24015 (N_24015,N_23596,N_22612);
or U24016 (N_24016,N_22711,N_23644);
nand U24017 (N_24017,N_22202,N_23608);
nor U24018 (N_24018,N_22858,N_23257);
or U24019 (N_24019,N_23360,N_23233);
nor U24020 (N_24020,N_23759,N_22672);
and U24021 (N_24021,N_23224,N_22349);
or U24022 (N_24022,N_22306,N_22397);
xnor U24023 (N_24023,N_23873,N_23686);
nand U24024 (N_24024,N_22889,N_23882);
or U24025 (N_24025,N_23348,N_23653);
and U24026 (N_24026,N_23019,N_23690);
xor U24027 (N_24027,N_22989,N_23112);
nand U24028 (N_24028,N_22922,N_22490);
nor U24029 (N_24029,N_22186,N_23420);
nand U24030 (N_24030,N_22847,N_23404);
or U24031 (N_24031,N_23743,N_22731);
and U24032 (N_24032,N_22749,N_23130);
nor U24033 (N_24033,N_23026,N_23063);
or U24034 (N_24034,N_23168,N_23095);
xor U24035 (N_24035,N_22603,N_23062);
or U24036 (N_24036,N_22511,N_22302);
nand U24037 (N_24037,N_23500,N_23713);
xor U24038 (N_24038,N_23048,N_23210);
and U24039 (N_24039,N_23290,N_22232);
nor U24040 (N_24040,N_23734,N_22789);
and U24041 (N_24041,N_23736,N_22801);
and U24042 (N_24042,N_22403,N_22367);
and U24043 (N_24043,N_22866,N_22300);
xor U24044 (N_24044,N_23140,N_22588);
nand U24045 (N_24045,N_23192,N_22558);
xnor U24046 (N_24046,N_23909,N_23856);
nand U24047 (N_24047,N_22193,N_23568);
and U24048 (N_24048,N_23643,N_23011);
xor U24049 (N_24049,N_22802,N_22914);
nor U24050 (N_24050,N_22919,N_23179);
xnor U24051 (N_24051,N_23370,N_22336);
nand U24052 (N_24052,N_23945,N_23213);
or U24053 (N_24053,N_22138,N_23116);
or U24054 (N_24054,N_23247,N_22319);
xor U24055 (N_24055,N_23927,N_22518);
or U24056 (N_24056,N_23835,N_23515);
xnor U24057 (N_24057,N_22695,N_22572);
and U24058 (N_24058,N_22087,N_23479);
nor U24059 (N_24059,N_22975,N_23359);
xor U24060 (N_24060,N_22345,N_22410);
or U24061 (N_24061,N_23305,N_23226);
xnor U24062 (N_24062,N_23947,N_23833);
and U24063 (N_24063,N_22983,N_23913);
or U24064 (N_24064,N_23763,N_23096);
nor U24065 (N_24065,N_22875,N_23390);
or U24066 (N_24066,N_23920,N_23100);
and U24067 (N_24067,N_23214,N_23142);
and U24068 (N_24068,N_23351,N_22150);
and U24069 (N_24069,N_23950,N_22548);
or U24070 (N_24070,N_23342,N_22222);
and U24071 (N_24071,N_23667,N_22824);
nand U24072 (N_24072,N_23468,N_22192);
and U24073 (N_24073,N_23242,N_23151);
nor U24074 (N_24074,N_23992,N_22303);
xor U24075 (N_24075,N_22358,N_23366);
nand U24076 (N_24076,N_22465,N_23990);
nand U24077 (N_24077,N_23782,N_23204);
or U24078 (N_24078,N_23004,N_22630);
nand U24079 (N_24079,N_22917,N_22284);
nand U24080 (N_24080,N_23519,N_22826);
or U24081 (N_24081,N_23921,N_23633);
xnor U24082 (N_24082,N_22174,N_22476);
xor U24083 (N_24083,N_23944,N_22813);
nand U24084 (N_24084,N_23382,N_23041);
nand U24085 (N_24085,N_23306,N_22162);
nor U24086 (N_24086,N_23691,N_22433);
xnor U24087 (N_24087,N_22398,N_22442);
nor U24088 (N_24088,N_23929,N_23170);
xnor U24089 (N_24089,N_23013,N_23783);
nor U24090 (N_24090,N_22415,N_23528);
xnor U24091 (N_24091,N_22609,N_23769);
nand U24092 (N_24092,N_23294,N_23578);
and U24093 (N_24093,N_22843,N_22329);
or U24094 (N_24094,N_23732,N_22120);
or U24095 (N_24095,N_22873,N_23613);
xor U24096 (N_24096,N_22706,N_22987);
or U24097 (N_24097,N_22363,N_23006);
or U24098 (N_24098,N_23745,N_23387);
nor U24099 (N_24099,N_22468,N_23791);
nor U24100 (N_24100,N_22269,N_22708);
and U24101 (N_24101,N_22109,N_23017);
xor U24102 (N_24102,N_22633,N_22301);
and U24103 (N_24103,N_23349,N_23655);
nand U24104 (N_24104,N_23815,N_22154);
nor U24105 (N_24105,N_23138,N_23730);
xor U24106 (N_24106,N_22309,N_23275);
and U24107 (N_24107,N_22064,N_22126);
or U24108 (N_24108,N_23900,N_22215);
nand U24109 (N_24109,N_23163,N_22788);
nor U24110 (N_24110,N_22510,N_22435);
nand U24111 (N_24111,N_22728,N_22751);
or U24112 (N_24112,N_23657,N_23735);
nor U24113 (N_24113,N_23535,N_22496);
nand U24114 (N_24114,N_23804,N_23796);
nor U24115 (N_24115,N_22057,N_22485);
or U24116 (N_24116,N_23180,N_23482);
or U24117 (N_24117,N_23493,N_23631);
xor U24118 (N_24118,N_22187,N_22430);
or U24119 (N_24119,N_22602,N_22935);
or U24120 (N_24120,N_22456,N_22599);
xor U24121 (N_24121,N_22070,N_23339);
and U24122 (N_24122,N_23392,N_22778);
or U24123 (N_24123,N_22231,N_22979);
and U24124 (N_24124,N_22136,N_22635);
or U24125 (N_24125,N_23523,N_23716);
nor U24126 (N_24126,N_22277,N_22412);
or U24127 (N_24127,N_23039,N_22692);
and U24128 (N_24128,N_22893,N_23037);
nand U24129 (N_24129,N_22304,N_22876);
xnor U24130 (N_24130,N_22481,N_22295);
nor U24131 (N_24131,N_22921,N_22075);
and U24132 (N_24132,N_22455,N_23543);
nor U24133 (N_24133,N_22253,N_22111);
and U24134 (N_24134,N_23637,N_22153);
nand U24135 (N_24135,N_23032,N_22591);
nor U24136 (N_24136,N_22330,N_23396);
nor U24137 (N_24137,N_22952,N_23984);
xnor U24138 (N_24138,N_22394,N_23787);
xor U24139 (N_24139,N_23975,N_22560);
and U24140 (N_24140,N_22988,N_22125);
or U24141 (N_24141,N_22950,N_23453);
and U24142 (N_24142,N_22170,N_23647);
nor U24143 (N_24143,N_22369,N_22738);
or U24144 (N_24144,N_22758,N_23808);
or U24145 (N_24145,N_22513,N_22252);
and U24146 (N_24146,N_23181,N_23939);
or U24147 (N_24147,N_22242,N_22827);
and U24148 (N_24148,N_22529,N_22821);
nand U24149 (N_24149,N_23276,N_23252);
nor U24150 (N_24150,N_22947,N_23982);
nor U24151 (N_24151,N_22288,N_22595);
nor U24152 (N_24152,N_23271,N_22332);
and U24153 (N_24153,N_22981,N_23943);
nor U24154 (N_24154,N_22608,N_22164);
nor U24155 (N_24155,N_23255,N_23309);
xnor U24156 (N_24156,N_23948,N_22933);
and U24157 (N_24157,N_23172,N_23991);
nand U24158 (N_24158,N_23976,N_22770);
nand U24159 (N_24159,N_23002,N_22908);
and U24160 (N_24160,N_23332,N_22487);
or U24161 (N_24161,N_23418,N_22258);
and U24162 (N_24162,N_22948,N_23709);
xnor U24163 (N_24163,N_22857,N_22763);
xor U24164 (N_24164,N_22765,N_22058);
nand U24165 (N_24165,N_22026,N_23220);
nor U24166 (N_24166,N_23588,N_22573);
or U24167 (N_24167,N_22799,N_22268);
nand U24168 (N_24168,N_22168,N_23639);
or U24169 (N_24169,N_22411,N_23788);
or U24170 (N_24170,N_22634,N_22619);
nand U24171 (N_24171,N_22382,N_22484);
nand U24172 (N_24172,N_22088,N_23614);
nor U24173 (N_24173,N_22836,N_22526);
xor U24174 (N_24174,N_23187,N_22912);
nand U24175 (N_24175,N_22003,N_23521);
nand U24176 (N_24176,N_23999,N_22899);
nor U24177 (N_24177,N_23166,N_23406);
xnor U24178 (N_24178,N_22920,N_23258);
and U24179 (N_24179,N_23353,N_22974);
nor U24180 (N_24180,N_23288,N_22698);
nand U24181 (N_24181,N_23956,N_22477);
nor U24182 (N_24182,N_23823,N_23560);
or U24183 (N_24183,N_23864,N_23818);
xnor U24184 (N_24184,N_23968,N_22308);
nand U24185 (N_24185,N_22533,N_23610);
nand U24186 (N_24186,N_23520,N_22766);
nor U24187 (N_24187,N_22185,N_22915);
nor U24188 (N_24188,N_23946,N_23137);
or U24189 (N_24189,N_23737,N_22531);
nor U24190 (N_24190,N_22149,N_22822);
nand U24191 (N_24191,N_22495,N_22173);
nor U24192 (N_24192,N_22144,N_23300);
nand U24193 (N_24193,N_23705,N_23099);
xor U24194 (N_24194,N_23419,N_23394);
nor U24195 (N_24195,N_23399,N_22094);
nand U24196 (N_24196,N_23652,N_23295);
xnor U24197 (N_24197,N_22502,N_22462);
and U24198 (N_24198,N_23451,N_23001);
or U24199 (N_24199,N_23888,N_23025);
and U24200 (N_24200,N_22916,N_22217);
or U24201 (N_24201,N_23518,N_23113);
and U24202 (N_24202,N_22236,N_22965);
nand U24203 (N_24203,N_22527,N_22687);
xor U24204 (N_24204,N_22507,N_23376);
nor U24205 (N_24205,N_22072,N_23860);
nor U24206 (N_24206,N_23282,N_22571);
nor U24207 (N_24207,N_22506,N_23317);
xnor U24208 (N_24208,N_22761,N_23671);
nor U24209 (N_24209,N_23849,N_23491);
or U24210 (N_24210,N_22638,N_22171);
or U24211 (N_24211,N_22275,N_22867);
nand U24212 (N_24212,N_23768,N_23169);
and U24213 (N_24213,N_23741,N_22498);
xor U24214 (N_24214,N_23908,N_23502);
and U24215 (N_24215,N_23278,N_22311);
xor U24216 (N_24216,N_23775,N_23703);
and U24217 (N_24217,N_23374,N_23325);
xnor U24218 (N_24218,N_23758,N_23827);
xor U24219 (N_24219,N_22872,N_23051);
xor U24220 (N_24220,N_22928,N_23906);
and U24221 (N_24221,N_23426,N_23158);
xnor U24222 (N_24222,N_23156,N_22943);
xnor U24223 (N_24223,N_22605,N_22264);
or U24224 (N_24224,N_23102,N_22239);
and U24225 (N_24225,N_22113,N_23280);
nand U24226 (N_24226,N_23486,N_23701);
or U24227 (N_24227,N_22830,N_23831);
nor U24228 (N_24228,N_23403,N_22444);
or U24229 (N_24229,N_23429,N_23119);
xnor U24230 (N_24230,N_22354,N_22265);
nor U24231 (N_24231,N_23718,N_22971);
and U24232 (N_24232,N_23668,N_22800);
and U24233 (N_24233,N_23662,N_23915);
and U24234 (N_24234,N_22840,N_22520);
nor U24235 (N_24235,N_23965,N_23246);
nor U24236 (N_24236,N_23884,N_22715);
xor U24237 (N_24237,N_22169,N_22624);
nor U24238 (N_24238,N_23425,N_22771);
nor U24239 (N_24239,N_23766,N_22639);
or U24240 (N_24240,N_22229,N_22844);
nand U24241 (N_24241,N_23128,N_23423);
nor U24242 (N_24242,N_22133,N_22885);
nor U24243 (N_24243,N_22936,N_22175);
and U24244 (N_24244,N_23802,N_23072);
nand U24245 (N_24245,N_22563,N_23338);
and U24246 (N_24246,N_23196,N_23961);
nand U24247 (N_24247,N_22365,N_23503);
and U24248 (N_24248,N_22562,N_23885);
nor U24249 (N_24249,N_23589,N_22048);
nor U24250 (N_24250,N_23414,N_23512);
or U24251 (N_24251,N_23564,N_22969);
or U24252 (N_24252,N_23283,N_23424);
and U24253 (N_24253,N_22768,N_23053);
xor U24254 (N_24254,N_22420,N_23987);
nor U24255 (N_24255,N_22559,N_22240);
or U24256 (N_24256,N_22655,N_23682);
nand U24257 (N_24257,N_23822,N_23846);
nor U24258 (N_24258,N_22419,N_22748);
and U24259 (N_24259,N_22331,N_22880);
and U24260 (N_24260,N_22226,N_23244);
nand U24261 (N_24261,N_22790,N_22046);
or U24262 (N_24262,N_22680,N_22029);
or U24263 (N_24263,N_22500,N_22341);
or U24264 (N_24264,N_22964,N_22584);
and U24265 (N_24265,N_23061,N_22347);
xnor U24266 (N_24266,N_22654,N_22135);
and U24267 (N_24267,N_22862,N_22219);
and U24268 (N_24268,N_22315,N_22597);
nand U24269 (N_24269,N_23485,N_23940);
xnor U24270 (N_24270,N_22414,N_22156);
and U24271 (N_24271,N_23889,N_23391);
and U24272 (N_24272,N_22927,N_23186);
nand U24273 (N_24273,N_23807,N_23206);
nand U24274 (N_24274,N_23058,N_22205);
nor U24275 (N_24275,N_23925,N_22593);
nor U24276 (N_24276,N_23607,N_23498);
nand U24277 (N_24277,N_23141,N_22587);
nor U24278 (N_24278,N_23816,N_23316);
nand U24279 (N_24279,N_23297,N_22614);
nor U24280 (N_24280,N_23262,N_22626);
or U24281 (N_24281,N_22176,N_23974);
nand U24282 (N_24282,N_22353,N_23836);
and U24283 (N_24283,N_22877,N_22723);
nor U24284 (N_24284,N_22632,N_22036);
or U24285 (N_24285,N_22716,N_23462);
xor U24286 (N_24286,N_23739,N_22503);
xor U24287 (N_24287,N_23337,N_23164);
or U24288 (N_24288,N_22776,N_22069);
and U24289 (N_24289,N_22409,N_23334);
nor U24290 (N_24290,N_22116,N_23937);
and U24291 (N_24291,N_22960,N_23380);
nor U24292 (N_24292,N_23555,N_22184);
and U24293 (N_24293,N_22678,N_22196);
nand U24294 (N_24294,N_23042,N_23695);
and U24295 (N_24295,N_22677,N_22926);
or U24296 (N_24296,N_23875,N_22181);
and U24297 (N_24297,N_23202,N_22640);
nor U24298 (N_24298,N_23761,N_22213);
nor U24299 (N_24299,N_22710,N_22041);
nand U24300 (N_24300,N_22071,N_22390);
xor U24301 (N_24301,N_23484,N_23794);
or U24302 (N_24302,N_23757,N_23448);
nand U24303 (N_24303,N_22567,N_23932);
and U24304 (N_24304,N_23707,N_23412);
or U24305 (N_24305,N_23447,N_22977);
nand U24306 (N_24306,N_22472,N_23477);
nand U24307 (N_24307,N_23779,N_22247);
and U24308 (N_24308,N_22137,N_22452);
xnor U24309 (N_24309,N_23372,N_22134);
nor U24310 (N_24310,N_23413,N_22543);
or U24311 (N_24311,N_22610,N_22729);
nand U24312 (N_24312,N_23840,N_22249);
and U24313 (N_24313,N_22243,N_23160);
xor U24314 (N_24314,N_23291,N_22483);
or U24315 (N_24315,N_22643,N_22266);
nand U24316 (N_24316,N_23356,N_22463);
nand U24317 (N_24317,N_22155,N_22600);
xor U24318 (N_24318,N_22179,N_23812);
xor U24319 (N_24319,N_22703,N_22777);
nand U24320 (N_24320,N_23383,N_23872);
and U24321 (N_24321,N_23729,N_23236);
and U24322 (N_24322,N_23362,N_22359);
nand U24323 (N_24323,N_22868,N_23641);
and U24324 (N_24324,N_22882,N_23431);
or U24325 (N_24325,N_23393,N_23223);
xor U24326 (N_24326,N_22084,N_23941);
nand U24327 (N_24327,N_22489,N_23702);
nand U24328 (N_24328,N_23587,N_23760);
and U24329 (N_24329,N_23828,N_23517);
nor U24330 (N_24330,N_22248,N_23243);
xor U24331 (N_24331,N_22114,N_22180);
or U24332 (N_24332,N_22719,N_22225);
nor U24333 (N_24333,N_23120,N_22376);
and U24334 (N_24334,N_23862,N_23361);
or U24335 (N_24335,N_22049,N_23774);
nor U24336 (N_24336,N_22956,N_22244);
and U24337 (N_24337,N_23126,N_23470);
nor U24338 (N_24338,N_22002,N_23959);
nor U24339 (N_24339,N_23865,N_23472);
or U24340 (N_24340,N_23661,N_23003);
nor U24341 (N_24341,N_23191,N_22387);
and U24342 (N_24342,N_23781,N_22725);
and U24343 (N_24343,N_23537,N_22890);
nor U24344 (N_24344,N_22019,N_22413);
xnor U24345 (N_24345,N_23844,N_22054);
and U24346 (N_24346,N_22523,N_23416);
nand U24347 (N_24347,N_23918,N_22340);
xor U24348 (N_24348,N_23617,N_23134);
xnor U24349 (N_24349,N_22539,N_23153);
nand U24350 (N_24350,N_23952,N_22661);
xnor U24351 (N_24351,N_22393,N_23509);
nor U24352 (N_24352,N_23964,N_22322);
nor U24353 (N_24353,N_23103,N_22980);
and U24354 (N_24354,N_23422,N_22707);
or U24355 (N_24355,N_22596,N_23955);
and U24356 (N_24356,N_23131,N_22383);
xor U24357 (N_24357,N_22092,N_23684);
and U24358 (N_24358,N_23710,N_23998);
nor U24359 (N_24359,N_22611,N_23645);
nand U24360 (N_24360,N_22177,N_22546);
xor U24361 (N_24361,N_23465,N_22620);
nor U24362 (N_24362,N_23752,N_23566);
or U24363 (N_24363,N_22110,N_23049);
nand U24364 (N_24364,N_23497,N_23154);
nand U24365 (N_24365,N_23594,N_23365);
xnor U24366 (N_24366,N_23327,N_23089);
and U24367 (N_24367,N_23616,N_22902);
nor U24368 (N_24368,N_23586,N_23241);
or U24369 (N_24369,N_23886,N_22212);
and U24370 (N_24370,N_23685,N_22894);
nand U24371 (N_24371,N_23516,N_22165);
nor U24372 (N_24372,N_22431,N_23328);
or U24373 (N_24373,N_23966,N_22128);
nor U24374 (N_24374,N_22755,N_23970);
nor U24375 (N_24375,N_23436,N_22080);
or U24376 (N_24376,N_23459,N_23307);
or U24377 (N_24377,N_22649,N_23274);
nor U24378 (N_24378,N_22741,N_22705);
and U24379 (N_24379,N_23367,N_22499);
or U24380 (N_24380,N_22853,N_23625);
and U24381 (N_24381,N_22424,N_22117);
and U24382 (N_24382,N_23091,N_23868);
nor U24383 (N_24383,N_22625,N_22550);
and U24384 (N_24384,N_22845,N_23531);
xnor U24385 (N_24385,N_22101,N_23678);
or U24386 (N_24386,N_22470,N_22407);
nand U24387 (N_24387,N_23540,N_22962);
nor U24388 (N_24388,N_22994,N_23666);
xor U24389 (N_24389,N_23973,N_22001);
nand U24390 (N_24390,N_23469,N_22547);
or U24391 (N_24391,N_22395,N_23722);
and U24392 (N_24392,N_23762,N_23087);
or U24393 (N_24393,N_23824,N_22321);
and U24394 (N_24394,N_22786,N_23912);
and U24395 (N_24395,N_23415,N_23162);
nor U24396 (N_24396,N_22760,N_22955);
or U24397 (N_24397,N_23237,N_23504);
xor U24398 (N_24398,N_22355,N_23660);
nor U24399 (N_24399,N_22050,N_22565);
and U24400 (N_24400,N_22287,N_22191);
nand U24401 (N_24401,N_23793,N_23178);
nand U24402 (N_24402,N_22835,N_22271);
or U24403 (N_24403,N_23304,N_23487);
or U24404 (N_24404,N_22934,N_23373);
or U24405 (N_24405,N_23215,N_22147);
and U24406 (N_24406,N_22474,N_22024);
or U24407 (N_24407,N_23183,N_22833);
xnor U24408 (N_24408,N_23917,N_23452);
xnor U24409 (N_24409,N_22296,N_22579);
and U24410 (N_24410,N_22891,N_22645);
and U24411 (N_24411,N_22000,N_23114);
nand U24412 (N_24412,N_23747,N_22682);
nor U24413 (N_24413,N_22348,N_22743);
nor U24414 (N_24414,N_23738,N_22097);
nor U24415 (N_24415,N_23301,N_23993);
and U24416 (N_24416,N_23123,N_22959);
nor U24417 (N_24417,N_23277,N_22528);
or U24418 (N_24418,N_23907,N_22005);
and U24419 (N_24419,N_23090,N_22525);
nor U24420 (N_24420,N_23958,N_22090);
nor U24421 (N_24421,N_23953,N_23024);
or U24422 (N_24422,N_23819,N_23047);
xor U24423 (N_24423,N_22973,N_22011);
nor U24424 (N_24424,N_22371,N_23539);
nor U24425 (N_24425,N_22190,N_22976);
nand U24426 (N_24426,N_23583,N_23298);
or U24427 (N_24427,N_22273,N_22052);
xnor U24428 (N_24428,N_22542,N_22556);
xor U24429 (N_24429,N_23038,N_23942);
and U24430 (N_24430,N_23995,N_22122);
nor U24431 (N_24431,N_23411,N_22929);
or U24432 (N_24432,N_22404,N_23044);
nand U24433 (N_24433,N_23933,N_23863);
xnor U24434 (N_24434,N_23358,N_22530);
and U24435 (N_24435,N_22014,N_22025);
nand U24436 (N_24436,N_23176,N_22792);
nor U24437 (N_24437,N_22820,N_22178);
xor U24438 (N_24438,N_22869,N_22425);
xnor U24439 (N_24439,N_22667,N_23855);
xor U24440 (N_24440,N_23859,N_23963);
nor U24441 (N_24441,N_22439,N_23867);
or U24442 (N_24442,N_22954,N_22063);
xor U24443 (N_24443,N_22028,N_22482);
nand U24444 (N_24444,N_23731,N_23629);
nor U24445 (N_24445,N_22860,N_22022);
xor U24446 (N_24446,N_22441,N_22004);
or U24447 (N_24447,N_22683,N_22132);
or U24448 (N_24448,N_22781,N_23630);
nor U24449 (N_24449,N_22228,N_23877);
or U24450 (N_24450,N_22290,N_22158);
or U24451 (N_24451,N_23626,N_23673);
and U24452 (N_24452,N_22582,N_22607);
xnor U24453 (N_24453,N_23852,N_22754);
or U24454 (N_24454,N_22453,N_23461);
and U24455 (N_24455,N_22123,N_22457);
and U24456 (N_24456,N_22042,N_23980);
xor U24457 (N_24457,N_22522,N_23597);
nor U24458 (N_24458,N_22131,N_22871);
nor U24459 (N_24459,N_23664,N_23847);
nand U24460 (N_24460,N_23445,N_23585);
nand U24461 (N_24461,N_22888,N_23430);
or U24462 (N_24462,N_23772,N_22993);
and U24463 (N_24463,N_22316,N_22617);
nand U24464 (N_24464,N_22750,N_22372);
nor U24465 (N_24465,N_23656,N_23075);
xnor U24466 (N_24466,N_22580,N_22037);
xor U24467 (N_24467,N_22031,N_23199);
nand U24468 (N_24468,N_23989,N_23245);
or U24469 (N_24469,N_23728,N_23104);
xor U24470 (N_24470,N_23533,N_23005);
and U24471 (N_24471,N_23997,N_23417);
nand U24472 (N_24472,N_22370,N_23525);
xnor U24473 (N_24473,N_23773,N_23746);
nand U24474 (N_24474,N_23511,N_22327);
and U24475 (N_24475,N_23279,N_22906);
nand U24476 (N_24476,N_22756,N_23478);
nand U24477 (N_24477,N_23015,N_22516);
or U24478 (N_24478,N_22554,N_23118);
or U24479 (N_24479,N_22245,N_22129);
nand U24480 (N_24480,N_23742,N_22333);
or U24481 (N_24481,N_23441,N_22021);
nand U24482 (N_24482,N_22378,N_22015);
or U24483 (N_24483,N_23067,N_23712);
xor U24484 (N_24484,N_23088,N_23129);
xor U24485 (N_24485,N_22590,N_23324);
nand U24486 (N_24486,N_22918,N_23771);
nand U24487 (N_24487,N_23527,N_22045);
or U24488 (N_24488,N_23251,N_22195);
nand U24489 (N_24489,N_23209,N_23217);
xnor U24490 (N_24490,N_22068,N_22328);
nor U24491 (N_24491,N_22183,N_22604);
nand U24492 (N_24492,N_22062,N_23018);
or U24493 (N_24493,N_22027,N_22712);
and U24494 (N_24494,N_22938,N_23810);
or U24495 (N_24495,N_23266,N_23801);
or U24496 (N_24496,N_23322,N_22825);
nor U24497 (N_24497,N_22839,N_22818);
xnor U24498 (N_24498,N_23029,N_22188);
nand U24499 (N_24499,N_23542,N_22552);
or U24500 (N_24500,N_23615,N_22944);
nand U24501 (N_24501,N_22142,N_23369);
or U24502 (N_24502,N_22995,N_23876);
nor U24503 (N_24503,N_22996,N_23845);
xor U24504 (N_24504,N_23008,N_22400);
nand U24505 (N_24505,N_22257,N_22901);
or U24506 (N_24506,N_22233,N_23046);
and U24507 (N_24507,N_23800,N_22681);
or U24508 (N_24508,N_23219,N_23972);
xor U24509 (N_24509,N_22318,N_22757);
xor U24510 (N_24510,N_23620,N_22594);
nor U24511 (N_24511,N_22656,N_23287);
xor U24512 (N_24512,N_22951,N_22998);
nor U24513 (N_24513,N_22020,N_23727);
xor U24514 (N_24514,N_22197,N_23159);
or U24515 (N_24515,N_22342,N_22985);
xor U24516 (N_24516,N_22535,N_23398);
or U24517 (N_24517,N_22855,N_22224);
nor U24518 (N_24518,N_22357,N_23981);
or U24519 (N_24519,N_22008,N_23234);
and U24520 (N_24520,N_22704,N_23534);
nand U24521 (N_24521,N_22443,N_22784);
nor U24522 (N_24522,N_22445,N_22544);
nor U24523 (N_24523,N_23805,N_23105);
and U24524 (N_24524,N_22809,N_22429);
or U24525 (N_24525,N_22083,N_23699);
xnor U24526 (N_24526,N_22796,N_23593);
nand U24527 (N_24527,N_23127,N_23592);
xor U24528 (N_24528,N_22966,N_22160);
nand U24529 (N_24529,N_23207,N_23601);
nand U24530 (N_24530,N_23834,N_22234);
nor U24531 (N_24531,N_23405,N_22782);
nor U24532 (N_24532,N_23572,N_23700);
nor U24533 (N_24533,N_23598,N_22689);
and U24534 (N_24534,N_23045,N_22972);
and U24535 (N_24535,N_23284,N_23433);
and U24536 (N_24536,N_22436,N_23971);
nand U24537 (N_24537,N_22702,N_23954);
xor U24538 (N_24538,N_23554,N_22812);
xor U24539 (N_24539,N_22752,N_23345);
nand U24540 (N_24540,N_23122,N_23386);
xnor U24541 (N_24541,N_23510,N_22053);
xor U24542 (N_24542,N_23221,N_23432);
or U24543 (N_24543,N_23326,N_22615);
nand U24544 (N_24544,N_23609,N_23216);
xor U24545 (N_24545,N_23488,N_22911);
xnor U24546 (N_24546,N_22787,N_23364);
xor U24547 (N_24547,N_23789,N_22854);
or U24548 (N_24548,N_23343,N_22446);
or U24549 (N_24549,N_22105,N_22892);
and U24550 (N_24550,N_22067,N_23150);
nand U24551 (N_24551,N_23513,N_22541);
or U24552 (N_24552,N_22256,N_23559);
nand U24553 (N_24553,N_23591,N_23155);
xnor U24554 (N_24554,N_23402,N_22684);
nand U24555 (N_24555,N_22406,N_23926);
or U24556 (N_24556,N_22281,N_23681);
nor U24557 (N_24557,N_22032,N_22870);
xnor U24558 (N_24558,N_23692,N_23079);
or U24559 (N_24559,N_23292,N_23194);
nand U24560 (N_24560,N_22200,N_22722);
nor U24561 (N_24561,N_22086,N_23421);
or U24562 (N_24562,N_22313,N_23674);
and U24563 (N_24563,N_23632,N_23696);
nand U24564 (N_24564,N_23460,N_23635);
xnor U24565 (N_24565,N_23407,N_22235);
nand U24566 (N_24566,N_23121,N_22402);
or U24567 (N_24567,N_23725,N_22167);
nor U24568 (N_24568,N_23967,N_22837);
or U24569 (N_24569,N_23780,N_22618);
or U24570 (N_24570,N_23795,N_22794);
xnor U24571 (N_24571,N_23060,N_22613);
or U24572 (N_24572,N_22904,N_22059);
nor U24573 (N_24573,N_23035,N_22759);
xor U24574 (N_24574,N_22671,N_23253);
or U24575 (N_24575,N_22356,N_23922);
nor U24576 (N_24576,N_22283,N_22381);
nor U24577 (N_24577,N_22691,N_22968);
and U24578 (N_24578,N_23286,N_22060);
or U24579 (N_24579,N_22039,N_22753);
nor U24580 (N_24580,N_22343,N_23951);
nand U24581 (N_24581,N_23851,N_23624);
nor U24582 (N_24582,N_23021,N_22564);
or U24583 (N_24583,N_22505,N_23443);
nand U24584 (N_24584,N_22713,N_23033);
xor U24585 (N_24585,N_23201,N_23385);
xnor U24586 (N_24586,N_22650,N_22467);
xnor U24587 (N_24587,N_23936,N_23077);
or U24588 (N_24588,N_22066,N_23841);
nor U24589 (N_24589,N_22740,N_23384);
and U24590 (N_24590,N_22970,N_23683);
and U24591 (N_24591,N_23861,N_23010);
nor U24592 (N_24592,N_22747,N_22307);
xor U24593 (N_24593,N_23858,N_23463);
or U24594 (N_24594,N_22538,N_22785);
nand U24595 (N_24595,N_22082,N_22646);
xnor U24596 (N_24596,N_23059,N_22574);
nand U24597 (N_24597,N_23371,N_23410);
or U24598 (N_24598,N_22978,N_23232);
nor U24599 (N_24599,N_23636,N_23832);
xnor U24600 (N_24600,N_23093,N_22673);
xor U24601 (N_24601,N_22335,N_22013);
xor U24602 (N_24602,N_22923,N_22578);
nand U24603 (N_24603,N_23606,N_22686);
xnor U24604 (N_24604,N_23268,N_23996);
and U24605 (N_24605,N_22797,N_22380);
nor U24606 (N_24606,N_22992,N_22368);
nor U24607 (N_24607,N_22990,N_23016);
xnor U24608 (N_24608,N_22422,N_23329);
or U24609 (N_24609,N_22194,N_22953);
and U24610 (N_24610,N_22720,N_22035);
nor U24611 (N_24611,N_22391,N_22846);
nor U24612 (N_24612,N_23080,N_22570);
and U24613 (N_24613,N_22112,N_23658);
or U24614 (N_24614,N_22221,N_23428);
and U24615 (N_24615,N_23281,N_23892);
nor U24616 (N_24616,N_23689,N_23108);
and U24617 (N_24617,N_23273,N_22669);
xnor U24618 (N_24618,N_23474,N_23466);
nor U24619 (N_24619,N_23960,N_23838);
or U24620 (N_24620,N_23544,N_23481);
and U24621 (N_24621,N_22515,N_22984);
or U24622 (N_24622,N_23218,N_23879);
xor U24623 (N_24623,N_22808,N_23748);
and U24624 (N_24624,N_23238,N_22724);
nor U24625 (N_24625,N_22272,N_23785);
and U24626 (N_24626,N_22851,N_22658);
or U24627 (N_24627,N_22206,N_23935);
nor U24628 (N_24628,N_22454,N_22601);
nor U24629 (N_24629,N_22732,N_22831);
or U24630 (N_24630,N_22621,N_23117);
or U24631 (N_24631,N_22945,N_23983);
nand U24632 (N_24632,N_23715,N_22883);
xor U24633 (N_24633,N_23270,N_22375);
nand U24634 (N_24634,N_23612,N_22805);
nor U24635 (N_24635,N_22700,N_23552);
nand U24636 (N_24636,N_22803,N_23663);
nor U24637 (N_24637,N_22159,N_23222);
and U24638 (N_24638,N_23496,N_22497);
nand U24639 (N_24639,N_23189,N_23924);
and U24640 (N_24640,N_23694,N_23211);
nand U24641 (N_24641,N_23697,N_23400);
or U24642 (N_24642,N_23074,N_23321);
nand U24643 (N_24643,N_22937,N_22282);
and U24644 (N_24644,N_22085,N_23427);
and U24645 (N_24645,N_22773,N_22076);
or U24646 (N_24646,N_23719,N_23299);
or U24647 (N_24647,N_22440,N_22958);
nand U24648 (N_24648,N_23148,N_23866);
xnor U24649 (N_24649,N_23249,N_22762);
xor U24650 (N_24650,N_22540,N_23577);
and U24651 (N_24651,N_23319,N_22775);
nand U24652 (N_24652,N_23870,N_23526);
nand U24653 (N_24653,N_23165,N_23634);
nor U24654 (N_24654,N_22685,N_22850);
and U24655 (N_24655,N_23092,N_23229);
or U24656 (N_24656,N_23826,N_22104);
and U24657 (N_24657,N_23084,N_23881);
nor U24658 (N_24658,N_23446,N_22545);
xor U24659 (N_24659,N_23009,N_22628);
or U24660 (N_24660,N_23902,N_22910);
nand U24661 (N_24661,N_23638,N_23669);
and U24662 (N_24662,N_23340,N_22997);
and U24663 (N_24663,N_23778,N_23809);
nor U24664 (N_24664,N_22652,N_23890);
and U24665 (N_24665,N_22093,N_23227);
nand U24666 (N_24666,N_23395,N_22298);
nor U24667 (N_24667,N_23581,N_23930);
xor U24668 (N_24668,N_23489,N_23579);
nand U24669 (N_24669,N_23659,N_23622);
xnor U24670 (N_24670,N_23052,N_22668);
and U24671 (N_24671,N_23028,N_22146);
nand U24672 (N_24672,N_22925,N_22718);
and U24673 (N_24673,N_23388,N_22448);
nor U24674 (N_24674,N_22469,N_22073);
or U24675 (N_24675,N_22007,N_23708);
or U24676 (N_24676,N_23897,N_23375);
nor U24677 (N_24677,N_23471,N_23231);
nand U24678 (N_24678,N_23901,N_22676);
or U24679 (N_24679,N_23354,N_22293);
and U24680 (N_24680,N_22930,N_22898);
nand U24681 (N_24681,N_23144,N_22512);
or U24682 (N_24682,N_22018,N_23157);
and U24683 (N_24683,N_22262,N_23318);
and U24684 (N_24684,N_22881,N_23750);
nor U24685 (N_24685,N_22636,N_23880);
or U24686 (N_24686,N_22647,N_23265);
or U24687 (N_24687,N_22494,N_22532);
xnor U24688 (N_24688,N_22317,N_22895);
or U24689 (N_24689,N_22434,N_23260);
nor U24690 (N_24690,N_22807,N_23721);
xor U24691 (N_24691,N_22172,N_23646);
and U24692 (N_24692,N_23714,N_22696);
and U24693 (N_24693,N_23904,N_23303);
nand U24694 (N_24694,N_22932,N_22447);
or U24695 (N_24695,N_22207,N_23195);
nand U24696 (N_24696,N_22863,N_22451);
nor U24697 (N_24697,N_23514,N_22246);
and U24698 (N_24698,N_22764,N_23650);
nand U24699 (N_24699,N_23027,N_22373);
xnor U24700 (N_24700,N_22897,N_22100);
nor U24701 (N_24701,N_22569,N_23272);
and U24702 (N_24702,N_23698,N_23056);
nor U24703 (N_24703,N_23330,N_23347);
xnor U24704 (N_24704,N_23557,N_22961);
nand U24705 (N_24705,N_22709,N_23031);
xnor U24706 (N_24706,N_23086,N_23379);
xnor U24707 (N_24707,N_22806,N_22816);
and U24708 (N_24708,N_22586,N_23254);
and U24709 (N_24709,N_22783,N_23854);
xor U24710 (N_24710,N_23171,N_23784);
and U24711 (N_24711,N_23023,N_23672);
or U24712 (N_24712,N_23628,N_23580);
or U24713 (N_24713,N_22819,N_23569);
nor U24714 (N_24714,N_23070,N_23444);
or U24715 (N_24715,N_23576,N_23057);
xnor U24716 (N_24716,N_22227,N_22940);
xor U24717 (N_24717,N_22665,N_23055);
and U24718 (N_24718,N_22338,N_23136);
xnor U24719 (N_24719,N_23110,N_22737);
and U24720 (N_24720,N_22464,N_23071);
nand U24721 (N_24721,N_22734,N_23050);
or U24722 (N_24722,N_23546,N_23225);
nand U24723 (N_24723,N_22774,N_22362);
xor U24724 (N_24724,N_23065,N_23723);
or U24725 (N_24725,N_22674,N_23352);
nor U24726 (N_24726,N_22903,N_22606);
nand U24727 (N_24727,N_23250,N_23235);
or U24728 (N_24728,N_22098,N_23505);
nor U24729 (N_24729,N_23007,N_22449);
and U24730 (N_24730,N_23097,N_22012);
xor U24731 (N_24731,N_23536,N_23916);
nor U24732 (N_24732,N_22874,N_22657);
or U24733 (N_24733,N_22061,N_22946);
nor U24734 (N_24734,N_23677,N_23455);
and U24735 (N_24735,N_23524,N_23985);
and U24736 (N_24736,N_22701,N_22585);
and U24737 (N_24737,N_23792,N_23302);
xor U24738 (N_24738,N_23435,N_22670);
nor U24739 (N_24739,N_23132,N_22056);
or U24740 (N_24740,N_23740,N_22210);
or U24741 (N_24741,N_22218,N_23814);
or U24742 (N_24742,N_22622,N_23848);
and U24743 (N_24743,N_23256,N_22714);
or U24744 (N_24744,N_22623,N_23570);
nand U24745 (N_24745,N_22384,N_23567);
nand U24746 (N_24746,N_23458,N_23454);
nor U24747 (N_24747,N_23175,N_22690);
xnor U24748 (N_24748,N_23602,N_22157);
nand U24749 (N_24749,N_22038,N_22009);
or U24750 (N_24750,N_23377,N_22099);
or U24751 (N_24751,N_23850,N_22553);
and U24752 (N_24752,N_22849,N_23820);
and U24753 (N_24753,N_22079,N_23957);
or U24754 (N_24754,N_22450,N_23776);
nand U24755 (N_24755,N_22346,N_23263);
xnor U24756 (N_24756,N_22237,N_22838);
or U24757 (N_24757,N_23786,N_22479);
nor U24758 (N_24758,N_23621,N_23177);
and U24759 (N_24759,N_23853,N_22473);
nor U24760 (N_24760,N_22865,N_23575);
nand U24761 (N_24761,N_23887,N_22524);
nor U24762 (N_24762,N_22566,N_22379);
or U24763 (N_24763,N_23618,N_22418);
nand U24764 (N_24764,N_23934,N_23548);
or U24765 (N_24765,N_23595,N_23507);
and U24766 (N_24766,N_22033,N_23437);
nor U24767 (N_24767,N_22742,N_22220);
and U24768 (N_24768,N_23931,N_22828);
nand U24769 (N_24769,N_22991,N_23565);
or U24770 (N_24770,N_22461,N_22203);
or U24771 (N_24771,N_23193,N_22896);
nand U24772 (N_24772,N_22859,N_23817);
or U24773 (N_24773,N_22458,N_23874);
nor U24774 (N_24774,N_23806,N_23147);
or U24775 (N_24775,N_23871,N_22583);
or U24776 (N_24776,N_22161,N_23098);
and U24777 (N_24777,N_23336,N_23693);
xor U24778 (N_24778,N_22405,N_22878);
or U24779 (N_24779,N_23054,N_22145);
or U24780 (N_24780,N_22314,N_22679);
nor U24781 (N_24781,N_22312,N_22351);
xor U24782 (N_24782,N_23676,N_22366);
nand U24783 (N_24783,N_23473,N_22377);
nor U24784 (N_24784,N_22337,N_23267);
xor U24785 (N_24785,N_22793,N_23409);
xnor U24786 (N_24786,N_23022,N_23651);
xor U24787 (N_24787,N_22267,N_23030);
xnor U24788 (N_24788,N_23000,N_22492);
nor U24789 (N_24789,N_22259,N_23962);
and U24790 (N_24790,N_23230,N_22040);
nor U24791 (N_24791,N_23556,N_22189);
and U24792 (N_24792,N_23239,N_22659);
nor U24793 (N_24793,N_22124,N_23726);
or U24794 (N_24794,N_23604,N_22396);
or U24795 (N_24795,N_22660,N_23891);
or U24796 (N_24796,N_22148,N_22141);
nand U24797 (N_24797,N_23969,N_22392);
and U24798 (N_24798,N_22592,N_23083);
nor U24799 (N_24799,N_22493,N_23293);
nor U24800 (N_24800,N_22096,N_22664);
nor U24801 (N_24801,N_22561,N_22089);
xnor U24802 (N_24802,N_22310,N_23799);
and U24803 (N_24803,N_22204,N_22517);
xor U24804 (N_24804,N_23530,N_23363);
and U24805 (N_24805,N_23182,N_23605);
and U24806 (N_24806,N_23640,N_22491);
or U24807 (N_24807,N_23457,N_23034);
nand U24808 (N_24808,N_22651,N_23476);
xor U24809 (N_24809,N_22091,N_23894);
xnor U24810 (N_24810,N_23751,N_22519);
xnor U24811 (N_24811,N_22401,N_23344);
nand U24812 (N_24812,N_23152,N_22907);
or U24813 (N_24813,N_22642,N_23797);
nor U24814 (N_24814,N_23688,N_22577);
and U24815 (N_24815,N_23938,N_23197);
or U24816 (N_24816,N_22118,N_23563);
nand U24817 (N_24817,N_23495,N_23081);
or U24818 (N_24818,N_23550,N_23571);
or U24819 (N_24819,N_22198,N_23381);
or U24820 (N_24820,N_22043,N_23494);
nor U24821 (N_24821,N_22374,N_23085);
nor U24822 (N_24822,N_22140,N_23314);
and U24823 (N_24823,N_22251,N_23821);
or U24824 (N_24824,N_22804,N_22417);
nor U24825 (N_24825,N_23623,N_23064);
nand U24826 (N_24826,N_23310,N_22772);
xor U24827 (N_24827,N_23145,N_23135);
xnor U24828 (N_24828,N_23670,N_22841);
nand U24829 (N_24829,N_23562,N_22924);
or U24830 (N_24830,N_22361,N_22285);
nand U24831 (N_24831,N_22488,N_23333);
xnor U24832 (N_24832,N_22077,N_23143);
and U24833 (N_24833,N_23149,N_22102);
nor U24834 (N_24834,N_22127,N_23717);
and U24835 (N_24835,N_22900,N_22823);
xnor U24836 (N_24836,N_22209,N_22339);
nor U24837 (N_24837,N_22051,N_23408);
or U24838 (N_24838,N_22416,N_23895);
and U24839 (N_24839,N_22201,N_22886);
and U24840 (N_24840,N_22982,N_22270);
or U24841 (N_24841,N_22663,N_23590);
and U24842 (N_24842,N_23665,N_23680);
xnor U24843 (N_24843,N_22931,N_22278);
or U24844 (N_24844,N_22627,N_23248);
xnor U24845 (N_24845,N_23167,N_22581);
nand U24846 (N_24846,N_23101,N_22662);
or U24847 (N_24847,N_23014,N_23811);
xor U24848 (N_24848,N_22814,N_23133);
xnor U24849 (N_24849,N_23350,N_22121);
nor U24850 (N_24850,N_22727,N_22736);
and U24851 (N_24851,N_23704,N_22408);
xnor U24852 (N_24852,N_23755,N_23320);
nand U24853 (N_24853,N_23756,N_22967);
nand U24854 (N_24854,N_22795,N_23076);
nand U24855 (N_24855,N_23724,N_22427);
nand U24856 (N_24856,N_23475,N_23790);
nand U24857 (N_24857,N_23869,N_23899);
nor U24858 (N_24858,N_23798,N_22726);
and U24859 (N_24859,N_22913,N_23401);
xnor U24860 (N_24860,N_23341,N_23261);
nand U24861 (N_24861,N_23036,N_23124);
or U24862 (N_24862,N_23289,N_23600);
xor U24863 (N_24863,N_23311,N_22815);
xnor U24864 (N_24864,N_23378,N_23012);
or U24865 (N_24865,N_23107,N_23857);
nor U24866 (N_24866,N_23109,N_23205);
and U24867 (N_24867,N_22034,N_23979);
nor U24868 (N_24868,N_22299,N_23883);
nor U24869 (N_24869,N_22279,N_22286);
and U24870 (N_24870,N_22095,N_22119);
nor U24871 (N_24871,N_23977,N_23720);
and U24872 (N_24872,N_22675,N_22471);
and U24873 (N_24873,N_23069,N_22388);
xnor U24874 (N_24874,N_22842,N_22130);
xor U24875 (N_24875,N_23346,N_22323);
nor U24876 (N_24876,N_23335,N_22432);
or U24877 (N_24877,N_22963,N_22856);
nor U24878 (N_24878,N_22108,N_23619);
nand U24879 (N_24879,N_22733,N_23492);
xor U24880 (N_24880,N_23020,N_22884);
nor U24881 (N_24881,N_23910,N_23825);
xor U24882 (N_24882,N_22644,N_22941);
xnor U24883 (N_24883,N_23264,N_22999);
nor U24884 (N_24884,N_22631,N_23066);
and U24885 (N_24885,N_22017,N_22023);
xnor U24886 (N_24886,N_22260,N_23919);
and U24887 (N_24887,N_22735,N_23082);
nor U24888 (N_24888,N_22746,N_23603);
and U24889 (N_24889,N_22721,N_23679);
and U24890 (N_24890,N_23558,N_22389);
nand U24891 (N_24891,N_23464,N_23777);
xnor U24892 (N_24892,N_23842,N_22274);
nand U24893 (N_24893,N_23749,N_22238);
xor U24894 (N_24894,N_22325,N_22065);
or U24895 (N_24895,N_23285,N_22666);
and U24896 (N_24896,N_23068,N_23094);
xnor U24897 (N_24897,N_22939,N_22334);
nand U24898 (N_24898,N_23240,N_22294);
nor U24899 (N_24899,N_23450,N_22852);
and U24900 (N_24900,N_22791,N_22261);
or U24901 (N_24901,N_22501,N_23903);
nand U24902 (N_24902,N_23648,N_22861);
and U24903 (N_24903,N_23574,N_23599);
and U24904 (N_24904,N_23185,N_22697);
nor U24905 (N_24905,N_22811,N_22438);
xnor U24906 (N_24906,N_23582,N_22589);
and U24907 (N_24907,N_22637,N_23161);
xnor U24908 (N_24908,N_23173,N_22810);
nand U24909 (N_24909,N_22350,N_23188);
nand U24910 (N_24910,N_22139,N_23994);
nand U24911 (N_24911,N_23115,N_22834);
and U24912 (N_24912,N_22717,N_22568);
or U24913 (N_24913,N_22103,N_23198);
or U24914 (N_24914,N_22905,N_23483);
nand U24915 (N_24915,N_23923,N_22694);
or U24916 (N_24916,N_22730,N_22428);
xnor U24917 (N_24917,N_22509,N_22909);
or U24918 (N_24918,N_22514,N_22230);
xnor U24919 (N_24919,N_22297,N_23896);
or U24920 (N_24920,N_23767,N_23125);
or U24921 (N_24921,N_22305,N_23296);
nor U24922 (N_24922,N_22016,N_22769);
xor U24923 (N_24923,N_23184,N_22423);
and U24924 (N_24924,N_22276,N_23442);
nand U24925 (N_24925,N_23898,N_23043);
nand U24926 (N_24926,N_23893,N_23545);
nor U24927 (N_24927,N_22475,N_22166);
and U24928 (N_24928,N_23911,N_22575);
nand U24929 (N_24929,N_22344,N_23687);
xor U24930 (N_24930,N_22555,N_22291);
xnor U24931 (N_24931,N_23228,N_22106);
nand U24932 (N_24932,N_23269,N_23368);
nor U24933 (N_24933,N_22739,N_22352);
nand U24934 (N_24934,N_22779,N_22211);
or U24935 (N_24935,N_23501,N_22486);
nor U24936 (N_24936,N_23312,N_22986);
nand U24937 (N_24937,N_22047,N_23843);
nand U24938 (N_24938,N_23208,N_23541);
nor U24939 (N_24939,N_22044,N_22744);
nand U24940 (N_24940,N_23146,N_22653);
and U24941 (N_24941,N_22223,N_22254);
and U24942 (N_24942,N_23928,N_22957);
or U24943 (N_24943,N_23308,N_23315);
and U24944 (N_24944,N_23949,N_22848);
nand U24945 (N_24945,N_22055,N_22460);
or U24946 (N_24946,N_22386,N_23259);
or U24947 (N_24947,N_22326,N_22508);
xor U24948 (N_24948,N_22199,N_23440);
nand U24949 (N_24949,N_22549,N_22421);
nand U24950 (N_24950,N_23878,N_23649);
nand U24951 (N_24951,N_22699,N_22536);
or U24952 (N_24952,N_22182,N_23549);
nor U24953 (N_24953,N_22107,N_23905);
xnor U24954 (N_24954,N_23733,N_22949);
xnor U24955 (N_24955,N_23754,N_23200);
and U24956 (N_24956,N_22426,N_23313);
or U24957 (N_24957,N_23551,N_23978);
and U24958 (N_24958,N_22437,N_23480);
and U24959 (N_24959,N_22214,N_22152);
nand U24960 (N_24960,N_23389,N_23449);
and U24961 (N_24961,N_22767,N_23355);
and U24962 (N_24962,N_22292,N_23803);
and U24963 (N_24963,N_23506,N_22360);
nor U24964 (N_24964,N_23357,N_23073);
or U24965 (N_24965,N_23203,N_22780);
or U24966 (N_24966,N_22521,N_23813);
nand U24967 (N_24967,N_23538,N_23467);
nor U24968 (N_24968,N_22466,N_23174);
nand U24969 (N_24969,N_22030,N_23627);
nand U24970 (N_24970,N_23642,N_23561);
nand U24971 (N_24971,N_23829,N_23190);
or U24972 (N_24972,N_22078,N_23553);
nand U24973 (N_24973,N_22320,N_23764);
or U24974 (N_24974,N_22693,N_22832);
nand U24975 (N_24975,N_22576,N_23839);
or U24976 (N_24976,N_23830,N_22074);
or U24977 (N_24977,N_23753,N_23438);
and U24978 (N_24978,N_23654,N_22250);
nor U24979 (N_24979,N_22537,N_22942);
or U24980 (N_24980,N_23490,N_22887);
and U24981 (N_24981,N_22817,N_22534);
or U24982 (N_24982,N_22551,N_23040);
nor U24983 (N_24983,N_23212,N_22629);
nor U24984 (N_24984,N_22399,N_22241);
or U24985 (N_24985,N_22216,N_22289);
nand U24986 (N_24986,N_22163,N_23508);
or U24987 (N_24987,N_23522,N_22598);
and U24988 (N_24988,N_22208,N_23706);
nor U24989 (N_24989,N_23547,N_23914);
or U24990 (N_24990,N_23711,N_23584);
nand U24991 (N_24991,N_23986,N_23331);
nand U24992 (N_24992,N_22459,N_23765);
xor U24993 (N_24993,N_23078,N_23499);
or U24994 (N_24994,N_22641,N_23770);
and U24995 (N_24995,N_22263,N_22280);
and U24996 (N_24996,N_23675,N_22864);
nor U24997 (N_24997,N_23611,N_22616);
nand U24998 (N_24998,N_23439,N_22478);
and U24999 (N_24999,N_22385,N_23397);
and U25000 (N_25000,N_23826,N_23092);
or U25001 (N_25001,N_22009,N_23064);
nor U25002 (N_25002,N_23222,N_23268);
nand U25003 (N_25003,N_23841,N_22953);
and U25004 (N_25004,N_22831,N_22798);
nor U25005 (N_25005,N_22117,N_23977);
xnor U25006 (N_25006,N_23224,N_23463);
nand U25007 (N_25007,N_22145,N_23217);
nor U25008 (N_25008,N_22780,N_23582);
nand U25009 (N_25009,N_23927,N_22081);
and U25010 (N_25010,N_23907,N_22706);
xnor U25011 (N_25011,N_23224,N_22544);
xor U25012 (N_25012,N_22391,N_23939);
and U25013 (N_25013,N_22156,N_23537);
or U25014 (N_25014,N_22996,N_23161);
or U25015 (N_25015,N_22540,N_23247);
and U25016 (N_25016,N_23761,N_22823);
nor U25017 (N_25017,N_22718,N_22147);
and U25018 (N_25018,N_22149,N_22467);
xnor U25019 (N_25019,N_23683,N_22923);
nor U25020 (N_25020,N_22211,N_22551);
and U25021 (N_25021,N_22937,N_23700);
nand U25022 (N_25022,N_22700,N_23132);
or U25023 (N_25023,N_23404,N_23147);
xnor U25024 (N_25024,N_22640,N_22755);
and U25025 (N_25025,N_22200,N_23499);
nor U25026 (N_25026,N_23020,N_23988);
nor U25027 (N_25027,N_22962,N_22536);
and U25028 (N_25028,N_22895,N_23158);
nand U25029 (N_25029,N_23737,N_23842);
or U25030 (N_25030,N_22669,N_23180);
nor U25031 (N_25031,N_23878,N_23056);
xor U25032 (N_25032,N_23569,N_22774);
nand U25033 (N_25033,N_22494,N_22063);
xor U25034 (N_25034,N_22147,N_22520);
nand U25035 (N_25035,N_22842,N_22414);
or U25036 (N_25036,N_23046,N_22226);
nor U25037 (N_25037,N_22513,N_23461);
and U25038 (N_25038,N_23749,N_22826);
nor U25039 (N_25039,N_22654,N_23409);
nor U25040 (N_25040,N_22909,N_22571);
nand U25041 (N_25041,N_22409,N_22122);
nor U25042 (N_25042,N_23092,N_22328);
or U25043 (N_25043,N_22133,N_22234);
nor U25044 (N_25044,N_23448,N_22659);
xnor U25045 (N_25045,N_23484,N_22911);
xor U25046 (N_25046,N_23978,N_23255);
or U25047 (N_25047,N_22592,N_23308);
and U25048 (N_25048,N_22867,N_23458);
nand U25049 (N_25049,N_22134,N_22689);
xnor U25050 (N_25050,N_22833,N_22868);
and U25051 (N_25051,N_22971,N_23891);
xnor U25052 (N_25052,N_23667,N_22769);
nor U25053 (N_25053,N_23672,N_22048);
nand U25054 (N_25054,N_23415,N_22780);
and U25055 (N_25055,N_23846,N_22958);
xnor U25056 (N_25056,N_22102,N_23407);
and U25057 (N_25057,N_22078,N_22768);
nand U25058 (N_25058,N_23821,N_22460);
and U25059 (N_25059,N_23061,N_23430);
nand U25060 (N_25060,N_23705,N_22005);
nand U25061 (N_25061,N_23642,N_22153);
nor U25062 (N_25062,N_22481,N_22137);
and U25063 (N_25063,N_23037,N_22975);
xnor U25064 (N_25064,N_23497,N_23428);
and U25065 (N_25065,N_23807,N_22178);
and U25066 (N_25066,N_22311,N_23977);
xnor U25067 (N_25067,N_22055,N_23112);
nand U25068 (N_25068,N_23068,N_23723);
nor U25069 (N_25069,N_23098,N_23563);
or U25070 (N_25070,N_22027,N_22721);
nand U25071 (N_25071,N_22417,N_23408);
nor U25072 (N_25072,N_22191,N_23986);
nor U25073 (N_25073,N_23804,N_23584);
nor U25074 (N_25074,N_22652,N_23864);
nand U25075 (N_25075,N_22952,N_23207);
nand U25076 (N_25076,N_23398,N_23679);
or U25077 (N_25077,N_23475,N_22557);
nor U25078 (N_25078,N_22799,N_23509);
or U25079 (N_25079,N_23179,N_22676);
nor U25080 (N_25080,N_23617,N_23177);
and U25081 (N_25081,N_22523,N_22340);
or U25082 (N_25082,N_22142,N_23498);
or U25083 (N_25083,N_22608,N_22531);
or U25084 (N_25084,N_22340,N_22243);
nor U25085 (N_25085,N_23743,N_22215);
xor U25086 (N_25086,N_23730,N_23883);
and U25087 (N_25087,N_23399,N_22274);
and U25088 (N_25088,N_23776,N_22497);
xnor U25089 (N_25089,N_22016,N_23215);
xor U25090 (N_25090,N_23893,N_23666);
xor U25091 (N_25091,N_23868,N_22016);
xor U25092 (N_25092,N_22310,N_23472);
or U25093 (N_25093,N_23726,N_22764);
nand U25094 (N_25094,N_23478,N_23602);
and U25095 (N_25095,N_22951,N_23168);
and U25096 (N_25096,N_23126,N_22474);
nand U25097 (N_25097,N_23957,N_22572);
nand U25098 (N_25098,N_23042,N_23961);
xor U25099 (N_25099,N_23833,N_22447);
nor U25100 (N_25100,N_23845,N_23663);
xor U25101 (N_25101,N_23517,N_22742);
nor U25102 (N_25102,N_22214,N_22992);
xnor U25103 (N_25103,N_23779,N_22900);
and U25104 (N_25104,N_22589,N_22547);
and U25105 (N_25105,N_22670,N_22733);
or U25106 (N_25106,N_23433,N_23206);
and U25107 (N_25107,N_22916,N_23700);
and U25108 (N_25108,N_23499,N_23112);
or U25109 (N_25109,N_22857,N_22310);
nand U25110 (N_25110,N_22419,N_23804);
xor U25111 (N_25111,N_22109,N_23234);
nor U25112 (N_25112,N_23687,N_23928);
and U25113 (N_25113,N_23235,N_22027);
or U25114 (N_25114,N_23034,N_23325);
nor U25115 (N_25115,N_22426,N_22324);
and U25116 (N_25116,N_22063,N_22932);
or U25117 (N_25117,N_22468,N_22513);
and U25118 (N_25118,N_22830,N_22952);
nor U25119 (N_25119,N_22764,N_22584);
and U25120 (N_25120,N_23248,N_23074);
and U25121 (N_25121,N_22731,N_22984);
and U25122 (N_25122,N_22854,N_22434);
or U25123 (N_25123,N_22525,N_22889);
and U25124 (N_25124,N_22335,N_22508);
nor U25125 (N_25125,N_23693,N_23281);
or U25126 (N_25126,N_22452,N_22223);
or U25127 (N_25127,N_22113,N_23067);
or U25128 (N_25128,N_22336,N_22992);
nand U25129 (N_25129,N_23276,N_22507);
or U25130 (N_25130,N_23811,N_23648);
and U25131 (N_25131,N_23643,N_23412);
or U25132 (N_25132,N_23888,N_23186);
and U25133 (N_25133,N_22985,N_22632);
and U25134 (N_25134,N_23730,N_23680);
nor U25135 (N_25135,N_23919,N_23094);
xor U25136 (N_25136,N_23828,N_22275);
xnor U25137 (N_25137,N_23070,N_23762);
and U25138 (N_25138,N_22498,N_22674);
nand U25139 (N_25139,N_22063,N_23619);
or U25140 (N_25140,N_22166,N_22696);
xnor U25141 (N_25141,N_22842,N_23590);
or U25142 (N_25142,N_23834,N_23749);
nand U25143 (N_25143,N_22601,N_23120);
nor U25144 (N_25144,N_22419,N_22816);
nor U25145 (N_25145,N_23972,N_23756);
or U25146 (N_25146,N_23833,N_23604);
and U25147 (N_25147,N_23070,N_22895);
nor U25148 (N_25148,N_22619,N_22546);
xor U25149 (N_25149,N_23827,N_23451);
and U25150 (N_25150,N_22490,N_23846);
and U25151 (N_25151,N_23386,N_23785);
nand U25152 (N_25152,N_22351,N_23121);
xnor U25153 (N_25153,N_23960,N_23335);
xor U25154 (N_25154,N_22122,N_23331);
nor U25155 (N_25155,N_23809,N_23326);
and U25156 (N_25156,N_22807,N_22149);
and U25157 (N_25157,N_23164,N_23214);
nand U25158 (N_25158,N_23438,N_22357);
and U25159 (N_25159,N_23369,N_23719);
nand U25160 (N_25160,N_22258,N_22570);
or U25161 (N_25161,N_23917,N_22584);
or U25162 (N_25162,N_22185,N_22191);
or U25163 (N_25163,N_22650,N_23534);
nand U25164 (N_25164,N_23386,N_23917);
or U25165 (N_25165,N_23629,N_23720);
xnor U25166 (N_25166,N_23817,N_22443);
or U25167 (N_25167,N_23465,N_22763);
xor U25168 (N_25168,N_22246,N_22101);
and U25169 (N_25169,N_23883,N_22778);
and U25170 (N_25170,N_22711,N_22323);
nand U25171 (N_25171,N_22694,N_23320);
or U25172 (N_25172,N_23641,N_23248);
nor U25173 (N_25173,N_22038,N_22153);
or U25174 (N_25174,N_23520,N_23359);
xnor U25175 (N_25175,N_23329,N_22207);
nor U25176 (N_25176,N_23259,N_22458);
nand U25177 (N_25177,N_22299,N_22032);
nand U25178 (N_25178,N_22256,N_23250);
and U25179 (N_25179,N_23321,N_23186);
xnor U25180 (N_25180,N_23006,N_22696);
or U25181 (N_25181,N_22622,N_22235);
nor U25182 (N_25182,N_23297,N_22490);
and U25183 (N_25183,N_23204,N_22212);
and U25184 (N_25184,N_22904,N_23007);
xnor U25185 (N_25185,N_22523,N_22675);
nor U25186 (N_25186,N_23301,N_22430);
nand U25187 (N_25187,N_22277,N_22181);
and U25188 (N_25188,N_22611,N_22895);
nor U25189 (N_25189,N_23428,N_23286);
xor U25190 (N_25190,N_23780,N_22470);
nor U25191 (N_25191,N_22681,N_23614);
or U25192 (N_25192,N_23018,N_23512);
nand U25193 (N_25193,N_22759,N_23066);
nor U25194 (N_25194,N_23482,N_22407);
nor U25195 (N_25195,N_22175,N_22829);
nand U25196 (N_25196,N_23131,N_22969);
and U25197 (N_25197,N_22211,N_22472);
and U25198 (N_25198,N_23003,N_23228);
nand U25199 (N_25199,N_23649,N_23725);
or U25200 (N_25200,N_23223,N_23935);
nor U25201 (N_25201,N_23109,N_23293);
nor U25202 (N_25202,N_22963,N_22585);
xnor U25203 (N_25203,N_22422,N_23758);
nand U25204 (N_25204,N_23948,N_23190);
nor U25205 (N_25205,N_23464,N_22280);
or U25206 (N_25206,N_22434,N_22341);
nand U25207 (N_25207,N_23326,N_23335);
and U25208 (N_25208,N_23768,N_23372);
nor U25209 (N_25209,N_22001,N_22370);
or U25210 (N_25210,N_22063,N_22025);
xnor U25211 (N_25211,N_23479,N_22055);
or U25212 (N_25212,N_22185,N_23512);
and U25213 (N_25213,N_22098,N_23155);
and U25214 (N_25214,N_22689,N_22007);
nand U25215 (N_25215,N_22640,N_22340);
and U25216 (N_25216,N_23580,N_22495);
xnor U25217 (N_25217,N_22187,N_23980);
or U25218 (N_25218,N_22865,N_22116);
and U25219 (N_25219,N_22847,N_23580);
and U25220 (N_25220,N_22145,N_22041);
and U25221 (N_25221,N_23101,N_23070);
nand U25222 (N_25222,N_23843,N_22452);
nand U25223 (N_25223,N_23023,N_22478);
and U25224 (N_25224,N_22781,N_22540);
and U25225 (N_25225,N_23755,N_23355);
nand U25226 (N_25226,N_23169,N_23654);
nand U25227 (N_25227,N_22009,N_23409);
xor U25228 (N_25228,N_23928,N_22236);
and U25229 (N_25229,N_23252,N_23639);
or U25230 (N_25230,N_22180,N_23500);
nor U25231 (N_25231,N_23438,N_22593);
nand U25232 (N_25232,N_23608,N_23585);
xor U25233 (N_25233,N_22708,N_23482);
nand U25234 (N_25234,N_23637,N_23434);
xnor U25235 (N_25235,N_22046,N_23489);
nand U25236 (N_25236,N_23171,N_23793);
xnor U25237 (N_25237,N_22008,N_23557);
nand U25238 (N_25238,N_22111,N_23849);
nor U25239 (N_25239,N_22359,N_22207);
and U25240 (N_25240,N_22334,N_22446);
and U25241 (N_25241,N_22526,N_22290);
nor U25242 (N_25242,N_22629,N_23163);
and U25243 (N_25243,N_23004,N_22923);
xnor U25244 (N_25244,N_22339,N_23334);
nor U25245 (N_25245,N_23905,N_22270);
or U25246 (N_25246,N_23108,N_22297);
or U25247 (N_25247,N_23503,N_23023);
or U25248 (N_25248,N_22349,N_23779);
and U25249 (N_25249,N_23919,N_22244);
or U25250 (N_25250,N_23990,N_22812);
and U25251 (N_25251,N_22206,N_23027);
and U25252 (N_25252,N_22917,N_23273);
nor U25253 (N_25253,N_22184,N_22043);
nand U25254 (N_25254,N_22956,N_22226);
or U25255 (N_25255,N_23827,N_22306);
xor U25256 (N_25256,N_23226,N_23483);
and U25257 (N_25257,N_22464,N_23050);
nand U25258 (N_25258,N_22868,N_22158);
nand U25259 (N_25259,N_22378,N_23297);
and U25260 (N_25260,N_22962,N_22649);
xor U25261 (N_25261,N_23148,N_23273);
or U25262 (N_25262,N_23209,N_22832);
nand U25263 (N_25263,N_22136,N_23355);
nand U25264 (N_25264,N_22709,N_22933);
nand U25265 (N_25265,N_22543,N_22616);
nor U25266 (N_25266,N_22759,N_22637);
nand U25267 (N_25267,N_23640,N_22798);
nand U25268 (N_25268,N_22833,N_23632);
nor U25269 (N_25269,N_22855,N_23011);
and U25270 (N_25270,N_23867,N_23163);
xnor U25271 (N_25271,N_22597,N_22909);
and U25272 (N_25272,N_23997,N_22973);
xor U25273 (N_25273,N_22728,N_23962);
nor U25274 (N_25274,N_22520,N_23756);
and U25275 (N_25275,N_22525,N_23502);
and U25276 (N_25276,N_23953,N_23177);
or U25277 (N_25277,N_23449,N_23274);
or U25278 (N_25278,N_23713,N_22838);
or U25279 (N_25279,N_23374,N_23471);
xor U25280 (N_25280,N_23370,N_22762);
nor U25281 (N_25281,N_22583,N_22614);
xnor U25282 (N_25282,N_22275,N_23855);
and U25283 (N_25283,N_23492,N_22255);
nand U25284 (N_25284,N_23178,N_23870);
nor U25285 (N_25285,N_22458,N_23547);
xor U25286 (N_25286,N_23340,N_22686);
nand U25287 (N_25287,N_22377,N_22003);
xor U25288 (N_25288,N_22578,N_22514);
nand U25289 (N_25289,N_23043,N_23969);
nand U25290 (N_25290,N_23367,N_22836);
xor U25291 (N_25291,N_22291,N_23155);
or U25292 (N_25292,N_22533,N_22949);
nand U25293 (N_25293,N_22902,N_23651);
xnor U25294 (N_25294,N_22089,N_23831);
nor U25295 (N_25295,N_23463,N_23179);
nand U25296 (N_25296,N_23174,N_22855);
xor U25297 (N_25297,N_23036,N_22751);
xor U25298 (N_25298,N_22538,N_23702);
nor U25299 (N_25299,N_22964,N_22760);
nor U25300 (N_25300,N_22580,N_22986);
nor U25301 (N_25301,N_23457,N_23479);
or U25302 (N_25302,N_23652,N_23690);
nor U25303 (N_25303,N_22836,N_22741);
nor U25304 (N_25304,N_22983,N_23108);
nor U25305 (N_25305,N_23750,N_22398);
and U25306 (N_25306,N_22716,N_23465);
and U25307 (N_25307,N_23075,N_23052);
nand U25308 (N_25308,N_22828,N_22055);
nor U25309 (N_25309,N_23336,N_23816);
xor U25310 (N_25310,N_23560,N_23608);
or U25311 (N_25311,N_23994,N_22255);
xor U25312 (N_25312,N_22975,N_23630);
or U25313 (N_25313,N_22951,N_23627);
and U25314 (N_25314,N_22459,N_23410);
or U25315 (N_25315,N_23451,N_22998);
nand U25316 (N_25316,N_23040,N_22431);
nand U25317 (N_25317,N_23978,N_23110);
xnor U25318 (N_25318,N_22619,N_22413);
or U25319 (N_25319,N_23685,N_23016);
nor U25320 (N_25320,N_22571,N_22821);
and U25321 (N_25321,N_23390,N_22044);
nand U25322 (N_25322,N_22792,N_23231);
or U25323 (N_25323,N_22734,N_23125);
nor U25324 (N_25324,N_23880,N_22669);
and U25325 (N_25325,N_22620,N_23399);
nor U25326 (N_25326,N_22186,N_22664);
nand U25327 (N_25327,N_23975,N_22859);
and U25328 (N_25328,N_23384,N_22050);
and U25329 (N_25329,N_22328,N_22541);
xnor U25330 (N_25330,N_23221,N_22856);
and U25331 (N_25331,N_23130,N_23385);
nor U25332 (N_25332,N_23167,N_22735);
xor U25333 (N_25333,N_23297,N_23686);
xnor U25334 (N_25334,N_22489,N_22922);
nor U25335 (N_25335,N_22579,N_23901);
nand U25336 (N_25336,N_22286,N_22596);
nor U25337 (N_25337,N_23308,N_23052);
and U25338 (N_25338,N_22148,N_23655);
nor U25339 (N_25339,N_22843,N_22185);
or U25340 (N_25340,N_23614,N_22365);
and U25341 (N_25341,N_23013,N_23909);
xnor U25342 (N_25342,N_23024,N_23542);
and U25343 (N_25343,N_22879,N_23598);
nor U25344 (N_25344,N_23404,N_23311);
nor U25345 (N_25345,N_22857,N_23156);
or U25346 (N_25346,N_23689,N_23815);
nand U25347 (N_25347,N_23821,N_23787);
and U25348 (N_25348,N_23221,N_23899);
and U25349 (N_25349,N_22064,N_22982);
xnor U25350 (N_25350,N_23410,N_22366);
or U25351 (N_25351,N_23380,N_22385);
xnor U25352 (N_25352,N_22864,N_22296);
or U25353 (N_25353,N_22247,N_23527);
nor U25354 (N_25354,N_22593,N_22068);
and U25355 (N_25355,N_22996,N_22096);
xnor U25356 (N_25356,N_22540,N_23482);
or U25357 (N_25357,N_22552,N_23582);
and U25358 (N_25358,N_23300,N_23783);
or U25359 (N_25359,N_23445,N_23999);
nand U25360 (N_25360,N_22389,N_23227);
nor U25361 (N_25361,N_22742,N_23648);
nor U25362 (N_25362,N_22709,N_22785);
nor U25363 (N_25363,N_23500,N_23764);
or U25364 (N_25364,N_23217,N_22322);
nand U25365 (N_25365,N_22062,N_23368);
or U25366 (N_25366,N_22513,N_22297);
and U25367 (N_25367,N_22882,N_23585);
or U25368 (N_25368,N_22922,N_22638);
nor U25369 (N_25369,N_22963,N_23176);
nand U25370 (N_25370,N_22837,N_22728);
and U25371 (N_25371,N_23955,N_23950);
xnor U25372 (N_25372,N_23945,N_23138);
nand U25373 (N_25373,N_23787,N_22089);
nor U25374 (N_25374,N_22112,N_23670);
nor U25375 (N_25375,N_22184,N_22348);
and U25376 (N_25376,N_23667,N_22467);
or U25377 (N_25377,N_22383,N_22170);
nand U25378 (N_25378,N_23522,N_23862);
or U25379 (N_25379,N_23126,N_22133);
nor U25380 (N_25380,N_22344,N_22094);
nand U25381 (N_25381,N_22609,N_23219);
nor U25382 (N_25382,N_23043,N_22909);
nor U25383 (N_25383,N_22523,N_23940);
nor U25384 (N_25384,N_23747,N_23192);
nor U25385 (N_25385,N_23955,N_23538);
and U25386 (N_25386,N_23990,N_23674);
or U25387 (N_25387,N_22627,N_22133);
xnor U25388 (N_25388,N_23810,N_23274);
xor U25389 (N_25389,N_22846,N_23369);
and U25390 (N_25390,N_22989,N_22113);
and U25391 (N_25391,N_22901,N_22403);
and U25392 (N_25392,N_22910,N_23164);
xor U25393 (N_25393,N_22054,N_22698);
xnor U25394 (N_25394,N_22589,N_23737);
or U25395 (N_25395,N_23564,N_22137);
xnor U25396 (N_25396,N_22964,N_22020);
xnor U25397 (N_25397,N_22930,N_23912);
and U25398 (N_25398,N_22365,N_23187);
nand U25399 (N_25399,N_22658,N_22627);
nor U25400 (N_25400,N_23517,N_22913);
nand U25401 (N_25401,N_22158,N_22933);
xnor U25402 (N_25402,N_22255,N_23507);
xnor U25403 (N_25403,N_22307,N_22978);
and U25404 (N_25404,N_23075,N_23796);
and U25405 (N_25405,N_22045,N_23654);
or U25406 (N_25406,N_23441,N_23099);
and U25407 (N_25407,N_23134,N_22598);
and U25408 (N_25408,N_23151,N_23287);
and U25409 (N_25409,N_22620,N_22039);
nor U25410 (N_25410,N_22421,N_23881);
or U25411 (N_25411,N_23064,N_23630);
nor U25412 (N_25412,N_23610,N_23729);
nand U25413 (N_25413,N_23394,N_23389);
nand U25414 (N_25414,N_23201,N_23681);
xnor U25415 (N_25415,N_23921,N_22792);
xnor U25416 (N_25416,N_23776,N_23984);
nor U25417 (N_25417,N_22322,N_23783);
and U25418 (N_25418,N_23473,N_22510);
or U25419 (N_25419,N_23026,N_23948);
xor U25420 (N_25420,N_22719,N_22363);
xor U25421 (N_25421,N_22509,N_22588);
or U25422 (N_25422,N_22166,N_22717);
and U25423 (N_25423,N_23054,N_22157);
or U25424 (N_25424,N_22793,N_23947);
and U25425 (N_25425,N_23287,N_23828);
xor U25426 (N_25426,N_22499,N_23920);
or U25427 (N_25427,N_22832,N_23530);
nand U25428 (N_25428,N_22951,N_23550);
and U25429 (N_25429,N_22267,N_23247);
xor U25430 (N_25430,N_22669,N_22969);
nand U25431 (N_25431,N_22388,N_23395);
xnor U25432 (N_25432,N_22376,N_23549);
and U25433 (N_25433,N_23289,N_22304);
and U25434 (N_25434,N_23028,N_23949);
or U25435 (N_25435,N_22058,N_22187);
and U25436 (N_25436,N_22804,N_23132);
nand U25437 (N_25437,N_22069,N_22088);
xor U25438 (N_25438,N_22082,N_23552);
and U25439 (N_25439,N_22046,N_23830);
nand U25440 (N_25440,N_22946,N_22797);
xnor U25441 (N_25441,N_23036,N_23632);
xor U25442 (N_25442,N_23529,N_22666);
xnor U25443 (N_25443,N_22425,N_23012);
nand U25444 (N_25444,N_23016,N_23463);
and U25445 (N_25445,N_23827,N_22771);
and U25446 (N_25446,N_23800,N_23903);
nand U25447 (N_25447,N_23221,N_22994);
nand U25448 (N_25448,N_22073,N_22782);
xor U25449 (N_25449,N_23205,N_22126);
or U25450 (N_25450,N_23579,N_22488);
nor U25451 (N_25451,N_22650,N_23702);
or U25452 (N_25452,N_22691,N_23530);
nor U25453 (N_25453,N_22927,N_23316);
nand U25454 (N_25454,N_23170,N_22931);
xor U25455 (N_25455,N_22401,N_23115);
xor U25456 (N_25456,N_23271,N_23401);
nor U25457 (N_25457,N_22382,N_23563);
nor U25458 (N_25458,N_23805,N_22563);
xor U25459 (N_25459,N_22917,N_23146);
xnor U25460 (N_25460,N_22874,N_22082);
xor U25461 (N_25461,N_23324,N_23267);
and U25462 (N_25462,N_22869,N_22510);
nand U25463 (N_25463,N_23316,N_23689);
nor U25464 (N_25464,N_23729,N_23549);
nor U25465 (N_25465,N_22794,N_23166);
and U25466 (N_25466,N_23462,N_23302);
or U25467 (N_25467,N_22300,N_22613);
xor U25468 (N_25468,N_23804,N_22856);
or U25469 (N_25469,N_23889,N_22233);
and U25470 (N_25470,N_22741,N_23617);
xor U25471 (N_25471,N_22511,N_23509);
nor U25472 (N_25472,N_22415,N_23800);
nor U25473 (N_25473,N_23950,N_22243);
nor U25474 (N_25474,N_23356,N_23058);
or U25475 (N_25475,N_23344,N_22188);
and U25476 (N_25476,N_22629,N_23230);
xnor U25477 (N_25477,N_23842,N_23237);
nand U25478 (N_25478,N_22550,N_23724);
nand U25479 (N_25479,N_23098,N_23606);
nand U25480 (N_25480,N_22672,N_23781);
and U25481 (N_25481,N_23960,N_23581);
nand U25482 (N_25482,N_22525,N_23281);
nand U25483 (N_25483,N_22612,N_22118);
xor U25484 (N_25484,N_23282,N_22666);
nand U25485 (N_25485,N_23002,N_22045);
xnor U25486 (N_25486,N_23441,N_23423);
xnor U25487 (N_25487,N_22590,N_23393);
nor U25488 (N_25488,N_22399,N_23251);
or U25489 (N_25489,N_22816,N_23973);
nor U25490 (N_25490,N_23179,N_23553);
nor U25491 (N_25491,N_22331,N_22295);
and U25492 (N_25492,N_23154,N_22456);
or U25493 (N_25493,N_22316,N_22048);
xor U25494 (N_25494,N_23205,N_22393);
or U25495 (N_25495,N_22135,N_22073);
nor U25496 (N_25496,N_23788,N_23219);
or U25497 (N_25497,N_22238,N_22718);
nor U25498 (N_25498,N_23013,N_22771);
xor U25499 (N_25499,N_23188,N_23835);
xor U25500 (N_25500,N_22054,N_22562);
nor U25501 (N_25501,N_23204,N_22650);
or U25502 (N_25502,N_23063,N_22881);
nand U25503 (N_25503,N_23900,N_22578);
or U25504 (N_25504,N_23948,N_23465);
or U25505 (N_25505,N_23494,N_22963);
or U25506 (N_25506,N_23871,N_22293);
nor U25507 (N_25507,N_23163,N_22821);
or U25508 (N_25508,N_22047,N_22690);
or U25509 (N_25509,N_23399,N_23780);
xor U25510 (N_25510,N_22582,N_23921);
or U25511 (N_25511,N_22055,N_22130);
or U25512 (N_25512,N_22357,N_22601);
xor U25513 (N_25513,N_23729,N_22391);
and U25514 (N_25514,N_23984,N_23508);
nor U25515 (N_25515,N_22980,N_22647);
and U25516 (N_25516,N_23615,N_23175);
nand U25517 (N_25517,N_23275,N_23133);
nor U25518 (N_25518,N_23465,N_22868);
xnor U25519 (N_25519,N_22753,N_23014);
or U25520 (N_25520,N_23591,N_23280);
and U25521 (N_25521,N_22714,N_22581);
and U25522 (N_25522,N_23076,N_23634);
or U25523 (N_25523,N_22195,N_22092);
xnor U25524 (N_25524,N_23836,N_22345);
nand U25525 (N_25525,N_23270,N_23813);
and U25526 (N_25526,N_23138,N_22773);
nor U25527 (N_25527,N_23133,N_22746);
nand U25528 (N_25528,N_22582,N_23999);
nor U25529 (N_25529,N_22811,N_23296);
and U25530 (N_25530,N_22942,N_23999);
or U25531 (N_25531,N_22705,N_23995);
nor U25532 (N_25532,N_23767,N_23499);
nor U25533 (N_25533,N_23355,N_23126);
nor U25534 (N_25534,N_23005,N_23573);
nand U25535 (N_25535,N_23123,N_22361);
nand U25536 (N_25536,N_23703,N_22955);
and U25537 (N_25537,N_22092,N_22488);
or U25538 (N_25538,N_22161,N_23533);
and U25539 (N_25539,N_23081,N_23370);
xnor U25540 (N_25540,N_22043,N_22472);
nor U25541 (N_25541,N_23316,N_22531);
nor U25542 (N_25542,N_22062,N_23113);
nor U25543 (N_25543,N_23542,N_22475);
nor U25544 (N_25544,N_23169,N_23168);
or U25545 (N_25545,N_23846,N_22265);
xor U25546 (N_25546,N_22751,N_22101);
or U25547 (N_25547,N_23496,N_23105);
nand U25548 (N_25548,N_23447,N_23825);
nand U25549 (N_25549,N_23171,N_22663);
or U25550 (N_25550,N_22862,N_23663);
xnor U25551 (N_25551,N_23613,N_23375);
and U25552 (N_25552,N_23686,N_22656);
xor U25553 (N_25553,N_22301,N_22883);
xnor U25554 (N_25554,N_22385,N_22550);
xor U25555 (N_25555,N_23054,N_23923);
or U25556 (N_25556,N_22032,N_22974);
nor U25557 (N_25557,N_22701,N_23011);
xnor U25558 (N_25558,N_23448,N_22868);
nand U25559 (N_25559,N_22215,N_23376);
nor U25560 (N_25560,N_22018,N_23643);
nand U25561 (N_25561,N_22993,N_23516);
and U25562 (N_25562,N_23134,N_22050);
xor U25563 (N_25563,N_23757,N_22348);
and U25564 (N_25564,N_23493,N_22265);
and U25565 (N_25565,N_23321,N_23088);
xnor U25566 (N_25566,N_22625,N_23309);
xor U25567 (N_25567,N_23255,N_22729);
and U25568 (N_25568,N_22488,N_23925);
nor U25569 (N_25569,N_23146,N_22280);
and U25570 (N_25570,N_22897,N_22478);
xor U25571 (N_25571,N_22931,N_23585);
xor U25572 (N_25572,N_23260,N_23016);
or U25573 (N_25573,N_22767,N_23063);
and U25574 (N_25574,N_22111,N_23223);
nand U25575 (N_25575,N_23607,N_22077);
or U25576 (N_25576,N_22591,N_22201);
or U25577 (N_25577,N_22041,N_23720);
nor U25578 (N_25578,N_23947,N_22731);
nand U25579 (N_25579,N_22799,N_23488);
nor U25580 (N_25580,N_22594,N_22854);
nand U25581 (N_25581,N_22750,N_23072);
and U25582 (N_25582,N_23714,N_23961);
and U25583 (N_25583,N_22183,N_22124);
xor U25584 (N_25584,N_23256,N_22175);
nand U25585 (N_25585,N_23985,N_23166);
nor U25586 (N_25586,N_23377,N_22421);
xnor U25587 (N_25587,N_23933,N_22273);
xnor U25588 (N_25588,N_22461,N_23607);
nor U25589 (N_25589,N_23515,N_23589);
or U25590 (N_25590,N_23210,N_23120);
and U25591 (N_25591,N_23576,N_23009);
nand U25592 (N_25592,N_23855,N_22674);
or U25593 (N_25593,N_23657,N_23413);
xor U25594 (N_25594,N_23713,N_22847);
and U25595 (N_25595,N_23627,N_23574);
xor U25596 (N_25596,N_23537,N_23055);
or U25597 (N_25597,N_23940,N_23428);
nand U25598 (N_25598,N_23223,N_23285);
nand U25599 (N_25599,N_22763,N_23342);
nor U25600 (N_25600,N_23653,N_22022);
nand U25601 (N_25601,N_22501,N_22097);
and U25602 (N_25602,N_22417,N_23841);
nand U25603 (N_25603,N_22724,N_23465);
nor U25604 (N_25604,N_22868,N_22223);
nor U25605 (N_25605,N_23026,N_23586);
nand U25606 (N_25606,N_23612,N_23700);
nor U25607 (N_25607,N_22117,N_22328);
or U25608 (N_25608,N_22779,N_22253);
nand U25609 (N_25609,N_23442,N_22147);
nor U25610 (N_25610,N_23590,N_22023);
xor U25611 (N_25611,N_22222,N_22207);
xnor U25612 (N_25612,N_22567,N_22617);
nor U25613 (N_25613,N_23379,N_23537);
nand U25614 (N_25614,N_22498,N_22094);
or U25615 (N_25615,N_22038,N_22811);
or U25616 (N_25616,N_22796,N_22430);
or U25617 (N_25617,N_22221,N_23597);
xor U25618 (N_25618,N_23269,N_22338);
and U25619 (N_25619,N_23615,N_22704);
nand U25620 (N_25620,N_22082,N_22483);
or U25621 (N_25621,N_22302,N_22462);
and U25622 (N_25622,N_23864,N_23508);
and U25623 (N_25623,N_22896,N_22417);
nand U25624 (N_25624,N_22405,N_22235);
and U25625 (N_25625,N_22431,N_22330);
and U25626 (N_25626,N_23642,N_23401);
xor U25627 (N_25627,N_23043,N_23504);
and U25628 (N_25628,N_22404,N_23465);
xor U25629 (N_25629,N_22521,N_22201);
or U25630 (N_25630,N_22698,N_23053);
nor U25631 (N_25631,N_22946,N_23487);
or U25632 (N_25632,N_23812,N_23068);
or U25633 (N_25633,N_23417,N_22439);
nand U25634 (N_25634,N_23849,N_23934);
nor U25635 (N_25635,N_23879,N_23513);
or U25636 (N_25636,N_23441,N_22886);
nand U25637 (N_25637,N_22379,N_22744);
nand U25638 (N_25638,N_22877,N_22476);
nor U25639 (N_25639,N_22678,N_23884);
or U25640 (N_25640,N_22464,N_22821);
and U25641 (N_25641,N_22721,N_22370);
or U25642 (N_25642,N_23908,N_22024);
or U25643 (N_25643,N_23773,N_23286);
nor U25644 (N_25644,N_23853,N_22253);
or U25645 (N_25645,N_23842,N_23077);
and U25646 (N_25646,N_22120,N_22360);
nand U25647 (N_25647,N_23002,N_22479);
xnor U25648 (N_25648,N_23394,N_23561);
nor U25649 (N_25649,N_22806,N_22138);
nand U25650 (N_25650,N_22212,N_23330);
and U25651 (N_25651,N_22074,N_22366);
xor U25652 (N_25652,N_22420,N_23544);
or U25653 (N_25653,N_23361,N_23477);
nand U25654 (N_25654,N_23948,N_23483);
nand U25655 (N_25655,N_23927,N_23787);
xnor U25656 (N_25656,N_22580,N_22140);
and U25657 (N_25657,N_22285,N_22192);
and U25658 (N_25658,N_22718,N_23560);
or U25659 (N_25659,N_23099,N_23150);
nor U25660 (N_25660,N_22153,N_22179);
or U25661 (N_25661,N_23594,N_22026);
nand U25662 (N_25662,N_22612,N_22847);
xnor U25663 (N_25663,N_23442,N_23985);
xnor U25664 (N_25664,N_23565,N_22141);
nor U25665 (N_25665,N_22378,N_23234);
nor U25666 (N_25666,N_23544,N_23406);
or U25667 (N_25667,N_22335,N_22952);
and U25668 (N_25668,N_22019,N_23721);
nor U25669 (N_25669,N_22969,N_22355);
xnor U25670 (N_25670,N_22101,N_23727);
nor U25671 (N_25671,N_22661,N_22905);
nand U25672 (N_25672,N_23496,N_22840);
nor U25673 (N_25673,N_23521,N_23541);
xnor U25674 (N_25674,N_22224,N_22148);
or U25675 (N_25675,N_22286,N_22151);
and U25676 (N_25676,N_23118,N_22704);
nand U25677 (N_25677,N_22965,N_23409);
and U25678 (N_25678,N_22526,N_23488);
or U25679 (N_25679,N_23669,N_23361);
xnor U25680 (N_25680,N_23393,N_22796);
nor U25681 (N_25681,N_23576,N_23803);
nand U25682 (N_25682,N_22261,N_22877);
xnor U25683 (N_25683,N_23571,N_22333);
and U25684 (N_25684,N_22009,N_23599);
nor U25685 (N_25685,N_23398,N_22135);
xor U25686 (N_25686,N_22912,N_22818);
nor U25687 (N_25687,N_23584,N_23093);
and U25688 (N_25688,N_22386,N_22418);
or U25689 (N_25689,N_23461,N_23895);
nand U25690 (N_25690,N_22989,N_22254);
xnor U25691 (N_25691,N_22857,N_23363);
nor U25692 (N_25692,N_23636,N_22296);
nor U25693 (N_25693,N_23849,N_22375);
xnor U25694 (N_25694,N_22422,N_23572);
nor U25695 (N_25695,N_22118,N_22789);
and U25696 (N_25696,N_22733,N_23264);
or U25697 (N_25697,N_22707,N_23145);
and U25698 (N_25698,N_22965,N_22939);
nand U25699 (N_25699,N_23342,N_23897);
and U25700 (N_25700,N_23759,N_22748);
xor U25701 (N_25701,N_23993,N_23034);
and U25702 (N_25702,N_23799,N_22903);
xor U25703 (N_25703,N_23943,N_22272);
nand U25704 (N_25704,N_22917,N_23424);
nor U25705 (N_25705,N_23732,N_22210);
nor U25706 (N_25706,N_22580,N_23434);
and U25707 (N_25707,N_22655,N_22881);
and U25708 (N_25708,N_22783,N_23047);
nor U25709 (N_25709,N_23077,N_22770);
or U25710 (N_25710,N_22657,N_22918);
xnor U25711 (N_25711,N_23275,N_22277);
xor U25712 (N_25712,N_23838,N_22106);
nor U25713 (N_25713,N_22263,N_23876);
xnor U25714 (N_25714,N_23091,N_22109);
xor U25715 (N_25715,N_22552,N_22874);
or U25716 (N_25716,N_22757,N_23901);
or U25717 (N_25717,N_23013,N_22988);
or U25718 (N_25718,N_23209,N_23821);
xor U25719 (N_25719,N_23930,N_23447);
and U25720 (N_25720,N_22558,N_23672);
nand U25721 (N_25721,N_23493,N_23412);
nand U25722 (N_25722,N_23015,N_22538);
xor U25723 (N_25723,N_22549,N_23181);
xnor U25724 (N_25724,N_23921,N_23778);
xnor U25725 (N_25725,N_22214,N_22630);
and U25726 (N_25726,N_23903,N_22238);
nor U25727 (N_25727,N_22702,N_23606);
or U25728 (N_25728,N_22094,N_23941);
nand U25729 (N_25729,N_22490,N_22034);
or U25730 (N_25730,N_22579,N_23365);
or U25731 (N_25731,N_23949,N_22086);
xor U25732 (N_25732,N_22578,N_22874);
or U25733 (N_25733,N_22944,N_22109);
nand U25734 (N_25734,N_22017,N_22681);
or U25735 (N_25735,N_23525,N_22947);
xnor U25736 (N_25736,N_22408,N_23029);
nand U25737 (N_25737,N_22768,N_22904);
nand U25738 (N_25738,N_22882,N_23682);
nand U25739 (N_25739,N_22908,N_22599);
nor U25740 (N_25740,N_22895,N_22984);
or U25741 (N_25741,N_22177,N_22439);
and U25742 (N_25742,N_23148,N_23334);
nor U25743 (N_25743,N_23811,N_23730);
nor U25744 (N_25744,N_22474,N_22313);
nor U25745 (N_25745,N_23009,N_22920);
nor U25746 (N_25746,N_22986,N_23344);
nor U25747 (N_25747,N_23911,N_22752);
nor U25748 (N_25748,N_23423,N_22196);
nand U25749 (N_25749,N_23790,N_23968);
and U25750 (N_25750,N_23679,N_22871);
or U25751 (N_25751,N_23837,N_22908);
and U25752 (N_25752,N_23013,N_23787);
xor U25753 (N_25753,N_22545,N_23274);
and U25754 (N_25754,N_22135,N_22860);
nand U25755 (N_25755,N_22437,N_22592);
nor U25756 (N_25756,N_23098,N_23015);
nor U25757 (N_25757,N_23703,N_22075);
and U25758 (N_25758,N_23624,N_22764);
or U25759 (N_25759,N_23087,N_23838);
xnor U25760 (N_25760,N_23582,N_22465);
nor U25761 (N_25761,N_22635,N_23905);
xor U25762 (N_25762,N_22866,N_22315);
nor U25763 (N_25763,N_23127,N_23538);
and U25764 (N_25764,N_22134,N_22911);
nor U25765 (N_25765,N_22126,N_23401);
nand U25766 (N_25766,N_22638,N_22836);
nand U25767 (N_25767,N_22219,N_23980);
or U25768 (N_25768,N_23414,N_23721);
and U25769 (N_25769,N_22364,N_23990);
nand U25770 (N_25770,N_22531,N_23155);
and U25771 (N_25771,N_23288,N_23095);
xor U25772 (N_25772,N_22596,N_23545);
xor U25773 (N_25773,N_22093,N_22135);
nor U25774 (N_25774,N_23990,N_23320);
nor U25775 (N_25775,N_22510,N_22011);
nand U25776 (N_25776,N_22774,N_22411);
nand U25777 (N_25777,N_23394,N_23535);
nand U25778 (N_25778,N_22571,N_23263);
nand U25779 (N_25779,N_23663,N_22264);
nor U25780 (N_25780,N_23023,N_22347);
and U25781 (N_25781,N_23475,N_23832);
xor U25782 (N_25782,N_22674,N_23870);
xnor U25783 (N_25783,N_23173,N_23362);
nand U25784 (N_25784,N_23518,N_22584);
or U25785 (N_25785,N_23573,N_22243);
nor U25786 (N_25786,N_22801,N_22012);
and U25787 (N_25787,N_22860,N_22157);
and U25788 (N_25788,N_22254,N_22269);
xor U25789 (N_25789,N_22233,N_23876);
or U25790 (N_25790,N_22019,N_23450);
nor U25791 (N_25791,N_23554,N_23301);
or U25792 (N_25792,N_22918,N_22986);
nor U25793 (N_25793,N_23598,N_22274);
nor U25794 (N_25794,N_23100,N_22289);
or U25795 (N_25795,N_23601,N_22012);
nor U25796 (N_25796,N_23257,N_23418);
xnor U25797 (N_25797,N_22032,N_22160);
xor U25798 (N_25798,N_22233,N_22293);
and U25799 (N_25799,N_23774,N_23654);
or U25800 (N_25800,N_23398,N_22422);
and U25801 (N_25801,N_22258,N_23431);
and U25802 (N_25802,N_22904,N_23320);
nand U25803 (N_25803,N_23930,N_22997);
or U25804 (N_25804,N_22892,N_22074);
or U25805 (N_25805,N_22750,N_23348);
and U25806 (N_25806,N_23894,N_23544);
nand U25807 (N_25807,N_23995,N_22231);
nor U25808 (N_25808,N_22931,N_22566);
or U25809 (N_25809,N_23873,N_22334);
nor U25810 (N_25810,N_23653,N_23866);
or U25811 (N_25811,N_23226,N_22986);
nand U25812 (N_25812,N_22737,N_22792);
xor U25813 (N_25813,N_22437,N_23655);
nor U25814 (N_25814,N_22604,N_23616);
or U25815 (N_25815,N_22558,N_22204);
and U25816 (N_25816,N_22820,N_23214);
xor U25817 (N_25817,N_23937,N_23677);
nor U25818 (N_25818,N_23140,N_22927);
or U25819 (N_25819,N_22429,N_22154);
nor U25820 (N_25820,N_23184,N_23927);
nand U25821 (N_25821,N_22084,N_22771);
and U25822 (N_25822,N_22298,N_23872);
or U25823 (N_25823,N_23958,N_22281);
and U25824 (N_25824,N_22160,N_22141);
xnor U25825 (N_25825,N_23660,N_23805);
and U25826 (N_25826,N_22126,N_23797);
and U25827 (N_25827,N_22997,N_23469);
xor U25828 (N_25828,N_22734,N_23484);
nand U25829 (N_25829,N_22502,N_22070);
xor U25830 (N_25830,N_22554,N_23016);
xnor U25831 (N_25831,N_23451,N_23624);
or U25832 (N_25832,N_23901,N_23741);
nor U25833 (N_25833,N_22818,N_23610);
nor U25834 (N_25834,N_22664,N_23897);
or U25835 (N_25835,N_22192,N_22661);
nand U25836 (N_25836,N_22102,N_23378);
xnor U25837 (N_25837,N_23848,N_23620);
or U25838 (N_25838,N_23786,N_22489);
or U25839 (N_25839,N_22796,N_22966);
xor U25840 (N_25840,N_23482,N_22629);
xor U25841 (N_25841,N_22514,N_23857);
nor U25842 (N_25842,N_23272,N_22375);
nand U25843 (N_25843,N_23104,N_22730);
nor U25844 (N_25844,N_23734,N_22578);
nor U25845 (N_25845,N_23735,N_23090);
and U25846 (N_25846,N_22606,N_23858);
xnor U25847 (N_25847,N_23462,N_23592);
nand U25848 (N_25848,N_22750,N_22093);
nand U25849 (N_25849,N_22479,N_22747);
nand U25850 (N_25850,N_22778,N_22688);
and U25851 (N_25851,N_23753,N_23724);
or U25852 (N_25852,N_23424,N_22141);
xnor U25853 (N_25853,N_23856,N_23499);
xnor U25854 (N_25854,N_23799,N_23725);
or U25855 (N_25855,N_23165,N_22752);
and U25856 (N_25856,N_23138,N_22001);
nor U25857 (N_25857,N_22594,N_22402);
or U25858 (N_25858,N_23310,N_22740);
nor U25859 (N_25859,N_23578,N_23172);
and U25860 (N_25860,N_22755,N_23083);
and U25861 (N_25861,N_23588,N_22874);
or U25862 (N_25862,N_22898,N_22709);
xor U25863 (N_25863,N_23749,N_23123);
nor U25864 (N_25864,N_23890,N_23658);
nor U25865 (N_25865,N_23548,N_22890);
and U25866 (N_25866,N_22566,N_22584);
or U25867 (N_25867,N_22188,N_23080);
nand U25868 (N_25868,N_23990,N_22968);
and U25869 (N_25869,N_22685,N_22833);
nand U25870 (N_25870,N_22782,N_22512);
nand U25871 (N_25871,N_22493,N_23967);
or U25872 (N_25872,N_22039,N_22575);
or U25873 (N_25873,N_23111,N_22483);
and U25874 (N_25874,N_23381,N_23140);
xor U25875 (N_25875,N_23282,N_22977);
nand U25876 (N_25876,N_23926,N_22607);
and U25877 (N_25877,N_23633,N_22789);
and U25878 (N_25878,N_22970,N_22188);
nor U25879 (N_25879,N_23593,N_22944);
or U25880 (N_25880,N_22582,N_23423);
nand U25881 (N_25881,N_22518,N_23558);
nor U25882 (N_25882,N_22855,N_23375);
nor U25883 (N_25883,N_23664,N_22200);
and U25884 (N_25884,N_23062,N_22479);
nand U25885 (N_25885,N_23292,N_22950);
xor U25886 (N_25886,N_23879,N_23031);
or U25887 (N_25887,N_23280,N_23012);
nor U25888 (N_25888,N_22216,N_23523);
nand U25889 (N_25889,N_23765,N_23961);
nand U25890 (N_25890,N_22291,N_22686);
nor U25891 (N_25891,N_22414,N_23721);
and U25892 (N_25892,N_23547,N_23646);
nor U25893 (N_25893,N_22627,N_22432);
or U25894 (N_25894,N_23546,N_23961);
nand U25895 (N_25895,N_22599,N_23495);
and U25896 (N_25896,N_22220,N_23379);
nor U25897 (N_25897,N_23032,N_22746);
nand U25898 (N_25898,N_23626,N_23267);
xor U25899 (N_25899,N_22834,N_22854);
or U25900 (N_25900,N_23881,N_22864);
and U25901 (N_25901,N_23567,N_23633);
nor U25902 (N_25902,N_23764,N_23798);
xor U25903 (N_25903,N_22703,N_22459);
xor U25904 (N_25904,N_23226,N_22780);
xnor U25905 (N_25905,N_23965,N_23319);
nand U25906 (N_25906,N_23424,N_23852);
nor U25907 (N_25907,N_23923,N_23999);
nor U25908 (N_25908,N_22389,N_23092);
and U25909 (N_25909,N_22629,N_23660);
or U25910 (N_25910,N_22710,N_22855);
or U25911 (N_25911,N_23764,N_22326);
nand U25912 (N_25912,N_22375,N_22582);
nor U25913 (N_25913,N_22909,N_22273);
nand U25914 (N_25914,N_23975,N_23247);
nor U25915 (N_25915,N_23060,N_23097);
xnor U25916 (N_25916,N_22543,N_23226);
nor U25917 (N_25917,N_22334,N_23257);
xnor U25918 (N_25918,N_23492,N_23702);
and U25919 (N_25919,N_22445,N_23387);
xor U25920 (N_25920,N_23631,N_22148);
nand U25921 (N_25921,N_23647,N_22982);
or U25922 (N_25922,N_22928,N_23486);
and U25923 (N_25923,N_22799,N_22150);
nand U25924 (N_25924,N_23177,N_22449);
nor U25925 (N_25925,N_22931,N_22975);
xnor U25926 (N_25926,N_22320,N_22214);
xnor U25927 (N_25927,N_22571,N_22806);
nor U25928 (N_25928,N_22360,N_23114);
nand U25929 (N_25929,N_23050,N_23082);
and U25930 (N_25930,N_22640,N_23775);
nor U25931 (N_25931,N_22249,N_23087);
or U25932 (N_25932,N_22094,N_22625);
and U25933 (N_25933,N_22297,N_23922);
nor U25934 (N_25934,N_23929,N_23903);
nand U25935 (N_25935,N_23264,N_22295);
xor U25936 (N_25936,N_23123,N_22698);
and U25937 (N_25937,N_23459,N_23255);
nand U25938 (N_25938,N_22954,N_22738);
nor U25939 (N_25939,N_22224,N_23401);
nand U25940 (N_25940,N_23173,N_23929);
and U25941 (N_25941,N_22905,N_23441);
and U25942 (N_25942,N_23269,N_22859);
nand U25943 (N_25943,N_23061,N_23425);
nor U25944 (N_25944,N_23379,N_22996);
nor U25945 (N_25945,N_22318,N_22305);
nor U25946 (N_25946,N_23003,N_22380);
and U25947 (N_25947,N_23725,N_23905);
or U25948 (N_25948,N_22683,N_22226);
xnor U25949 (N_25949,N_23609,N_23694);
or U25950 (N_25950,N_22527,N_23737);
or U25951 (N_25951,N_23570,N_23676);
nand U25952 (N_25952,N_22739,N_22272);
or U25953 (N_25953,N_22974,N_23937);
and U25954 (N_25954,N_22846,N_23748);
nand U25955 (N_25955,N_23317,N_22003);
nand U25956 (N_25956,N_22378,N_23350);
nand U25957 (N_25957,N_22093,N_23918);
xor U25958 (N_25958,N_23120,N_23742);
nand U25959 (N_25959,N_23413,N_22836);
nand U25960 (N_25960,N_22876,N_22714);
or U25961 (N_25961,N_23776,N_23045);
or U25962 (N_25962,N_22133,N_22385);
nor U25963 (N_25963,N_23105,N_22266);
nor U25964 (N_25964,N_22429,N_22126);
nor U25965 (N_25965,N_22622,N_23011);
or U25966 (N_25966,N_22029,N_23522);
nor U25967 (N_25967,N_22245,N_23539);
or U25968 (N_25968,N_22737,N_23083);
xor U25969 (N_25969,N_23626,N_23124);
xor U25970 (N_25970,N_23731,N_22426);
nor U25971 (N_25971,N_22972,N_23612);
nand U25972 (N_25972,N_22200,N_22256);
nor U25973 (N_25973,N_22302,N_22932);
nor U25974 (N_25974,N_23755,N_22400);
or U25975 (N_25975,N_23252,N_23769);
and U25976 (N_25976,N_23967,N_23164);
nor U25977 (N_25977,N_23171,N_23134);
xor U25978 (N_25978,N_23300,N_22025);
nand U25979 (N_25979,N_22725,N_22493);
nor U25980 (N_25980,N_22314,N_23378);
and U25981 (N_25981,N_22714,N_22861);
or U25982 (N_25982,N_22300,N_22924);
nor U25983 (N_25983,N_23798,N_22087);
nor U25984 (N_25984,N_22720,N_22057);
or U25985 (N_25985,N_22868,N_22283);
or U25986 (N_25986,N_23526,N_23485);
nor U25987 (N_25987,N_22563,N_22150);
nand U25988 (N_25988,N_23407,N_22476);
or U25989 (N_25989,N_23078,N_23660);
nand U25990 (N_25990,N_22343,N_23706);
nand U25991 (N_25991,N_22112,N_23030);
nand U25992 (N_25992,N_23622,N_23853);
or U25993 (N_25993,N_23118,N_23005);
nand U25994 (N_25994,N_22966,N_22771);
and U25995 (N_25995,N_23698,N_22564);
xnor U25996 (N_25996,N_23490,N_22786);
and U25997 (N_25997,N_23109,N_22208);
nand U25998 (N_25998,N_22283,N_22183);
or U25999 (N_25999,N_23535,N_22399);
xnor U26000 (N_26000,N_25217,N_25696);
nand U26001 (N_26001,N_25590,N_24239);
xor U26002 (N_26002,N_24629,N_25798);
xor U26003 (N_26003,N_24904,N_25693);
xor U26004 (N_26004,N_24879,N_25716);
xor U26005 (N_26005,N_25632,N_25496);
nand U26006 (N_26006,N_25109,N_24832);
or U26007 (N_26007,N_25244,N_25376);
nand U26008 (N_26008,N_25873,N_24459);
and U26009 (N_26009,N_25541,N_24698);
nor U26010 (N_26010,N_25200,N_25897);
xor U26011 (N_26011,N_24678,N_25165);
or U26012 (N_26012,N_24840,N_24173);
and U26013 (N_26013,N_25099,N_24383);
xor U26014 (N_26014,N_25146,N_25457);
xnor U26015 (N_26015,N_25345,N_24405);
or U26016 (N_26016,N_24863,N_25233);
and U26017 (N_26017,N_25446,N_24739);
xor U26018 (N_26018,N_24509,N_25971);
or U26019 (N_26019,N_24030,N_24649);
xnor U26020 (N_26020,N_25239,N_25451);
nor U26021 (N_26021,N_25121,N_24848);
and U26022 (N_26022,N_24265,N_25566);
nor U26023 (N_26023,N_24395,N_24429);
and U26024 (N_26024,N_24465,N_24836);
xor U26025 (N_26025,N_25319,N_25361);
and U26026 (N_26026,N_25374,N_24216);
or U26027 (N_26027,N_24112,N_25096);
and U26028 (N_26028,N_24387,N_24727);
or U26029 (N_26029,N_24307,N_24577);
xnor U26030 (N_26030,N_25282,N_24165);
and U26031 (N_26031,N_24224,N_24500);
nand U26032 (N_26032,N_25092,N_25279);
nand U26033 (N_26033,N_24343,N_24448);
nor U26034 (N_26034,N_24772,N_24450);
xor U26035 (N_26035,N_24281,N_25934);
or U26036 (N_26036,N_24236,N_25932);
nor U26037 (N_26037,N_25117,N_25245);
nand U26038 (N_26038,N_25802,N_24267);
nand U26039 (N_26039,N_24285,N_25445);
nand U26040 (N_26040,N_25366,N_24133);
and U26041 (N_26041,N_25722,N_24699);
xnor U26042 (N_26042,N_25562,N_24347);
and U26043 (N_26043,N_25638,N_24110);
nand U26044 (N_26044,N_24306,N_24948);
nand U26045 (N_26045,N_24378,N_25699);
xor U26046 (N_26046,N_24080,N_24147);
xor U26047 (N_26047,N_24135,N_25786);
nand U26048 (N_26048,N_24303,N_24501);
nand U26049 (N_26049,N_24017,N_24161);
and U26050 (N_26050,N_24547,N_25054);
nor U26051 (N_26051,N_25154,N_25019);
nor U26052 (N_26052,N_25704,N_24619);
xor U26053 (N_26053,N_25461,N_25213);
nor U26054 (N_26054,N_25964,N_24985);
xnor U26055 (N_26055,N_24601,N_25959);
or U26056 (N_26056,N_24978,N_24758);
or U26057 (N_26057,N_25483,N_25236);
or U26058 (N_26058,N_24116,N_24624);
and U26059 (N_26059,N_24205,N_25998);
nor U26060 (N_26060,N_24872,N_25202);
or U26061 (N_26061,N_24851,N_25066);
xor U26062 (N_26062,N_25384,N_24591);
xnor U26063 (N_26063,N_24578,N_25396);
nand U26064 (N_26064,N_24003,N_25424);
or U26065 (N_26065,N_25620,N_25878);
and U26066 (N_26066,N_25967,N_24167);
xnor U26067 (N_26067,N_25501,N_25455);
or U26068 (N_26068,N_25063,N_25456);
nor U26069 (N_26069,N_25460,N_24573);
nor U26070 (N_26070,N_24873,N_25194);
nand U26071 (N_26071,N_24249,N_25556);
and U26072 (N_26072,N_25883,N_25206);
nand U26073 (N_26073,N_25776,N_25125);
and U26074 (N_26074,N_25310,N_24934);
xnor U26075 (N_26075,N_24084,N_25104);
and U26076 (N_26076,N_25685,N_25952);
or U26077 (N_26077,N_25865,N_24548);
and U26078 (N_26078,N_24790,N_24476);
xnor U26079 (N_26079,N_24046,N_25951);
and U26080 (N_26080,N_25133,N_25037);
xnor U26081 (N_26081,N_24055,N_24291);
and U26082 (N_26082,N_24217,N_24759);
or U26083 (N_26083,N_24109,N_25264);
or U26084 (N_26084,N_25588,N_24953);
and U26085 (N_26085,N_24066,N_24685);
nand U26086 (N_26086,N_25612,N_24036);
nor U26087 (N_26087,N_25403,N_25508);
and U26088 (N_26088,N_25850,N_24855);
nor U26089 (N_26089,N_24014,N_25559);
nand U26090 (N_26090,N_24566,N_24033);
xor U26091 (N_26091,N_25695,N_25475);
nand U26092 (N_26092,N_25675,N_24958);
or U26093 (N_26093,N_25933,N_24766);
xnor U26094 (N_26094,N_24241,N_24233);
or U26095 (N_26095,N_24426,N_25163);
xnor U26096 (N_26096,N_24326,N_25809);
and U26097 (N_26097,N_24364,N_24568);
and U26098 (N_26098,N_24527,N_25619);
or U26099 (N_26099,N_25986,N_24882);
nand U26100 (N_26100,N_24164,N_24918);
xor U26101 (N_26101,N_24104,N_25022);
or U26102 (N_26102,N_24632,N_24775);
nand U26103 (N_26103,N_25315,N_24345);
nand U26104 (N_26104,N_24599,N_24681);
nand U26105 (N_26105,N_25118,N_24746);
nand U26106 (N_26106,N_24246,N_24102);
and U26107 (N_26107,N_24461,N_25758);
or U26108 (N_26108,N_25771,N_24410);
or U26109 (N_26109,N_24447,N_24021);
and U26110 (N_26110,N_24412,N_24451);
nor U26111 (N_26111,N_25956,N_24034);
nor U26112 (N_26112,N_24423,N_25819);
nand U26113 (N_26113,N_25907,N_24397);
nor U26114 (N_26114,N_25751,N_25683);
nor U26115 (N_26115,N_25868,N_25304);
xor U26116 (N_26116,N_24234,N_24835);
or U26117 (N_26117,N_25831,N_24594);
xor U26118 (N_26118,N_25308,N_24314);
and U26119 (N_26119,N_25357,N_25631);
or U26120 (N_26120,N_24063,N_24422);
nor U26121 (N_26121,N_25654,N_24433);
nand U26122 (N_26122,N_25923,N_24089);
nand U26123 (N_26123,N_24489,N_25199);
xnor U26124 (N_26124,N_24714,N_24270);
xnor U26125 (N_26125,N_24440,N_24574);
xor U26126 (N_26126,N_25145,N_24081);
nand U26127 (N_26127,N_25237,N_24590);
nand U26128 (N_26128,N_25792,N_25979);
and U26129 (N_26129,N_24644,N_25225);
nor U26130 (N_26130,N_25368,N_25207);
nor U26131 (N_26131,N_25656,N_25925);
and U26132 (N_26132,N_25415,N_25625);
nor U26133 (N_26133,N_24959,N_24386);
xor U26134 (N_26134,N_25116,N_25313);
or U26135 (N_26135,N_24235,N_25431);
nor U26136 (N_26136,N_25421,N_25557);
xnor U26137 (N_26137,N_24930,N_24262);
and U26138 (N_26138,N_24750,N_24610);
nand U26139 (N_26139,N_24210,N_25487);
and U26140 (N_26140,N_25746,N_24976);
nor U26141 (N_26141,N_24616,N_25673);
or U26142 (N_26142,N_24126,N_25161);
nor U26143 (N_26143,N_25263,N_25734);
nand U26144 (N_26144,N_25135,N_24850);
nand U26145 (N_26145,N_25482,N_25587);
nor U26146 (N_26146,N_24881,N_24809);
nor U26147 (N_26147,N_25079,N_24458);
xnor U26148 (N_26148,N_25278,N_25769);
and U26149 (N_26149,N_25558,N_24979);
or U26150 (N_26150,N_25807,N_24226);
nand U26151 (N_26151,N_25427,N_25533);
xnor U26152 (N_26152,N_24705,N_24263);
and U26153 (N_26153,N_24582,N_25834);
or U26154 (N_26154,N_24981,N_24402);
and U26155 (N_26155,N_25682,N_25276);
xnor U26156 (N_26156,N_25314,N_24097);
nand U26157 (N_26157,N_25929,N_25597);
and U26158 (N_26158,N_25780,N_24277);
and U26159 (N_26159,N_24951,N_24301);
or U26160 (N_26160,N_24514,N_25546);
nor U26161 (N_26161,N_24354,N_25908);
or U26162 (N_26162,N_24803,N_24741);
nand U26163 (N_26163,N_24572,N_24592);
xnor U26164 (N_26164,N_24288,N_24072);
or U26165 (N_26165,N_24630,N_25761);
nor U26166 (N_26166,N_24519,N_25754);
and U26167 (N_26167,N_25000,N_25863);
xor U26168 (N_26168,N_24670,N_24571);
or U26169 (N_26169,N_24039,N_24861);
xnor U26170 (N_26170,N_24789,N_24128);
nand U26171 (N_26171,N_24119,N_25611);
or U26172 (N_26172,N_25589,N_25380);
nand U26173 (N_26173,N_25718,N_25791);
or U26174 (N_26174,N_25574,N_25895);
xor U26175 (N_26175,N_25339,N_25347);
xnor U26176 (N_26176,N_24980,N_24122);
xor U26177 (N_26177,N_24598,N_24731);
xnor U26178 (N_26178,N_25976,N_25367);
or U26179 (N_26179,N_25195,N_25355);
nor U26180 (N_26180,N_25586,N_24642);
and U26181 (N_26181,N_24986,N_24550);
or U26182 (N_26182,N_24087,N_24579);
xnor U26183 (N_26183,N_24196,N_25797);
or U26184 (N_26184,N_24316,N_24664);
xor U26185 (N_26185,N_25666,N_24048);
nand U26186 (N_26186,N_24323,N_25226);
or U26187 (N_26187,N_24657,N_24770);
xor U26188 (N_26188,N_24812,N_24340);
or U26189 (N_26189,N_25606,N_24283);
or U26190 (N_26190,N_24889,N_24963);
nor U26191 (N_26191,N_25604,N_24192);
xnor U26192 (N_26192,N_24600,N_25261);
nor U26193 (N_26193,N_24893,N_24862);
or U26194 (N_26194,N_24666,N_25227);
nand U26195 (N_26195,N_25193,N_25982);
nand U26196 (N_26196,N_24074,N_25476);
nor U26197 (N_26197,N_25515,N_24182);
or U26198 (N_26198,N_25253,N_25062);
nand U26199 (N_26199,N_25958,N_25886);
nor U26200 (N_26200,N_25548,N_24427);
and U26201 (N_26201,N_24774,N_25039);
nor U26202 (N_26202,N_24010,N_24208);
and U26203 (N_26203,N_25273,N_24655);
nor U26204 (N_26204,N_24361,N_24312);
xor U26205 (N_26205,N_24520,N_24073);
nor U26206 (N_26206,N_24810,N_25223);
or U26207 (N_26207,N_25905,N_25488);
nand U26208 (N_26208,N_24016,N_25267);
nor U26209 (N_26209,N_24299,N_24031);
nor U26210 (N_26210,N_25720,N_24682);
nor U26211 (N_26211,N_25745,N_25494);
and U26212 (N_26212,N_25983,N_24901);
xor U26213 (N_26213,N_24141,N_25749);
xnor U26214 (N_26214,N_25860,N_24227);
nand U26215 (N_26215,N_25793,N_24778);
nand U26216 (N_26216,N_24996,N_25406);
or U26217 (N_26217,N_25107,N_25038);
nor U26218 (N_26218,N_24777,N_24908);
nor U26219 (N_26219,N_24223,N_24732);
nand U26220 (N_26220,N_24178,N_25531);
and U26221 (N_26221,N_25600,N_24172);
nand U26222 (N_26222,N_25535,N_24138);
nand U26223 (N_26223,N_25605,N_24114);
or U26224 (N_26224,N_24026,N_25286);
xnor U26225 (N_26225,N_24555,N_25766);
nand U26226 (N_26226,N_24379,N_25829);
and U26227 (N_26227,N_25156,N_25861);
nand U26228 (N_26228,N_24987,N_25473);
nor U26229 (N_26229,N_25744,N_25658);
and U26230 (N_26230,N_24310,N_25081);
nand U26231 (N_26231,N_25428,N_25763);
and U26232 (N_26232,N_25256,N_24139);
xor U26233 (N_26233,N_25034,N_24372);
nor U26234 (N_26234,N_24738,N_25452);
or U26235 (N_26235,N_24703,N_24059);
nor U26236 (N_26236,N_25065,N_24942);
or U26237 (N_26237,N_25218,N_25235);
nor U26238 (N_26238,N_24069,N_25180);
nor U26239 (N_26239,N_24043,N_25901);
or U26240 (N_26240,N_24931,N_25700);
nand U26241 (N_26241,N_25220,N_25184);
xnor U26242 (N_26242,N_24160,N_25914);
nand U26243 (N_26243,N_25375,N_24845);
nand U26244 (N_26244,N_25325,N_24020);
and U26245 (N_26245,N_25166,N_25527);
nand U26246 (N_26246,N_24919,N_25513);
nand U26247 (N_26247,N_24169,N_24502);
xnor U26248 (N_26248,N_25930,N_25516);
nor U26249 (N_26249,N_24710,N_24654);
nor U26250 (N_26250,N_24240,N_25972);
and U26251 (N_26251,N_24174,N_24067);
nand U26252 (N_26252,N_25813,N_24825);
xnor U26253 (N_26253,N_24330,N_24242);
nor U26254 (N_26254,N_24858,N_25708);
and U26255 (N_26255,N_24508,N_24800);
nand U26256 (N_26256,N_24415,N_24480);
nand U26257 (N_26257,N_25551,N_25290);
nor U26258 (N_26258,N_24284,N_24822);
and U26259 (N_26259,N_25271,N_25651);
or U26260 (N_26260,N_25041,N_24757);
nand U26261 (N_26261,N_25035,N_24311);
nand U26262 (N_26262,N_25316,N_24209);
nand U26263 (N_26263,N_24785,N_25836);
xor U26264 (N_26264,N_25894,N_25690);
nand U26265 (N_26265,N_24761,N_25067);
or U26266 (N_26266,N_25387,N_24878);
and U26267 (N_26267,N_24237,N_24085);
nor U26268 (N_26268,N_25594,N_24317);
nand U26269 (N_26269,N_25337,N_24042);
and U26270 (N_26270,N_25134,N_25843);
xnor U26271 (N_26271,N_24793,N_25214);
xor U26272 (N_26272,N_25961,N_25444);
xnor U26273 (N_26273,N_25162,N_24683);
and U26274 (N_26274,N_24620,N_25300);
or U26275 (N_26275,N_25911,N_24200);
nor U26276 (N_26276,N_25856,N_24045);
nand U26277 (N_26277,N_25664,N_24184);
or U26278 (N_26278,N_24635,N_24542);
nand U26279 (N_26279,N_25921,N_24896);
nand U26280 (N_26280,N_25910,N_25497);
nor U26281 (N_26281,N_24539,N_25917);
and U26282 (N_26282,N_25505,N_25634);
or U26283 (N_26283,N_24193,N_24337);
xor U26284 (N_26284,N_24887,N_24814);
nor U26285 (N_26285,N_25191,N_25047);
xnor U26286 (N_26286,N_25639,N_25999);
or U26287 (N_26287,N_25944,N_24168);
nor U26288 (N_26288,N_25420,N_24499);
nor U26289 (N_26289,N_24211,N_25719);
xnor U26290 (N_26290,N_24818,N_25434);
nand U26291 (N_26291,N_24298,N_24890);
nand U26292 (N_26292,N_24910,N_25411);
and U26293 (N_26293,N_24222,N_25143);
nand U26294 (N_26294,N_25224,N_24324);
nor U26295 (N_26295,N_25867,N_24622);
nor U26296 (N_26296,N_25647,N_25108);
and U26297 (N_26297,N_24396,N_24843);
or U26298 (N_26298,N_24556,N_25371);
xnor U26299 (N_26299,N_25024,N_25378);
nand U26300 (N_26300,N_25928,N_25847);
or U26301 (N_26301,N_25111,N_25692);
xnor U26302 (N_26302,N_25565,N_24454);
or U26303 (N_26303,N_25234,N_24342);
and U26304 (N_26304,N_25138,N_25948);
xnor U26305 (N_26305,N_24320,N_25215);
and U26306 (N_26306,N_24570,N_24231);
nand U26307 (N_26307,N_24100,N_24170);
and U26308 (N_26308,N_25728,N_24005);
or U26309 (N_26309,N_25168,N_25004);
or U26310 (N_26310,N_24481,N_24701);
and U26311 (N_26311,N_24892,N_25528);
or U26312 (N_26312,N_24035,N_25201);
or U26313 (N_26313,N_24864,N_25462);
xor U26314 (N_26314,N_25825,N_25447);
or U26315 (N_26315,N_24078,N_24689);
xor U26316 (N_26316,N_24584,N_25269);
or U26317 (N_26317,N_25128,N_25975);
xor U26318 (N_26318,N_24972,N_24743);
nor U26319 (N_26319,N_25796,N_25386);
and U26320 (N_26320,N_25257,N_24968);
or U26321 (N_26321,N_24521,N_25080);
and U26322 (N_26322,N_25167,N_25474);
nand U26323 (N_26323,N_24712,N_25677);
or U26324 (N_26324,N_25866,N_24004);
or U26325 (N_26325,N_24421,N_25794);
or U26326 (N_26326,N_24029,N_24051);
nand U26327 (N_26327,N_24515,N_25610);
xnor U26328 (N_26328,N_24561,N_25430);
and U26329 (N_26329,N_24054,N_24365);
nand U26330 (N_26330,N_25830,N_24745);
nor U26331 (N_26331,N_24401,N_24124);
xor U26332 (N_26332,N_24916,N_24728);
xnor U26333 (N_26333,N_25703,N_25429);
and U26334 (N_26334,N_25552,N_24470);
or U26335 (N_26335,N_24297,N_24513);
and U26336 (N_26336,N_24482,N_24965);
or U26337 (N_26337,N_24282,N_25326);
and U26338 (N_26338,N_24735,N_25741);
xor U26339 (N_26339,N_24961,N_24279);
nor U26340 (N_26340,N_25906,N_25500);
nor U26341 (N_26341,N_25196,N_25721);
and U26342 (N_26342,N_25989,N_25105);
or U26343 (N_26343,N_24407,N_25209);
xor U26344 (N_26344,N_24129,N_25119);
xor U26345 (N_26345,N_25575,N_25857);
nand U26346 (N_26346,N_25808,N_25727);
xnor U26347 (N_26347,N_24001,N_25896);
xor U26348 (N_26348,N_25301,N_25828);
xor U26349 (N_26349,N_25726,N_25186);
or U26350 (N_26350,N_25110,N_25027);
or U26351 (N_26351,N_25169,N_25084);
nor U26352 (N_26352,N_25289,N_24773);
and U26353 (N_26353,N_24469,N_24537);
or U26354 (N_26354,N_24175,N_24937);
nor U26355 (N_26355,N_25203,N_25918);
or U26356 (N_26356,N_24273,N_25188);
nand U26357 (N_26357,N_25083,N_24441);
and U26358 (N_26358,N_24729,N_25013);
xnor U26359 (N_26359,N_25942,N_25077);
xor U26360 (N_26360,N_25064,N_24013);
and U26361 (N_26361,N_25132,N_24704);
and U26362 (N_26362,N_25120,N_24844);
or U26363 (N_26363,N_25748,N_25032);
nand U26364 (N_26364,N_24417,N_25846);
xor U26365 (N_26365,N_25576,N_25171);
nand U26366 (N_26366,N_25787,N_25628);
xor U26367 (N_26367,N_25635,N_24212);
nand U26368 (N_26368,N_25876,N_25822);
or U26369 (N_26369,N_25299,N_24531);
xnor U26370 (N_26370,N_25141,N_25757);
nand U26371 (N_26371,N_25385,N_24885);
nor U26372 (N_26372,N_25103,N_25592);
xor U26373 (N_26373,N_24319,N_24510);
nand U26374 (N_26374,N_25030,N_25981);
nand U26375 (N_26375,N_24115,N_25800);
nand U26376 (N_26376,N_24251,N_24204);
or U26377 (N_26377,N_24841,N_24260);
and U26378 (N_26378,N_25210,N_25147);
and U26379 (N_26379,N_25593,N_25595);
nor U26380 (N_26380,N_24296,N_24506);
xor U26381 (N_26381,N_25775,N_24797);
xor U26382 (N_26382,N_25753,N_25176);
nand U26383 (N_26383,N_25855,N_25520);
nand U26384 (N_26384,N_24406,N_25835);
nand U26385 (N_26385,N_25075,N_25493);
nand U26386 (N_26386,N_25662,N_24891);
xor U26387 (N_26387,N_24015,N_25614);
and U26388 (N_26388,N_24829,N_25106);
xnor U26389 (N_26389,N_25288,N_24232);
nand U26390 (N_26390,N_25676,N_24111);
xnor U26391 (N_26391,N_24389,N_25543);
nand U26392 (N_26392,N_24875,N_24593);
or U26393 (N_26393,N_25879,N_25060);
nand U26394 (N_26394,N_25644,N_24612);
nand U26395 (N_26395,N_25724,N_24162);
nor U26396 (N_26396,N_24802,N_24998);
xnor U26397 (N_26397,N_25441,N_24952);
nand U26398 (N_26398,N_24022,N_24424);
xor U26399 (N_26399,N_24467,N_25569);
xnor U26400 (N_26400,N_25920,N_24127);
and U26401 (N_26401,N_25890,N_25490);
or U26402 (N_26402,N_24357,N_24473);
xor U26403 (N_26403,N_25713,N_25335);
nand U26404 (N_26404,N_24061,N_25139);
or U26405 (N_26405,N_24189,N_25737);
nor U26406 (N_26406,N_25657,N_25837);
and U26407 (N_26407,N_25481,N_25102);
nand U26408 (N_26408,N_25115,N_24912);
nand U26409 (N_26409,N_24854,N_25182);
xor U26410 (N_26410,N_25284,N_24544);
xnor U26411 (N_26411,N_24762,N_24245);
and U26412 (N_26412,N_24322,N_25479);
nand U26413 (N_26413,N_24276,N_24826);
nor U26414 (N_26414,N_25463,N_25653);
or U26415 (N_26415,N_25327,N_25328);
xnor U26416 (N_26416,N_25016,N_24557);
nor U26417 (N_26417,N_24795,N_25158);
and U26418 (N_26418,N_24463,N_25701);
nand U26419 (N_26419,N_24487,N_24253);
nand U26420 (N_26420,N_24101,N_24768);
or U26421 (N_26421,N_24538,N_25502);
nand U26422 (N_26422,N_25400,N_24852);
or U26423 (N_26423,N_24618,N_24497);
nand U26424 (N_26424,N_24603,N_25272);
xor U26425 (N_26425,N_24157,N_24356);
or U26426 (N_26426,N_24070,N_24446);
xnor U26427 (N_26427,N_25507,N_25097);
nand U26428 (N_26428,N_24631,N_24229);
or U26429 (N_26429,N_24915,N_24414);
and U26430 (N_26430,N_24989,N_25408);
and U26431 (N_26431,N_24369,N_25965);
or U26432 (N_26432,N_24079,N_24975);
nor U26433 (N_26433,N_24966,N_25179);
xor U26434 (N_26434,N_25159,N_25842);
or U26435 (N_26435,N_24117,N_25439);
and U26436 (N_26436,N_25880,N_25491);
or U26437 (N_26437,N_24723,N_25354);
nand U26438 (N_26438,N_24302,N_24740);
nand U26439 (N_26439,N_25648,N_25804);
or U26440 (N_26440,N_25583,N_25511);
nor U26441 (N_26441,N_24028,N_25613);
nand U26442 (N_26442,N_25629,N_25093);
or U26443 (N_26443,N_25599,N_25872);
nor U26444 (N_26444,N_25137,N_24536);
xnor U26445 (N_26445,N_24847,N_25715);
xor U26446 (N_26446,N_24432,N_24702);
and U26447 (N_26447,N_25003,N_24394);
or U26448 (N_26448,N_25033,N_24286);
nor U26449 (N_26449,N_24837,N_25853);
nand U26450 (N_26450,N_25448,N_24661);
or U26451 (N_26451,N_25694,N_25888);
xnor U26452 (N_26452,N_25801,N_25324);
nor U26453 (N_26453,N_25529,N_25514);
and U26454 (N_26454,N_24195,N_24694);
or U26455 (N_26455,N_24056,N_25329);
xnor U26456 (N_26456,N_24477,N_25449);
and U26457 (N_26457,N_25711,N_25440);
nand U26458 (N_26458,N_24883,N_24567);
or U26459 (N_26459,N_24783,N_24156);
or U26460 (N_26460,N_24849,N_24041);
nand U26461 (N_26461,N_24250,N_25545);
and U26462 (N_26462,N_24874,N_25509);
or U26463 (N_26463,N_24425,N_25001);
or U26464 (N_26464,N_25011,N_24988);
or U26465 (N_26465,N_25839,N_24788);
nand U26466 (N_26466,N_25887,N_25344);
nor U26467 (N_26467,N_25450,N_25416);
and U26468 (N_26468,N_25687,N_25009);
nor U26469 (N_26469,N_25740,N_25208);
or U26470 (N_26470,N_24511,N_24094);
xor U26471 (N_26471,N_24518,N_25752);
or U26472 (N_26472,N_24688,N_25250);
and U26473 (N_26473,N_24280,N_24428);
or U26474 (N_26474,N_24219,N_25155);
or U26475 (N_26475,N_24190,N_24484);
nor U26476 (N_26476,N_24636,N_24530);
or U26477 (N_26477,N_25229,N_25221);
or U26478 (N_26478,N_24742,N_24651);
or U26479 (N_26479,N_24569,N_25020);
nor U26480 (N_26480,N_24154,N_25841);
nand U26481 (N_26481,N_24724,N_24201);
nor U26482 (N_26482,N_25294,N_24782);
and U26483 (N_26483,N_24384,N_25885);
nand U26484 (N_26484,N_25517,N_24786);
and U26485 (N_26485,N_25173,N_25418);
or U26486 (N_26486,N_25759,N_24920);
xnor U26487 (N_26487,N_24827,N_25698);
and U26488 (N_26488,N_25777,N_25542);
xor U26489 (N_26489,N_25309,N_25818);
nor U26490 (N_26490,N_24318,N_25938);
nand U26491 (N_26491,N_24650,N_24335);
xor U26492 (N_26492,N_24679,N_25992);
or U26493 (N_26493,N_25052,N_25691);
or U26494 (N_26494,N_25725,N_24082);
nor U26495 (N_26495,N_24880,N_25303);
or U26496 (N_26496,N_25012,N_24225);
xor U26497 (N_26497,N_25358,N_24617);
or U26498 (N_26498,N_25671,N_25636);
or U26499 (N_26499,N_25002,N_25098);
xor U26500 (N_26500,N_24504,N_25164);
or U26501 (N_26501,N_25774,N_24816);
and U26502 (N_26502,N_24420,N_25123);
nand U26503 (N_26503,N_25410,N_25277);
and U26504 (N_26504,N_24971,N_24491);
xnor U26505 (N_26505,N_24341,N_25784);
nor U26506 (N_26506,N_25402,N_25391);
nand U26507 (N_26507,N_24171,N_24581);
and U26508 (N_26508,N_25506,N_25526);
and U26509 (N_26509,N_25874,N_24464);
xor U26510 (N_26510,N_25338,N_24922);
nor U26511 (N_26511,N_25779,N_24751);
xnor U26512 (N_26512,N_24674,N_25823);
nor U26513 (N_26513,N_25070,N_24294);
nand U26514 (N_26514,N_24062,N_25425);
and U26515 (N_26515,N_24468,N_24687);
nor U26516 (N_26516,N_24604,N_25190);
xor U26517 (N_26517,N_25519,N_24533);
nand U26518 (N_26518,N_24646,N_25995);
nor U26519 (N_26519,N_25684,N_25438);
xnor U26520 (N_26520,N_24027,N_24437);
nand U26521 (N_26521,N_25977,N_24289);
nor U26522 (N_26522,N_25302,N_24091);
xor U26523 (N_26523,N_24024,N_25031);
or U26524 (N_26524,N_24939,N_25074);
or U26525 (N_26525,N_25609,N_24643);
nor U26526 (N_26526,N_24479,N_24040);
and U26527 (N_26527,N_24137,N_24970);
or U26528 (N_26528,N_24552,N_24776);
and U26529 (N_26529,N_24360,N_24551);
nor U26530 (N_26530,N_25401,N_25650);
or U26531 (N_26531,N_24404,N_24991);
nor U26532 (N_26532,N_24149,N_25927);
nand U26533 (N_26533,N_24833,N_25772);
nand U26534 (N_26534,N_24718,N_25322);
or U26535 (N_26535,N_25663,N_25521);
xor U26536 (N_26536,N_24186,N_25767);
nand U26537 (N_26537,N_24867,N_24392);
and U26538 (N_26538,N_25988,N_25788);
or U26539 (N_26539,N_24870,N_24707);
xor U26540 (N_26540,N_25243,N_25187);
nor U26541 (N_26541,N_24416,N_25926);
xor U26542 (N_26542,N_25765,N_24823);
nor U26543 (N_26543,N_25317,N_25398);
and U26544 (N_26544,N_24131,N_25466);
and U26545 (N_26545,N_25352,N_24456);
and U26546 (N_26546,N_25803,N_25045);
nor U26547 (N_26547,N_25197,N_24371);
and U26548 (N_26548,N_24462,N_25283);
xnor U26549 (N_26549,N_25585,N_25810);
nand U26550 (N_26550,N_24188,N_24668);
nor U26551 (N_26551,N_24486,N_24512);
or U26552 (N_26552,N_25572,N_25549);
and U26553 (N_26553,N_25573,N_25530);
xor U26554 (N_26554,N_24653,N_25710);
and U26555 (N_26555,N_25382,N_24206);
xor U26556 (N_26556,N_24691,N_25731);
or U26557 (N_26557,N_24749,N_25086);
and U26558 (N_26558,N_25730,N_24676);
and U26559 (N_26559,N_25963,N_24564);
nand U26560 (N_26560,N_24220,N_24057);
and U26561 (N_26561,N_25471,N_25127);
xnor U26562 (N_26562,N_24907,N_25265);
or U26563 (N_26563,N_24143,N_24838);
nand U26564 (N_26564,N_24380,N_25395);
nand U26565 (N_26565,N_25555,N_24271);
and U26566 (N_26566,N_25377,N_25820);
xor U26567 (N_26567,N_24820,N_24693);
and U26568 (N_26568,N_24944,N_25939);
and U26569 (N_26569,N_24008,N_24123);
or U26570 (N_26570,N_25414,N_24492);
and U26571 (N_26571,N_24355,N_24438);
nor U26572 (N_26572,N_24752,N_24268);
xnor U26573 (N_26573,N_24628,N_24753);
nand U26574 (N_26574,N_24673,N_24525);
or U26575 (N_26575,N_25305,N_24605);
or U26576 (N_26576,N_25185,N_24248);
or U26577 (N_26577,N_25006,N_24607);
and U26578 (N_26578,N_25478,N_24197);
and U26579 (N_26579,N_24546,N_25140);
nor U26580 (N_26580,N_25089,N_25570);
nand U26581 (N_26581,N_24103,N_24120);
or U26582 (N_26582,N_25623,N_25889);
xor U26583 (N_26583,N_24583,N_25626);
nor U26584 (N_26584,N_25900,N_25768);
nor U26585 (N_26585,N_25172,N_24244);
and U26586 (N_26586,N_24373,N_25348);
xor U26587 (N_26587,N_24905,N_24860);
nand U26588 (N_26588,N_25817,N_24313);
or U26589 (N_26589,N_24614,N_25902);
nand U26590 (N_26590,N_25238,N_24152);
and U26591 (N_26591,N_24215,N_25157);
nand U26592 (N_26592,N_25390,N_25667);
xor U26593 (N_26593,N_24866,N_25966);
and U26594 (N_26594,N_25762,N_24060);
or U26595 (N_26595,N_25435,N_24247);
and U26596 (N_26596,N_25144,N_24807);
and U26597 (N_26597,N_24767,N_24736);
and U26598 (N_26598,N_25373,N_24052);
nand U26599 (N_26599,N_24903,N_25399);
nor U26600 (N_26600,N_25346,N_24025);
nand U26601 (N_26601,N_24439,N_25312);
nor U26602 (N_26602,N_25287,N_25242);
or U26603 (N_26603,N_25845,N_24199);
nor U26604 (N_26604,N_24293,N_24338);
and U26605 (N_26605,N_25706,N_25170);
nand U26606 (N_26606,N_24259,N_24696);
or U26607 (N_26607,N_25360,N_24960);
and U26608 (N_26608,N_25640,N_25912);
nor U26609 (N_26609,N_25498,N_24997);
and U26610 (N_26610,N_24792,N_25756);
nand U26611 (N_26611,N_24096,N_25298);
nand U26612 (N_26612,N_25524,N_24308);
or U26613 (N_26613,N_25838,N_24747);
nand U26614 (N_26614,N_24076,N_25670);
or U26615 (N_26615,N_24523,N_24485);
xor U26616 (N_26616,N_24478,N_24136);
nand U26617 (N_26617,N_25783,N_24325);
and U26618 (N_26618,N_24933,N_25292);
and U26619 (N_26619,N_24419,N_24488);
nor U26620 (N_26620,N_24012,N_24064);
xnor U26621 (N_26621,N_25073,N_25078);
xnor U26622 (N_26622,N_24333,N_24000);
and U26623 (N_26623,N_25122,N_24058);
nand U26624 (N_26624,N_25655,N_24621);
and U26625 (N_26625,N_24580,N_24911);
or U26626 (N_26626,N_25903,N_25058);
nor U26627 (N_26627,N_24183,N_25212);
nand U26628 (N_26628,N_25262,N_25055);
or U26629 (N_26629,N_24381,N_24637);
xnor U26630 (N_26630,N_25547,N_25090);
nand U26631 (N_26631,N_25806,N_25652);
nor U26632 (N_26632,N_24824,N_24522);
nor U26633 (N_26633,N_24348,N_24708);
nor U26634 (N_26634,N_24798,N_24411);
and U26635 (N_26635,N_25616,N_24007);
or U26636 (N_26636,N_24949,N_25379);
and U26637 (N_26637,N_25954,N_24956);
and U26638 (N_26638,N_25124,N_25567);
and U26639 (N_26639,N_24207,N_25844);
xor U26640 (N_26640,N_25633,N_25241);
nor U26641 (N_26641,N_25014,N_25459);
nor U26642 (N_26642,N_24181,N_24529);
and U26643 (N_26643,N_24309,N_24460);
nand U26644 (N_26644,N_24779,N_25413);
nand U26645 (N_26645,N_24494,N_24507);
or U26646 (N_26646,N_24769,N_25432);
and U26647 (N_26647,N_24967,N_25858);
and U26648 (N_26648,N_25056,N_25702);
and U26649 (N_26649,N_24606,N_25381);
or U26650 (N_26650,N_24092,N_25343);
and U26651 (N_26651,N_24926,N_24813);
xor U26652 (N_26652,N_24558,N_25827);
and U26653 (N_26653,N_25617,N_25018);
or U26654 (N_26654,N_24142,N_24686);
xnor U26655 (N_26655,N_24083,N_25160);
nand U26656 (N_26656,N_24121,N_25909);
or U26657 (N_26657,N_24819,N_24938);
and U26658 (N_26658,N_25364,N_25537);
nor U26659 (N_26659,N_24927,N_25525);
or U26660 (N_26660,N_25306,N_25222);
and U26661 (N_26661,N_24706,N_24932);
or U26662 (N_26662,N_25805,N_25356);
or U26663 (N_26663,N_24993,N_25072);
and U26664 (N_26664,N_24400,N_25240);
xnor U26665 (N_26665,N_24213,N_25915);
and U26666 (N_26666,N_24158,N_24349);
nor U26667 (N_26667,N_24053,N_24794);
nand U26668 (N_26668,N_24009,N_25869);
nand U26669 (N_26669,N_24408,N_24943);
and U26670 (N_26670,N_24897,N_25152);
nor U26671 (N_26671,N_25936,N_25814);
nand U26672 (N_26672,N_25993,N_25870);
nand U26673 (N_26673,N_24471,N_24159);
or U26674 (N_26674,N_25584,N_24198);
nand U26675 (N_26675,N_24925,N_25486);
and U26676 (N_26676,N_24817,N_25532);
xnor U26677 (N_26677,N_24719,N_25705);
and U26678 (N_26678,N_25404,N_24884);
nand U26679 (N_26679,N_25602,N_25940);
xnor U26680 (N_26680,N_24490,N_24266);
xnor U26681 (N_26681,N_24955,N_24962);
nand U26682 (N_26682,N_24711,N_24238);
nor U26683 (N_26683,N_24254,N_25174);
xor U26684 (N_26684,N_25630,N_24528);
nand U26685 (N_26685,N_24436,N_24608);
nor U26686 (N_26686,N_25443,N_25028);
or U26687 (N_26687,N_24272,N_24726);
nand U26688 (N_26688,N_24334,N_25578);
nor U26689 (N_26689,N_24452,N_24638);
nand U26690 (N_26690,N_24388,N_24941);
nor U26691 (N_26691,N_25862,N_25540);
nand U26692 (N_26692,N_24516,N_25736);
or U26693 (N_26693,N_25260,N_24936);
xnor U26694 (N_26694,N_25598,N_24295);
nor U26695 (N_26695,N_25742,N_25252);
nor U26696 (N_26696,N_24145,N_25816);
nand U26697 (N_26697,N_25997,N_25919);
or U26698 (N_26698,N_25884,N_24663);
xnor U26699 (N_26699,N_24842,N_25149);
and U26700 (N_26700,N_24214,N_24615);
nand U26701 (N_26701,N_24924,N_24586);
xnor U26702 (N_26702,N_24992,N_25503);
and U26703 (N_26703,N_25563,N_24275);
and U26704 (N_26704,N_24830,N_24393);
and U26705 (N_26705,N_24144,N_25681);
or U26706 (N_26706,N_25353,N_25579);
nand U26707 (N_26707,N_24900,N_24756);
nor U26708 (N_26708,N_24641,N_25898);
and U26709 (N_26709,N_24560,N_24535);
and U26710 (N_26710,N_25249,N_24700);
or U26711 (N_26711,N_24697,N_24744);
nor U26712 (N_26712,N_24543,N_24898);
xnor U26713 (N_26713,N_25351,N_25922);
and U26714 (N_26714,N_24304,N_25848);
nand U26715 (N_26715,N_24665,N_25051);
nor U26716 (N_26716,N_24194,N_25495);
xnor U26717 (N_26717,N_25522,N_25945);
nor U26718 (N_26718,N_24559,N_25943);
and U26719 (N_26719,N_25659,N_25359);
and U26720 (N_26720,N_25023,N_25181);
nor U26721 (N_26721,N_24541,N_25258);
or U26722 (N_26722,N_25405,N_25469);
and U26723 (N_26723,N_24787,N_25596);
nand U26724 (N_26724,N_25336,N_24090);
nor U26725 (N_26725,N_25082,N_25333);
and U26726 (N_26726,N_25550,N_25875);
and U26727 (N_26727,N_24274,N_25949);
xor U26728 (N_26728,N_24669,N_24713);
or U26729 (N_26729,N_24804,N_25423);
nand U26730 (N_26730,N_25518,N_25464);
nand U26731 (N_26731,N_24375,N_25069);
nor U26732 (N_26732,N_24113,N_24565);
xnor U26733 (N_26733,N_24909,N_25334);
nor U26734 (N_26734,N_25935,N_24398);
nand U26735 (N_26735,N_25465,N_24877);
nand U26736 (N_26736,N_24095,N_24362);
and U26737 (N_26737,N_24554,N_25365);
xnor U26738 (N_26738,N_25068,N_25645);
and U26739 (N_26739,N_25057,N_25646);
nor U26740 (N_26740,N_24264,N_25970);
nand U26741 (N_26741,N_24562,N_24765);
and U26742 (N_26742,N_24385,N_25821);
and U26743 (N_26743,N_24929,N_24645);
nor U26744 (N_26744,N_24894,N_24935);
nand U26745 (N_26745,N_24493,N_25293);
and U26746 (N_26746,N_25026,N_25729);
xor U26747 (N_26747,N_25733,N_25955);
or U26748 (N_26748,N_24639,N_25247);
xnor U26749 (N_26749,N_25059,N_25864);
xnor U26750 (N_26750,N_24917,N_24382);
nor U26751 (N_26751,N_25130,N_24148);
nand U26752 (N_26752,N_24640,N_24140);
or U26753 (N_26753,N_25177,N_25849);
nand U26754 (N_26754,N_24453,N_24023);
xnor U26755 (N_26755,N_24660,N_24576);
nor U26756 (N_26756,N_24805,N_24588);
or U26757 (N_26757,N_25994,N_24166);
nor U26758 (N_26758,N_24019,N_24075);
and U26759 (N_26759,N_24946,N_25990);
nor U26760 (N_26760,N_24950,N_24886);
xnor U26761 (N_26761,N_24107,N_24764);
or U26762 (N_26762,N_24002,N_24821);
or U26763 (N_26763,N_24784,N_24185);
and U26764 (N_26764,N_25852,N_25877);
xnor U26765 (N_26765,N_25770,N_25388);
nor U26766 (N_26766,N_25076,N_24466);
nand U26767 (N_26767,N_24134,N_25142);
and U26768 (N_26768,N_25580,N_24692);
xor U26769 (N_26769,N_25008,N_25991);
or U26770 (N_26770,N_24037,N_25296);
and U26771 (N_26771,N_24376,N_25280);
xnor U26772 (N_26772,N_25832,N_25622);
and U26773 (N_26773,N_24044,N_25040);
nor U26774 (N_26774,N_25781,N_24359);
or U26775 (N_26775,N_24626,N_24258);
and U26776 (N_26776,N_25150,N_24475);
or U26777 (N_26777,N_24146,N_24763);
nand U26778 (N_26778,N_25680,N_25175);
xnor U26779 (N_26779,N_25916,N_24613);
nand U26780 (N_26780,N_25178,N_25492);
xnor U26781 (N_26781,N_25591,N_25467);
or U26782 (N_26782,N_25615,N_24990);
nor U26783 (N_26783,N_25112,N_25007);
and U26784 (N_26784,N_24625,N_24964);
or U26785 (N_26785,N_25601,N_24049);
or U26786 (N_26786,N_24940,N_25815);
or U26787 (N_26787,N_25707,N_25297);
or U26788 (N_26788,N_24634,N_24018);
and U26789 (N_26789,N_24099,N_24652);
nand U26790 (N_26790,N_25735,N_24086);
or U26791 (N_26791,N_25458,N_24352);
or U26792 (N_26792,N_25369,N_25017);
xnor U26793 (N_26793,N_24647,N_24358);
nor U26794 (N_26794,N_25738,N_24984);
nor U26795 (N_26795,N_24609,N_25088);
nor U26796 (N_26796,N_25363,N_25968);
xor U26797 (N_26797,N_25561,N_25036);
or U26798 (N_26798,N_24755,N_24068);
nor U26799 (N_26799,N_25230,N_25442);
or U26800 (N_26800,N_25709,N_24722);
or U26801 (N_26801,N_25285,N_24370);
nor U26802 (N_26802,N_25755,N_25219);
xor U26803 (N_26803,N_24331,N_25953);
xor U26804 (N_26804,N_24733,N_25050);
nor U26805 (N_26805,N_24667,N_25129);
nor U26806 (N_26806,N_25544,N_25510);
or U26807 (N_26807,N_25087,N_25723);
or U26808 (N_26808,N_24895,N_25679);
nand U26809 (N_26809,N_25960,N_25231);
nand U26810 (N_26810,N_24973,N_24483);
and U26811 (N_26811,N_25136,N_25248);
or U26812 (N_26812,N_25582,N_25372);
nor U26813 (N_26813,N_25409,N_24954);
or U26814 (N_26814,N_25621,N_25470);
nand U26815 (N_26815,N_25042,N_24627);
and U26816 (N_26816,N_24716,N_25362);
or U26817 (N_26817,N_25349,N_25383);
nor U26818 (N_26818,N_25393,N_25624);
xor U26819 (N_26819,N_24585,N_25904);
nor U26820 (N_26820,N_25198,N_25350);
and U26821 (N_26821,N_25618,N_25950);
or U26822 (N_26822,N_24399,N_25859);
or U26823 (N_26823,N_24315,N_24065);
and U26824 (N_26824,N_24754,N_24888);
nand U26825 (N_26825,N_24503,N_24346);
xor U26826 (N_26826,N_25778,N_25672);
nor U26827 (N_26827,N_24902,N_24125);
nand U26828 (N_26828,N_24391,N_25669);
and U26829 (N_26829,N_24921,N_25318);
nor U26830 (N_26830,N_25661,N_25113);
xor U26831 (N_26831,N_25947,N_25044);
nor U26832 (N_26832,N_25049,N_24457);
and U26833 (N_26833,N_25126,N_24526);
and U26834 (N_26834,N_25397,N_25697);
nand U26835 (N_26835,N_24596,N_24549);
nand U26836 (N_26836,N_24252,N_25512);
xor U26837 (N_26837,N_25607,N_24430);
and U26838 (N_26838,N_25192,N_25892);
nor U26839 (N_26839,N_25504,N_25882);
or U26840 (N_26840,N_24524,N_24730);
xnor U26841 (N_26841,N_25571,N_24077);
or U26842 (N_26842,N_25996,N_24859);
nand U26843 (N_26843,N_24455,N_24602);
xor U26844 (N_26844,N_24105,N_24339);
xnor U26845 (N_26845,N_25029,N_25739);
or U26846 (N_26846,N_25937,N_24725);
and U26847 (N_26847,N_25005,N_24221);
nor U26848 (N_26848,N_24720,N_24801);
and U26849 (N_26849,N_24808,N_25275);
nand U26850 (N_26850,N_24228,N_24292);
or U26851 (N_26851,N_24218,N_25969);
or U26852 (N_26852,N_25712,N_25422);
or U26853 (N_26853,N_24680,N_25984);
or U26854 (N_26854,N_24906,N_24869);
nor U26855 (N_26855,N_25281,N_25931);
or U26856 (N_26856,N_25295,N_25307);
or U26857 (N_26857,N_24715,N_25538);
nand U26858 (N_26858,N_25660,N_24656);
and U26859 (N_26859,N_25523,N_25568);
or U26860 (N_26860,N_25259,N_25254);
nand U26861 (N_26861,N_24517,N_24709);
nand U26862 (N_26862,N_25534,N_25826);
and U26863 (N_26863,N_24868,N_24180);
or U26864 (N_26864,N_25812,N_24982);
or U26865 (N_26865,N_25987,N_24799);
xnor U26866 (N_26866,N_25114,N_24366);
or U26867 (N_26867,N_25924,N_24305);
xnor U26868 (N_26868,N_25419,N_24098);
nand U26869 (N_26869,N_24781,N_24151);
or U26870 (N_26870,N_24672,N_24328);
or U26871 (N_26871,N_25554,N_24327);
nand U26872 (N_26872,N_25553,N_24300);
or U26873 (N_26873,N_24623,N_24505);
nand U26874 (N_26874,N_24038,N_25560);
or U26875 (N_26875,N_25795,N_25204);
nor U26876 (N_26876,N_24431,N_24857);
nand U26877 (N_26877,N_25010,N_24815);
and U26878 (N_26878,N_24118,N_24999);
nor U26879 (N_26879,N_24353,N_24443);
and U26880 (N_26880,N_25957,N_24671);
nand U26881 (N_26881,N_25714,N_24032);
or U26882 (N_26882,N_25151,N_24575);
xor U26883 (N_26883,N_25101,N_25131);
or U26884 (N_26884,N_24957,N_25426);
and U26885 (N_26885,N_24472,N_25477);
or U26886 (N_26886,N_25581,N_25342);
or U26887 (N_26887,N_24974,N_24540);
or U26888 (N_26888,N_25750,N_25085);
nor U26889 (N_26889,N_24684,N_24418);
or U26890 (N_26890,N_25913,N_25851);
and U26891 (N_26891,N_24163,N_25091);
and U26892 (N_26892,N_24865,N_25642);
nor U26893 (N_26893,N_24695,N_25674);
nor U26894 (N_26894,N_25799,N_24287);
nor U26895 (N_26895,N_24945,N_25811);
and U26896 (N_26896,N_25608,N_25094);
and U26897 (N_26897,N_25389,N_24050);
nor U26898 (N_26898,N_24332,N_25015);
or U26899 (N_26899,N_24914,N_24871);
nand U26900 (N_26900,N_25228,N_24321);
nand U26901 (N_26901,N_24994,N_24923);
or U26902 (N_26902,N_25747,N_25251);
or U26903 (N_26903,N_24846,N_24368);
and U26904 (N_26904,N_24155,N_24737);
nor U26905 (N_26905,N_25341,N_24899);
or U26906 (N_26906,N_25649,N_25603);
nand U26907 (N_26907,N_25686,N_24434);
nor U26908 (N_26908,N_24658,N_24278);
nor U26909 (N_26909,N_25941,N_25472);
and U26910 (N_26910,N_24344,N_24363);
nor U26911 (N_26911,N_24106,N_25291);
or U26912 (N_26912,N_25717,N_24648);
nor U26913 (N_26913,N_24806,N_25370);
and U26914 (N_26914,N_24675,N_25046);
nand U26915 (N_26915,N_24257,N_25833);
nand U26916 (N_26916,N_25899,N_24071);
nor U26917 (N_26917,N_24444,N_24717);
or U26918 (N_26918,N_25436,N_24721);
or U26919 (N_26919,N_25484,N_24659);
or U26920 (N_26920,N_25760,N_24969);
nand U26921 (N_26921,N_24498,N_24132);
and U26922 (N_26922,N_25980,N_25871);
or U26923 (N_26923,N_24203,N_25789);
nor U26924 (N_26924,N_25678,N_25637);
and U26925 (N_26925,N_25974,N_24495);
or U26926 (N_26926,N_25392,N_24409);
and U26927 (N_26927,N_25320,N_24390);
xor U26928 (N_26928,N_25255,N_24047);
nand U26929 (N_26929,N_25773,N_25095);
and U26930 (N_26930,N_24351,N_24261);
nor U26931 (N_26931,N_25891,N_24374);
or U26932 (N_26932,N_25332,N_24006);
nand U26933 (N_26933,N_24811,N_25266);
and U26934 (N_26934,N_24377,N_24191);
nand U26935 (N_26935,N_25205,N_25183);
and U26936 (N_26936,N_25412,N_24088);
or U26937 (N_26937,N_24256,N_24153);
nand U26938 (N_26938,N_24336,N_25407);
nand U26939 (N_26939,N_24435,N_25468);
nand U26940 (N_26940,N_25043,N_25485);
xor U26941 (N_26941,N_24587,N_24839);
nand U26942 (N_26942,N_25274,N_25232);
nor U26943 (N_26943,N_25433,N_25480);
nor U26944 (N_26944,N_24176,N_24662);
and U26945 (N_26945,N_25053,N_24496);
or U26946 (N_26946,N_24928,N_24011);
nor U26947 (N_26947,N_24445,N_24553);
nand U26948 (N_26948,N_24442,N_24202);
nor U26949 (N_26949,N_24403,N_25973);
and U26950 (N_26950,N_25331,N_25071);
xor U26951 (N_26951,N_24995,N_25216);
nor U26952 (N_26952,N_25189,N_25417);
or U26953 (N_26953,N_25061,N_24269);
nand U26954 (N_26954,N_24834,N_25689);
xor U26955 (N_26955,N_25270,N_25321);
or U26956 (N_26956,N_24597,N_24780);
or U26957 (N_26957,N_24828,N_25539);
or U26958 (N_26958,N_25330,N_25627);
xnor U26959 (N_26959,N_24611,N_25643);
or U26960 (N_26960,N_24290,N_25048);
nand U26961 (N_26961,N_25824,N_25577);
xnor U26962 (N_26962,N_24771,N_24474);
nor U26963 (N_26963,N_24150,N_24449);
nand U26964 (N_26964,N_24748,N_24595);
or U26965 (N_26965,N_25893,N_25246);
nand U26966 (N_26966,N_25153,N_24367);
xor U26967 (N_26967,N_25323,N_25489);
nand U26968 (N_26968,N_24532,N_25985);
xnor U26969 (N_26969,N_25840,N_25732);
nand U26970 (N_26970,N_25437,N_24255);
xor U26971 (N_26971,N_25453,N_25268);
and U26972 (N_26972,N_25100,N_25454);
nand U26973 (N_26973,N_24690,N_25962);
and U26974 (N_26974,N_25881,N_25764);
and U26975 (N_26975,N_25665,N_24633);
nand U26976 (N_26976,N_24853,N_24983);
nand U26977 (N_26977,N_24545,N_25641);
and U26978 (N_26978,N_24734,N_24329);
or U26979 (N_26979,N_25668,N_25211);
nor U26980 (N_26980,N_24534,N_24179);
nor U26981 (N_26981,N_24093,N_24796);
xor U26982 (N_26982,N_24856,N_25536);
nor U26983 (N_26983,N_25311,N_25394);
and U26984 (N_26984,N_24677,N_25148);
nand U26985 (N_26985,N_24977,N_25782);
xnor U26986 (N_26986,N_24177,N_24563);
nor U26987 (N_26987,N_25854,N_25564);
or U26988 (N_26988,N_25946,N_25025);
nor U26989 (N_26989,N_25021,N_24243);
or U26990 (N_26990,N_24413,N_24589);
or U26991 (N_26991,N_24876,N_25499);
xor U26992 (N_26992,N_24187,N_24760);
xor U26993 (N_26993,N_24108,N_25340);
nor U26994 (N_26994,N_24350,N_25743);
or U26995 (N_26995,N_25688,N_24791);
xor U26996 (N_26996,N_25978,N_24230);
nor U26997 (N_26997,N_24130,N_24947);
xor U26998 (N_26998,N_24913,N_25790);
nor U26999 (N_26999,N_25785,N_24831);
or U27000 (N_27000,N_24964,N_24130);
nand U27001 (N_27001,N_25968,N_25640);
nand U27002 (N_27002,N_24265,N_24490);
and U27003 (N_27003,N_24811,N_24023);
or U27004 (N_27004,N_24810,N_25148);
and U27005 (N_27005,N_24227,N_25056);
or U27006 (N_27006,N_24738,N_24414);
nor U27007 (N_27007,N_25768,N_25501);
or U27008 (N_27008,N_25760,N_25192);
and U27009 (N_27009,N_25252,N_24681);
xor U27010 (N_27010,N_24179,N_24927);
or U27011 (N_27011,N_24073,N_25562);
xnor U27012 (N_27012,N_25543,N_24292);
nor U27013 (N_27013,N_25876,N_24732);
and U27014 (N_27014,N_25671,N_25379);
nor U27015 (N_27015,N_25136,N_25852);
nand U27016 (N_27016,N_24213,N_24809);
or U27017 (N_27017,N_25877,N_25332);
xnor U27018 (N_27018,N_24144,N_25809);
nand U27019 (N_27019,N_25207,N_25415);
or U27020 (N_27020,N_25412,N_25226);
or U27021 (N_27021,N_25993,N_25423);
nand U27022 (N_27022,N_24429,N_24606);
and U27023 (N_27023,N_24515,N_24418);
nor U27024 (N_27024,N_24423,N_25594);
xnor U27025 (N_27025,N_25967,N_24750);
nor U27026 (N_27026,N_25010,N_24319);
nand U27027 (N_27027,N_25404,N_25279);
nor U27028 (N_27028,N_25260,N_25187);
or U27029 (N_27029,N_24625,N_25113);
or U27030 (N_27030,N_24411,N_24725);
nor U27031 (N_27031,N_24942,N_25163);
nand U27032 (N_27032,N_24080,N_24652);
nor U27033 (N_27033,N_25772,N_25742);
nand U27034 (N_27034,N_25728,N_24480);
nor U27035 (N_27035,N_25307,N_24659);
and U27036 (N_27036,N_24012,N_24662);
and U27037 (N_27037,N_24317,N_25189);
nand U27038 (N_27038,N_24030,N_24455);
and U27039 (N_27039,N_25401,N_25375);
xnor U27040 (N_27040,N_25610,N_25390);
xor U27041 (N_27041,N_24118,N_25314);
nand U27042 (N_27042,N_25668,N_25904);
xnor U27043 (N_27043,N_25258,N_25403);
nor U27044 (N_27044,N_25177,N_25644);
xnor U27045 (N_27045,N_24214,N_24258);
and U27046 (N_27046,N_24069,N_25580);
xnor U27047 (N_27047,N_24228,N_24805);
or U27048 (N_27048,N_24363,N_24540);
nor U27049 (N_27049,N_25146,N_24431);
nand U27050 (N_27050,N_24701,N_25984);
nor U27051 (N_27051,N_25136,N_24982);
and U27052 (N_27052,N_25321,N_25977);
and U27053 (N_27053,N_25899,N_24537);
xnor U27054 (N_27054,N_24984,N_25961);
nor U27055 (N_27055,N_25179,N_25715);
xnor U27056 (N_27056,N_25175,N_25900);
and U27057 (N_27057,N_25459,N_25402);
or U27058 (N_27058,N_24080,N_25216);
or U27059 (N_27059,N_25413,N_24167);
xor U27060 (N_27060,N_24242,N_24022);
or U27061 (N_27061,N_24158,N_24155);
nand U27062 (N_27062,N_24821,N_24662);
and U27063 (N_27063,N_24634,N_25728);
xnor U27064 (N_27064,N_25356,N_25526);
xnor U27065 (N_27065,N_25842,N_24750);
xor U27066 (N_27066,N_25969,N_24921);
nand U27067 (N_27067,N_24366,N_25133);
xnor U27068 (N_27068,N_24619,N_24971);
nor U27069 (N_27069,N_24111,N_24732);
xnor U27070 (N_27070,N_24101,N_25703);
and U27071 (N_27071,N_25877,N_25910);
and U27072 (N_27072,N_25682,N_24116);
nand U27073 (N_27073,N_25589,N_24359);
nor U27074 (N_27074,N_25698,N_25874);
or U27075 (N_27075,N_24595,N_25810);
and U27076 (N_27076,N_25882,N_24642);
nor U27077 (N_27077,N_25961,N_25740);
or U27078 (N_27078,N_24189,N_25196);
and U27079 (N_27079,N_25811,N_25561);
or U27080 (N_27080,N_24456,N_25905);
and U27081 (N_27081,N_25512,N_25457);
nand U27082 (N_27082,N_25680,N_24188);
nor U27083 (N_27083,N_25428,N_25208);
nor U27084 (N_27084,N_25112,N_24686);
xor U27085 (N_27085,N_24973,N_25532);
nand U27086 (N_27086,N_25564,N_24372);
and U27087 (N_27087,N_25501,N_25752);
nor U27088 (N_27088,N_25819,N_25988);
or U27089 (N_27089,N_25150,N_24815);
nand U27090 (N_27090,N_25136,N_24546);
xnor U27091 (N_27091,N_24533,N_24416);
nand U27092 (N_27092,N_24082,N_24900);
and U27093 (N_27093,N_24152,N_25242);
nand U27094 (N_27094,N_24890,N_25231);
and U27095 (N_27095,N_24467,N_24349);
nand U27096 (N_27096,N_24521,N_25032);
nor U27097 (N_27097,N_25284,N_24568);
xnor U27098 (N_27098,N_24305,N_25241);
and U27099 (N_27099,N_24936,N_25299);
and U27100 (N_27100,N_24585,N_25564);
or U27101 (N_27101,N_24775,N_24129);
xnor U27102 (N_27102,N_24470,N_25280);
or U27103 (N_27103,N_24138,N_25459);
and U27104 (N_27104,N_24908,N_25087);
or U27105 (N_27105,N_24113,N_25957);
xor U27106 (N_27106,N_25415,N_24645);
nor U27107 (N_27107,N_24178,N_25451);
xnor U27108 (N_27108,N_25785,N_25213);
nor U27109 (N_27109,N_24496,N_25343);
and U27110 (N_27110,N_24358,N_24141);
nor U27111 (N_27111,N_24341,N_25922);
and U27112 (N_27112,N_24244,N_25273);
or U27113 (N_27113,N_25859,N_24554);
and U27114 (N_27114,N_25867,N_24419);
xor U27115 (N_27115,N_25324,N_24762);
or U27116 (N_27116,N_25289,N_24947);
nand U27117 (N_27117,N_25875,N_24717);
or U27118 (N_27118,N_24461,N_25066);
and U27119 (N_27119,N_24499,N_25847);
nor U27120 (N_27120,N_25283,N_25959);
nor U27121 (N_27121,N_25661,N_24709);
nor U27122 (N_27122,N_25766,N_24047);
xor U27123 (N_27123,N_25134,N_24394);
and U27124 (N_27124,N_25023,N_25390);
nand U27125 (N_27125,N_25377,N_25382);
and U27126 (N_27126,N_24472,N_25548);
nand U27127 (N_27127,N_24960,N_25543);
nand U27128 (N_27128,N_25132,N_25330);
and U27129 (N_27129,N_24255,N_24032);
and U27130 (N_27130,N_24845,N_24787);
or U27131 (N_27131,N_25542,N_24308);
nand U27132 (N_27132,N_24516,N_25737);
or U27133 (N_27133,N_24438,N_25979);
or U27134 (N_27134,N_25590,N_24160);
nand U27135 (N_27135,N_24748,N_24173);
and U27136 (N_27136,N_25835,N_24700);
or U27137 (N_27137,N_24637,N_24351);
xnor U27138 (N_27138,N_24649,N_24100);
or U27139 (N_27139,N_24779,N_24153);
xnor U27140 (N_27140,N_25692,N_24755);
or U27141 (N_27141,N_25831,N_25108);
or U27142 (N_27142,N_25976,N_25995);
nor U27143 (N_27143,N_24073,N_24770);
nor U27144 (N_27144,N_25893,N_24189);
and U27145 (N_27145,N_24851,N_24427);
nand U27146 (N_27146,N_24923,N_24194);
xnor U27147 (N_27147,N_24771,N_25822);
xor U27148 (N_27148,N_25396,N_25818);
and U27149 (N_27149,N_24651,N_24896);
xnor U27150 (N_27150,N_25167,N_24145);
nand U27151 (N_27151,N_25211,N_24332);
or U27152 (N_27152,N_24493,N_25167);
nor U27153 (N_27153,N_25959,N_25264);
nor U27154 (N_27154,N_24496,N_25807);
nor U27155 (N_27155,N_24360,N_25206);
xnor U27156 (N_27156,N_24881,N_24504);
xnor U27157 (N_27157,N_25783,N_24357);
and U27158 (N_27158,N_25987,N_24981);
and U27159 (N_27159,N_25451,N_24209);
nand U27160 (N_27160,N_25251,N_25295);
nand U27161 (N_27161,N_24565,N_24586);
and U27162 (N_27162,N_24925,N_24151);
nand U27163 (N_27163,N_24567,N_24552);
xor U27164 (N_27164,N_25145,N_25328);
and U27165 (N_27165,N_24514,N_24885);
nor U27166 (N_27166,N_25913,N_25646);
nor U27167 (N_27167,N_25646,N_25273);
nand U27168 (N_27168,N_25652,N_25747);
nor U27169 (N_27169,N_24731,N_25225);
or U27170 (N_27170,N_24466,N_25517);
nor U27171 (N_27171,N_24115,N_25111);
or U27172 (N_27172,N_25518,N_25319);
or U27173 (N_27173,N_25613,N_24360);
and U27174 (N_27174,N_25418,N_25147);
xnor U27175 (N_27175,N_25417,N_25048);
nor U27176 (N_27176,N_24854,N_25789);
xnor U27177 (N_27177,N_25531,N_25185);
xnor U27178 (N_27178,N_25873,N_24606);
nor U27179 (N_27179,N_25376,N_24718);
nand U27180 (N_27180,N_24640,N_24697);
xor U27181 (N_27181,N_25774,N_25323);
nand U27182 (N_27182,N_24035,N_24523);
nand U27183 (N_27183,N_25854,N_25593);
nor U27184 (N_27184,N_25780,N_24561);
and U27185 (N_27185,N_24281,N_25655);
nand U27186 (N_27186,N_25965,N_25142);
xor U27187 (N_27187,N_24144,N_24234);
and U27188 (N_27188,N_25969,N_24159);
nand U27189 (N_27189,N_25417,N_25156);
nand U27190 (N_27190,N_24503,N_24354);
nand U27191 (N_27191,N_25330,N_24070);
or U27192 (N_27192,N_24992,N_24467);
or U27193 (N_27193,N_24701,N_25932);
and U27194 (N_27194,N_24896,N_24333);
nor U27195 (N_27195,N_24897,N_25664);
or U27196 (N_27196,N_24182,N_24265);
nand U27197 (N_27197,N_25447,N_25686);
and U27198 (N_27198,N_24014,N_25577);
nand U27199 (N_27199,N_24651,N_25542);
or U27200 (N_27200,N_25647,N_24356);
nor U27201 (N_27201,N_25120,N_25586);
and U27202 (N_27202,N_25678,N_24790);
and U27203 (N_27203,N_25863,N_25682);
or U27204 (N_27204,N_24634,N_24778);
xnor U27205 (N_27205,N_24203,N_24269);
nor U27206 (N_27206,N_25096,N_25471);
or U27207 (N_27207,N_24175,N_24239);
xor U27208 (N_27208,N_24166,N_24864);
and U27209 (N_27209,N_25236,N_24756);
and U27210 (N_27210,N_24246,N_25406);
and U27211 (N_27211,N_25220,N_24988);
and U27212 (N_27212,N_24876,N_24180);
or U27213 (N_27213,N_25205,N_25635);
and U27214 (N_27214,N_24943,N_24035);
or U27215 (N_27215,N_25658,N_24019);
and U27216 (N_27216,N_25143,N_25035);
xor U27217 (N_27217,N_25026,N_25943);
nor U27218 (N_27218,N_24057,N_25698);
and U27219 (N_27219,N_24052,N_25678);
or U27220 (N_27220,N_25455,N_24280);
or U27221 (N_27221,N_25387,N_25960);
nor U27222 (N_27222,N_24940,N_24962);
nor U27223 (N_27223,N_25666,N_25251);
nand U27224 (N_27224,N_25681,N_25616);
and U27225 (N_27225,N_25714,N_25716);
nand U27226 (N_27226,N_24952,N_24069);
xor U27227 (N_27227,N_25901,N_24057);
and U27228 (N_27228,N_25191,N_24275);
and U27229 (N_27229,N_24661,N_25781);
xor U27230 (N_27230,N_25254,N_24714);
xnor U27231 (N_27231,N_24114,N_25567);
nor U27232 (N_27232,N_25642,N_25016);
nand U27233 (N_27233,N_25544,N_25409);
and U27234 (N_27234,N_25617,N_24603);
and U27235 (N_27235,N_25205,N_25372);
or U27236 (N_27236,N_24943,N_24876);
nor U27237 (N_27237,N_24255,N_25728);
or U27238 (N_27238,N_25164,N_25887);
and U27239 (N_27239,N_24245,N_24502);
and U27240 (N_27240,N_24432,N_24935);
nand U27241 (N_27241,N_24172,N_25057);
nand U27242 (N_27242,N_24938,N_24223);
and U27243 (N_27243,N_25248,N_24356);
and U27244 (N_27244,N_25021,N_24094);
nand U27245 (N_27245,N_24705,N_24127);
and U27246 (N_27246,N_24032,N_24660);
or U27247 (N_27247,N_25121,N_24505);
nor U27248 (N_27248,N_24277,N_25553);
nand U27249 (N_27249,N_24145,N_25112);
xor U27250 (N_27250,N_24463,N_25699);
nand U27251 (N_27251,N_25720,N_25741);
nand U27252 (N_27252,N_24424,N_24426);
or U27253 (N_27253,N_24536,N_25232);
or U27254 (N_27254,N_25309,N_25390);
and U27255 (N_27255,N_24702,N_25664);
and U27256 (N_27256,N_24895,N_24021);
nand U27257 (N_27257,N_24731,N_24782);
nor U27258 (N_27258,N_25636,N_24614);
and U27259 (N_27259,N_25270,N_25249);
and U27260 (N_27260,N_24470,N_25127);
xor U27261 (N_27261,N_24701,N_24124);
xor U27262 (N_27262,N_24501,N_25689);
and U27263 (N_27263,N_25056,N_24733);
nand U27264 (N_27264,N_25285,N_24260);
nor U27265 (N_27265,N_24604,N_24839);
nand U27266 (N_27266,N_25078,N_25018);
nor U27267 (N_27267,N_24668,N_25847);
and U27268 (N_27268,N_25407,N_25979);
nor U27269 (N_27269,N_24313,N_24909);
or U27270 (N_27270,N_24729,N_25136);
xor U27271 (N_27271,N_25491,N_25713);
or U27272 (N_27272,N_24675,N_24071);
and U27273 (N_27273,N_24954,N_24353);
and U27274 (N_27274,N_24952,N_25656);
nor U27275 (N_27275,N_24296,N_25110);
and U27276 (N_27276,N_24432,N_24717);
nor U27277 (N_27277,N_25459,N_25869);
or U27278 (N_27278,N_24381,N_25181);
nand U27279 (N_27279,N_25888,N_25301);
and U27280 (N_27280,N_25831,N_25464);
and U27281 (N_27281,N_25645,N_24499);
nand U27282 (N_27282,N_25196,N_25646);
nor U27283 (N_27283,N_24782,N_25580);
nand U27284 (N_27284,N_24353,N_25676);
and U27285 (N_27285,N_25287,N_24795);
xor U27286 (N_27286,N_24998,N_24294);
nand U27287 (N_27287,N_25524,N_24075);
nand U27288 (N_27288,N_25331,N_24730);
nor U27289 (N_27289,N_25778,N_24759);
and U27290 (N_27290,N_24091,N_24946);
or U27291 (N_27291,N_24763,N_25122);
and U27292 (N_27292,N_25391,N_25980);
xnor U27293 (N_27293,N_24328,N_25126);
and U27294 (N_27294,N_25041,N_24767);
nand U27295 (N_27295,N_24554,N_25567);
or U27296 (N_27296,N_24872,N_24315);
or U27297 (N_27297,N_24075,N_24740);
nor U27298 (N_27298,N_25109,N_25965);
or U27299 (N_27299,N_24835,N_25222);
nand U27300 (N_27300,N_24209,N_25939);
nor U27301 (N_27301,N_25947,N_25281);
nand U27302 (N_27302,N_24477,N_25923);
xnor U27303 (N_27303,N_24952,N_25969);
nand U27304 (N_27304,N_24580,N_24204);
nand U27305 (N_27305,N_25013,N_24817);
and U27306 (N_27306,N_24176,N_25687);
or U27307 (N_27307,N_24010,N_25501);
and U27308 (N_27308,N_25791,N_24870);
and U27309 (N_27309,N_24542,N_25736);
and U27310 (N_27310,N_25899,N_25352);
and U27311 (N_27311,N_25123,N_25611);
xnor U27312 (N_27312,N_24304,N_24375);
nor U27313 (N_27313,N_25385,N_24370);
nor U27314 (N_27314,N_24403,N_24494);
and U27315 (N_27315,N_24579,N_25699);
and U27316 (N_27316,N_24803,N_25661);
nand U27317 (N_27317,N_25276,N_25125);
or U27318 (N_27318,N_25257,N_24586);
or U27319 (N_27319,N_25118,N_24591);
xor U27320 (N_27320,N_24725,N_24314);
xor U27321 (N_27321,N_24753,N_25926);
or U27322 (N_27322,N_24521,N_25739);
xor U27323 (N_27323,N_25997,N_24680);
or U27324 (N_27324,N_25178,N_25477);
and U27325 (N_27325,N_24244,N_25605);
and U27326 (N_27326,N_24577,N_25825);
nor U27327 (N_27327,N_25001,N_24543);
nand U27328 (N_27328,N_24920,N_25694);
nor U27329 (N_27329,N_25063,N_25122);
nand U27330 (N_27330,N_24792,N_24128);
or U27331 (N_27331,N_24782,N_25003);
nand U27332 (N_27332,N_24534,N_25994);
and U27333 (N_27333,N_24333,N_24535);
nor U27334 (N_27334,N_24322,N_24812);
nor U27335 (N_27335,N_25061,N_24902);
xnor U27336 (N_27336,N_24993,N_25825);
xnor U27337 (N_27337,N_24193,N_25603);
or U27338 (N_27338,N_25438,N_24149);
and U27339 (N_27339,N_24123,N_25328);
or U27340 (N_27340,N_25249,N_25959);
nand U27341 (N_27341,N_25209,N_25744);
or U27342 (N_27342,N_25405,N_24527);
nor U27343 (N_27343,N_24507,N_24718);
and U27344 (N_27344,N_24082,N_24661);
xnor U27345 (N_27345,N_25705,N_24205);
or U27346 (N_27346,N_25550,N_25104);
nor U27347 (N_27347,N_24430,N_24522);
and U27348 (N_27348,N_25884,N_25708);
xor U27349 (N_27349,N_24864,N_24199);
or U27350 (N_27350,N_25896,N_24211);
xor U27351 (N_27351,N_25570,N_25345);
xor U27352 (N_27352,N_24858,N_25931);
xor U27353 (N_27353,N_24183,N_25565);
or U27354 (N_27354,N_25915,N_24190);
nor U27355 (N_27355,N_25270,N_25392);
nor U27356 (N_27356,N_24390,N_25706);
and U27357 (N_27357,N_25720,N_24141);
nor U27358 (N_27358,N_24303,N_25578);
or U27359 (N_27359,N_25799,N_25615);
or U27360 (N_27360,N_25201,N_25768);
nor U27361 (N_27361,N_25785,N_24280);
and U27362 (N_27362,N_24179,N_24492);
and U27363 (N_27363,N_25813,N_25503);
xor U27364 (N_27364,N_25277,N_25832);
xor U27365 (N_27365,N_25603,N_24421);
xor U27366 (N_27366,N_24290,N_25691);
xnor U27367 (N_27367,N_25990,N_25250);
xnor U27368 (N_27368,N_24571,N_24295);
nand U27369 (N_27369,N_24416,N_25776);
xnor U27370 (N_27370,N_24180,N_24499);
or U27371 (N_27371,N_24415,N_24589);
nand U27372 (N_27372,N_24294,N_24134);
xnor U27373 (N_27373,N_24191,N_24209);
nand U27374 (N_27374,N_25584,N_24744);
nand U27375 (N_27375,N_25497,N_24350);
nor U27376 (N_27376,N_24206,N_25293);
or U27377 (N_27377,N_25360,N_24282);
nor U27378 (N_27378,N_25146,N_24642);
or U27379 (N_27379,N_24371,N_25961);
and U27380 (N_27380,N_25317,N_24329);
xnor U27381 (N_27381,N_25746,N_24574);
nand U27382 (N_27382,N_24641,N_24697);
xor U27383 (N_27383,N_25668,N_25443);
nand U27384 (N_27384,N_24818,N_24082);
and U27385 (N_27385,N_25608,N_24314);
nand U27386 (N_27386,N_25569,N_25842);
nor U27387 (N_27387,N_24640,N_25736);
xor U27388 (N_27388,N_24675,N_24355);
nor U27389 (N_27389,N_24655,N_25579);
and U27390 (N_27390,N_24389,N_24608);
or U27391 (N_27391,N_25137,N_25262);
xnor U27392 (N_27392,N_25314,N_24742);
and U27393 (N_27393,N_25303,N_24865);
nor U27394 (N_27394,N_24914,N_24447);
nor U27395 (N_27395,N_25070,N_24210);
nand U27396 (N_27396,N_24926,N_25542);
and U27397 (N_27397,N_25391,N_25316);
or U27398 (N_27398,N_25468,N_25965);
or U27399 (N_27399,N_25501,N_25990);
nor U27400 (N_27400,N_24024,N_25909);
nand U27401 (N_27401,N_25704,N_24198);
nand U27402 (N_27402,N_24616,N_24065);
and U27403 (N_27403,N_25930,N_25830);
nand U27404 (N_27404,N_25206,N_25222);
or U27405 (N_27405,N_25703,N_24805);
nor U27406 (N_27406,N_25754,N_25227);
or U27407 (N_27407,N_24761,N_25491);
nor U27408 (N_27408,N_25573,N_25654);
nor U27409 (N_27409,N_24915,N_25120);
xnor U27410 (N_27410,N_24022,N_24339);
xor U27411 (N_27411,N_25451,N_25623);
or U27412 (N_27412,N_24578,N_24894);
nor U27413 (N_27413,N_25319,N_24735);
and U27414 (N_27414,N_24878,N_24178);
xor U27415 (N_27415,N_24907,N_24416);
and U27416 (N_27416,N_24390,N_25992);
and U27417 (N_27417,N_25608,N_25809);
xnor U27418 (N_27418,N_25512,N_24883);
and U27419 (N_27419,N_24450,N_25234);
or U27420 (N_27420,N_25204,N_24618);
and U27421 (N_27421,N_24325,N_24785);
and U27422 (N_27422,N_24470,N_25648);
nor U27423 (N_27423,N_24876,N_24574);
xor U27424 (N_27424,N_24098,N_24601);
and U27425 (N_27425,N_25819,N_25312);
xnor U27426 (N_27426,N_24662,N_25622);
nand U27427 (N_27427,N_25636,N_24139);
nor U27428 (N_27428,N_25765,N_24197);
xor U27429 (N_27429,N_24874,N_24246);
nand U27430 (N_27430,N_24868,N_25865);
or U27431 (N_27431,N_24300,N_24248);
nand U27432 (N_27432,N_25033,N_25061);
xnor U27433 (N_27433,N_25388,N_24333);
nor U27434 (N_27434,N_24903,N_24650);
and U27435 (N_27435,N_25449,N_25863);
xnor U27436 (N_27436,N_24379,N_24440);
or U27437 (N_27437,N_25625,N_25528);
nor U27438 (N_27438,N_24378,N_24168);
and U27439 (N_27439,N_24104,N_25819);
and U27440 (N_27440,N_24602,N_24637);
nor U27441 (N_27441,N_25967,N_24057);
nand U27442 (N_27442,N_25523,N_25383);
nor U27443 (N_27443,N_25776,N_24727);
xor U27444 (N_27444,N_25675,N_24964);
nand U27445 (N_27445,N_24589,N_24419);
and U27446 (N_27446,N_25673,N_24030);
or U27447 (N_27447,N_24236,N_24369);
nand U27448 (N_27448,N_25725,N_25922);
nand U27449 (N_27449,N_25087,N_24605);
nor U27450 (N_27450,N_24097,N_24584);
nand U27451 (N_27451,N_24236,N_24107);
nand U27452 (N_27452,N_25372,N_25287);
nand U27453 (N_27453,N_24792,N_25504);
nand U27454 (N_27454,N_24986,N_25351);
and U27455 (N_27455,N_25855,N_24656);
xnor U27456 (N_27456,N_25960,N_25681);
nand U27457 (N_27457,N_24165,N_24285);
or U27458 (N_27458,N_24369,N_24621);
nand U27459 (N_27459,N_24776,N_24936);
and U27460 (N_27460,N_24570,N_25986);
or U27461 (N_27461,N_25251,N_24766);
nand U27462 (N_27462,N_24039,N_24172);
or U27463 (N_27463,N_25756,N_24830);
or U27464 (N_27464,N_25670,N_25748);
nor U27465 (N_27465,N_25779,N_24563);
or U27466 (N_27466,N_24770,N_25903);
or U27467 (N_27467,N_25375,N_25186);
nand U27468 (N_27468,N_24221,N_25039);
and U27469 (N_27469,N_24866,N_25441);
and U27470 (N_27470,N_24316,N_25810);
and U27471 (N_27471,N_25812,N_24355);
nor U27472 (N_27472,N_25564,N_24414);
and U27473 (N_27473,N_24182,N_24544);
or U27474 (N_27474,N_25309,N_24012);
and U27475 (N_27475,N_24825,N_24925);
nand U27476 (N_27476,N_24740,N_24579);
or U27477 (N_27477,N_24770,N_25463);
nor U27478 (N_27478,N_24548,N_25766);
nor U27479 (N_27479,N_24821,N_24365);
or U27480 (N_27480,N_24720,N_24697);
or U27481 (N_27481,N_24835,N_25174);
nand U27482 (N_27482,N_24357,N_24196);
or U27483 (N_27483,N_25676,N_24794);
nor U27484 (N_27484,N_24335,N_25263);
nor U27485 (N_27485,N_25055,N_24232);
or U27486 (N_27486,N_24592,N_25988);
and U27487 (N_27487,N_25457,N_25692);
or U27488 (N_27488,N_25588,N_24471);
nand U27489 (N_27489,N_24945,N_25512);
and U27490 (N_27490,N_24599,N_25324);
xor U27491 (N_27491,N_25545,N_25750);
xor U27492 (N_27492,N_24380,N_24954);
and U27493 (N_27493,N_24357,N_25589);
or U27494 (N_27494,N_24666,N_24627);
xnor U27495 (N_27495,N_25899,N_25103);
or U27496 (N_27496,N_25528,N_24860);
xnor U27497 (N_27497,N_25284,N_24409);
and U27498 (N_27498,N_25744,N_24522);
or U27499 (N_27499,N_25513,N_24855);
and U27500 (N_27500,N_25849,N_24198);
xnor U27501 (N_27501,N_25382,N_24872);
and U27502 (N_27502,N_24678,N_24453);
xnor U27503 (N_27503,N_25615,N_25913);
and U27504 (N_27504,N_25709,N_25518);
and U27505 (N_27505,N_24687,N_25752);
or U27506 (N_27506,N_24002,N_24256);
or U27507 (N_27507,N_24592,N_24658);
xor U27508 (N_27508,N_24671,N_25836);
xnor U27509 (N_27509,N_24387,N_24121);
and U27510 (N_27510,N_24076,N_25909);
and U27511 (N_27511,N_25372,N_25204);
nand U27512 (N_27512,N_24725,N_24864);
xor U27513 (N_27513,N_25113,N_24645);
nor U27514 (N_27514,N_25688,N_25034);
or U27515 (N_27515,N_24578,N_24853);
nand U27516 (N_27516,N_24003,N_24125);
nor U27517 (N_27517,N_24139,N_24720);
xor U27518 (N_27518,N_24207,N_25685);
and U27519 (N_27519,N_24351,N_24281);
nand U27520 (N_27520,N_25073,N_25613);
xor U27521 (N_27521,N_25372,N_24367);
and U27522 (N_27522,N_24131,N_25863);
nand U27523 (N_27523,N_25577,N_24813);
nor U27524 (N_27524,N_25551,N_25251);
xor U27525 (N_27525,N_24708,N_24559);
nor U27526 (N_27526,N_25232,N_25198);
nand U27527 (N_27527,N_24800,N_24596);
nor U27528 (N_27528,N_24293,N_25767);
nor U27529 (N_27529,N_24833,N_24203);
xor U27530 (N_27530,N_25361,N_25657);
and U27531 (N_27531,N_25822,N_24139);
nand U27532 (N_27532,N_24173,N_24015);
nand U27533 (N_27533,N_25487,N_24724);
xnor U27534 (N_27534,N_25408,N_24388);
nand U27535 (N_27535,N_24763,N_25104);
xnor U27536 (N_27536,N_24585,N_25108);
nor U27537 (N_27537,N_24003,N_24020);
nor U27538 (N_27538,N_24933,N_25186);
nand U27539 (N_27539,N_25598,N_25278);
and U27540 (N_27540,N_25589,N_24212);
or U27541 (N_27541,N_24767,N_25663);
nor U27542 (N_27542,N_25619,N_24337);
xnor U27543 (N_27543,N_24080,N_25283);
and U27544 (N_27544,N_25455,N_24225);
and U27545 (N_27545,N_25757,N_24752);
nand U27546 (N_27546,N_25156,N_24228);
or U27547 (N_27547,N_25344,N_24120);
and U27548 (N_27548,N_24641,N_24356);
nor U27549 (N_27549,N_24292,N_24396);
nor U27550 (N_27550,N_25392,N_24553);
xor U27551 (N_27551,N_24561,N_24867);
or U27552 (N_27552,N_25693,N_25211);
xor U27553 (N_27553,N_24862,N_25266);
and U27554 (N_27554,N_25639,N_24710);
nor U27555 (N_27555,N_25199,N_25204);
nand U27556 (N_27556,N_24074,N_24494);
nor U27557 (N_27557,N_25829,N_24517);
xnor U27558 (N_27558,N_24469,N_25388);
nand U27559 (N_27559,N_25209,N_25636);
nand U27560 (N_27560,N_24055,N_25481);
xnor U27561 (N_27561,N_24945,N_24524);
xnor U27562 (N_27562,N_25127,N_25502);
nor U27563 (N_27563,N_24087,N_24854);
nand U27564 (N_27564,N_24807,N_25191);
nand U27565 (N_27565,N_24225,N_24030);
xnor U27566 (N_27566,N_25910,N_25950);
nand U27567 (N_27567,N_25855,N_24872);
and U27568 (N_27568,N_24476,N_24983);
and U27569 (N_27569,N_25375,N_25146);
and U27570 (N_27570,N_25423,N_24128);
and U27571 (N_27571,N_25579,N_24171);
nand U27572 (N_27572,N_25453,N_25820);
and U27573 (N_27573,N_25170,N_24444);
nand U27574 (N_27574,N_24092,N_24645);
and U27575 (N_27575,N_24471,N_25489);
xnor U27576 (N_27576,N_24404,N_24728);
xnor U27577 (N_27577,N_24045,N_25124);
nand U27578 (N_27578,N_25553,N_24184);
nand U27579 (N_27579,N_25329,N_24575);
and U27580 (N_27580,N_25782,N_25198);
nand U27581 (N_27581,N_24284,N_24731);
nand U27582 (N_27582,N_25972,N_25735);
and U27583 (N_27583,N_24069,N_24284);
and U27584 (N_27584,N_24264,N_24638);
and U27585 (N_27585,N_24883,N_24137);
nor U27586 (N_27586,N_24021,N_25332);
nor U27587 (N_27587,N_24709,N_24084);
or U27588 (N_27588,N_24216,N_25608);
nor U27589 (N_27589,N_25826,N_25082);
or U27590 (N_27590,N_25045,N_24431);
xnor U27591 (N_27591,N_24225,N_24509);
or U27592 (N_27592,N_24170,N_24696);
nand U27593 (N_27593,N_25323,N_24889);
or U27594 (N_27594,N_24379,N_25057);
nor U27595 (N_27595,N_25913,N_25156);
nand U27596 (N_27596,N_24575,N_24097);
nor U27597 (N_27597,N_25268,N_25990);
and U27598 (N_27598,N_24517,N_25405);
nor U27599 (N_27599,N_25972,N_24276);
nand U27600 (N_27600,N_25453,N_24246);
or U27601 (N_27601,N_25501,N_25827);
and U27602 (N_27602,N_25994,N_24170);
or U27603 (N_27603,N_25598,N_24277);
xnor U27604 (N_27604,N_25054,N_25398);
or U27605 (N_27605,N_24171,N_25147);
nor U27606 (N_27606,N_25103,N_25302);
or U27607 (N_27607,N_24210,N_24142);
xnor U27608 (N_27608,N_25235,N_24226);
xor U27609 (N_27609,N_24991,N_25314);
nand U27610 (N_27610,N_24369,N_25618);
xor U27611 (N_27611,N_24497,N_25729);
xnor U27612 (N_27612,N_25410,N_25325);
or U27613 (N_27613,N_25138,N_24757);
xor U27614 (N_27614,N_25697,N_24265);
and U27615 (N_27615,N_25521,N_25920);
nor U27616 (N_27616,N_25361,N_24995);
and U27617 (N_27617,N_25272,N_24235);
or U27618 (N_27618,N_24029,N_24645);
nand U27619 (N_27619,N_24939,N_25734);
or U27620 (N_27620,N_25273,N_25840);
or U27621 (N_27621,N_25762,N_25721);
and U27622 (N_27622,N_24728,N_24400);
nor U27623 (N_27623,N_24175,N_25096);
nand U27624 (N_27624,N_24396,N_25035);
xnor U27625 (N_27625,N_24423,N_24033);
and U27626 (N_27626,N_24271,N_25773);
and U27627 (N_27627,N_25748,N_24590);
xnor U27628 (N_27628,N_25482,N_24355);
nand U27629 (N_27629,N_24468,N_25316);
nand U27630 (N_27630,N_25386,N_24597);
and U27631 (N_27631,N_25044,N_24910);
and U27632 (N_27632,N_24731,N_24109);
nand U27633 (N_27633,N_24514,N_24635);
or U27634 (N_27634,N_25821,N_24701);
nand U27635 (N_27635,N_24181,N_24422);
or U27636 (N_27636,N_25270,N_25740);
nand U27637 (N_27637,N_25278,N_24332);
nor U27638 (N_27638,N_24165,N_25830);
xnor U27639 (N_27639,N_24643,N_24310);
and U27640 (N_27640,N_24735,N_25166);
nor U27641 (N_27641,N_25466,N_25722);
nand U27642 (N_27642,N_24937,N_25318);
and U27643 (N_27643,N_24537,N_24099);
nand U27644 (N_27644,N_24349,N_24075);
or U27645 (N_27645,N_25744,N_25822);
nand U27646 (N_27646,N_25541,N_25812);
nor U27647 (N_27647,N_25879,N_25381);
and U27648 (N_27648,N_24442,N_25413);
xor U27649 (N_27649,N_25303,N_24336);
xnor U27650 (N_27650,N_25052,N_25621);
nand U27651 (N_27651,N_25227,N_25824);
or U27652 (N_27652,N_24472,N_24332);
or U27653 (N_27653,N_24417,N_25979);
nor U27654 (N_27654,N_24413,N_25109);
and U27655 (N_27655,N_24768,N_24666);
nand U27656 (N_27656,N_25469,N_24731);
nor U27657 (N_27657,N_24857,N_24094);
nor U27658 (N_27658,N_24279,N_25705);
nand U27659 (N_27659,N_24773,N_24992);
nor U27660 (N_27660,N_25965,N_25844);
and U27661 (N_27661,N_25202,N_24135);
nor U27662 (N_27662,N_25246,N_25201);
nor U27663 (N_27663,N_25077,N_24024);
nand U27664 (N_27664,N_25814,N_24852);
nor U27665 (N_27665,N_25975,N_24374);
nor U27666 (N_27666,N_24519,N_24001);
and U27667 (N_27667,N_25351,N_25496);
xor U27668 (N_27668,N_25372,N_25977);
nor U27669 (N_27669,N_24072,N_25540);
nand U27670 (N_27670,N_24488,N_24404);
xor U27671 (N_27671,N_24417,N_24863);
nand U27672 (N_27672,N_25245,N_24681);
or U27673 (N_27673,N_24654,N_24604);
or U27674 (N_27674,N_24863,N_25353);
xor U27675 (N_27675,N_24016,N_25666);
nor U27676 (N_27676,N_25204,N_24802);
nand U27677 (N_27677,N_25938,N_24982);
nand U27678 (N_27678,N_24910,N_24060);
nor U27679 (N_27679,N_25048,N_24501);
nor U27680 (N_27680,N_25184,N_25941);
nor U27681 (N_27681,N_24653,N_24007);
nor U27682 (N_27682,N_24204,N_25299);
and U27683 (N_27683,N_24206,N_25202);
or U27684 (N_27684,N_24527,N_24108);
nand U27685 (N_27685,N_25172,N_25199);
and U27686 (N_27686,N_24996,N_25879);
xor U27687 (N_27687,N_25725,N_24542);
nand U27688 (N_27688,N_24940,N_25269);
nor U27689 (N_27689,N_24949,N_24118);
nor U27690 (N_27690,N_24901,N_25993);
nand U27691 (N_27691,N_24708,N_24920);
nand U27692 (N_27692,N_25393,N_25251);
nand U27693 (N_27693,N_24772,N_24444);
nand U27694 (N_27694,N_24292,N_24802);
nand U27695 (N_27695,N_24513,N_25500);
xnor U27696 (N_27696,N_24621,N_24556);
and U27697 (N_27697,N_25863,N_25974);
or U27698 (N_27698,N_24867,N_25537);
xnor U27699 (N_27699,N_25704,N_24242);
nand U27700 (N_27700,N_25004,N_24733);
nor U27701 (N_27701,N_24406,N_25329);
and U27702 (N_27702,N_24043,N_24195);
xnor U27703 (N_27703,N_24777,N_25221);
nand U27704 (N_27704,N_25326,N_25774);
nand U27705 (N_27705,N_24678,N_24152);
nand U27706 (N_27706,N_25056,N_24389);
nand U27707 (N_27707,N_24203,N_25471);
nor U27708 (N_27708,N_24919,N_25240);
nand U27709 (N_27709,N_25325,N_24899);
or U27710 (N_27710,N_24484,N_24184);
nor U27711 (N_27711,N_25831,N_24119);
or U27712 (N_27712,N_25895,N_24158);
or U27713 (N_27713,N_25450,N_25587);
xor U27714 (N_27714,N_25788,N_25486);
xnor U27715 (N_27715,N_24877,N_25777);
xnor U27716 (N_27716,N_25777,N_24361);
nand U27717 (N_27717,N_24007,N_25046);
and U27718 (N_27718,N_24260,N_24914);
xor U27719 (N_27719,N_25994,N_24916);
and U27720 (N_27720,N_25600,N_25421);
or U27721 (N_27721,N_24261,N_24292);
nand U27722 (N_27722,N_24695,N_25911);
nand U27723 (N_27723,N_25898,N_24917);
and U27724 (N_27724,N_25868,N_24440);
nand U27725 (N_27725,N_25394,N_24196);
nor U27726 (N_27726,N_25763,N_25818);
and U27727 (N_27727,N_24337,N_25658);
and U27728 (N_27728,N_25363,N_25434);
nand U27729 (N_27729,N_25354,N_25842);
xor U27730 (N_27730,N_25762,N_25517);
xnor U27731 (N_27731,N_25769,N_25979);
nand U27732 (N_27732,N_25560,N_25580);
or U27733 (N_27733,N_25944,N_25393);
nand U27734 (N_27734,N_25276,N_24136);
nand U27735 (N_27735,N_25028,N_24723);
xor U27736 (N_27736,N_24127,N_25181);
nand U27737 (N_27737,N_24886,N_24058);
nor U27738 (N_27738,N_25356,N_24201);
nor U27739 (N_27739,N_24816,N_25317);
nor U27740 (N_27740,N_25593,N_25036);
or U27741 (N_27741,N_25967,N_25333);
nor U27742 (N_27742,N_24482,N_25143);
xor U27743 (N_27743,N_24734,N_24692);
or U27744 (N_27744,N_25479,N_24670);
xnor U27745 (N_27745,N_25282,N_25146);
nor U27746 (N_27746,N_24294,N_25855);
nor U27747 (N_27747,N_25707,N_24327);
nor U27748 (N_27748,N_24331,N_24437);
nor U27749 (N_27749,N_25485,N_25187);
xor U27750 (N_27750,N_25755,N_24224);
and U27751 (N_27751,N_25415,N_24965);
nor U27752 (N_27752,N_25490,N_25963);
nand U27753 (N_27753,N_25122,N_25806);
nand U27754 (N_27754,N_24298,N_24590);
or U27755 (N_27755,N_25670,N_24764);
nand U27756 (N_27756,N_24781,N_25591);
and U27757 (N_27757,N_24840,N_24559);
nand U27758 (N_27758,N_25203,N_24639);
and U27759 (N_27759,N_24332,N_25037);
and U27760 (N_27760,N_25226,N_25710);
and U27761 (N_27761,N_24549,N_24670);
xnor U27762 (N_27762,N_25878,N_25633);
nor U27763 (N_27763,N_25870,N_24870);
or U27764 (N_27764,N_24681,N_24634);
or U27765 (N_27765,N_25071,N_24663);
nand U27766 (N_27766,N_25279,N_24566);
nor U27767 (N_27767,N_24939,N_24678);
and U27768 (N_27768,N_25091,N_25883);
and U27769 (N_27769,N_25662,N_25525);
nor U27770 (N_27770,N_25394,N_25957);
nand U27771 (N_27771,N_25441,N_25542);
and U27772 (N_27772,N_25404,N_25105);
nor U27773 (N_27773,N_25856,N_24265);
nor U27774 (N_27774,N_25614,N_25856);
or U27775 (N_27775,N_24824,N_25501);
and U27776 (N_27776,N_25612,N_25554);
xnor U27777 (N_27777,N_24736,N_24965);
and U27778 (N_27778,N_24708,N_24038);
and U27779 (N_27779,N_24254,N_25771);
nand U27780 (N_27780,N_25062,N_25408);
and U27781 (N_27781,N_25692,N_25684);
and U27782 (N_27782,N_24854,N_24419);
xnor U27783 (N_27783,N_24045,N_25494);
xnor U27784 (N_27784,N_24943,N_25404);
and U27785 (N_27785,N_25067,N_24850);
or U27786 (N_27786,N_25611,N_25818);
nand U27787 (N_27787,N_24669,N_25983);
or U27788 (N_27788,N_25097,N_24156);
xnor U27789 (N_27789,N_25286,N_24861);
and U27790 (N_27790,N_25787,N_25000);
nor U27791 (N_27791,N_24473,N_25253);
or U27792 (N_27792,N_25425,N_24264);
nand U27793 (N_27793,N_24235,N_24124);
nor U27794 (N_27794,N_25505,N_24977);
and U27795 (N_27795,N_25917,N_25882);
nor U27796 (N_27796,N_25901,N_25173);
xor U27797 (N_27797,N_24330,N_24084);
nor U27798 (N_27798,N_25237,N_25470);
nor U27799 (N_27799,N_24921,N_25860);
nand U27800 (N_27800,N_24718,N_25015);
and U27801 (N_27801,N_24449,N_25544);
nand U27802 (N_27802,N_25261,N_24133);
or U27803 (N_27803,N_24758,N_24329);
or U27804 (N_27804,N_24836,N_24071);
and U27805 (N_27805,N_25176,N_24736);
and U27806 (N_27806,N_25304,N_24780);
nor U27807 (N_27807,N_24296,N_25337);
nand U27808 (N_27808,N_24817,N_25057);
and U27809 (N_27809,N_24138,N_24981);
nor U27810 (N_27810,N_25986,N_24678);
or U27811 (N_27811,N_24085,N_24469);
nand U27812 (N_27812,N_24297,N_24855);
nor U27813 (N_27813,N_25842,N_25882);
or U27814 (N_27814,N_24840,N_25121);
or U27815 (N_27815,N_24297,N_25649);
and U27816 (N_27816,N_24436,N_24021);
xnor U27817 (N_27817,N_24698,N_24960);
nor U27818 (N_27818,N_25836,N_25502);
and U27819 (N_27819,N_24101,N_25111);
nor U27820 (N_27820,N_25801,N_25805);
nor U27821 (N_27821,N_24808,N_25155);
and U27822 (N_27822,N_25182,N_24463);
nor U27823 (N_27823,N_24947,N_24878);
or U27824 (N_27824,N_24449,N_24798);
and U27825 (N_27825,N_24331,N_25359);
nand U27826 (N_27826,N_25993,N_25115);
or U27827 (N_27827,N_25798,N_24970);
and U27828 (N_27828,N_24471,N_25635);
or U27829 (N_27829,N_25946,N_25401);
nand U27830 (N_27830,N_25104,N_25649);
nor U27831 (N_27831,N_24641,N_24744);
nor U27832 (N_27832,N_25808,N_25449);
and U27833 (N_27833,N_25571,N_25514);
or U27834 (N_27834,N_25195,N_25484);
nor U27835 (N_27835,N_24493,N_25776);
nand U27836 (N_27836,N_25583,N_24527);
or U27837 (N_27837,N_25967,N_24602);
nor U27838 (N_27838,N_25855,N_25543);
xnor U27839 (N_27839,N_24063,N_24323);
or U27840 (N_27840,N_24665,N_25296);
and U27841 (N_27841,N_25364,N_24411);
nor U27842 (N_27842,N_25349,N_24893);
and U27843 (N_27843,N_24784,N_25733);
and U27844 (N_27844,N_24652,N_25004);
xor U27845 (N_27845,N_24682,N_24306);
nand U27846 (N_27846,N_25193,N_24119);
nand U27847 (N_27847,N_24925,N_24990);
or U27848 (N_27848,N_24797,N_24485);
nor U27849 (N_27849,N_24462,N_25425);
or U27850 (N_27850,N_25305,N_25185);
nor U27851 (N_27851,N_24134,N_25941);
nand U27852 (N_27852,N_24465,N_24641);
nor U27853 (N_27853,N_25635,N_24362);
and U27854 (N_27854,N_24029,N_25510);
or U27855 (N_27855,N_24076,N_24542);
and U27856 (N_27856,N_25281,N_25650);
and U27857 (N_27857,N_24273,N_25126);
nor U27858 (N_27858,N_25449,N_24499);
nor U27859 (N_27859,N_25395,N_24361);
or U27860 (N_27860,N_25516,N_24415);
xnor U27861 (N_27861,N_25162,N_24130);
or U27862 (N_27862,N_24188,N_24728);
nand U27863 (N_27863,N_25948,N_25029);
or U27864 (N_27864,N_24821,N_25163);
xor U27865 (N_27865,N_24688,N_24240);
and U27866 (N_27866,N_24662,N_25243);
xnor U27867 (N_27867,N_25308,N_24439);
and U27868 (N_27868,N_24116,N_25941);
or U27869 (N_27869,N_24591,N_24927);
nand U27870 (N_27870,N_24932,N_25023);
and U27871 (N_27871,N_24861,N_25020);
nand U27872 (N_27872,N_24068,N_25941);
nand U27873 (N_27873,N_24295,N_25365);
and U27874 (N_27874,N_25414,N_25620);
or U27875 (N_27875,N_24555,N_25391);
and U27876 (N_27876,N_25847,N_24916);
nand U27877 (N_27877,N_25676,N_25471);
nor U27878 (N_27878,N_24919,N_24044);
nor U27879 (N_27879,N_25425,N_24595);
and U27880 (N_27880,N_25247,N_24281);
or U27881 (N_27881,N_24491,N_25700);
xor U27882 (N_27882,N_24776,N_25519);
nor U27883 (N_27883,N_25249,N_24595);
and U27884 (N_27884,N_24758,N_25219);
or U27885 (N_27885,N_25967,N_25461);
nand U27886 (N_27886,N_25519,N_24993);
xnor U27887 (N_27887,N_25587,N_24393);
and U27888 (N_27888,N_25867,N_24542);
and U27889 (N_27889,N_25681,N_25120);
xor U27890 (N_27890,N_25314,N_25394);
nand U27891 (N_27891,N_25202,N_24689);
nand U27892 (N_27892,N_24542,N_25477);
nor U27893 (N_27893,N_24848,N_24582);
or U27894 (N_27894,N_25322,N_25908);
and U27895 (N_27895,N_25833,N_25735);
xnor U27896 (N_27896,N_24338,N_24113);
xor U27897 (N_27897,N_24954,N_24989);
nand U27898 (N_27898,N_24002,N_24912);
nand U27899 (N_27899,N_25797,N_24649);
or U27900 (N_27900,N_25118,N_25154);
and U27901 (N_27901,N_25073,N_24278);
or U27902 (N_27902,N_25798,N_25849);
and U27903 (N_27903,N_25930,N_25965);
nand U27904 (N_27904,N_24153,N_24477);
or U27905 (N_27905,N_24942,N_24064);
nor U27906 (N_27906,N_24561,N_25768);
nand U27907 (N_27907,N_24572,N_24947);
xnor U27908 (N_27908,N_25878,N_25527);
xor U27909 (N_27909,N_25815,N_24059);
or U27910 (N_27910,N_25882,N_25643);
nor U27911 (N_27911,N_24728,N_24464);
and U27912 (N_27912,N_25312,N_24860);
nor U27913 (N_27913,N_25852,N_24674);
nand U27914 (N_27914,N_25395,N_24994);
and U27915 (N_27915,N_25956,N_25488);
nand U27916 (N_27916,N_25205,N_25005);
nand U27917 (N_27917,N_24253,N_24860);
xnor U27918 (N_27918,N_25232,N_25428);
and U27919 (N_27919,N_24134,N_25822);
nor U27920 (N_27920,N_25966,N_25447);
or U27921 (N_27921,N_25554,N_25353);
or U27922 (N_27922,N_24327,N_24374);
and U27923 (N_27923,N_25386,N_25652);
nor U27924 (N_27924,N_25763,N_25444);
or U27925 (N_27925,N_25598,N_24932);
nor U27926 (N_27926,N_25708,N_25230);
and U27927 (N_27927,N_25971,N_24386);
and U27928 (N_27928,N_24578,N_24864);
xnor U27929 (N_27929,N_24824,N_25954);
and U27930 (N_27930,N_24321,N_25720);
nor U27931 (N_27931,N_25704,N_25856);
nor U27932 (N_27932,N_24192,N_25255);
or U27933 (N_27933,N_25308,N_25766);
or U27934 (N_27934,N_24540,N_25294);
or U27935 (N_27935,N_25764,N_25279);
nor U27936 (N_27936,N_24348,N_25182);
nor U27937 (N_27937,N_25405,N_25277);
xnor U27938 (N_27938,N_25947,N_24373);
nand U27939 (N_27939,N_25570,N_24776);
xor U27940 (N_27940,N_24337,N_25981);
or U27941 (N_27941,N_25798,N_24972);
and U27942 (N_27942,N_24532,N_25491);
and U27943 (N_27943,N_25164,N_24472);
and U27944 (N_27944,N_24762,N_25837);
nor U27945 (N_27945,N_24505,N_25339);
and U27946 (N_27946,N_25010,N_25844);
and U27947 (N_27947,N_24390,N_24767);
and U27948 (N_27948,N_25190,N_25375);
or U27949 (N_27949,N_24530,N_25900);
and U27950 (N_27950,N_25371,N_25633);
or U27951 (N_27951,N_25388,N_24832);
and U27952 (N_27952,N_25579,N_24057);
xnor U27953 (N_27953,N_24371,N_25129);
nand U27954 (N_27954,N_24681,N_25638);
xor U27955 (N_27955,N_24359,N_25383);
and U27956 (N_27956,N_25762,N_25820);
nand U27957 (N_27957,N_25881,N_25298);
xor U27958 (N_27958,N_24379,N_24771);
nor U27959 (N_27959,N_24331,N_24312);
or U27960 (N_27960,N_24698,N_25825);
nor U27961 (N_27961,N_25273,N_24413);
and U27962 (N_27962,N_24455,N_25883);
nor U27963 (N_27963,N_25228,N_25432);
nor U27964 (N_27964,N_25266,N_24658);
nor U27965 (N_27965,N_24367,N_24046);
xnor U27966 (N_27966,N_25048,N_24930);
xor U27967 (N_27967,N_25173,N_25930);
and U27968 (N_27968,N_24565,N_25874);
nor U27969 (N_27969,N_24480,N_25369);
or U27970 (N_27970,N_25606,N_24426);
nor U27971 (N_27971,N_25937,N_24830);
nor U27972 (N_27972,N_24519,N_25408);
nand U27973 (N_27973,N_25474,N_24100);
or U27974 (N_27974,N_24321,N_25376);
or U27975 (N_27975,N_24942,N_24219);
nor U27976 (N_27976,N_24814,N_25623);
and U27977 (N_27977,N_24750,N_24788);
nor U27978 (N_27978,N_25381,N_25852);
or U27979 (N_27979,N_24655,N_25886);
xnor U27980 (N_27980,N_25944,N_24490);
and U27981 (N_27981,N_25381,N_24904);
xor U27982 (N_27982,N_25912,N_25033);
nor U27983 (N_27983,N_24494,N_24833);
nor U27984 (N_27984,N_25228,N_25167);
nand U27985 (N_27985,N_25919,N_25093);
nand U27986 (N_27986,N_24888,N_25299);
or U27987 (N_27987,N_25961,N_25761);
and U27988 (N_27988,N_24690,N_25260);
nand U27989 (N_27989,N_25353,N_24701);
and U27990 (N_27990,N_24666,N_24963);
nand U27991 (N_27991,N_25392,N_24941);
nor U27992 (N_27992,N_24079,N_24033);
nor U27993 (N_27993,N_25239,N_24691);
xor U27994 (N_27994,N_24176,N_25676);
nand U27995 (N_27995,N_24704,N_25104);
nor U27996 (N_27996,N_24046,N_24904);
nor U27997 (N_27997,N_24744,N_24471);
or U27998 (N_27998,N_25781,N_24656);
or U27999 (N_27999,N_24782,N_25894);
or U28000 (N_28000,N_26275,N_26132);
nand U28001 (N_28001,N_27719,N_26459);
xnor U28002 (N_28002,N_27024,N_26196);
nor U28003 (N_28003,N_27178,N_26591);
nor U28004 (N_28004,N_27105,N_27126);
nor U28005 (N_28005,N_27334,N_26256);
or U28006 (N_28006,N_27367,N_26614);
xnor U28007 (N_28007,N_27897,N_27400);
or U28008 (N_28008,N_26126,N_27220);
xnor U28009 (N_28009,N_26220,N_27412);
nand U28010 (N_28010,N_27085,N_26321);
nand U28011 (N_28011,N_26695,N_27317);
nand U28012 (N_28012,N_26341,N_27210);
nor U28013 (N_28013,N_27653,N_27003);
and U28014 (N_28014,N_26508,N_27724);
nand U28015 (N_28015,N_27411,N_26288);
and U28016 (N_28016,N_27685,N_26381);
or U28017 (N_28017,N_27114,N_27982);
xor U28018 (N_28018,N_27993,N_27592);
nor U28019 (N_28019,N_26465,N_27505);
and U28020 (N_28020,N_27465,N_26129);
nor U28021 (N_28021,N_27185,N_27845);
xnor U28022 (N_28022,N_26812,N_26332);
xor U28023 (N_28023,N_26215,N_27347);
nand U28024 (N_28024,N_26680,N_26647);
nor U28025 (N_28025,N_26474,N_27824);
nor U28026 (N_28026,N_27459,N_27738);
nor U28027 (N_28027,N_27774,N_27103);
xnor U28028 (N_28028,N_26350,N_26443);
xnor U28029 (N_28029,N_26995,N_27856);
and U28030 (N_28030,N_27663,N_27839);
or U28031 (N_28031,N_27504,N_27167);
and U28032 (N_28032,N_26011,N_27966);
nor U28033 (N_28033,N_27299,N_26391);
or U28034 (N_28034,N_27564,N_26127);
nand U28035 (N_28035,N_26344,N_27475);
xnor U28036 (N_28036,N_26472,N_26273);
nand U28037 (N_28037,N_27528,N_27526);
or U28038 (N_28038,N_27550,N_26518);
and U28039 (N_28039,N_27182,N_26179);
and U28040 (N_28040,N_27760,N_27232);
xnor U28041 (N_28041,N_27454,N_26879);
nor U28042 (N_28042,N_26401,N_26022);
and U28043 (N_28043,N_27370,N_26062);
xor U28044 (N_28044,N_26525,N_27518);
nand U28045 (N_28045,N_26934,N_26621);
or U28046 (N_28046,N_26742,N_26663);
nor U28047 (N_28047,N_26703,N_27890);
nand U28048 (N_28048,N_27609,N_26191);
nor U28049 (N_28049,N_27779,N_26312);
and U28050 (N_28050,N_27937,N_27977);
and U28051 (N_28051,N_27493,N_26377);
nand U28052 (N_28052,N_27339,N_27762);
or U28053 (N_28053,N_27580,N_27260);
nand U28054 (N_28054,N_26067,N_26863);
or U28055 (N_28055,N_26039,N_26826);
nor U28056 (N_28056,N_27610,N_26837);
nand U28057 (N_28057,N_27576,N_27758);
xnor U28058 (N_28058,N_27695,N_26648);
nor U28059 (N_28059,N_26493,N_26760);
xnor U28060 (N_28060,N_27674,N_26726);
nand U28061 (N_28061,N_27583,N_26492);
nor U28062 (N_28062,N_27233,N_27643);
xor U28063 (N_28063,N_27739,N_26274);
xnor U28064 (N_28064,N_27679,N_27136);
xnor U28065 (N_28065,N_27457,N_26977);
nand U28066 (N_28066,N_26659,N_27945);
nor U28067 (N_28067,N_26357,N_27050);
or U28068 (N_28068,N_27778,N_26537);
and U28069 (N_28069,N_27115,N_27353);
and U28070 (N_28070,N_26666,N_27892);
nand U28071 (N_28071,N_26636,N_27924);
or U28072 (N_28072,N_27468,N_27780);
nand U28073 (N_28073,N_26951,N_26932);
and U28074 (N_28074,N_26478,N_26319);
nand U28075 (N_28075,N_26853,N_26107);
and U28076 (N_28076,N_27763,N_27512);
nand U28077 (N_28077,N_27259,N_27731);
or U28078 (N_28078,N_26326,N_27480);
nand U28079 (N_28079,N_27263,N_27219);
xor U28080 (N_28080,N_27531,N_27179);
xor U28081 (N_28081,N_26119,N_26419);
or U28082 (N_28082,N_26148,N_27656);
nand U28083 (N_28083,N_26491,N_26436);
or U28084 (N_28084,N_27020,N_26014);
xnor U28085 (N_28085,N_27336,N_26918);
and U28086 (N_28086,N_26009,N_26780);
and U28087 (N_28087,N_27713,N_26475);
and U28088 (N_28088,N_26969,N_26200);
nor U28089 (N_28089,N_26059,N_27437);
nor U28090 (N_28090,N_26967,N_27959);
or U28091 (N_28091,N_26248,N_27062);
nor U28092 (N_28092,N_26163,N_26923);
nand U28093 (N_28093,N_26035,N_26555);
and U28094 (N_28094,N_27511,N_26868);
and U28095 (N_28095,N_27539,N_27968);
and U28096 (N_28096,N_27056,N_27556);
nor U28097 (N_28097,N_26403,N_27923);
nor U28098 (N_28098,N_26487,N_27326);
nor U28099 (N_28099,N_27417,N_26392);
nor U28100 (N_28100,N_26158,N_26856);
and U28101 (N_28101,N_27686,N_26700);
and U28102 (N_28102,N_27360,N_27201);
xnor U28103 (N_28103,N_27542,N_27080);
nor U28104 (N_28104,N_27358,N_26396);
nor U28105 (N_28105,N_26414,N_26084);
or U28106 (N_28106,N_26723,N_26207);
and U28107 (N_28107,N_27549,N_27588);
nand U28108 (N_28108,N_26060,N_27883);
nand U28109 (N_28109,N_27055,N_27031);
and U28110 (N_28110,N_27106,N_27585);
nor U28111 (N_28111,N_26910,N_27757);
or U28112 (N_28112,N_26115,N_26224);
nand U28113 (N_28113,N_26547,N_26762);
and U28114 (N_28114,N_27172,N_26042);
nor U28115 (N_28115,N_26485,N_27163);
or U28116 (N_28116,N_26779,N_26108);
and U28117 (N_28117,N_26363,N_27869);
nand U28118 (N_28118,N_26330,N_26552);
nor U28119 (N_28119,N_26184,N_26267);
xnor U28120 (N_28120,N_27913,N_27865);
or U28121 (N_28121,N_26820,N_27122);
xnor U28122 (N_28122,N_27994,N_27377);
nand U28123 (N_28123,N_27217,N_26778);
and U28124 (N_28124,N_27906,N_26875);
nand U28125 (N_28125,N_27754,N_27327);
and U28126 (N_28126,N_27218,N_27683);
or U28127 (N_28127,N_27064,N_26586);
nor U28128 (N_28128,N_27271,N_27809);
nor U28129 (N_28129,N_26811,N_26506);
nand U28130 (N_28130,N_27440,N_27642);
or U28131 (N_28131,N_27245,N_26175);
xor U28132 (N_28132,N_26739,N_26583);
xnor U28133 (N_28133,N_27407,N_26291);
xnor U28134 (N_28134,N_27775,N_27519);
and U28135 (N_28135,N_27714,N_27551);
nand U28136 (N_28136,N_27045,N_26888);
xnor U28137 (N_28137,N_26705,N_27503);
nand U28138 (N_28138,N_27972,N_27699);
nor U28139 (N_28139,N_27269,N_26304);
nand U28140 (N_28140,N_27666,N_27971);
nand U28141 (N_28141,N_27169,N_26343);
nor U28142 (N_28142,N_27759,N_26861);
nor U28143 (N_28143,N_26140,N_27230);
and U28144 (N_28144,N_26893,N_27221);
nand U28145 (N_28145,N_26266,N_27433);
and U28146 (N_28146,N_27662,N_26120);
nor U28147 (N_28147,N_26323,N_27051);
and U28148 (N_28148,N_27250,N_27072);
and U28149 (N_28149,N_27578,N_27535);
xnor U28150 (N_28150,N_26997,N_26437);
or U28151 (N_28151,N_27036,N_27229);
and U28152 (N_28152,N_26584,N_27956);
or U28153 (N_28153,N_27522,N_27744);
or U28154 (N_28154,N_27768,N_27595);
nor U28155 (N_28155,N_26962,N_27351);
and U28156 (N_28156,N_27575,N_26305);
xnor U28157 (N_28157,N_27543,N_26989);
or U28158 (N_28158,N_26041,N_27037);
or U28159 (N_28159,N_27704,N_27851);
nor U28160 (N_28160,N_26830,N_26633);
xnor U28161 (N_28161,N_27962,N_26295);
and U28162 (N_28162,N_26483,N_26806);
nand U28163 (N_28163,N_27319,N_26069);
and U28164 (N_28164,N_27111,N_26423);
xor U28165 (N_28165,N_26573,N_26921);
nor U28166 (N_28166,N_26610,N_27429);
nor U28167 (N_28167,N_27767,N_27730);
nor U28168 (N_28168,N_26089,N_27290);
nand U28169 (N_28169,N_27307,N_27008);
xnor U28170 (N_28170,N_26664,N_26049);
and U28171 (N_28171,N_27277,N_27690);
nor U28172 (N_28172,N_27577,N_26113);
nand U28173 (N_28173,N_26829,N_26539);
nand U28174 (N_28174,N_27227,N_26745);
nand U28175 (N_28175,N_26605,N_26956);
nor U28176 (N_28176,N_27732,N_27131);
and U28177 (N_28177,N_27948,N_26681);
or U28178 (N_28178,N_26418,N_26821);
nand U28179 (N_28179,N_26892,N_26557);
xnor U28180 (N_28180,N_27190,N_26153);
nand U28181 (N_28181,N_26917,N_26192);
or U28182 (N_28182,N_27668,N_27902);
nand U28183 (N_28183,N_26625,N_27280);
nand U28184 (N_28184,N_26029,N_26709);
xnor U28185 (N_28185,N_26137,N_27047);
or U28186 (N_28186,N_26637,N_27618);
xnor U28187 (N_28187,N_26138,N_26390);
nand U28188 (N_28188,N_26792,N_26412);
nor U28189 (N_28189,N_26499,N_27860);
or U28190 (N_28190,N_26168,N_27622);
and U28191 (N_28191,N_26691,N_26817);
xnor U28192 (N_28192,N_27027,N_26670);
xnor U28193 (N_28193,N_27435,N_27660);
and U28194 (N_28194,N_27041,N_27193);
xor U28195 (N_28195,N_26789,N_27019);
and U28196 (N_28196,N_26241,N_26898);
nand U28197 (N_28197,N_26674,N_27084);
or U28198 (N_28198,N_26983,N_27991);
nor U28199 (N_28199,N_27381,N_27238);
xor U28200 (N_28200,N_26818,N_26984);
or U28201 (N_28201,N_27887,N_27999);
xor U28202 (N_28202,N_26704,N_26259);
nor U28203 (N_28203,N_27162,N_26914);
and U28204 (N_28204,N_27586,N_26653);
and U28205 (N_28205,N_27946,N_26206);
or U28206 (N_28206,N_26193,N_27239);
nor U28207 (N_28207,N_26835,N_26415);
and U28208 (N_28208,N_27687,N_26699);
or U28209 (N_28209,N_27895,N_26566);
and U28210 (N_28210,N_26247,N_26397);
nor U28211 (N_28211,N_26535,N_26534);
nor U28212 (N_28212,N_26225,N_26630);
nor U28213 (N_28213,N_27615,N_27188);
or U28214 (N_28214,N_26567,N_27752);
nor U28215 (N_28215,N_26968,N_26971);
xnor U28216 (N_28216,N_27667,N_26121);
or U28217 (N_28217,N_26366,N_26144);
nand U28218 (N_28218,N_26514,N_26787);
or U28219 (N_28219,N_26420,N_26000);
nor U28220 (N_28220,N_27311,N_26574);
or U28221 (N_28221,N_27840,N_27444);
nand U28222 (N_28222,N_27806,N_26667);
nor U28223 (N_28223,N_27127,N_27125);
nor U28224 (N_28224,N_27678,N_26135);
xnor U28225 (N_28225,N_27949,N_26590);
or U28226 (N_28226,N_26136,N_26913);
nand U28227 (N_28227,N_26854,N_27645);
or U28228 (N_28228,N_27741,N_26092);
or U28229 (N_28229,N_26719,N_26816);
or U28230 (N_28230,N_27248,N_27349);
nand U28231 (N_28231,N_27694,N_26793);
nand U28232 (N_28232,N_26445,N_26301);
and U28233 (N_28233,N_27710,N_26318);
nor U28234 (N_28234,N_26505,N_27517);
nand U28235 (N_28235,N_26587,N_27723);
and U28236 (N_28236,N_26024,N_26199);
or U28237 (N_28237,N_26016,N_27054);
xnor U28238 (N_28238,N_27282,N_26497);
and U28239 (N_28239,N_27152,N_27029);
or U28240 (N_28240,N_27212,N_27487);
nand U28241 (N_28241,N_27960,N_27788);
nand U28242 (N_28242,N_26204,N_27074);
nand U28243 (N_28243,N_27396,N_26687);
nand U28244 (N_28244,N_26572,N_27346);
nor U28245 (N_28245,N_27011,N_26568);
nand U28246 (N_28246,N_26645,N_27315);
nand U28247 (N_28247,N_26994,N_26407);
xor U28248 (N_28248,N_27142,N_27933);
and U28249 (N_28249,N_26008,N_27533);
nor U28250 (N_28250,N_26966,N_27641);
and U28251 (N_28251,N_27734,N_26481);
or U28252 (N_28252,N_27529,N_27623);
nand U28253 (N_28253,N_26683,N_27120);
and U28254 (N_28254,N_27886,N_27509);
or U28255 (N_28255,N_26188,N_26894);
nand U28256 (N_28256,N_27350,N_26870);
nor U28257 (N_28257,N_26713,N_27006);
nand U28258 (N_28258,N_26790,N_27208);
xnor U28259 (N_28259,N_27273,N_26015);
or U28260 (N_28260,N_26733,N_26752);
or U28261 (N_28261,N_26309,N_27825);
xnor U28262 (N_28262,N_27793,N_26227);
or U28263 (N_28263,N_27325,N_27743);
or U28264 (N_28264,N_26424,N_26617);
or U28265 (N_28265,N_27159,N_27375);
and U28266 (N_28266,N_27415,N_27117);
and U28267 (N_28267,N_26027,N_26882);
or U28268 (N_28268,N_26198,N_26251);
xor U28269 (N_28269,N_26513,N_26285);
nand U28270 (N_28270,N_27146,N_27344);
nand U28271 (N_28271,N_26622,N_26554);
nor U28272 (N_28272,N_26161,N_26538);
xnor U28273 (N_28273,N_26374,N_26012);
or U28274 (N_28274,N_26579,N_27057);
xor U28275 (N_28275,N_26624,N_26523);
and U28276 (N_28276,N_27010,N_27394);
or U28277 (N_28277,N_26839,N_27499);
nand U28278 (N_28278,N_26991,N_26571);
and U28279 (N_28279,N_27464,N_27414);
nor U28280 (N_28280,N_26222,N_26873);
or U28281 (N_28281,N_26010,N_26577);
nand U28282 (N_28282,N_27655,N_27471);
and U28283 (N_28283,N_27613,N_27822);
xor U28284 (N_28284,N_27261,N_26949);
nor U28285 (N_28285,N_26233,N_26734);
xor U28286 (N_28286,N_27288,N_26197);
nor U28287 (N_28287,N_26280,N_26930);
nor U28288 (N_28288,N_27249,N_27878);
xnor U28289 (N_28289,N_26150,N_26306);
xnor U28290 (N_28290,N_26846,N_26243);
xnor U28291 (N_28291,N_26398,N_27821);
nor U28292 (N_28292,N_27022,N_26157);
xor U28293 (N_28293,N_27861,N_27721);
and U28294 (N_28294,N_26048,N_27448);
xor U28295 (N_28295,N_27872,N_27804);
nand U28296 (N_28296,N_27070,N_27102);
and U28297 (N_28297,N_26827,N_26869);
and U28298 (N_28298,N_26720,N_26980);
and U28299 (N_28299,N_26046,N_26928);
or U28300 (N_28300,N_27606,N_26771);
nand U28301 (N_28301,N_26400,N_27134);
xnor U28302 (N_28302,N_26682,N_27039);
xor U28303 (N_28303,N_27997,N_26651);
nor U28304 (N_28304,N_26620,N_26242);
nor U28305 (N_28305,N_26348,N_26946);
xor U28306 (N_28306,N_27552,N_27756);
or U28307 (N_28307,N_27124,N_26074);
and U28308 (N_28308,N_27781,N_26335);
nand U28309 (N_28309,N_27943,N_27581);
and U28310 (N_28310,N_27461,N_27737);
xor U28311 (N_28311,N_26228,N_27443);
nand U28312 (N_28312,N_27755,N_26214);
or U28313 (N_28313,N_26948,N_27604);
nand U28314 (N_28314,N_27525,N_26026);
nor U28315 (N_28315,N_27130,N_27633);
xnor U28316 (N_28316,N_27005,N_27491);
and U28317 (N_28317,N_26336,N_27289);
nand U28318 (N_28318,N_27107,N_26230);
xor U28319 (N_28319,N_26844,N_27110);
and U28320 (N_28320,N_26263,N_27281);
nor U28321 (N_28321,N_27534,N_27980);
and U28322 (N_28322,N_26495,N_26749);
nand U28323 (N_28323,N_26105,N_27398);
or U28324 (N_28324,N_26100,N_27403);
or U28325 (N_28325,N_27244,N_27191);
nor U28326 (N_28326,N_27940,N_26410);
nand U28327 (N_28327,N_26471,N_26342);
xor U28328 (N_28328,N_27482,N_26281);
or U28329 (N_28329,N_27366,N_26447);
nand U28330 (N_28330,N_27870,N_27380);
nand U28331 (N_28331,N_27242,N_27386);
xnor U28332 (N_28332,N_26833,N_26441);
nor U28333 (N_28333,N_27888,N_27452);
nor U28334 (N_28334,N_27287,N_26402);
nand U28335 (N_28335,N_27555,N_27657);
xor U28336 (N_28336,N_26520,N_26382);
nand U28337 (N_28337,N_27270,N_26676);
nor U28338 (N_28338,N_26735,N_27602);
nor U28339 (N_28339,N_26900,N_26096);
nor U28340 (N_28340,N_27922,N_27450);
nand U28341 (N_28341,N_26708,N_26784);
nor U28342 (N_28342,N_26025,N_27896);
nand U28343 (N_28343,N_27745,N_27619);
or U28344 (N_28344,N_27082,N_27941);
nor U28345 (N_28345,N_27352,N_27173);
xnor U28346 (N_28346,N_26809,N_27203);
nor U28347 (N_28347,N_27376,N_27337);
nand U28348 (N_28348,N_26619,N_27279);
nor U28349 (N_28349,N_27097,N_27969);
nor U28350 (N_28350,N_26961,N_27796);
nand U28351 (N_28351,N_27021,N_26880);
and U28352 (N_28352,N_26627,N_26313);
nor U28353 (N_28353,N_27880,N_27761);
and U28354 (N_28354,N_26031,N_27200);
nor U28355 (N_28355,N_26417,N_27930);
xnor U28356 (N_28356,N_26152,N_27389);
nor U28357 (N_28357,N_27144,N_26594);
xnor U28358 (N_28358,N_26072,N_27331);
nor U28359 (N_28359,N_27365,N_26367);
and U28360 (N_28360,N_27506,N_27086);
or U28361 (N_28361,N_26075,N_27803);
nor U28362 (N_28362,N_27850,N_26102);
or U28363 (N_28363,N_26795,N_27799);
xnor U28364 (N_28364,N_27357,N_26600);
and U28365 (N_28365,N_27729,N_26270);
and U28366 (N_28366,N_26339,N_26775);
or U28367 (N_28367,N_26669,N_27540);
nand U28368 (N_28368,N_27301,N_27648);
nand U28369 (N_28369,N_27129,N_27026);
or U28370 (N_28370,N_27541,N_27369);
and U28371 (N_28371,N_26284,N_27765);
or U28372 (N_28372,N_27338,N_26299);
xnor U28373 (N_28373,N_26797,N_26353);
or U28374 (N_28374,N_27195,N_27640);
and U28375 (N_28375,N_27700,N_26020);
nor U28376 (N_28376,N_27296,N_27079);
xor U28377 (N_28377,N_26599,N_27364);
nor U28378 (N_28378,N_27516,N_26229);
nor U28379 (N_28379,N_26741,N_26783);
nand U28380 (N_28380,N_26987,N_27236);
or U28381 (N_28381,N_27841,N_27866);
nand U28382 (N_28382,N_26316,N_26467);
and U28383 (N_28383,N_26232,N_26328);
nand U28384 (N_28384,N_27286,N_26964);
and U28385 (N_28385,N_27740,N_26209);
xnor U28386 (N_28386,N_27626,N_27794);
xor U28387 (N_28387,N_26159,N_26068);
or U28388 (N_28388,N_27356,N_27785);
and U28389 (N_28389,N_27463,N_26975);
nor U28390 (N_28390,N_26548,N_27884);
or U28391 (N_28391,N_26738,N_26433);
and U28392 (N_28392,N_26383,N_26889);
and U28393 (N_28393,N_26927,N_27829);
and U28394 (N_28394,N_26289,N_27145);
or U28395 (N_28395,N_26810,N_27876);
or U28396 (N_28396,N_27198,N_27953);
and U28397 (N_28397,N_27790,N_26265);
and U28398 (N_28398,N_26576,N_27328);
nand U28399 (N_28399,N_27693,N_26439);
and U28400 (N_28400,N_27314,N_27661);
xnor U28401 (N_28401,N_26920,N_26464);
xor U28402 (N_28402,N_27976,N_27671);
nand U28403 (N_28403,N_26307,N_26389);
and U28404 (N_28404,N_27255,N_26457);
nor U28405 (N_28405,N_27777,N_26688);
xor U28406 (N_28406,N_26678,N_27816);
and U28407 (N_28407,N_26824,N_27702);
nor U28408 (N_28408,N_27772,N_26768);
nor U28409 (N_28409,N_27215,N_27449);
nor U28410 (N_28410,N_27165,N_26761);
nor U28411 (N_28411,N_27954,N_27044);
nand U28412 (N_28412,N_27362,N_26038);
xor U28413 (N_28413,N_27858,N_26271);
nand U28414 (N_28414,N_26940,N_27189);
or U28415 (N_28415,N_26634,N_26832);
nand U28416 (N_28416,N_27109,N_26171);
or U28417 (N_28417,N_26314,N_27749);
or U28418 (N_28418,N_27789,N_26327);
nor U28419 (N_28419,N_26529,N_26325);
xor U28420 (N_28420,N_27625,N_26843);
nor U28421 (N_28421,N_27566,N_27567);
nand U28422 (N_28422,N_26729,N_26502);
or U28423 (N_28423,N_26244,N_26231);
nand U28424 (N_28424,N_26580,N_27494);
nand U28425 (N_28425,N_27116,N_26300);
nor U28426 (N_28426,N_26386,N_27974);
or U28427 (N_28427,N_26945,N_26823);
and U28428 (N_28428,N_26292,N_27392);
or U28429 (N_28429,N_26311,N_27597);
or U28430 (N_28430,N_27514,N_26394);
nor U28431 (N_28431,N_26489,N_27470);
and U28432 (N_28432,N_27907,N_27893);
nor U28433 (N_28433,N_26550,N_27701);
or U28434 (N_28434,N_27716,N_26358);
xor U28435 (N_28435,N_27554,N_26006);
nor U28436 (N_28436,N_26702,N_26250);
nand U28437 (N_28437,N_27262,N_27784);
xor U28438 (N_28438,N_26086,N_27458);
xnor U28439 (N_28439,N_27206,N_27591);
or U28440 (N_28440,N_27706,N_26650);
xnor U28441 (N_28441,N_27620,N_27171);
xnor U28442 (N_28442,N_26924,N_26114);
nor U28443 (N_28443,N_26799,N_26162);
nor U28444 (N_28444,N_27634,N_26017);
xor U28445 (N_28445,N_27069,N_26836);
xnor U28446 (N_28446,N_26303,N_27676);
and U28447 (N_28447,N_27278,N_27497);
nor U28448 (N_28448,N_26044,N_27835);
or U28449 (N_28449,N_26895,N_26262);
nand U28450 (N_28450,N_26473,N_26758);
nor U28451 (N_28451,N_27899,N_27406);
xor U28452 (N_28452,N_26543,N_26510);
and U28453 (N_28453,N_26395,N_27063);
nor U28454 (N_28454,N_27033,N_27717);
xor U28455 (N_28455,N_27553,N_26909);
or U28456 (N_28456,N_26116,N_27207);
or U28457 (N_28457,N_27978,N_26208);
and U28458 (N_28458,N_27987,N_26246);
or U28459 (N_28459,N_26334,N_27828);
or U28460 (N_28460,N_27644,N_27532);
nand U28461 (N_28461,N_26542,N_27486);
and U28462 (N_28462,N_27510,N_27472);
nand U28463 (N_28463,N_26449,N_27646);
xor U28464 (N_28464,N_26957,N_27569);
nand U28465 (N_28465,N_26461,N_27548);
nor U28466 (N_28466,N_26684,N_26950);
and U28467 (N_28467,N_27333,N_27926);
nor U28468 (N_28468,N_27254,N_26689);
xor U28469 (N_28469,N_26373,N_26287);
and U28470 (N_28470,N_27688,N_26532);
nand U28471 (N_28471,N_26364,N_27708);
nand U28472 (N_28472,N_26455,N_27931);
or U28473 (N_28473,N_26857,N_27920);
nand U28474 (N_28474,N_26180,N_26052);
nand U28475 (N_28475,N_27986,N_26845);
nand U28476 (N_28476,N_27485,N_27722);
and U28477 (N_28477,N_26562,N_27800);
or U28478 (N_28478,N_26970,N_27842);
nand U28479 (N_28479,N_26871,N_27970);
xnor U28480 (N_28480,N_26588,N_26149);
or U28481 (N_28481,N_26859,N_27908);
xor U28482 (N_28482,N_27300,N_26446);
xnor U28483 (N_28483,N_26759,N_27343);
nor U28484 (N_28484,N_26123,N_26254);
nor U28485 (N_28485,N_27698,N_26142);
or U28486 (N_28486,N_27378,N_26352);
xnor U28487 (N_28487,N_27783,N_27984);
xor U28488 (N_28488,N_26782,N_27133);
xor U28489 (N_28489,N_26602,N_27579);
nand U28490 (N_28490,N_26903,N_26718);
and U28491 (N_28491,N_27294,N_26444);
xnor U28492 (N_28492,N_26393,N_26380);
and U28493 (N_28493,N_26626,N_26643);
or U28494 (N_28494,N_27481,N_26376);
nor U28495 (N_28495,N_27612,N_26090);
and U28496 (N_28496,N_26076,N_26279);
xor U28497 (N_28497,N_26053,N_26324);
or U28498 (N_28498,N_27515,N_27513);
nor U28499 (N_28499,N_26531,N_26901);
or U28500 (N_28500,N_27932,N_26176);
nand U28501 (N_28501,N_26876,N_27002);
xor U28502 (N_28502,N_26177,N_27222);
xor U28503 (N_28503,N_27501,N_27335);
xnor U28504 (N_28504,N_26887,N_26103);
and U28505 (N_28505,N_27049,N_26612);
or U28506 (N_28506,N_26050,N_27846);
xnor U28507 (N_28507,N_26595,N_27368);
xor U28508 (N_28508,N_27150,N_26297);
or U28509 (N_28509,N_27427,N_27638);
nor U28510 (N_28510,N_27409,N_26831);
xor U28511 (N_28511,N_26872,N_26737);
and U28512 (N_28512,N_26698,N_26933);
or U28513 (N_28513,N_26819,N_26238);
and U28514 (N_28514,N_26104,N_27979);
nor U28515 (N_28515,N_26519,N_27393);
and U28516 (N_28516,N_26960,N_26988);
or U28517 (N_28517,N_27187,N_26611);
nand U28518 (N_28518,N_27175,N_27934);
and U28519 (N_28519,N_26286,N_26173);
nand U28520 (N_28520,N_26165,N_27958);
xor U28521 (N_28521,N_26346,N_26786);
nor U28522 (N_28522,N_26714,N_27628);
xor U28523 (N_28523,N_27753,N_26710);
nand U28524 (N_28524,N_27882,N_26249);
or U28525 (N_28525,N_26462,N_26355);
nor U28526 (N_28526,N_27894,N_27305);
nand U28527 (N_28527,N_26582,N_27961);
nor U28528 (N_28528,N_27827,N_26855);
nor U28529 (N_28529,N_27402,N_26753);
nor U28530 (N_28530,N_26701,N_27138);
nor U28531 (N_28531,N_26805,N_27166);
nand U28532 (N_28532,N_27696,N_27891);
nand U28533 (N_28533,N_26772,N_26609);
nor U28534 (N_28534,N_27170,N_27149);
nand U28535 (N_28535,N_26706,N_27659);
or U28536 (N_28536,N_27771,N_27076);
and U28537 (N_28537,N_27235,N_26884);
and U28538 (N_28538,N_27616,N_27466);
xnor U28539 (N_28539,N_27423,N_27214);
nor U28540 (N_28540,N_26511,N_27705);
or U28541 (N_28541,N_26986,N_27373);
and U28542 (N_28542,N_27012,N_27176);
nor U28543 (N_28543,N_26106,N_26767);
or U28544 (N_28544,N_26186,N_26294);
nand U28545 (N_28545,N_26018,N_27834);
and U28546 (N_28546,N_26133,N_27359);
nor U28547 (N_28547,N_26890,N_26754);
and U28548 (N_28548,N_27537,N_27787);
nor U28549 (N_28549,N_26507,N_26834);
nand U28550 (N_28550,N_27769,N_27438);
nand U28551 (N_28551,N_27395,N_26458);
and U28552 (N_28552,N_26375,N_27536);
xnor U28553 (N_28553,N_27837,N_26435);
nand U28554 (N_28554,N_27139,N_27559);
and U28555 (N_28555,N_26094,N_26456);
xor U28556 (N_28556,N_26672,N_26007);
and U28557 (N_28557,N_26866,N_27318);
and U28558 (N_28558,N_26858,N_27766);
nor U28559 (N_28559,N_27241,N_26711);
xnor U28560 (N_28560,N_26631,N_26240);
xor U28561 (N_28561,N_27614,N_26796);
nor U28562 (N_28562,N_26925,N_26213);
nor U28563 (N_28563,N_27158,N_27649);
nor U28564 (N_28564,N_26959,N_26891);
nand U28565 (N_28565,N_27007,N_27252);
nand U28566 (N_28566,N_27297,N_26030);
or U28567 (N_28567,N_26993,N_27565);
and U28568 (N_28568,N_26524,N_27684);
xnor U28569 (N_28569,N_27025,N_27092);
nand U28570 (N_28570,N_26278,N_27264);
or U28571 (N_28571,N_27652,N_27345);
and U28572 (N_28572,N_27099,N_27205);
or U28573 (N_28573,N_26183,N_26902);
and U28574 (N_28574,N_27726,N_26365);
and U28575 (N_28575,N_26237,N_26218);
or U28576 (N_28576,N_26952,N_26131);
and U28577 (N_28577,N_26635,N_27322);
nand U28578 (N_28578,N_26033,N_27900);
nor U28579 (N_28579,N_26765,N_26088);
and U28580 (N_28580,N_26744,N_26581);
or U28581 (N_28581,N_27813,N_27015);
xor U28582 (N_28582,N_27975,N_27881);
nand U28583 (N_28583,N_26504,N_27546);
or U28584 (N_28584,N_27830,N_26569);
or U28585 (N_28585,N_27184,N_27808);
or U28586 (N_28586,N_27177,N_27736);
nor U28587 (N_28587,N_26345,N_27060);
xor U28588 (N_28588,N_26814,N_26878);
nor U28589 (N_28589,N_27384,N_27607);
or U28590 (N_28590,N_26947,N_27293);
nand U28591 (N_28591,N_26066,N_26079);
nor U28592 (N_28592,N_27313,N_27283);
nor U28593 (N_28593,N_27157,N_26174);
and U28594 (N_28594,N_27942,N_26656);
xnor U28595 (N_28595,N_26838,N_27568);
nand U28596 (N_28596,N_26883,N_26110);
nand U28597 (N_28597,N_26662,N_26788);
nand U28598 (N_28598,N_27174,N_26360);
or U28599 (N_28599,N_27715,N_26623);
nand U28600 (N_28600,N_26261,N_26530);
and U28601 (N_28601,N_27764,N_27303);
xnor U28602 (N_28602,N_26276,N_27843);
xnor U28603 (N_28603,N_27520,N_27247);
xnor U28604 (N_28604,N_26146,N_26660);
xor U28605 (N_28605,N_26451,N_26516);
xor U28606 (N_28606,N_27868,N_26646);
or U28607 (N_28607,N_27879,N_27196);
nand U28608 (N_28608,N_26468,N_27446);
nor U28609 (N_28609,N_27391,N_26860);
nor U28610 (N_28610,N_27964,N_26001);
nand U28611 (N_28611,N_26794,N_27087);
or U28612 (N_28612,N_26329,N_26773);
nand U28613 (N_28613,N_27034,N_26082);
xor U28614 (N_28614,N_26755,N_26411);
xor U28615 (N_28615,N_27140,N_27043);
nand U28616 (N_28616,N_26540,N_26652);
or U28617 (N_28617,N_27995,N_27088);
nand U28618 (N_28618,N_26978,N_27792);
nor U28619 (N_28619,N_26731,N_27584);
or U28620 (N_28620,N_26430,N_26351);
or U28621 (N_28621,N_27014,N_26750);
or U28622 (N_28622,N_27664,N_27996);
and U28623 (N_28623,N_26097,N_27308);
nand U28624 (N_28624,N_27089,N_26427);
nor U28625 (N_28625,N_27728,N_26118);
nor U28626 (N_28626,N_26558,N_26541);
nor U28627 (N_28627,N_27910,N_26850);
nand U28628 (N_28628,N_26434,N_26867);
or U28629 (N_28629,N_26221,N_26585);
nor U28630 (N_28630,N_26955,N_26460);
nand U28631 (N_28631,N_27077,N_26852);
xor U28632 (N_28632,N_26618,N_26766);
xor U28633 (N_28633,N_26777,N_26362);
and U28634 (N_28634,N_26725,N_26322);
xnor U28635 (N_28635,N_27434,N_27681);
xor U28636 (N_28636,N_27682,N_27593);
nor U28637 (N_28637,N_27500,N_26912);
and U28638 (N_28638,N_27707,N_26640);
nor U28639 (N_28639,N_26675,N_26421);
or U28640 (N_28640,N_26649,N_26748);
and U28641 (N_28641,N_26981,N_26613);
xor U28642 (N_28642,N_26716,N_27153);
and U28643 (N_28643,N_27951,N_27673);
and U28644 (N_28644,N_26058,N_26503);
or U28645 (N_28645,N_26615,N_27387);
nor U28646 (N_28646,N_27831,N_26219);
nand U28647 (N_28647,N_27197,N_27818);
xor U28648 (N_28648,N_26657,N_27611);
nand U28649 (N_28649,N_27441,N_26440);
or U28650 (N_28650,N_27276,N_27489);
xnor U28651 (N_28651,N_27950,N_26549);
and U28652 (N_28652,N_26992,N_27091);
nand U28653 (N_28653,N_26747,N_27914);
or U28654 (N_28654,N_27119,N_26258);
xor U28655 (N_28655,N_27560,N_27257);
nand U28656 (N_28656,N_26825,N_27823);
xnor U28657 (N_28657,N_26372,N_26340);
or U28658 (N_28658,N_27670,N_27864);
and U28659 (N_28659,N_27456,N_27329);
or U28660 (N_28660,N_26098,N_27137);
and U28661 (N_28661,N_26283,N_27001);
or U28662 (N_28662,N_27801,N_27944);
xor U28663 (N_28663,N_26201,N_26848);
and U28664 (N_28664,N_26606,N_26563);
or U28665 (N_28665,N_26781,N_26071);
nand U28666 (N_28666,N_27621,N_26093);
and U28667 (N_28667,N_27405,N_27453);
and U28668 (N_28668,N_26906,N_27038);
and U28669 (N_28669,N_27256,N_27164);
nor U28670 (N_28670,N_27524,N_26239);
nand U28671 (N_28671,N_27291,N_27371);
and U28672 (N_28672,N_27905,N_27413);
or U28673 (N_28673,N_26939,N_27669);
or U28674 (N_28674,N_27009,N_27939);
nand U28675 (N_28675,N_26037,N_26190);
xor U28676 (N_28676,N_27320,N_26528);
or U28677 (N_28677,N_26272,N_27430);
or U28678 (N_28678,N_26774,N_26802);
and U28679 (N_28679,N_27811,N_26963);
or U28680 (N_28680,N_27797,N_26919);
xor U28681 (N_28681,N_27000,N_26936);
nor U28682 (N_28682,N_26592,N_26632);
nor U28683 (N_28683,N_26776,N_26601);
nand U28684 (N_28684,N_26712,N_27981);
or U28685 (N_28685,N_26211,N_26371);
nor U28686 (N_28686,N_27285,N_27680);
nand U28687 (N_28687,N_27316,N_26454);
nand U28688 (N_28688,N_26628,N_27627);
xnor U28689 (N_28689,N_26607,N_27410);
and U28690 (N_28690,N_27770,N_27935);
xor U28691 (N_28691,N_27004,N_27385);
or U28692 (N_28692,N_26578,N_26315);
or U28693 (N_28693,N_26840,N_26087);
or U28694 (N_28694,N_27479,N_27330);
xnor U28695 (N_28695,N_27904,N_27383);
nand U28696 (N_28696,N_27901,N_26021);
and U28697 (N_28697,N_27275,N_26141);
nor U28698 (N_28698,N_27052,N_27877);
xor U28699 (N_28699,N_26990,N_26736);
xnor U28700 (N_28700,N_26899,N_26679);
xnor U28701 (N_28701,N_27090,N_27637);
xor U28702 (N_28702,N_26399,N_27836);
nand U28703 (N_28703,N_27101,N_27557);
nor U28704 (N_28704,N_26556,N_26536);
and U28705 (N_28705,N_26501,N_26527);
and U28706 (N_28706,N_27268,N_27957);
or U28707 (N_28707,N_26470,N_26911);
or U28708 (N_28708,N_26694,N_26486);
or U28709 (N_28709,N_26938,N_27418);
nor U28710 (N_28710,N_26063,N_27601);
xor U28711 (N_28711,N_27928,N_27147);
xor U28712 (N_28712,N_26169,N_26996);
nor U28713 (N_28713,N_27725,N_27636);
xnor U28714 (N_28714,N_27938,N_27889);
nand U28715 (N_28715,N_27849,N_27989);
nand U28716 (N_28716,N_26083,N_26561);
nand U28717 (N_28717,N_26644,N_26269);
nor U28718 (N_28718,N_26488,N_26099);
and U28719 (N_28719,N_26686,N_26931);
or U28720 (N_28720,N_26944,N_27473);
and U28721 (N_28721,N_26051,N_26255);
xor U28722 (N_28722,N_27104,N_26156);
or U28723 (N_28723,N_26553,N_27067);
and U28724 (N_28724,N_26641,N_26974);
or U28725 (N_28725,N_26302,N_26122);
xor U28726 (N_28726,N_26808,N_26575);
or U28727 (N_28727,N_26170,N_27439);
nor U28728 (N_28728,N_26043,N_26143);
nand U28729 (N_28729,N_27477,N_26125);
nor U28730 (N_28730,N_27563,N_27424);
or U28731 (N_28731,N_26333,N_27302);
xor U28732 (N_28732,N_26166,N_27274);
nand U28733 (N_28733,N_27154,N_27672);
or U28734 (N_28734,N_26798,N_26028);
and U28735 (N_28735,N_26841,N_27258);
and U28736 (N_28736,N_26724,N_27068);
or U28737 (N_28737,N_27492,N_27113);
and U28738 (N_28738,N_27490,N_26203);
and U28739 (N_28739,N_26164,N_26361);
or U28740 (N_28740,N_26277,N_27404);
xnor U28741 (N_28741,N_27805,N_27231);
xor U28742 (N_28742,N_26597,N_27647);
and U28743 (N_28743,N_27058,N_27631);
or U28744 (N_28744,N_26896,N_27677);
xor U28745 (N_28745,N_26693,N_26565);
or U28746 (N_28746,N_27240,N_27862);
nor U28747 (N_28747,N_27284,N_27265);
or U28748 (N_28748,N_26842,N_26236);
nor U28749 (N_28749,N_27912,N_27748);
xnor U28750 (N_28750,N_27629,N_27915);
and U28751 (N_28751,N_27711,N_26849);
and U28752 (N_28752,N_27635,N_26509);
nor U28753 (N_28753,N_26661,N_27243);
nand U28754 (N_28754,N_26387,N_27075);
or U28755 (N_28755,N_26764,N_26056);
and U28756 (N_28756,N_27874,N_27310);
nand U28757 (N_28757,N_27018,N_27608);
nand U28758 (N_28758,N_26429,N_26257);
xor U28759 (N_28759,N_26639,N_26128);
xnor U28760 (N_28760,N_27712,N_26223);
nand U28761 (N_28761,N_26546,N_26828);
or U28762 (N_28762,N_27469,N_27312);
or U28763 (N_28763,N_26937,N_27544);
nor U28764 (N_28764,N_26642,N_27990);
and U28765 (N_28765,N_26655,N_26057);
and U28766 (N_28766,N_26134,N_27929);
xnor U28767 (N_28767,N_26915,N_27108);
or U28768 (N_28768,N_27573,N_26707);
xnor U28769 (N_28769,N_26178,N_26965);
or U28770 (N_28770,N_27428,N_27848);
and U28771 (N_28771,N_26973,N_26673);
and U28772 (N_28772,N_26379,N_27186);
xor U28773 (N_28773,N_26212,N_26210);
nand U28774 (N_28774,N_26751,N_27508);
nand U28775 (N_28775,N_26432,N_27630);
or U28776 (N_28776,N_26054,N_26260);
nand U28777 (N_28777,N_27909,N_27425);
nor U28778 (N_28778,N_26154,N_27332);
nor U28779 (N_28779,N_26359,N_26598);
or U28780 (N_28780,N_26109,N_26253);
or U28781 (N_28781,N_27654,N_26929);
and U28782 (N_28782,N_26147,N_27985);
xnor U28783 (N_28783,N_26690,N_27484);
and U28784 (N_28784,N_27582,N_26194);
xnor U28785 (N_28785,N_26078,N_27083);
nor U28786 (N_28786,N_27820,N_26999);
and U28787 (N_28787,N_27709,N_27650);
xor U28788 (N_28788,N_27545,N_27885);
nand U28789 (N_28789,N_27852,N_27570);
nor U28790 (N_28790,N_27445,N_27128);
and U28791 (N_28791,N_26953,N_27455);
nor U28792 (N_28792,N_27199,N_26985);
nand U28793 (N_28793,N_26732,N_27750);
or U28794 (N_28794,N_27059,N_26160);
nor U28795 (N_28795,N_27507,N_27735);
nor U28796 (N_28796,N_27161,N_27298);
nor U28797 (N_28797,N_27703,N_27355);
nor U28798 (N_28798,N_27589,N_26181);
nor U28799 (N_28799,N_26864,N_26453);
or U28800 (N_28800,N_27562,N_27955);
or U28801 (N_28801,N_27689,N_27095);
nor U28802 (N_28802,N_27802,N_27156);
xnor U28803 (N_28803,N_27028,N_27304);
xor U28804 (N_28804,N_27844,N_26055);
and U28805 (N_28805,N_26908,N_27992);
xor U28806 (N_28806,N_27100,N_27053);
xor U28807 (N_28807,N_26151,N_26526);
and U28808 (N_28808,N_27382,N_27898);
and U28809 (N_28809,N_27918,N_26422);
nand U28810 (N_28810,N_27223,N_27925);
nand U28811 (N_28811,N_27798,N_27030);
nor U28812 (N_28812,N_27594,N_26293);
nor U28813 (N_28813,N_26596,N_27571);
xnor U28814 (N_28814,N_27810,N_26822);
or U28815 (N_28815,N_27812,N_27061);
and U28816 (N_28816,N_26448,N_26065);
nand U28817 (N_28817,N_26378,N_27786);
nand U28818 (N_28818,N_27967,N_27527);
nor U28819 (N_28819,N_27016,N_27639);
and U28820 (N_28820,N_26172,N_27447);
or U28821 (N_28821,N_26264,N_26282);
xnor U28822 (N_28822,N_26111,N_27658);
and U28823 (N_28823,N_27747,N_27155);
nand U28824 (N_28824,N_26073,N_27746);
xor U28825 (N_28825,N_27372,N_26182);
nor U28826 (N_28826,N_27081,N_26217);
or U28827 (N_28827,N_26885,N_26490);
nand U28828 (N_28828,N_26874,N_26638);
nor U28829 (N_28829,N_26466,N_27094);
or U28830 (N_28830,N_27952,N_26479);
xor U28831 (N_28831,N_27947,N_26851);
and U28832 (N_28832,N_26205,N_26308);
nor U28833 (N_28833,N_27460,N_26226);
xor U28834 (N_28834,N_26545,N_27065);
xnor U28835 (N_28835,N_26943,N_27374);
nand U28836 (N_28836,N_27988,N_27873);
nor U28837 (N_28837,N_26298,N_26080);
nand U28838 (N_28838,N_27574,N_26406);
xor U28839 (N_28839,N_26498,N_26337);
and U28840 (N_28840,N_26185,N_27875);
and U28841 (N_28841,N_27599,N_27042);
nand U28842 (N_28842,N_27632,N_26654);
xor U28843 (N_28843,N_26728,N_27867);
nor U28844 (N_28844,N_26791,N_26746);
or U28845 (N_28845,N_27547,N_27983);
or U28846 (N_28846,N_26155,N_26942);
nor U28847 (N_28847,N_26847,N_27854);
and U28848 (N_28848,N_27432,N_26091);
or U28849 (N_28849,N_27963,N_27720);
nand U28850 (N_28850,N_27776,N_26560);
and U28851 (N_28851,N_27181,N_26559);
or U28852 (N_28852,N_26717,N_26763);
and U28853 (N_28853,N_27251,N_26070);
xor U28854 (N_28854,N_26310,N_26331);
nand U28855 (N_28855,N_26954,N_26047);
nand U28856 (N_28856,N_27936,N_27272);
nor U28857 (N_28857,N_27596,N_26034);
nand U28858 (N_28858,N_27998,N_27348);
and U28859 (N_28859,N_27379,N_26494);
or U28860 (N_28860,N_27488,N_27826);
and U28861 (N_28861,N_26426,N_27590);
xnor U28862 (N_28862,N_27342,N_27204);
xor U28863 (N_28863,N_27474,N_27066);
nand U28864 (N_28864,N_27921,N_27253);
nand U28865 (N_28865,N_27558,N_27692);
nand U28866 (N_28866,N_26916,N_26500);
and U28867 (N_28867,N_27267,N_27420);
or U28868 (N_28868,N_27431,N_26517);
xnor U28869 (N_28869,N_27209,N_26368);
and U28870 (N_28870,N_27224,N_26603);
and U28871 (N_28871,N_26800,N_27598);
nor U28872 (N_28872,N_27927,N_27467);
xor U28873 (N_28873,N_27853,N_27073);
and U28874 (N_28874,N_27476,N_27572);
nand U28875 (N_28875,N_27442,N_27399);
nand U28876 (N_28876,N_26404,N_26665);
or U28877 (N_28877,N_27093,N_26408);
nand U28878 (N_28878,N_26167,N_27436);
and U28879 (N_28879,N_26003,N_26245);
nand U28880 (N_28880,N_26347,N_27815);
or U28881 (N_28881,N_27225,N_26482);
nand U28882 (N_28882,N_27132,N_27151);
nor U28883 (N_28883,N_26469,N_26036);
and U28884 (N_28884,N_27141,N_27919);
nand U28885 (N_28885,N_26668,N_27587);
and U28886 (N_28886,N_26976,N_27226);
or U28887 (N_28887,N_26804,N_27462);
nor U28888 (N_28888,N_26101,N_27246);
nor U28889 (N_28889,N_27098,N_27817);
nand U28890 (N_28890,N_27795,N_26972);
nor U28891 (N_28891,N_27321,N_26905);
or U28892 (N_28892,N_26477,N_27017);
nand U28893 (N_28893,N_27211,N_26384);
nor U28894 (N_28894,N_26081,N_27651);
or U28895 (N_28895,N_27624,N_26616);
xor U28896 (N_28896,N_27751,N_26354);
or U28897 (N_28897,N_26019,N_26005);
nor U28898 (N_28898,N_26388,N_26320);
and U28899 (N_28899,N_27135,N_27814);
xor U28900 (N_28900,N_26290,N_27421);
xor U28901 (N_28901,N_27180,N_26604);
or U28902 (N_28902,N_26189,N_27408);
or U28903 (N_28903,N_27306,N_26608);
nor U28904 (N_28904,N_27416,N_26564);
or U28905 (N_28905,N_27194,N_27143);
nor U28906 (N_28906,N_26815,N_26715);
nand U28907 (N_28907,N_26139,N_27859);
nand U28908 (N_28908,N_26907,N_26533);
nor U28909 (N_28909,N_27727,N_27309);
xor U28910 (N_28910,N_27871,N_27478);
or U28911 (N_28911,N_27401,N_26409);
nand U28912 (N_28912,N_27323,N_26629);
xnor U28913 (N_28913,N_26442,N_27916);
nand U28914 (N_28914,N_27451,N_26425);
or U28915 (N_28915,N_27148,N_26476);
xor U28916 (N_28916,N_26770,N_26480);
or U28917 (N_28917,N_26438,N_26496);
or U28918 (N_28918,N_26722,N_27341);
or U28919 (N_28919,N_27911,N_26202);
nand U28920 (N_28920,N_27422,N_27600);
and U28921 (N_28921,N_27032,N_27665);
or U28922 (N_28922,N_27295,N_27390);
or U28923 (N_28923,N_27035,N_27496);
xnor U28924 (N_28924,N_26095,N_26877);
or U28925 (N_28925,N_27419,N_27742);
nor U28926 (N_28926,N_27237,N_26740);
xor U28927 (N_28927,N_27340,N_27046);
and U28928 (N_28928,N_27118,N_26452);
and U28929 (N_28929,N_27903,N_26769);
nand U28930 (N_28930,N_27838,N_26117);
and U28931 (N_28931,N_26897,N_27234);
or U28932 (N_28932,N_27023,N_26431);
xnor U28933 (N_28933,N_26551,N_26982);
and U28934 (N_28934,N_27617,N_26216);
xnor U28935 (N_28935,N_26187,N_26002);
xnor U28936 (N_28936,N_26515,N_26727);
and U28937 (N_28937,N_26235,N_27819);
or U28938 (N_28938,N_27530,N_27096);
or U28939 (N_28939,N_27675,N_26338);
and U28940 (N_28940,N_26512,N_27213);
or U28941 (N_28941,N_27718,N_26032);
and U28942 (N_28942,N_26004,N_26130);
xnor U28943 (N_28943,N_26045,N_27857);
nor U28944 (N_28944,N_26317,N_26405);
or U28945 (N_28945,N_26484,N_26658);
and U28946 (N_28946,N_26544,N_26349);
xor U28947 (N_28947,N_26671,N_26807);
nand U28948 (N_28948,N_27216,N_26941);
and U28949 (N_28949,N_27502,N_27228);
and U28950 (N_28950,N_26085,N_26743);
xor U28951 (N_28951,N_27078,N_27791);
nand U28952 (N_28952,N_27361,N_27782);
xnor U28953 (N_28953,N_27483,N_26013);
nand U28954 (N_28954,N_26040,N_27691);
and U28955 (N_28955,N_27426,N_26370);
xor U28956 (N_28956,N_26112,N_27973);
xnor U28957 (N_28957,N_26589,N_27183);
nand U28958 (N_28958,N_27160,N_27603);
and U28959 (N_28959,N_26998,N_26886);
and U28960 (N_28960,N_27071,N_26696);
xnor U28961 (N_28961,N_27354,N_27523);
nor U28962 (N_28962,N_26813,N_26356);
nor U28963 (N_28963,N_26757,N_26904);
nor U28964 (N_28964,N_26268,N_27847);
nor U28965 (N_28965,N_26677,N_26935);
xor U28966 (N_28966,N_26077,N_27917);
nor U28967 (N_28967,N_27048,N_26922);
and U28968 (N_28968,N_26570,N_26785);
nor U28969 (N_28969,N_27202,N_27363);
nor U28970 (N_28970,N_27121,N_27605);
xnor U28971 (N_28971,N_27495,N_27863);
nor U28972 (N_28972,N_27807,N_27561);
nand U28973 (N_28973,N_27833,N_26413);
or U28974 (N_28974,N_26730,N_27832);
nand U28975 (N_28975,N_27168,N_26521);
or U28976 (N_28976,N_26803,N_26881);
xor U28977 (N_28977,N_27697,N_26428);
and U28978 (N_28978,N_26593,N_27292);
nand U28979 (N_28979,N_26369,N_26023);
and U28980 (N_28980,N_26801,N_26385);
or U28981 (N_28981,N_26145,N_27123);
xnor U28982 (N_28982,N_26061,N_26862);
xnor U28983 (N_28983,N_27521,N_27192);
and U28984 (N_28984,N_26416,N_26195);
or U28985 (N_28985,N_26450,N_27112);
nand U28986 (N_28986,N_26756,N_26958);
nand U28987 (N_28987,N_26234,N_27040);
or U28988 (N_28988,N_27324,N_26064);
or U28989 (N_28989,N_27397,N_26296);
or U28990 (N_28990,N_26124,N_27855);
xnor U28991 (N_28991,N_27498,N_27965);
or U28992 (N_28992,N_26522,N_26692);
and U28993 (N_28993,N_27733,N_26252);
nor U28994 (N_28994,N_26979,N_27773);
nand U28995 (N_28995,N_26697,N_26865);
xor U28996 (N_28996,N_26926,N_26463);
xor U28997 (N_28997,N_27266,N_27388);
nand U28998 (N_28998,N_27013,N_26685);
nor U28999 (N_28999,N_27538,N_26721);
xnor U29000 (N_29000,N_27609,N_27498);
nand U29001 (N_29001,N_27984,N_27724);
nor U29002 (N_29002,N_27773,N_26902);
or U29003 (N_29003,N_26689,N_27807);
and U29004 (N_29004,N_26427,N_27488);
nand U29005 (N_29005,N_26449,N_27891);
nand U29006 (N_29006,N_26337,N_26640);
or U29007 (N_29007,N_26875,N_26573);
nor U29008 (N_29008,N_26467,N_27570);
nand U29009 (N_29009,N_26731,N_27734);
or U29010 (N_29010,N_26338,N_27017);
nor U29011 (N_29011,N_26438,N_27563);
and U29012 (N_29012,N_26329,N_27901);
or U29013 (N_29013,N_27630,N_27697);
nand U29014 (N_29014,N_26280,N_26597);
and U29015 (N_29015,N_27971,N_27169);
nor U29016 (N_29016,N_26309,N_26367);
xor U29017 (N_29017,N_26106,N_26798);
xnor U29018 (N_29018,N_27324,N_26052);
and U29019 (N_29019,N_26542,N_26523);
nor U29020 (N_29020,N_26394,N_26294);
nand U29021 (N_29021,N_26465,N_26064);
xnor U29022 (N_29022,N_26691,N_27369);
nand U29023 (N_29023,N_26755,N_26082);
xnor U29024 (N_29024,N_26890,N_27862);
or U29025 (N_29025,N_27769,N_27775);
xnor U29026 (N_29026,N_27384,N_27082);
or U29027 (N_29027,N_26566,N_26693);
xnor U29028 (N_29028,N_26473,N_27034);
and U29029 (N_29029,N_26100,N_26817);
nand U29030 (N_29030,N_27957,N_27032);
or U29031 (N_29031,N_27682,N_27931);
or U29032 (N_29032,N_26745,N_26757);
xnor U29033 (N_29033,N_27844,N_27015);
or U29034 (N_29034,N_26039,N_27871);
and U29035 (N_29035,N_26550,N_26628);
or U29036 (N_29036,N_27699,N_26644);
nand U29037 (N_29037,N_26580,N_26104);
xnor U29038 (N_29038,N_27207,N_26377);
xnor U29039 (N_29039,N_26557,N_27195);
and U29040 (N_29040,N_27606,N_26878);
and U29041 (N_29041,N_27628,N_27859);
or U29042 (N_29042,N_26804,N_27806);
nand U29043 (N_29043,N_26888,N_26153);
xnor U29044 (N_29044,N_27300,N_27756);
xnor U29045 (N_29045,N_27399,N_26072);
or U29046 (N_29046,N_26028,N_27420);
nand U29047 (N_29047,N_27702,N_26662);
nand U29048 (N_29048,N_27605,N_27675);
nor U29049 (N_29049,N_27487,N_26679);
nand U29050 (N_29050,N_27391,N_26154);
and U29051 (N_29051,N_26688,N_26443);
and U29052 (N_29052,N_27174,N_27734);
xnor U29053 (N_29053,N_27084,N_26259);
nor U29054 (N_29054,N_26181,N_26404);
or U29055 (N_29055,N_27865,N_27625);
and U29056 (N_29056,N_27834,N_27999);
xnor U29057 (N_29057,N_26289,N_26642);
and U29058 (N_29058,N_26275,N_27274);
or U29059 (N_29059,N_26986,N_26970);
xnor U29060 (N_29060,N_26403,N_26697);
nand U29061 (N_29061,N_27536,N_26959);
nand U29062 (N_29062,N_27765,N_26005);
nor U29063 (N_29063,N_26979,N_26036);
or U29064 (N_29064,N_27973,N_27406);
or U29065 (N_29065,N_27304,N_26250);
and U29066 (N_29066,N_26316,N_27275);
xor U29067 (N_29067,N_26555,N_26659);
or U29068 (N_29068,N_26078,N_26786);
nor U29069 (N_29069,N_27818,N_26707);
nand U29070 (N_29070,N_26970,N_27020);
xor U29071 (N_29071,N_27384,N_26352);
nand U29072 (N_29072,N_26722,N_27216);
xor U29073 (N_29073,N_27562,N_26021);
or U29074 (N_29074,N_26078,N_27026);
or U29075 (N_29075,N_26380,N_26693);
nor U29076 (N_29076,N_26398,N_26242);
xor U29077 (N_29077,N_26044,N_26294);
xnor U29078 (N_29078,N_27099,N_27700);
and U29079 (N_29079,N_26559,N_27213);
or U29080 (N_29080,N_26055,N_27139);
nand U29081 (N_29081,N_26643,N_26119);
xnor U29082 (N_29082,N_26985,N_27447);
xor U29083 (N_29083,N_26137,N_26431);
and U29084 (N_29084,N_26453,N_27593);
xor U29085 (N_29085,N_26833,N_27078);
or U29086 (N_29086,N_26741,N_27452);
nand U29087 (N_29087,N_26657,N_27647);
and U29088 (N_29088,N_26629,N_27413);
nand U29089 (N_29089,N_27827,N_27023);
and U29090 (N_29090,N_27038,N_26800);
and U29091 (N_29091,N_26271,N_27608);
xnor U29092 (N_29092,N_26336,N_26627);
or U29093 (N_29093,N_27091,N_27908);
or U29094 (N_29094,N_27716,N_26545);
nand U29095 (N_29095,N_27677,N_26110);
nand U29096 (N_29096,N_26474,N_27025);
nand U29097 (N_29097,N_27612,N_26055);
nand U29098 (N_29098,N_26539,N_27238);
or U29099 (N_29099,N_26468,N_27442);
and U29100 (N_29100,N_27756,N_27451);
nor U29101 (N_29101,N_27155,N_26645);
xor U29102 (N_29102,N_27893,N_26701);
xor U29103 (N_29103,N_27439,N_27947);
nand U29104 (N_29104,N_26806,N_26136);
nand U29105 (N_29105,N_27525,N_27928);
nand U29106 (N_29106,N_26793,N_27814);
or U29107 (N_29107,N_26482,N_27658);
xor U29108 (N_29108,N_26130,N_26141);
or U29109 (N_29109,N_27140,N_27480);
or U29110 (N_29110,N_27355,N_26816);
nand U29111 (N_29111,N_27403,N_26803);
and U29112 (N_29112,N_26385,N_27774);
or U29113 (N_29113,N_27534,N_27582);
nand U29114 (N_29114,N_26343,N_26901);
and U29115 (N_29115,N_26970,N_27662);
nand U29116 (N_29116,N_27024,N_26936);
nand U29117 (N_29117,N_26263,N_26008);
nor U29118 (N_29118,N_26653,N_26667);
nor U29119 (N_29119,N_26196,N_26123);
and U29120 (N_29120,N_27108,N_26250);
nand U29121 (N_29121,N_27843,N_27003);
nand U29122 (N_29122,N_27300,N_26497);
nor U29123 (N_29123,N_26893,N_26684);
xnor U29124 (N_29124,N_26052,N_27430);
nand U29125 (N_29125,N_27750,N_27108);
xor U29126 (N_29126,N_26654,N_27834);
or U29127 (N_29127,N_27096,N_27819);
nand U29128 (N_29128,N_26649,N_27941);
nand U29129 (N_29129,N_27309,N_27218);
and U29130 (N_29130,N_26719,N_27159);
and U29131 (N_29131,N_26232,N_26944);
or U29132 (N_29132,N_26015,N_26123);
and U29133 (N_29133,N_26730,N_26565);
nor U29134 (N_29134,N_26625,N_27837);
xnor U29135 (N_29135,N_26365,N_26046);
or U29136 (N_29136,N_26195,N_26264);
nor U29137 (N_29137,N_27889,N_26559);
or U29138 (N_29138,N_27133,N_27130);
nor U29139 (N_29139,N_26152,N_27821);
xnor U29140 (N_29140,N_26686,N_27972);
or U29141 (N_29141,N_26983,N_27337);
nor U29142 (N_29142,N_27235,N_26634);
and U29143 (N_29143,N_26511,N_26914);
or U29144 (N_29144,N_27161,N_27568);
nor U29145 (N_29145,N_27213,N_26691);
nor U29146 (N_29146,N_26695,N_26681);
xor U29147 (N_29147,N_27721,N_27453);
nor U29148 (N_29148,N_27627,N_27354);
or U29149 (N_29149,N_27042,N_26855);
nor U29150 (N_29150,N_26660,N_27351);
nand U29151 (N_29151,N_26648,N_26806);
and U29152 (N_29152,N_26976,N_26908);
and U29153 (N_29153,N_27062,N_27470);
and U29154 (N_29154,N_27721,N_26712);
or U29155 (N_29155,N_27109,N_27370);
nand U29156 (N_29156,N_26377,N_26146);
and U29157 (N_29157,N_26828,N_27481);
nor U29158 (N_29158,N_26342,N_26827);
or U29159 (N_29159,N_27744,N_27138);
nor U29160 (N_29160,N_27699,N_27707);
nand U29161 (N_29161,N_27040,N_27744);
nand U29162 (N_29162,N_26305,N_26978);
and U29163 (N_29163,N_26088,N_26469);
or U29164 (N_29164,N_26157,N_27984);
or U29165 (N_29165,N_26031,N_26591);
xor U29166 (N_29166,N_26584,N_27300);
or U29167 (N_29167,N_26811,N_26784);
nor U29168 (N_29168,N_26189,N_27993);
and U29169 (N_29169,N_26069,N_26498);
nand U29170 (N_29170,N_27074,N_26802);
nand U29171 (N_29171,N_27294,N_26790);
and U29172 (N_29172,N_27853,N_26762);
or U29173 (N_29173,N_27728,N_26278);
and U29174 (N_29174,N_26847,N_26499);
nor U29175 (N_29175,N_27807,N_27565);
nand U29176 (N_29176,N_27824,N_27052);
and U29177 (N_29177,N_27609,N_26754);
nor U29178 (N_29178,N_27672,N_26570);
or U29179 (N_29179,N_27957,N_26205);
and U29180 (N_29180,N_27183,N_26904);
xor U29181 (N_29181,N_27254,N_26553);
xnor U29182 (N_29182,N_27181,N_26331);
nor U29183 (N_29183,N_26837,N_26168);
nor U29184 (N_29184,N_27703,N_26510);
nor U29185 (N_29185,N_26054,N_27559);
nand U29186 (N_29186,N_27375,N_27190);
or U29187 (N_29187,N_27081,N_26277);
or U29188 (N_29188,N_26242,N_27039);
xor U29189 (N_29189,N_27521,N_26712);
and U29190 (N_29190,N_26444,N_26871);
xor U29191 (N_29191,N_27040,N_27905);
or U29192 (N_29192,N_26189,N_27036);
and U29193 (N_29193,N_27736,N_26847);
and U29194 (N_29194,N_26923,N_27923);
nand U29195 (N_29195,N_27970,N_27385);
nand U29196 (N_29196,N_26054,N_27575);
nand U29197 (N_29197,N_27878,N_27180);
nor U29198 (N_29198,N_26134,N_26609);
and U29199 (N_29199,N_26681,N_26676);
nand U29200 (N_29200,N_27532,N_26992);
or U29201 (N_29201,N_26287,N_27422);
nand U29202 (N_29202,N_27564,N_27046);
and U29203 (N_29203,N_26830,N_26896);
xor U29204 (N_29204,N_27621,N_27666);
xor U29205 (N_29205,N_26083,N_26246);
xor U29206 (N_29206,N_27329,N_26272);
nand U29207 (N_29207,N_26375,N_27231);
and U29208 (N_29208,N_26079,N_26478);
xnor U29209 (N_29209,N_26475,N_26575);
xnor U29210 (N_29210,N_26673,N_26838);
and U29211 (N_29211,N_27507,N_26155);
nand U29212 (N_29212,N_26152,N_27498);
nand U29213 (N_29213,N_26186,N_26626);
xnor U29214 (N_29214,N_27036,N_27947);
nand U29215 (N_29215,N_26154,N_27881);
and U29216 (N_29216,N_27066,N_26367);
or U29217 (N_29217,N_26445,N_27274);
and U29218 (N_29218,N_26451,N_27246);
and U29219 (N_29219,N_26298,N_26256);
nor U29220 (N_29220,N_27467,N_27190);
xor U29221 (N_29221,N_27896,N_27285);
xor U29222 (N_29222,N_27057,N_27784);
nand U29223 (N_29223,N_26034,N_26310);
nor U29224 (N_29224,N_26514,N_26051);
and U29225 (N_29225,N_26159,N_27257);
or U29226 (N_29226,N_27005,N_27953);
nor U29227 (N_29227,N_27786,N_27681);
nor U29228 (N_29228,N_27699,N_26814);
and U29229 (N_29229,N_27345,N_27493);
or U29230 (N_29230,N_26339,N_26611);
xor U29231 (N_29231,N_27070,N_27023);
and U29232 (N_29232,N_27189,N_26725);
xnor U29233 (N_29233,N_26083,N_26394);
nor U29234 (N_29234,N_27144,N_26568);
xor U29235 (N_29235,N_26274,N_26091);
nor U29236 (N_29236,N_27709,N_26969);
or U29237 (N_29237,N_27576,N_26699);
xor U29238 (N_29238,N_26271,N_26784);
nand U29239 (N_29239,N_26564,N_26945);
and U29240 (N_29240,N_27613,N_27244);
and U29241 (N_29241,N_27504,N_26763);
xor U29242 (N_29242,N_27933,N_26061);
and U29243 (N_29243,N_26971,N_26868);
nand U29244 (N_29244,N_26147,N_26412);
nor U29245 (N_29245,N_27515,N_27170);
or U29246 (N_29246,N_26214,N_26475);
nand U29247 (N_29247,N_26430,N_27557);
nor U29248 (N_29248,N_27898,N_26650);
nand U29249 (N_29249,N_26022,N_27627);
and U29250 (N_29250,N_27199,N_27597);
and U29251 (N_29251,N_27559,N_27123);
xnor U29252 (N_29252,N_27502,N_27191);
and U29253 (N_29253,N_27694,N_27449);
nor U29254 (N_29254,N_27863,N_27116);
nor U29255 (N_29255,N_27351,N_26369);
or U29256 (N_29256,N_27951,N_27140);
nand U29257 (N_29257,N_27052,N_26709);
or U29258 (N_29258,N_27536,N_26674);
or U29259 (N_29259,N_26611,N_27508);
nor U29260 (N_29260,N_26954,N_27151);
nor U29261 (N_29261,N_27456,N_27634);
nand U29262 (N_29262,N_26350,N_26885);
xor U29263 (N_29263,N_27469,N_27515);
xor U29264 (N_29264,N_26907,N_27615);
or U29265 (N_29265,N_26391,N_26791);
nor U29266 (N_29266,N_26576,N_26361);
and U29267 (N_29267,N_26143,N_26514);
nand U29268 (N_29268,N_26977,N_27307);
xnor U29269 (N_29269,N_27920,N_27883);
or U29270 (N_29270,N_26707,N_26109);
nor U29271 (N_29271,N_26596,N_26633);
and U29272 (N_29272,N_26619,N_26298);
nor U29273 (N_29273,N_26034,N_27991);
or U29274 (N_29274,N_26438,N_27568);
nor U29275 (N_29275,N_27012,N_27571);
xor U29276 (N_29276,N_27327,N_27816);
nor U29277 (N_29277,N_26396,N_27226);
xor U29278 (N_29278,N_26040,N_27147);
or U29279 (N_29279,N_26655,N_27363);
nand U29280 (N_29280,N_27422,N_27651);
or U29281 (N_29281,N_26577,N_26793);
or U29282 (N_29282,N_26563,N_26543);
nand U29283 (N_29283,N_27043,N_27915);
and U29284 (N_29284,N_26659,N_26414);
nand U29285 (N_29285,N_26707,N_27157);
and U29286 (N_29286,N_27516,N_26098);
nor U29287 (N_29287,N_27435,N_26759);
nand U29288 (N_29288,N_26214,N_26890);
xor U29289 (N_29289,N_27777,N_26342);
nor U29290 (N_29290,N_26441,N_27115);
and U29291 (N_29291,N_27006,N_27588);
and U29292 (N_29292,N_26030,N_26472);
nor U29293 (N_29293,N_26519,N_26741);
xnor U29294 (N_29294,N_26325,N_27310);
or U29295 (N_29295,N_27246,N_26098);
xnor U29296 (N_29296,N_27100,N_27569);
nor U29297 (N_29297,N_26527,N_27694);
or U29298 (N_29298,N_27521,N_27399);
xor U29299 (N_29299,N_26258,N_26140);
nor U29300 (N_29300,N_27084,N_26990);
nand U29301 (N_29301,N_26380,N_26728);
or U29302 (N_29302,N_26378,N_27491);
nor U29303 (N_29303,N_26322,N_26252);
nand U29304 (N_29304,N_26551,N_26779);
xor U29305 (N_29305,N_26249,N_26988);
and U29306 (N_29306,N_27985,N_27698);
nor U29307 (N_29307,N_26951,N_26063);
xor U29308 (N_29308,N_27929,N_26504);
nor U29309 (N_29309,N_26514,N_26229);
nand U29310 (N_29310,N_27008,N_27191);
and U29311 (N_29311,N_27487,N_27223);
nor U29312 (N_29312,N_26931,N_26199);
nor U29313 (N_29313,N_26714,N_27367);
nand U29314 (N_29314,N_26772,N_27506);
xnor U29315 (N_29315,N_26259,N_26004);
or U29316 (N_29316,N_27116,N_26541);
and U29317 (N_29317,N_27305,N_26588);
nor U29318 (N_29318,N_26818,N_26897);
nand U29319 (N_29319,N_26718,N_26311);
or U29320 (N_29320,N_27516,N_26204);
nor U29321 (N_29321,N_27713,N_26634);
or U29322 (N_29322,N_26561,N_26442);
or U29323 (N_29323,N_26376,N_26848);
or U29324 (N_29324,N_26452,N_26776);
xnor U29325 (N_29325,N_27058,N_27627);
or U29326 (N_29326,N_26809,N_26608);
or U29327 (N_29327,N_27034,N_27869);
nand U29328 (N_29328,N_27574,N_26562);
xor U29329 (N_29329,N_26370,N_26950);
nor U29330 (N_29330,N_26255,N_26374);
nor U29331 (N_29331,N_26202,N_27800);
xnor U29332 (N_29332,N_27788,N_26390);
xor U29333 (N_29333,N_26181,N_27175);
nor U29334 (N_29334,N_27529,N_27511);
xnor U29335 (N_29335,N_27816,N_26049);
and U29336 (N_29336,N_26363,N_27475);
xnor U29337 (N_29337,N_27081,N_26570);
nor U29338 (N_29338,N_26024,N_27933);
or U29339 (N_29339,N_26555,N_27507);
xnor U29340 (N_29340,N_27730,N_26406);
and U29341 (N_29341,N_26277,N_26075);
and U29342 (N_29342,N_26579,N_26963);
nand U29343 (N_29343,N_26673,N_27549);
and U29344 (N_29344,N_27163,N_27864);
nor U29345 (N_29345,N_27194,N_26608);
xnor U29346 (N_29346,N_27203,N_26794);
or U29347 (N_29347,N_26322,N_26659);
xor U29348 (N_29348,N_27618,N_26984);
and U29349 (N_29349,N_27361,N_26259);
xnor U29350 (N_29350,N_27837,N_27912);
nand U29351 (N_29351,N_26587,N_26170);
and U29352 (N_29352,N_27570,N_26382);
xnor U29353 (N_29353,N_27842,N_27695);
nor U29354 (N_29354,N_26053,N_27854);
xnor U29355 (N_29355,N_27813,N_27748);
xnor U29356 (N_29356,N_27627,N_26877);
or U29357 (N_29357,N_27809,N_26671);
xnor U29358 (N_29358,N_27293,N_27933);
and U29359 (N_29359,N_26673,N_27630);
or U29360 (N_29360,N_27829,N_27693);
nand U29361 (N_29361,N_27591,N_26104);
nor U29362 (N_29362,N_27726,N_27772);
xnor U29363 (N_29363,N_26716,N_26006);
and U29364 (N_29364,N_27464,N_27740);
and U29365 (N_29365,N_26532,N_27917);
nor U29366 (N_29366,N_26159,N_27859);
nand U29367 (N_29367,N_26300,N_27067);
nand U29368 (N_29368,N_26181,N_26876);
and U29369 (N_29369,N_26362,N_26699);
nand U29370 (N_29370,N_26783,N_27084);
xnor U29371 (N_29371,N_27323,N_27597);
nor U29372 (N_29372,N_27149,N_27957);
or U29373 (N_29373,N_27423,N_26155);
xnor U29374 (N_29374,N_27379,N_26869);
xnor U29375 (N_29375,N_26484,N_27803);
or U29376 (N_29376,N_27872,N_27210);
nand U29377 (N_29377,N_27957,N_26334);
nand U29378 (N_29378,N_27418,N_27000);
nor U29379 (N_29379,N_26045,N_27484);
and U29380 (N_29380,N_27685,N_27621);
nor U29381 (N_29381,N_26073,N_26106);
nand U29382 (N_29382,N_26246,N_27513);
xnor U29383 (N_29383,N_27011,N_26169);
and U29384 (N_29384,N_26841,N_27862);
and U29385 (N_29385,N_27117,N_26337);
or U29386 (N_29386,N_26302,N_26523);
or U29387 (N_29387,N_26409,N_27257);
or U29388 (N_29388,N_27739,N_26116);
nor U29389 (N_29389,N_27127,N_26557);
nor U29390 (N_29390,N_26562,N_26889);
nand U29391 (N_29391,N_26569,N_27972);
xnor U29392 (N_29392,N_27251,N_26731);
or U29393 (N_29393,N_26023,N_26705);
xor U29394 (N_29394,N_26569,N_26165);
nand U29395 (N_29395,N_27953,N_27392);
and U29396 (N_29396,N_26342,N_26781);
nor U29397 (N_29397,N_26253,N_27800);
and U29398 (N_29398,N_27010,N_27881);
nand U29399 (N_29399,N_26787,N_26705);
xnor U29400 (N_29400,N_26031,N_26752);
or U29401 (N_29401,N_26724,N_27884);
or U29402 (N_29402,N_27485,N_27302);
and U29403 (N_29403,N_27069,N_26891);
nor U29404 (N_29404,N_26861,N_26104);
nand U29405 (N_29405,N_27529,N_26037);
and U29406 (N_29406,N_26550,N_27952);
xor U29407 (N_29407,N_27045,N_26615);
or U29408 (N_29408,N_26441,N_26935);
nor U29409 (N_29409,N_27333,N_27981);
or U29410 (N_29410,N_26807,N_26932);
and U29411 (N_29411,N_27566,N_26178);
nand U29412 (N_29412,N_27652,N_27072);
nand U29413 (N_29413,N_27280,N_27869);
xor U29414 (N_29414,N_26475,N_27488);
or U29415 (N_29415,N_27875,N_27098);
xor U29416 (N_29416,N_26049,N_26910);
and U29417 (N_29417,N_26598,N_26525);
and U29418 (N_29418,N_26655,N_27468);
nor U29419 (N_29419,N_27802,N_26870);
xor U29420 (N_29420,N_27548,N_26185);
and U29421 (N_29421,N_27155,N_27890);
and U29422 (N_29422,N_26633,N_27789);
or U29423 (N_29423,N_26443,N_26196);
or U29424 (N_29424,N_26262,N_27762);
and U29425 (N_29425,N_26637,N_26564);
and U29426 (N_29426,N_27848,N_27505);
and U29427 (N_29427,N_26871,N_26147);
nand U29428 (N_29428,N_27530,N_27374);
xnor U29429 (N_29429,N_26164,N_26123);
nor U29430 (N_29430,N_27673,N_27533);
xor U29431 (N_29431,N_27318,N_26427);
and U29432 (N_29432,N_27196,N_27357);
or U29433 (N_29433,N_26886,N_27578);
nor U29434 (N_29434,N_27564,N_26005);
or U29435 (N_29435,N_26255,N_27557);
and U29436 (N_29436,N_27092,N_26717);
or U29437 (N_29437,N_27979,N_26956);
or U29438 (N_29438,N_26931,N_26713);
xor U29439 (N_29439,N_26723,N_26732);
xnor U29440 (N_29440,N_27997,N_26664);
nand U29441 (N_29441,N_26489,N_27130);
xnor U29442 (N_29442,N_26478,N_26149);
xnor U29443 (N_29443,N_27714,N_27066);
nor U29444 (N_29444,N_27570,N_27456);
nor U29445 (N_29445,N_27481,N_27714);
nand U29446 (N_29446,N_26012,N_26710);
and U29447 (N_29447,N_26804,N_26461);
or U29448 (N_29448,N_26912,N_27376);
or U29449 (N_29449,N_26368,N_26937);
nor U29450 (N_29450,N_27117,N_27264);
nand U29451 (N_29451,N_26306,N_27095);
and U29452 (N_29452,N_27590,N_27173);
nand U29453 (N_29453,N_27975,N_26009);
or U29454 (N_29454,N_26037,N_26937);
and U29455 (N_29455,N_27728,N_27015);
or U29456 (N_29456,N_26862,N_27015);
or U29457 (N_29457,N_26158,N_26790);
nor U29458 (N_29458,N_26153,N_26316);
nand U29459 (N_29459,N_26150,N_27381);
and U29460 (N_29460,N_26646,N_26890);
nor U29461 (N_29461,N_26886,N_26933);
and U29462 (N_29462,N_27704,N_27645);
xor U29463 (N_29463,N_27158,N_26108);
nor U29464 (N_29464,N_26420,N_26537);
or U29465 (N_29465,N_26889,N_26488);
nor U29466 (N_29466,N_26657,N_26607);
nand U29467 (N_29467,N_27230,N_26633);
xor U29468 (N_29468,N_27110,N_26151);
and U29469 (N_29469,N_27743,N_26074);
nand U29470 (N_29470,N_26319,N_27269);
xnor U29471 (N_29471,N_27683,N_26063);
nor U29472 (N_29472,N_26242,N_26848);
nor U29473 (N_29473,N_26625,N_27943);
and U29474 (N_29474,N_26825,N_27091);
and U29475 (N_29475,N_26927,N_26446);
nand U29476 (N_29476,N_27597,N_26364);
nand U29477 (N_29477,N_26570,N_27246);
nor U29478 (N_29478,N_26297,N_27522);
nor U29479 (N_29479,N_26966,N_27843);
xor U29480 (N_29480,N_26039,N_27526);
or U29481 (N_29481,N_26864,N_27210);
and U29482 (N_29482,N_27006,N_27280);
or U29483 (N_29483,N_27485,N_26205);
xor U29484 (N_29484,N_26713,N_26029);
nand U29485 (N_29485,N_27389,N_27603);
and U29486 (N_29486,N_26172,N_27648);
or U29487 (N_29487,N_26054,N_27655);
xnor U29488 (N_29488,N_26779,N_27640);
and U29489 (N_29489,N_27414,N_26833);
or U29490 (N_29490,N_26136,N_27372);
xnor U29491 (N_29491,N_26459,N_27461);
nor U29492 (N_29492,N_26064,N_26721);
nand U29493 (N_29493,N_26917,N_26590);
xnor U29494 (N_29494,N_26690,N_26863);
or U29495 (N_29495,N_26569,N_27706);
and U29496 (N_29496,N_27893,N_27936);
or U29497 (N_29497,N_27370,N_27935);
nor U29498 (N_29498,N_27095,N_27040);
or U29499 (N_29499,N_26027,N_27566);
xor U29500 (N_29500,N_26762,N_26338);
nor U29501 (N_29501,N_27077,N_27301);
nor U29502 (N_29502,N_27093,N_26436);
nor U29503 (N_29503,N_26691,N_27917);
nor U29504 (N_29504,N_26156,N_27957);
or U29505 (N_29505,N_26822,N_26597);
and U29506 (N_29506,N_27129,N_26729);
nor U29507 (N_29507,N_27286,N_26582);
nor U29508 (N_29508,N_27515,N_26513);
nand U29509 (N_29509,N_26108,N_27719);
nand U29510 (N_29510,N_27725,N_26793);
nand U29511 (N_29511,N_26805,N_26178);
and U29512 (N_29512,N_26907,N_27540);
or U29513 (N_29513,N_26937,N_27478);
nor U29514 (N_29514,N_27540,N_27140);
nor U29515 (N_29515,N_26705,N_27699);
xor U29516 (N_29516,N_27542,N_27231);
nand U29517 (N_29517,N_27662,N_26621);
nand U29518 (N_29518,N_27812,N_26686);
nand U29519 (N_29519,N_26836,N_27358);
and U29520 (N_29520,N_26791,N_27633);
or U29521 (N_29521,N_27065,N_27652);
nand U29522 (N_29522,N_27335,N_27031);
or U29523 (N_29523,N_26372,N_26325);
nand U29524 (N_29524,N_26817,N_26464);
or U29525 (N_29525,N_26964,N_27639);
and U29526 (N_29526,N_26342,N_26407);
and U29527 (N_29527,N_26237,N_26239);
or U29528 (N_29528,N_26566,N_26711);
or U29529 (N_29529,N_26903,N_27035);
nor U29530 (N_29530,N_27216,N_27194);
nand U29531 (N_29531,N_26314,N_27493);
nand U29532 (N_29532,N_26482,N_26114);
xor U29533 (N_29533,N_27828,N_27914);
xnor U29534 (N_29534,N_26123,N_26429);
xnor U29535 (N_29535,N_27862,N_27861);
nand U29536 (N_29536,N_27665,N_26627);
xnor U29537 (N_29537,N_27150,N_27832);
nor U29538 (N_29538,N_26413,N_27102);
or U29539 (N_29539,N_27341,N_26093);
or U29540 (N_29540,N_27981,N_27291);
xnor U29541 (N_29541,N_27411,N_26482);
nor U29542 (N_29542,N_27417,N_26832);
nor U29543 (N_29543,N_26390,N_27023);
nand U29544 (N_29544,N_26697,N_26910);
xor U29545 (N_29545,N_27634,N_27327);
or U29546 (N_29546,N_26353,N_26656);
and U29547 (N_29547,N_26704,N_26789);
nand U29548 (N_29548,N_26096,N_26855);
and U29549 (N_29549,N_27968,N_26176);
nor U29550 (N_29550,N_26617,N_26940);
xor U29551 (N_29551,N_27395,N_27328);
or U29552 (N_29552,N_27302,N_26906);
nand U29553 (N_29553,N_26130,N_26871);
and U29554 (N_29554,N_26191,N_26177);
nand U29555 (N_29555,N_26134,N_27815);
xor U29556 (N_29556,N_26524,N_27671);
and U29557 (N_29557,N_27053,N_27016);
or U29558 (N_29558,N_26464,N_26123);
nand U29559 (N_29559,N_26308,N_27586);
nand U29560 (N_29560,N_27403,N_26368);
or U29561 (N_29561,N_27732,N_26623);
nand U29562 (N_29562,N_27495,N_26616);
and U29563 (N_29563,N_27315,N_26285);
nor U29564 (N_29564,N_26109,N_26228);
or U29565 (N_29565,N_26558,N_27989);
nor U29566 (N_29566,N_27968,N_26408);
nor U29567 (N_29567,N_27937,N_26192);
and U29568 (N_29568,N_26553,N_27557);
and U29569 (N_29569,N_27391,N_27264);
nand U29570 (N_29570,N_27014,N_27958);
and U29571 (N_29571,N_26392,N_26268);
nand U29572 (N_29572,N_27744,N_27941);
and U29573 (N_29573,N_27371,N_27716);
or U29574 (N_29574,N_26186,N_26228);
and U29575 (N_29575,N_27168,N_27307);
xor U29576 (N_29576,N_27462,N_27759);
or U29577 (N_29577,N_27291,N_26423);
and U29578 (N_29578,N_26297,N_26972);
or U29579 (N_29579,N_27703,N_27526);
and U29580 (N_29580,N_26677,N_27470);
xnor U29581 (N_29581,N_27424,N_26688);
or U29582 (N_29582,N_26991,N_26300);
xnor U29583 (N_29583,N_26137,N_27528);
nor U29584 (N_29584,N_26212,N_26621);
or U29585 (N_29585,N_27201,N_27761);
or U29586 (N_29586,N_26923,N_27960);
xor U29587 (N_29587,N_27302,N_27783);
xnor U29588 (N_29588,N_27033,N_26117);
or U29589 (N_29589,N_26168,N_26338);
xnor U29590 (N_29590,N_26975,N_27554);
or U29591 (N_29591,N_26181,N_27465);
nand U29592 (N_29592,N_27943,N_26284);
xnor U29593 (N_29593,N_27946,N_26276);
and U29594 (N_29594,N_27969,N_26610);
nand U29595 (N_29595,N_26209,N_27726);
and U29596 (N_29596,N_26161,N_27380);
or U29597 (N_29597,N_26945,N_26644);
xor U29598 (N_29598,N_26250,N_27478);
or U29599 (N_29599,N_27184,N_26957);
and U29600 (N_29600,N_26347,N_26196);
nor U29601 (N_29601,N_26207,N_27519);
nor U29602 (N_29602,N_26816,N_26433);
nor U29603 (N_29603,N_27138,N_26270);
and U29604 (N_29604,N_27151,N_27249);
or U29605 (N_29605,N_26969,N_27798);
nand U29606 (N_29606,N_27819,N_27008);
xnor U29607 (N_29607,N_26153,N_26862);
or U29608 (N_29608,N_26418,N_26679);
nand U29609 (N_29609,N_27265,N_26344);
nor U29610 (N_29610,N_26998,N_27317);
xor U29611 (N_29611,N_26550,N_26034);
xnor U29612 (N_29612,N_27419,N_26447);
nor U29613 (N_29613,N_26739,N_26888);
or U29614 (N_29614,N_26066,N_26723);
and U29615 (N_29615,N_26133,N_27149);
nand U29616 (N_29616,N_26614,N_27204);
or U29617 (N_29617,N_26320,N_26110);
and U29618 (N_29618,N_26271,N_26950);
xor U29619 (N_29619,N_26143,N_27392);
nand U29620 (N_29620,N_27767,N_27757);
or U29621 (N_29621,N_27196,N_27071);
nor U29622 (N_29622,N_27088,N_27970);
nor U29623 (N_29623,N_26940,N_27376);
or U29624 (N_29624,N_26485,N_27118);
nand U29625 (N_29625,N_26275,N_26940);
xnor U29626 (N_29626,N_27829,N_26464);
and U29627 (N_29627,N_26768,N_26349);
nand U29628 (N_29628,N_26302,N_26667);
nand U29629 (N_29629,N_26145,N_27882);
and U29630 (N_29630,N_27828,N_27667);
or U29631 (N_29631,N_27099,N_26349);
or U29632 (N_29632,N_26254,N_27423);
xor U29633 (N_29633,N_27780,N_26244);
or U29634 (N_29634,N_26073,N_26304);
and U29635 (N_29635,N_27298,N_26218);
nor U29636 (N_29636,N_27856,N_26174);
and U29637 (N_29637,N_26819,N_27269);
xor U29638 (N_29638,N_27726,N_26315);
nand U29639 (N_29639,N_26501,N_26077);
nand U29640 (N_29640,N_27226,N_26066);
and U29641 (N_29641,N_27773,N_27469);
xnor U29642 (N_29642,N_27690,N_26216);
xnor U29643 (N_29643,N_26296,N_27043);
and U29644 (N_29644,N_26712,N_27747);
or U29645 (N_29645,N_27099,N_26886);
or U29646 (N_29646,N_27086,N_26288);
nor U29647 (N_29647,N_26032,N_27992);
xor U29648 (N_29648,N_26842,N_27922);
nor U29649 (N_29649,N_26436,N_26208);
xor U29650 (N_29650,N_27286,N_27642);
nor U29651 (N_29651,N_27201,N_26038);
nor U29652 (N_29652,N_27748,N_26477);
and U29653 (N_29653,N_26455,N_26352);
or U29654 (N_29654,N_27791,N_26754);
nand U29655 (N_29655,N_27063,N_27600);
xnor U29656 (N_29656,N_26606,N_27747);
nor U29657 (N_29657,N_26349,N_27983);
and U29658 (N_29658,N_27177,N_27499);
nand U29659 (N_29659,N_27912,N_26652);
or U29660 (N_29660,N_26927,N_27064);
nand U29661 (N_29661,N_27393,N_27823);
or U29662 (N_29662,N_27584,N_26775);
xnor U29663 (N_29663,N_26526,N_27590);
and U29664 (N_29664,N_26935,N_27940);
or U29665 (N_29665,N_27881,N_27200);
xnor U29666 (N_29666,N_27338,N_27855);
nor U29667 (N_29667,N_26802,N_26758);
nor U29668 (N_29668,N_27238,N_26672);
or U29669 (N_29669,N_26955,N_27066);
nand U29670 (N_29670,N_27904,N_26160);
nand U29671 (N_29671,N_27573,N_26850);
xnor U29672 (N_29672,N_27629,N_26334);
or U29673 (N_29673,N_27693,N_26656);
xor U29674 (N_29674,N_27001,N_26837);
xnor U29675 (N_29675,N_26034,N_27076);
xnor U29676 (N_29676,N_26317,N_27962);
nor U29677 (N_29677,N_27817,N_27702);
nand U29678 (N_29678,N_26240,N_26357);
or U29679 (N_29679,N_26945,N_26321);
and U29680 (N_29680,N_27812,N_27760);
nand U29681 (N_29681,N_26175,N_26134);
nor U29682 (N_29682,N_26367,N_27820);
nand U29683 (N_29683,N_26204,N_26741);
or U29684 (N_29684,N_27543,N_27351);
xnor U29685 (N_29685,N_26275,N_27238);
nand U29686 (N_29686,N_26357,N_27684);
or U29687 (N_29687,N_26437,N_27099);
or U29688 (N_29688,N_26115,N_26389);
xnor U29689 (N_29689,N_26235,N_27152);
nand U29690 (N_29690,N_27150,N_26878);
or U29691 (N_29691,N_26432,N_26141);
nand U29692 (N_29692,N_26766,N_26331);
or U29693 (N_29693,N_27746,N_26244);
xnor U29694 (N_29694,N_27352,N_26465);
xnor U29695 (N_29695,N_26231,N_27688);
and U29696 (N_29696,N_27548,N_26723);
nand U29697 (N_29697,N_26017,N_27701);
nand U29698 (N_29698,N_26207,N_27120);
and U29699 (N_29699,N_26508,N_27402);
nand U29700 (N_29700,N_26667,N_27775);
nor U29701 (N_29701,N_26821,N_26932);
and U29702 (N_29702,N_27604,N_27555);
nand U29703 (N_29703,N_26030,N_27957);
nor U29704 (N_29704,N_27636,N_26640);
or U29705 (N_29705,N_27915,N_26003);
xnor U29706 (N_29706,N_26513,N_27164);
nand U29707 (N_29707,N_26391,N_26466);
or U29708 (N_29708,N_26363,N_26539);
xnor U29709 (N_29709,N_26575,N_26744);
nand U29710 (N_29710,N_26648,N_27795);
nor U29711 (N_29711,N_27050,N_26770);
and U29712 (N_29712,N_27721,N_27292);
or U29713 (N_29713,N_27787,N_27606);
xnor U29714 (N_29714,N_27494,N_27515);
nor U29715 (N_29715,N_27818,N_26334);
xor U29716 (N_29716,N_26601,N_26785);
or U29717 (N_29717,N_26375,N_27442);
xor U29718 (N_29718,N_26158,N_27136);
and U29719 (N_29719,N_27203,N_26481);
and U29720 (N_29720,N_27978,N_27535);
nor U29721 (N_29721,N_27610,N_26342);
nor U29722 (N_29722,N_27987,N_26695);
xnor U29723 (N_29723,N_27291,N_26351);
nand U29724 (N_29724,N_27036,N_27022);
or U29725 (N_29725,N_26363,N_26927);
xnor U29726 (N_29726,N_27678,N_27588);
xnor U29727 (N_29727,N_27313,N_27232);
nor U29728 (N_29728,N_27425,N_26576);
nor U29729 (N_29729,N_26164,N_26013);
or U29730 (N_29730,N_27404,N_26607);
nor U29731 (N_29731,N_26461,N_27686);
or U29732 (N_29732,N_26388,N_26037);
or U29733 (N_29733,N_26390,N_26295);
or U29734 (N_29734,N_27070,N_26755);
nand U29735 (N_29735,N_26149,N_27696);
and U29736 (N_29736,N_27079,N_26659);
nand U29737 (N_29737,N_26876,N_27861);
and U29738 (N_29738,N_27817,N_27587);
nand U29739 (N_29739,N_27341,N_27871);
nand U29740 (N_29740,N_27359,N_26908);
and U29741 (N_29741,N_26935,N_26661);
or U29742 (N_29742,N_26048,N_27754);
or U29743 (N_29743,N_26856,N_27675);
or U29744 (N_29744,N_26036,N_27948);
nand U29745 (N_29745,N_26330,N_26438);
nand U29746 (N_29746,N_27006,N_26693);
nand U29747 (N_29747,N_27052,N_27481);
and U29748 (N_29748,N_27933,N_26600);
nand U29749 (N_29749,N_27252,N_27963);
xnor U29750 (N_29750,N_27767,N_26271);
and U29751 (N_29751,N_26551,N_27809);
and U29752 (N_29752,N_27641,N_27894);
and U29753 (N_29753,N_27999,N_27264);
nand U29754 (N_29754,N_27430,N_26172);
nor U29755 (N_29755,N_27001,N_27998);
or U29756 (N_29756,N_26059,N_26235);
and U29757 (N_29757,N_26057,N_27153);
nor U29758 (N_29758,N_27411,N_26119);
nand U29759 (N_29759,N_27870,N_27930);
nand U29760 (N_29760,N_26620,N_27765);
xnor U29761 (N_29761,N_27701,N_27005);
or U29762 (N_29762,N_27770,N_26404);
and U29763 (N_29763,N_27128,N_26283);
nand U29764 (N_29764,N_26117,N_27426);
or U29765 (N_29765,N_26201,N_27459);
xor U29766 (N_29766,N_26404,N_27931);
or U29767 (N_29767,N_27268,N_26417);
nor U29768 (N_29768,N_27882,N_27104);
nor U29769 (N_29769,N_27894,N_27116);
nor U29770 (N_29770,N_26210,N_26382);
nor U29771 (N_29771,N_27308,N_26989);
xor U29772 (N_29772,N_27132,N_27979);
or U29773 (N_29773,N_26466,N_27814);
and U29774 (N_29774,N_27920,N_27247);
nand U29775 (N_29775,N_27986,N_27185);
and U29776 (N_29776,N_27086,N_27967);
nor U29777 (N_29777,N_26321,N_27393);
and U29778 (N_29778,N_26477,N_27239);
nor U29779 (N_29779,N_27812,N_27719);
nor U29780 (N_29780,N_26910,N_27495);
nor U29781 (N_29781,N_26507,N_26444);
nand U29782 (N_29782,N_26132,N_26715);
or U29783 (N_29783,N_27936,N_27531);
or U29784 (N_29784,N_27251,N_26257);
or U29785 (N_29785,N_26912,N_26446);
xor U29786 (N_29786,N_26275,N_26899);
and U29787 (N_29787,N_27185,N_26136);
nand U29788 (N_29788,N_27994,N_26564);
xnor U29789 (N_29789,N_26789,N_26878);
and U29790 (N_29790,N_26048,N_26694);
and U29791 (N_29791,N_27285,N_27288);
nor U29792 (N_29792,N_26627,N_27503);
or U29793 (N_29793,N_26520,N_26832);
xnor U29794 (N_29794,N_26047,N_26392);
or U29795 (N_29795,N_27702,N_26676);
or U29796 (N_29796,N_27238,N_27014);
nand U29797 (N_29797,N_27538,N_26331);
or U29798 (N_29798,N_27456,N_26248);
nor U29799 (N_29799,N_26268,N_26225);
nor U29800 (N_29800,N_26567,N_27545);
and U29801 (N_29801,N_27547,N_27200);
or U29802 (N_29802,N_27612,N_26972);
nand U29803 (N_29803,N_26516,N_27944);
nand U29804 (N_29804,N_26683,N_26138);
nand U29805 (N_29805,N_27427,N_26924);
or U29806 (N_29806,N_26379,N_26136);
nor U29807 (N_29807,N_27012,N_26217);
nor U29808 (N_29808,N_27274,N_26223);
xnor U29809 (N_29809,N_26114,N_27979);
nor U29810 (N_29810,N_27952,N_26841);
and U29811 (N_29811,N_27615,N_27504);
nor U29812 (N_29812,N_26362,N_26174);
nor U29813 (N_29813,N_27453,N_26186);
nor U29814 (N_29814,N_27587,N_26137);
or U29815 (N_29815,N_27771,N_26655);
nor U29816 (N_29816,N_27969,N_27288);
and U29817 (N_29817,N_27127,N_27012);
or U29818 (N_29818,N_26543,N_26227);
or U29819 (N_29819,N_26114,N_27117);
nand U29820 (N_29820,N_26064,N_26483);
and U29821 (N_29821,N_26234,N_27255);
nor U29822 (N_29822,N_26295,N_26516);
xor U29823 (N_29823,N_27297,N_26311);
nor U29824 (N_29824,N_27401,N_26466);
xor U29825 (N_29825,N_26611,N_27163);
nand U29826 (N_29826,N_27797,N_27070);
nor U29827 (N_29827,N_26452,N_26311);
nand U29828 (N_29828,N_27135,N_27795);
nor U29829 (N_29829,N_26189,N_27731);
nand U29830 (N_29830,N_27334,N_27624);
and U29831 (N_29831,N_26749,N_27090);
xnor U29832 (N_29832,N_27698,N_26082);
nor U29833 (N_29833,N_26015,N_27240);
nor U29834 (N_29834,N_27428,N_26863);
or U29835 (N_29835,N_27612,N_26880);
nand U29836 (N_29836,N_27966,N_26326);
nor U29837 (N_29837,N_27708,N_27767);
xnor U29838 (N_29838,N_27558,N_27786);
nor U29839 (N_29839,N_26288,N_27631);
nand U29840 (N_29840,N_27956,N_27763);
nand U29841 (N_29841,N_27254,N_26967);
nand U29842 (N_29842,N_26349,N_26753);
or U29843 (N_29843,N_27472,N_26639);
or U29844 (N_29844,N_26449,N_26739);
nand U29845 (N_29845,N_26684,N_26974);
nand U29846 (N_29846,N_27259,N_26975);
nor U29847 (N_29847,N_26373,N_27495);
xor U29848 (N_29848,N_26963,N_26815);
or U29849 (N_29849,N_26719,N_26110);
or U29850 (N_29850,N_26483,N_26364);
or U29851 (N_29851,N_26171,N_26913);
or U29852 (N_29852,N_27617,N_26792);
and U29853 (N_29853,N_27265,N_27385);
nor U29854 (N_29854,N_26641,N_26363);
or U29855 (N_29855,N_27829,N_27084);
xor U29856 (N_29856,N_27734,N_27860);
and U29857 (N_29857,N_26850,N_26577);
and U29858 (N_29858,N_27971,N_27106);
and U29859 (N_29859,N_26598,N_26837);
nand U29860 (N_29860,N_26925,N_27916);
xnor U29861 (N_29861,N_27435,N_27922);
nor U29862 (N_29862,N_27309,N_26197);
and U29863 (N_29863,N_27712,N_27266);
or U29864 (N_29864,N_27301,N_27559);
and U29865 (N_29865,N_27474,N_26251);
nor U29866 (N_29866,N_27865,N_27086);
or U29867 (N_29867,N_26773,N_27511);
nor U29868 (N_29868,N_26893,N_27117);
nand U29869 (N_29869,N_26289,N_26713);
or U29870 (N_29870,N_27594,N_27400);
nor U29871 (N_29871,N_26058,N_26665);
and U29872 (N_29872,N_26869,N_26267);
and U29873 (N_29873,N_26069,N_27988);
xnor U29874 (N_29874,N_26375,N_27732);
nor U29875 (N_29875,N_26899,N_26357);
nand U29876 (N_29876,N_27261,N_27082);
nor U29877 (N_29877,N_27106,N_27959);
nand U29878 (N_29878,N_27010,N_26959);
or U29879 (N_29879,N_27816,N_26224);
nor U29880 (N_29880,N_27017,N_26152);
or U29881 (N_29881,N_27853,N_27882);
xnor U29882 (N_29882,N_27992,N_26986);
xor U29883 (N_29883,N_27900,N_27755);
and U29884 (N_29884,N_27549,N_27004);
or U29885 (N_29885,N_26679,N_26471);
and U29886 (N_29886,N_26810,N_27953);
and U29887 (N_29887,N_27806,N_26028);
xnor U29888 (N_29888,N_26085,N_26893);
nand U29889 (N_29889,N_26108,N_26474);
and U29890 (N_29890,N_27972,N_27903);
xor U29891 (N_29891,N_26212,N_27014);
nor U29892 (N_29892,N_27441,N_26274);
nor U29893 (N_29893,N_26646,N_26747);
and U29894 (N_29894,N_27105,N_26393);
or U29895 (N_29895,N_26935,N_26768);
or U29896 (N_29896,N_26187,N_26443);
nor U29897 (N_29897,N_27922,N_26966);
and U29898 (N_29898,N_27436,N_26949);
nand U29899 (N_29899,N_27683,N_26555);
and U29900 (N_29900,N_26490,N_27976);
xor U29901 (N_29901,N_27619,N_26434);
nand U29902 (N_29902,N_27231,N_26241);
and U29903 (N_29903,N_26642,N_27647);
nor U29904 (N_29904,N_26881,N_27432);
nand U29905 (N_29905,N_26669,N_26939);
nand U29906 (N_29906,N_26699,N_26501);
and U29907 (N_29907,N_27900,N_26719);
or U29908 (N_29908,N_27044,N_27782);
nand U29909 (N_29909,N_27342,N_26614);
nor U29910 (N_29910,N_27916,N_27358);
xor U29911 (N_29911,N_27150,N_26779);
nand U29912 (N_29912,N_27097,N_27568);
xnor U29913 (N_29913,N_27402,N_26049);
nor U29914 (N_29914,N_27505,N_27503);
nor U29915 (N_29915,N_27923,N_27382);
xnor U29916 (N_29916,N_27986,N_27115);
or U29917 (N_29917,N_27485,N_26590);
xor U29918 (N_29918,N_27236,N_27039);
nand U29919 (N_29919,N_27215,N_26702);
or U29920 (N_29920,N_26637,N_27023);
or U29921 (N_29921,N_26571,N_26975);
and U29922 (N_29922,N_26962,N_26171);
or U29923 (N_29923,N_26345,N_26564);
or U29924 (N_29924,N_26979,N_27719);
and U29925 (N_29925,N_27719,N_27445);
and U29926 (N_29926,N_26806,N_26817);
nand U29927 (N_29927,N_27328,N_26743);
nor U29928 (N_29928,N_26248,N_26297);
or U29929 (N_29929,N_27298,N_26690);
nand U29930 (N_29930,N_27749,N_26088);
xor U29931 (N_29931,N_26407,N_26263);
nor U29932 (N_29932,N_27302,N_27368);
nand U29933 (N_29933,N_27132,N_27690);
xor U29934 (N_29934,N_26451,N_27389);
nand U29935 (N_29935,N_27799,N_27174);
nand U29936 (N_29936,N_27063,N_26818);
nand U29937 (N_29937,N_26341,N_26106);
nor U29938 (N_29938,N_26449,N_26488);
nand U29939 (N_29939,N_26019,N_26568);
and U29940 (N_29940,N_27585,N_27983);
and U29941 (N_29941,N_26805,N_27044);
and U29942 (N_29942,N_26513,N_27471);
nor U29943 (N_29943,N_26156,N_27956);
and U29944 (N_29944,N_27222,N_27177);
and U29945 (N_29945,N_26476,N_26993);
and U29946 (N_29946,N_27772,N_26981);
xnor U29947 (N_29947,N_26125,N_27956);
nand U29948 (N_29948,N_26035,N_27627);
nor U29949 (N_29949,N_27131,N_27468);
or U29950 (N_29950,N_27367,N_27552);
and U29951 (N_29951,N_27760,N_27764);
nand U29952 (N_29952,N_27614,N_27484);
or U29953 (N_29953,N_27754,N_26039);
and U29954 (N_29954,N_27560,N_27640);
and U29955 (N_29955,N_27471,N_27763);
and U29956 (N_29956,N_27857,N_27198);
nand U29957 (N_29957,N_27851,N_26361);
and U29958 (N_29958,N_26920,N_27349);
xnor U29959 (N_29959,N_26244,N_27125);
nand U29960 (N_29960,N_27404,N_27069);
nand U29961 (N_29961,N_26816,N_26836);
and U29962 (N_29962,N_26915,N_26780);
and U29963 (N_29963,N_26613,N_26688);
and U29964 (N_29964,N_26636,N_27856);
or U29965 (N_29965,N_27227,N_26528);
nand U29966 (N_29966,N_27271,N_26304);
nand U29967 (N_29967,N_26725,N_27460);
nor U29968 (N_29968,N_27913,N_27005);
xnor U29969 (N_29969,N_26520,N_26943);
nand U29970 (N_29970,N_27743,N_27779);
nor U29971 (N_29971,N_26339,N_26699);
or U29972 (N_29972,N_27513,N_27282);
xor U29973 (N_29973,N_27919,N_27975);
or U29974 (N_29974,N_27689,N_27968);
and U29975 (N_29975,N_27206,N_26071);
or U29976 (N_29976,N_26342,N_26722);
and U29977 (N_29977,N_26649,N_27312);
nand U29978 (N_29978,N_27855,N_27120);
and U29979 (N_29979,N_26303,N_26404);
nand U29980 (N_29980,N_26166,N_26130);
or U29981 (N_29981,N_26553,N_26696);
or U29982 (N_29982,N_26783,N_26493);
and U29983 (N_29983,N_26161,N_26075);
and U29984 (N_29984,N_26368,N_26262);
nor U29985 (N_29985,N_26923,N_26701);
and U29986 (N_29986,N_27581,N_26085);
or U29987 (N_29987,N_26660,N_26592);
nor U29988 (N_29988,N_27398,N_26329);
or U29989 (N_29989,N_27490,N_27391);
or U29990 (N_29990,N_26091,N_27265);
and U29991 (N_29991,N_26852,N_27769);
xnor U29992 (N_29992,N_26886,N_27396);
nand U29993 (N_29993,N_27999,N_27652);
nor U29994 (N_29994,N_26711,N_27055);
or U29995 (N_29995,N_27881,N_26500);
xnor U29996 (N_29996,N_26013,N_27116);
nand U29997 (N_29997,N_26310,N_27156);
xor U29998 (N_29998,N_27427,N_27822);
and U29999 (N_29999,N_26263,N_26616);
nand UO_0 (O_0,N_29487,N_29692);
or UO_1 (O_1,N_29925,N_29066);
nand UO_2 (O_2,N_29212,N_28470);
nand UO_3 (O_3,N_28443,N_29935);
xnor UO_4 (O_4,N_28397,N_29188);
nor UO_5 (O_5,N_29155,N_28826);
xor UO_6 (O_6,N_28413,N_29962);
xor UO_7 (O_7,N_29025,N_29742);
or UO_8 (O_8,N_29132,N_28921);
xnor UO_9 (O_9,N_28555,N_29289);
nor UO_10 (O_10,N_28900,N_29672);
xnor UO_11 (O_11,N_29712,N_28324);
nor UO_12 (O_12,N_28910,N_28014);
or UO_13 (O_13,N_28034,N_28290);
xnor UO_14 (O_14,N_28301,N_29717);
nor UO_15 (O_15,N_29825,N_28070);
and UO_16 (O_16,N_28552,N_29418);
and UO_17 (O_17,N_29785,N_29442);
or UO_18 (O_18,N_29529,N_29363);
xor UO_19 (O_19,N_29397,N_28458);
nand UO_20 (O_20,N_28556,N_29946);
and UO_21 (O_21,N_28386,N_28598);
or UO_22 (O_22,N_28948,N_29807);
or UO_23 (O_23,N_28908,N_28305);
and UO_24 (O_24,N_28756,N_29572);
nor UO_25 (O_25,N_28154,N_29608);
or UO_26 (O_26,N_28489,N_28614);
or UO_27 (O_27,N_29133,N_28090);
nor UO_28 (O_28,N_29857,N_29562);
nand UO_29 (O_29,N_28930,N_28449);
nand UO_30 (O_30,N_28485,N_28126);
nor UO_31 (O_31,N_28027,N_28459);
or UO_32 (O_32,N_28078,N_28742);
xor UO_33 (O_33,N_29837,N_28786);
nand UO_34 (O_34,N_28804,N_28822);
and UO_35 (O_35,N_28794,N_28717);
nor UO_36 (O_36,N_28279,N_29086);
or UO_37 (O_37,N_29854,N_29129);
nand UO_38 (O_38,N_29370,N_29765);
or UO_39 (O_39,N_29969,N_29364);
xnor UO_40 (O_40,N_29567,N_28241);
xnor UO_41 (O_41,N_29990,N_29172);
nor UO_42 (O_42,N_29213,N_28228);
xnor UO_43 (O_43,N_28438,N_29709);
or UO_44 (O_44,N_28807,N_28768);
nor UO_45 (O_45,N_29997,N_28419);
nor UO_46 (O_46,N_28145,N_29535);
or UO_47 (O_47,N_29094,N_28548);
xor UO_48 (O_48,N_29392,N_29910);
xor UO_49 (O_49,N_28295,N_29298);
nor UO_50 (O_50,N_28068,N_29210);
nor UO_51 (O_51,N_29582,N_28731);
nand UO_52 (O_52,N_28372,N_29506);
or UO_53 (O_53,N_29277,N_29992);
nor UO_54 (O_54,N_28551,N_29465);
or UO_55 (O_55,N_29773,N_29069);
nand UO_56 (O_56,N_29233,N_28170);
and UO_57 (O_57,N_28935,N_28480);
and UO_58 (O_58,N_29106,N_29116);
nand UO_59 (O_59,N_29326,N_29446);
nor UO_60 (O_60,N_28671,N_28907);
xor UO_61 (O_61,N_28106,N_29589);
nor UO_62 (O_62,N_28370,N_28361);
or UO_63 (O_63,N_29524,N_28718);
nand UO_64 (O_64,N_28680,N_28554);
nand UO_65 (O_65,N_28801,N_29552);
xor UO_66 (O_66,N_28193,N_28567);
or UO_67 (O_67,N_28882,N_29406);
xnor UO_68 (O_68,N_28783,N_28189);
nand UO_69 (O_69,N_28769,N_28772);
and UO_70 (O_70,N_28004,N_29369);
and UO_71 (O_71,N_29337,N_28841);
or UO_72 (O_72,N_28472,N_28119);
and UO_73 (O_73,N_29357,N_29647);
and UO_74 (O_74,N_28626,N_29372);
xnor UO_75 (O_75,N_28648,N_28481);
nor UO_76 (O_76,N_28562,N_28499);
nor UO_77 (O_77,N_29481,N_29901);
nor UO_78 (O_78,N_29830,N_29947);
or UO_79 (O_79,N_28906,N_29761);
nor UO_80 (O_80,N_29955,N_29559);
nor UO_81 (O_81,N_28961,N_29806);
nand UO_82 (O_82,N_29814,N_29686);
nand UO_83 (O_83,N_29045,N_29058);
nand UO_84 (O_84,N_28583,N_28590);
nand UO_85 (O_85,N_28162,N_28547);
xnor UO_86 (O_86,N_28057,N_29131);
or UO_87 (O_87,N_28748,N_28203);
nand UO_88 (O_88,N_29217,N_29417);
or UO_89 (O_89,N_28868,N_29952);
and UO_90 (O_90,N_29705,N_29262);
nor UO_91 (O_91,N_29751,N_28630);
or UO_92 (O_92,N_28277,N_29977);
nand UO_93 (O_93,N_29503,N_28858);
or UO_94 (O_94,N_28083,N_28166);
nor UO_95 (O_95,N_29564,N_28436);
and UO_96 (O_96,N_28694,N_29803);
nand UO_97 (O_97,N_28257,N_28011);
nand UO_98 (O_98,N_29579,N_28650);
and UO_99 (O_99,N_28433,N_29120);
nor UO_100 (O_100,N_28417,N_29226);
nand UO_101 (O_101,N_29024,N_28118);
xnor UO_102 (O_102,N_28254,N_29743);
and UO_103 (O_103,N_29159,N_29462);
nor UO_104 (O_104,N_28441,N_28950);
and UO_105 (O_105,N_29909,N_28710);
or UO_106 (O_106,N_29335,N_28494);
xnor UO_107 (O_107,N_28379,N_29605);
xnor UO_108 (O_108,N_28559,N_29278);
nor UO_109 (O_109,N_28952,N_29956);
and UO_110 (O_110,N_29143,N_28720);
or UO_111 (O_111,N_29333,N_28461);
or UO_112 (O_112,N_28116,N_28519);
or UO_113 (O_113,N_28751,N_29454);
nand UO_114 (O_114,N_29312,N_29078);
nor UO_115 (O_115,N_28408,N_29818);
nand UO_116 (O_116,N_29889,N_28052);
nor UO_117 (O_117,N_28577,N_29411);
xor UO_118 (O_118,N_28275,N_29254);
xor UO_119 (O_119,N_28043,N_28121);
nand UO_120 (O_120,N_29896,N_28545);
nor UO_121 (O_121,N_29306,N_29036);
nand UO_122 (O_122,N_28692,N_29911);
nand UO_123 (O_123,N_29198,N_29514);
xnor UO_124 (O_124,N_29016,N_28050);
or UO_125 (O_125,N_29474,N_28456);
nand UO_126 (O_126,N_28219,N_29802);
nand UO_127 (O_127,N_28155,N_29735);
nand UO_128 (O_128,N_28133,N_29520);
and UO_129 (O_129,N_28965,N_28482);
and UO_130 (O_130,N_29891,N_28610);
nor UO_131 (O_131,N_29434,N_28213);
nor UO_132 (O_132,N_29083,N_28007);
nand UO_133 (O_133,N_28670,N_28631);
nand UO_134 (O_134,N_29380,N_29917);
nor UO_135 (O_135,N_28374,N_28920);
or UO_136 (O_136,N_28281,N_28919);
xnor UO_137 (O_137,N_28345,N_28176);
nor UO_138 (O_138,N_29667,N_29122);
xnor UO_139 (O_139,N_29936,N_28503);
nand UO_140 (O_140,N_28396,N_29142);
nor UO_141 (O_141,N_29156,N_29511);
and UO_142 (O_142,N_29752,N_29930);
nor UO_143 (O_143,N_29195,N_28637);
or UO_144 (O_144,N_28899,N_28539);
nand UO_145 (O_145,N_29327,N_28869);
nor UO_146 (O_146,N_29076,N_28757);
nand UO_147 (O_147,N_28047,N_28025);
xnor UO_148 (O_148,N_28873,N_28411);
xnor UO_149 (O_149,N_29682,N_28838);
and UO_150 (O_150,N_28046,N_29883);
nor UO_151 (O_151,N_28513,N_29714);
nand UO_152 (O_152,N_28328,N_29477);
nand UO_153 (O_153,N_28561,N_28044);
or UO_154 (O_154,N_29102,N_28446);
or UO_155 (O_155,N_29887,N_28808);
and UO_156 (O_156,N_28495,N_28709);
or UO_157 (O_157,N_28420,N_28058);
nor UO_158 (O_158,N_29111,N_28914);
xor UO_159 (O_159,N_29443,N_29581);
xnor UO_160 (O_160,N_29680,N_28881);
or UO_161 (O_161,N_29407,N_28369);
nand UO_162 (O_162,N_29158,N_29671);
nor UO_163 (O_163,N_28988,N_29430);
nor UO_164 (O_164,N_29504,N_28278);
nor UO_165 (O_165,N_29878,N_29627);
and UO_166 (O_166,N_28165,N_29551);
nor UO_167 (O_167,N_28151,N_29770);
nand UO_168 (O_168,N_29147,N_29290);
and UO_169 (O_169,N_28476,N_28836);
and UO_170 (O_170,N_28287,N_29192);
nand UO_171 (O_171,N_28969,N_28973);
or UO_172 (O_172,N_28500,N_28898);
and UO_173 (O_173,N_29101,N_29252);
nor UO_174 (O_174,N_29341,N_29696);
and UO_175 (O_175,N_28553,N_28733);
or UO_176 (O_176,N_29745,N_29161);
xnor UO_177 (O_177,N_28284,N_29276);
nor UO_178 (O_178,N_28734,N_29833);
and UO_179 (O_179,N_29868,N_29852);
xnor UO_180 (O_180,N_29500,N_29820);
and UO_181 (O_181,N_28866,N_28477);
nor UO_182 (O_182,N_29483,N_29890);
and UO_183 (O_183,N_29166,N_29280);
nor UO_184 (O_184,N_28787,N_29618);
nand UO_185 (O_185,N_28421,N_28242);
xnor UO_186 (O_186,N_28887,N_28037);
nand UO_187 (O_187,N_28209,N_29377);
and UO_188 (O_188,N_28951,N_29261);
nor UO_189 (O_189,N_28222,N_29923);
nor UO_190 (O_190,N_28885,N_29757);
xnor UO_191 (O_191,N_28778,N_29173);
nor UO_192 (O_192,N_29000,N_29321);
or UO_193 (O_193,N_28888,N_29223);
or UO_194 (O_194,N_29248,N_28304);
or UO_195 (O_195,N_29848,N_28686);
xor UO_196 (O_196,N_28529,N_29685);
nor UO_197 (O_197,N_29112,N_29530);
nand UO_198 (O_198,N_29030,N_28507);
and UO_199 (O_199,N_29281,N_29292);
and UO_200 (O_200,N_28713,N_29642);
nand UO_201 (O_201,N_28375,N_29401);
and UO_202 (O_202,N_28855,N_28462);
and UO_203 (O_203,N_28272,N_28828);
and UO_204 (O_204,N_28049,N_29716);
and UO_205 (O_205,N_28829,N_28716);
and UO_206 (O_206,N_28352,N_28218);
or UO_207 (O_207,N_29623,N_29084);
and UO_208 (O_208,N_29697,N_28549);
nand UO_209 (O_209,N_28161,N_29836);
xor UO_210 (O_210,N_29580,N_29983);
nor UO_211 (O_211,N_28776,N_29609);
nor UO_212 (O_212,N_28138,N_29532);
or UO_213 (O_213,N_29275,N_28256);
or UO_214 (O_214,N_29272,N_28466);
nor UO_215 (O_215,N_28845,N_28200);
nor UO_216 (O_216,N_29221,N_28879);
nor UO_217 (O_217,N_29436,N_28152);
xnor UO_218 (O_218,N_29325,N_29468);
nor UO_219 (O_219,N_28764,N_28340);
xor UO_220 (O_220,N_28187,N_28619);
nand UO_221 (O_221,N_28488,N_29853);
nor UO_222 (O_222,N_28991,N_29387);
and UO_223 (O_223,N_29812,N_29362);
nand UO_224 (O_224,N_28010,N_29264);
xor UO_225 (O_225,N_28464,N_29413);
xor UO_226 (O_226,N_29209,N_29545);
and UO_227 (O_227,N_29404,N_29649);
nand UO_228 (O_228,N_28075,N_28115);
nand UO_229 (O_229,N_29867,N_28698);
nand UO_230 (O_230,N_29549,N_29031);
nor UO_231 (O_231,N_28915,N_29247);
nand UO_232 (O_232,N_28546,N_28707);
nand UO_233 (O_233,N_29469,N_28181);
nor UO_234 (O_234,N_28348,N_28163);
and UO_235 (O_235,N_29087,N_29653);
nor UO_236 (O_236,N_28026,N_28597);
or UO_237 (O_237,N_28678,N_29561);
xnor UO_238 (O_238,N_28414,N_29110);
and UO_239 (O_239,N_29660,N_28981);
xor UO_240 (O_240,N_29978,N_28179);
and UO_241 (O_241,N_29573,N_29073);
nor UO_242 (O_242,N_28825,N_28358);
or UO_243 (O_243,N_29228,N_28527);
and UO_244 (O_244,N_29669,N_29427);
and UO_245 (O_245,N_29144,N_28029);
or UO_246 (O_246,N_29656,N_29805);
and UO_247 (O_247,N_28629,N_29698);
nand UO_248 (O_248,N_28387,N_28434);
or UO_249 (O_249,N_28987,N_29738);
xor UO_250 (O_250,N_28585,N_28288);
nor UO_251 (O_251,N_29432,N_28066);
nor UO_252 (O_252,N_28308,N_28038);
xnor UO_253 (O_253,N_28782,N_28450);
and UO_254 (O_254,N_29493,N_29323);
and UO_255 (O_255,N_28839,N_28097);
nor UO_256 (O_256,N_28255,N_28112);
or UO_257 (O_257,N_28190,N_29934);
xnor UO_258 (O_258,N_29315,N_28139);
and UO_259 (O_259,N_28890,N_28602);
nand UO_260 (O_260,N_29300,N_29255);
nor UO_261 (O_261,N_28316,N_28262);
nor UO_262 (O_262,N_28440,N_28820);
nor UO_263 (O_263,N_28798,N_28940);
or UO_264 (O_264,N_28220,N_29117);
nand UO_265 (O_265,N_29350,N_29967);
and UO_266 (O_266,N_28834,N_29661);
and UO_267 (O_267,N_29190,N_29360);
or UO_268 (O_268,N_29488,N_28715);
nand UO_269 (O_269,N_29473,N_29140);
nand UO_270 (O_270,N_28221,N_29203);
and UO_271 (O_271,N_28964,N_29844);
nand UO_272 (O_272,N_29177,N_29965);
nor UO_273 (O_273,N_29668,N_29346);
and UO_274 (O_274,N_28140,N_28701);
or UO_275 (O_275,N_28966,N_29391);
xor UO_276 (O_276,N_29633,N_28410);
nand UO_277 (O_277,N_28122,N_28342);
nand UO_278 (O_278,N_29870,N_28889);
nand UO_279 (O_279,N_28060,N_29655);
or UO_280 (O_280,N_29639,N_29124);
and UO_281 (O_281,N_28194,N_28206);
and UO_282 (O_282,N_29594,N_28663);
nor UO_283 (O_283,N_28191,N_29885);
xnor UO_284 (O_284,N_29267,N_28978);
nor UO_285 (O_285,N_29314,N_28045);
nand UO_286 (O_286,N_28453,N_29957);
and UO_287 (O_287,N_29939,N_28917);
nor UO_288 (O_288,N_28697,N_28755);
nor UO_289 (O_289,N_28666,N_29246);
or UO_290 (O_290,N_28309,N_28282);
and UO_291 (O_291,N_29318,N_28473);
nor UO_292 (O_292,N_29239,N_28803);
nand UO_293 (O_293,N_28484,N_29585);
or UO_294 (O_294,N_28289,N_29577);
or UO_295 (O_295,N_29684,N_29271);
xnor UO_296 (O_296,N_29096,N_28674);
xnor UO_297 (O_297,N_29090,N_29948);
nand UO_298 (O_298,N_29658,N_28447);
or UO_299 (O_299,N_28028,N_28968);
nor UO_300 (O_300,N_28863,N_28550);
nor UO_301 (O_301,N_28124,N_29793);
nand UO_302 (O_302,N_28524,N_29553);
nand UO_303 (O_303,N_29951,N_29253);
and UO_304 (O_304,N_29393,N_29722);
xnor UO_305 (O_305,N_28265,N_29643);
nor UO_306 (O_306,N_29537,N_28336);
and UO_307 (O_307,N_29037,N_29527);
nor UO_308 (O_308,N_29376,N_29541);
and UO_309 (O_309,N_29826,N_29905);
and UO_310 (O_310,N_28051,N_29606);
or UO_311 (O_311,N_29512,N_28313);
nand UO_312 (O_312,N_28819,N_29448);
nand UO_313 (O_313,N_29548,N_29630);
nand UO_314 (O_314,N_28468,N_29006);
nand UO_315 (O_315,N_29074,N_28738);
xor UO_316 (O_316,N_29800,N_28832);
xnor UO_317 (O_317,N_29089,N_29165);
nor UO_318 (O_318,N_28248,N_28497);
xor UO_319 (O_319,N_29463,N_28022);
nor UO_320 (O_320,N_29498,N_28048);
or UO_321 (O_321,N_29183,N_29439);
xnor UO_322 (O_322,N_29624,N_29470);
and UO_323 (O_323,N_29798,N_28544);
xor UO_324 (O_324,N_28886,N_28791);
or UO_325 (O_325,N_29079,N_28283);
and UO_326 (O_326,N_29915,N_28185);
and UO_327 (O_327,N_28691,N_29508);
xor UO_328 (O_328,N_28019,N_29359);
and UO_329 (O_329,N_28065,N_29534);
xnor UO_330 (O_330,N_29813,N_28056);
nand UO_331 (O_331,N_28005,N_29931);
nor UO_332 (O_332,N_28003,N_29659);
and UO_333 (O_333,N_29790,N_29590);
and UO_334 (O_334,N_28745,N_28076);
or UO_335 (O_335,N_28537,N_29003);
nand UO_336 (O_336,N_28439,N_28905);
nor UO_337 (O_337,N_28393,N_28036);
xnor UO_338 (O_338,N_28658,N_29943);
or UO_339 (O_339,N_29816,N_28758);
nand UO_340 (O_340,N_28020,N_29544);
xor UO_341 (O_341,N_28327,N_28430);
or UO_342 (O_342,N_28231,N_29689);
and UO_343 (O_343,N_28586,N_28415);
or UO_344 (O_344,N_29789,N_29795);
nor UO_345 (O_345,N_28923,N_29232);
and UO_346 (O_346,N_28175,N_28291);
nand UO_347 (O_347,N_29693,N_29386);
or UO_348 (O_348,N_29240,N_29441);
nor UO_349 (O_349,N_29491,N_29942);
nor UO_350 (O_350,N_28243,N_29797);
nor UO_351 (O_351,N_29744,N_28508);
nor UO_352 (O_352,N_29061,N_29288);
or UO_353 (O_353,N_28897,N_29054);
or UO_354 (O_354,N_28662,N_28645);
and UO_355 (O_355,N_28759,N_28334);
xor UO_356 (O_356,N_28867,N_28303);
or UO_357 (O_357,N_29208,N_29274);
or UO_358 (O_358,N_28469,N_29841);
nor UO_359 (O_359,N_29851,N_29708);
and UO_360 (O_360,N_28672,N_29991);
nor UO_361 (O_361,N_29995,N_28814);
nor UO_362 (O_362,N_28687,N_28633);
nand UO_363 (O_363,N_29204,N_29625);
and UO_364 (O_364,N_29613,N_28850);
or UO_365 (O_365,N_28298,N_28041);
nand UO_366 (O_366,N_28895,N_29657);
nand UO_367 (O_367,N_28471,N_29619);
and UO_368 (O_368,N_29945,N_29381);
and UO_369 (O_369,N_29879,N_29695);
and UO_370 (O_370,N_28706,N_28398);
nand UO_371 (O_371,N_28103,N_29731);
or UO_372 (O_372,N_28605,N_29629);
nor UO_373 (O_373,N_29405,N_29718);
xor UO_374 (O_374,N_29041,N_28979);
and UO_375 (O_375,N_28296,N_29361);
and UO_376 (O_376,N_28937,N_29048);
or UO_377 (O_377,N_29847,N_28566);
nand UO_378 (O_378,N_28371,N_28958);
and UO_379 (O_379,N_29607,N_29842);
nor UO_380 (O_380,N_28800,N_29382);
or UO_381 (O_381,N_28205,N_29869);
and UO_382 (O_382,N_28074,N_28726);
and UO_383 (O_383,N_29196,N_29243);
nand UO_384 (O_384,N_29634,N_28306);
and UO_385 (O_385,N_29269,N_28012);
nor UO_386 (O_386,N_29666,N_28330);
xor UO_387 (O_387,N_28641,N_29876);
nand UO_388 (O_388,N_29701,N_29485);
xor UO_389 (O_389,N_29163,N_29395);
xor UO_390 (O_390,N_28040,N_28183);
and UO_391 (O_391,N_29916,N_28712);
nor UO_392 (O_392,N_29525,N_28942);
nor UO_393 (O_393,N_28840,N_28129);
and UO_394 (O_394,N_29308,N_28916);
nor UO_395 (O_395,N_29721,N_28541);
nor UO_396 (O_396,N_28315,N_29502);
xor UO_397 (O_397,N_28388,N_29164);
nand UO_398 (O_398,N_28267,N_29556);
nor UO_399 (O_399,N_29538,N_28523);
nor UO_400 (O_400,N_29831,N_28854);
nor UO_401 (O_401,N_29072,N_29961);
or UO_402 (O_402,N_28999,N_29332);
and UO_403 (O_403,N_29644,N_29622);
or UO_404 (O_404,N_29149,N_28409);
or UO_405 (O_405,N_28578,N_28232);
nand UO_406 (O_406,N_29145,N_28506);
nor UO_407 (O_407,N_29740,N_28269);
nand UO_408 (O_408,N_29871,N_29023);
nor UO_409 (O_409,N_28173,N_29415);
nor UO_410 (O_410,N_28927,N_29933);
nor UO_411 (O_411,N_29974,N_28568);
nor UO_412 (O_412,N_29645,N_29741);
xnor UO_413 (O_413,N_28842,N_28355);
and UO_414 (O_414,N_28399,N_28286);
nand UO_415 (O_415,N_28198,N_28487);
nor UO_416 (O_416,N_29047,N_29652);
and UO_417 (O_417,N_28130,N_28271);
or UO_418 (O_418,N_28613,N_28528);
and UO_419 (O_419,N_29777,N_29593);
xor UO_420 (O_420,N_28618,N_29595);
nor UO_421 (O_421,N_28735,N_28268);
nand UO_422 (O_422,N_28864,N_28107);
nor UO_423 (O_423,N_28402,N_29013);
xor UO_424 (O_424,N_28079,N_29467);
and UO_425 (O_425,N_29225,N_29231);
xor UO_426 (O_426,N_28463,N_28403);
and UO_427 (O_427,N_29151,N_29409);
nand UO_428 (O_428,N_28114,N_28394);
or UO_429 (O_429,N_29042,N_28857);
or UO_430 (O_430,N_28760,N_29766);
nand UO_431 (O_431,N_29104,N_29884);
nor UO_432 (O_432,N_28347,N_29328);
or UO_433 (O_433,N_29452,N_28069);
nand UO_434 (O_434,N_28490,N_28793);
or UO_435 (O_435,N_28238,N_28512);
nor UO_436 (O_436,N_29985,N_28244);
nor UO_437 (O_437,N_29109,N_29963);
or UO_438 (O_438,N_28592,N_29356);
nand UO_439 (O_439,N_29734,N_29260);
and UO_440 (O_440,N_28390,N_29338);
nor UO_441 (O_441,N_29707,N_28276);
or UO_442 (O_442,N_28703,N_29416);
nor UO_443 (O_443,N_28913,N_29703);
nor UO_444 (O_444,N_28928,N_29348);
and UO_445 (O_445,N_29250,N_29170);
nand UO_446 (O_446,N_29235,N_28784);
nor UO_447 (O_447,N_29732,N_28016);
and UO_448 (O_448,N_28249,N_28579);
nand UO_449 (O_449,N_29293,N_28606);
or UO_450 (O_450,N_29118,N_28178);
or UO_451 (O_451,N_29526,N_28156);
nor UO_452 (O_452,N_28071,N_28573);
or UO_453 (O_453,N_29566,N_28591);
nand UO_454 (O_454,N_28149,N_29829);
xnor UO_455 (O_455,N_28460,N_28360);
or UO_456 (O_456,N_28147,N_29460);
and UO_457 (O_457,N_28406,N_28581);
xor UO_458 (O_458,N_29039,N_28233);
and UO_459 (O_459,N_28227,N_29720);
and UO_460 (O_460,N_29057,N_29291);
nand UO_461 (O_461,N_29959,N_29762);
nand UO_462 (O_462,N_28754,N_28125);
nand UO_463 (O_463,N_28975,N_29154);
nor UO_464 (O_464,N_28013,N_29258);
or UO_465 (O_465,N_28113,N_28977);
nor UO_466 (O_466,N_29984,N_28024);
nor UO_467 (O_467,N_28947,N_28385);
xnor UO_468 (O_468,N_29082,N_29536);
nor UO_469 (O_469,N_29004,N_28363);
or UO_470 (O_470,N_29126,N_28261);
nand UO_471 (O_471,N_28167,N_28422);
and UO_472 (O_472,N_28426,N_28911);
xnor UO_473 (O_473,N_29850,N_29651);
nor UO_474 (O_474,N_29444,N_29388);
and UO_475 (O_475,N_29786,N_28063);
xnor UO_476 (O_476,N_28683,N_28682);
xor UO_477 (O_477,N_28376,N_29636);
xnor UO_478 (O_478,N_28412,N_29385);
and UO_479 (O_479,N_29543,N_28252);
xnor UO_480 (O_480,N_29309,N_28096);
nor UO_481 (O_481,N_28356,N_28962);
nand UO_482 (O_482,N_28753,N_28377);
nor UO_483 (O_483,N_29174,N_29772);
or UO_484 (O_484,N_28938,N_28770);
and UO_485 (O_485,N_28510,N_28699);
xnor UO_486 (O_486,N_29700,N_28815);
xnor UO_487 (O_487,N_29725,N_28643);
and UO_488 (O_488,N_29973,N_28883);
nor UO_489 (O_489,N_29914,N_28810);
and UO_490 (O_490,N_29032,N_29968);
or UO_491 (O_491,N_28540,N_28143);
nand UO_492 (O_492,N_28797,N_28542);
xor UO_493 (O_493,N_29085,N_28773);
nor UO_494 (O_494,N_29342,N_29496);
xnor UO_495 (O_495,N_28117,N_28903);
nand UO_496 (O_496,N_28516,N_28625);
nand UO_497 (O_497,N_28104,N_29139);
and UO_498 (O_498,N_28195,N_29399);
or UO_499 (O_499,N_28137,N_29938);
and UO_500 (O_500,N_28474,N_28996);
nand UO_501 (O_501,N_29200,N_29297);
xnor UO_502 (O_502,N_29224,N_29062);
xor UO_503 (O_503,N_29928,N_28201);
nand UO_504 (O_504,N_29302,N_29265);
and UO_505 (O_505,N_29480,N_29310);
and UO_506 (O_506,N_28844,N_28102);
nor UO_507 (O_507,N_29704,N_28690);
nor UO_508 (O_508,N_29431,N_29778);
nor UO_509 (O_509,N_29453,N_28714);
xor UO_510 (O_510,N_29877,N_29603);
nor UO_511 (O_511,N_28077,N_28362);
nor UO_512 (O_512,N_28722,N_29273);
nor UO_513 (O_513,N_29516,N_28777);
or UO_514 (O_514,N_28835,N_28314);
xnor UO_515 (O_515,N_28357,N_29419);
and UO_516 (O_516,N_28983,N_29378);
or UO_517 (O_517,N_28230,N_29191);
or UO_518 (O_518,N_28612,N_29365);
or UO_519 (O_519,N_28766,N_28444);
xor UO_520 (O_520,N_29123,N_28498);
or UO_521 (O_521,N_28294,N_29596);
nor UO_522 (O_522,N_29027,N_28665);
nor UO_523 (O_523,N_29810,N_29554);
xnor UO_524 (O_524,N_28627,N_29558);
and UO_525 (O_525,N_29105,N_29134);
xor UO_526 (O_526,N_29383,N_29989);
or UO_527 (O_527,N_28338,N_29403);
xor UO_528 (O_528,N_29906,N_29864);
or UO_529 (O_529,N_29095,N_29694);
or UO_530 (O_530,N_29412,N_28843);
nor UO_531 (O_531,N_28368,N_29303);
xor UO_532 (O_532,N_29597,N_29926);
nand UO_533 (O_533,N_29184,N_29550);
xor UO_534 (O_534,N_28719,N_28307);
or UO_535 (O_535,N_28171,N_29510);
nand UO_536 (O_536,N_28862,N_29616);
and UO_537 (O_537,N_29600,N_28936);
nor UO_538 (O_538,N_28653,N_28299);
nand UO_539 (O_539,N_29244,N_29187);
nand UO_540 (O_540,N_29621,N_28335);
or UO_541 (O_541,N_28945,N_29846);
xor UO_542 (O_542,N_28160,N_29242);
and UO_543 (O_543,N_29792,N_28587);
and UO_544 (O_544,N_29028,N_28002);
xnor UO_545 (O_545,N_28894,N_28604);
nor UO_546 (O_546,N_29455,N_28280);
and UO_547 (O_547,N_28234,N_28571);
xnor UO_548 (O_548,N_29307,N_28761);
nor UO_549 (O_549,N_29148,N_28405);
xnor UO_550 (O_550,N_29088,N_28711);
nor UO_551 (O_551,N_28608,N_29650);
nor UO_552 (O_552,N_28496,N_28861);
or UO_553 (O_553,N_28365,N_29533);
nor UO_554 (O_554,N_29970,N_28563);
nand UO_555 (O_555,N_29531,N_29044);
nand UO_556 (O_556,N_28332,N_29733);
or UO_557 (O_557,N_29033,N_29394);
or UO_558 (O_558,N_28639,N_28042);
xnor UO_559 (O_559,N_29903,N_29092);
xor UO_560 (O_560,N_28941,N_28144);
nor UO_561 (O_561,N_29097,N_28245);
and UO_562 (O_562,N_29893,N_29437);
nand UO_563 (O_563,N_28135,N_29501);
nor UO_564 (O_564,N_28728,N_29150);
nor UO_565 (O_565,N_29872,N_28407);
nor UO_566 (O_566,N_28235,N_29953);
xor UO_567 (O_567,N_28204,N_29216);
nand UO_568 (O_568,N_29449,N_29858);
or UO_569 (O_569,N_29282,N_29479);
and UO_570 (O_570,N_28557,N_29662);
xor UO_571 (O_571,N_29610,N_28132);
nand UO_572 (O_572,N_28454,N_29920);
nor UO_573 (O_573,N_28382,N_28317);
xnor UO_574 (O_574,N_29215,N_28628);
nand UO_575 (O_575,N_28891,N_29612);
xnor UO_576 (O_576,N_29002,N_29759);
nand UO_577 (O_577,N_29249,N_28681);
or UO_578 (O_578,N_29574,N_29426);
xor UO_579 (O_579,N_29690,N_28831);
xnor UO_580 (O_580,N_28081,N_28596);
or UO_581 (O_581,N_29902,N_28146);
xor UO_582 (O_582,N_28796,N_28811);
nand UO_583 (O_583,N_28724,N_28847);
nor UO_584 (O_584,N_29421,N_29472);
and UO_585 (O_585,N_28105,N_28343);
or UO_586 (O_586,N_29012,N_28830);
nand UO_587 (O_587,N_29547,N_29570);
and UO_588 (O_588,N_28212,N_29237);
and UO_589 (O_589,N_29010,N_29153);
and UO_590 (O_590,N_29351,N_29900);
and UO_591 (O_591,N_29598,N_29808);
xnor UO_592 (O_592,N_28871,N_29389);
or UO_593 (O_593,N_28727,N_28971);
or UO_594 (O_594,N_29726,N_28364);
xnor UO_595 (O_595,N_29202,N_28111);
nor UO_596 (O_596,N_29540,N_28901);
or UO_597 (O_597,N_28100,N_28188);
nor UO_598 (O_598,N_28088,N_29781);
nand UO_599 (O_599,N_29764,N_29285);
nor UO_600 (O_600,N_28326,N_28918);
nor UO_601 (O_601,N_29471,N_29782);
nor UO_602 (O_602,N_28428,N_29175);
nand UO_603 (O_603,N_28824,N_28424);
or UO_604 (O_604,N_28620,N_28452);
nand UO_605 (O_605,N_28635,N_28743);
nand UO_606 (O_606,N_28805,N_29687);
nand UO_607 (O_607,N_28263,N_28595);
xor UO_608 (O_608,N_28018,N_28264);
nand UO_609 (O_609,N_29823,N_29834);
xor UO_610 (O_610,N_29555,N_29051);
nor UO_611 (O_611,N_28491,N_28055);
xnor UO_612 (O_612,N_28084,N_28813);
and UO_613 (O_613,N_28685,N_28531);
and UO_614 (O_614,N_28158,N_28872);
nor UO_615 (O_615,N_28023,N_29560);
nor UO_616 (O_616,N_29211,N_28708);
nor UO_617 (O_617,N_28035,N_28932);
nand UO_618 (O_618,N_29575,N_29402);
nand UO_619 (O_619,N_29497,N_29017);
nand UO_620 (O_620,N_28127,N_29620);
nor UO_621 (O_621,N_29975,N_28391);
nand UO_622 (O_622,N_28792,N_28095);
xnor UO_623 (O_623,N_28101,N_28594);
xnor UO_624 (O_624,N_29352,N_29245);
and UO_625 (O_625,N_29422,N_29137);
xor UO_626 (O_626,N_28323,N_28445);
nor UO_627 (O_627,N_28827,N_29880);
and UO_628 (O_628,N_29100,N_29358);
and UO_629 (O_629,N_29679,N_29788);
or UO_630 (O_630,N_28990,N_29353);
and UO_631 (O_631,N_29710,N_29229);
nor UO_632 (O_632,N_29138,N_29034);
xnor UO_633 (O_633,N_29727,N_28818);
nand UO_634 (O_634,N_29676,N_28199);
nor UO_635 (O_635,N_28526,N_28632);
or UO_636 (O_636,N_29614,N_28504);
and UO_637 (O_637,N_28976,N_28781);
and UO_638 (O_638,N_29804,N_28211);
or UO_639 (O_639,N_28080,N_28634);
xor UO_640 (O_640,N_28790,N_29711);
or UO_641 (O_641,N_29638,N_29999);
xnor UO_642 (O_642,N_29040,N_28380);
or UO_643 (O_643,N_28253,N_29324);
or UO_644 (O_644,N_28478,N_28032);
and UO_645 (O_645,N_28142,N_29005);
nor UO_646 (O_646,N_28696,N_28763);
xor UO_647 (O_647,N_28944,N_28616);
or UO_648 (O_648,N_29811,N_28168);
nor UO_649 (O_649,N_28974,N_29026);
and UO_650 (O_650,N_29287,N_29998);
xor UO_651 (O_651,N_29912,N_29135);
nand UO_652 (O_652,N_29519,N_28479);
xor UO_653 (O_653,N_29583,N_29749);
or UO_654 (O_654,N_28015,N_29257);
nor UO_655 (O_655,N_29588,N_29699);
xnor UO_656 (O_656,N_29827,N_29179);
nor UO_657 (O_657,N_28837,N_29771);
nor UO_658 (O_658,N_29907,N_28437);
and UO_659 (O_659,N_29840,N_28558);
and UO_660 (O_660,N_28788,N_29832);
xnor UO_661 (O_661,N_28893,N_28902);
nor UO_662 (O_662,N_29319,N_29410);
or UO_663 (O_663,N_29728,N_29014);
or UO_664 (O_664,N_29919,N_29098);
and UO_665 (O_665,N_28465,N_29747);
or UO_666 (O_666,N_28404,N_28684);
nand UO_667 (O_667,N_28982,N_29571);
xor UO_668 (O_668,N_29263,N_29523);
nand UO_669 (O_669,N_28880,N_28350);
or UO_670 (O_670,N_29064,N_29492);
or UO_671 (O_671,N_28589,N_28789);
and UO_672 (O_672,N_28270,N_28483);
xor UO_673 (O_673,N_28986,N_29169);
or UO_674 (O_674,N_28615,N_29296);
nand UO_675 (O_675,N_29205,N_28543);
nand UO_676 (O_676,N_29119,N_28525);
nor UO_677 (O_677,N_29648,N_28522);
xnor UO_678 (O_678,N_29796,N_28749);
xor UO_679 (O_679,N_29591,N_28922);
or UO_680 (O_680,N_29982,N_28514);
xor UO_681 (O_681,N_28031,N_29366);
nor UO_682 (O_682,N_28723,N_29617);
or UO_683 (O_683,N_29892,N_28001);
nor UO_684 (O_684,N_29435,N_28878);
nor UO_685 (O_685,N_29713,N_28337);
or UO_686 (O_686,N_29882,N_28442);
nor UO_687 (O_687,N_29542,N_29071);
nor UO_688 (O_688,N_29528,N_28455);
nand UO_689 (O_689,N_28925,N_28120);
nand UO_690 (O_690,N_29099,N_28912);
or UO_691 (O_691,N_28416,N_29114);
xor UO_692 (O_692,N_29821,N_29322);
or UO_693 (O_693,N_28225,N_28182);
xor UO_694 (O_694,N_29509,N_29059);
xnor UO_695 (O_695,N_29230,N_28762);
nand UO_696 (O_696,N_28136,N_29972);
and UO_697 (O_697,N_28877,N_28197);
or UO_698 (O_698,N_29429,N_29301);
and UO_699 (O_699,N_29035,N_29665);
xor UO_700 (O_700,N_28644,N_29626);
nor UO_701 (O_701,N_29011,N_28574);
and UO_702 (O_702,N_29779,N_28226);
xor UO_703 (O_703,N_28780,N_29414);
xnor UO_704 (O_704,N_29344,N_28812);
xor UO_705 (O_705,N_29505,N_28515);
nor UO_706 (O_706,N_28876,N_28946);
and UO_707 (O_707,N_28030,N_28302);
nor UO_708 (O_708,N_28957,N_28993);
nand UO_709 (O_709,N_28846,N_29897);
nor UO_710 (O_710,N_28148,N_29865);
or UO_711 (O_711,N_28603,N_29753);
xnor UO_712 (O_712,N_28767,N_28972);
xor UO_713 (O_713,N_29628,N_28659);
nand UO_714 (O_714,N_28960,N_29937);
or UO_715 (O_715,N_29539,N_29576);
xor UO_716 (O_716,N_28849,N_29060);
and UO_717 (O_717,N_29688,N_28322);
and UO_718 (O_718,N_28833,N_28657);
xnor UO_719 (O_719,N_28207,N_28099);
xnor UO_720 (O_720,N_29259,N_28779);
and UO_721 (O_721,N_29769,N_28702);
nor UO_722 (O_722,N_29719,N_29881);
nor UO_723 (O_723,N_28909,N_28521);
xnor UO_724 (O_724,N_29018,N_29641);
nor UO_725 (O_725,N_28202,N_29199);
nand UO_726 (O_726,N_29664,N_28569);
and UO_727 (O_727,N_28669,N_28344);
or UO_728 (O_728,N_28180,N_28054);
nand UO_729 (O_729,N_28636,N_28852);
and UO_730 (O_730,N_29862,N_29125);
nor UO_731 (O_731,N_28802,N_29438);
or UO_732 (O_732,N_28351,N_28949);
xnor UO_733 (O_733,N_28128,N_28736);
nor UO_734 (O_734,N_28059,N_28401);
and UO_735 (O_735,N_29180,N_28565);
nor UO_736 (O_736,N_28418,N_28123);
or UO_737 (O_737,N_28259,N_28700);
nand UO_738 (O_738,N_29206,N_28943);
nor UO_739 (O_739,N_28530,N_28721);
and UO_740 (O_740,N_28739,N_28856);
xnor UO_741 (O_741,N_29081,N_28098);
or UO_742 (O_742,N_28572,N_29996);
nor UO_743 (O_743,N_28346,N_29838);
nor UO_744 (O_744,N_29478,N_28312);
and UO_745 (O_745,N_29855,N_29311);
and UO_746 (O_746,N_28033,N_29819);
xnor UO_747 (O_747,N_29065,N_29227);
and UO_748 (O_748,N_28310,N_29507);
nand UO_749 (O_749,N_29681,N_29932);
or UO_750 (O_750,N_28823,N_28955);
xnor UO_751 (O_751,N_28582,N_28593);
nand UO_752 (O_752,N_28646,N_28746);
xor UO_753 (O_753,N_28292,N_29675);
or UO_754 (O_754,N_28799,N_28229);
xnor UO_755 (O_755,N_28072,N_29739);
nand UO_756 (O_756,N_29093,N_28654);
nor UO_757 (O_757,N_29238,N_29964);
nor UO_758 (O_758,N_28963,N_28141);
nand UO_759 (O_759,N_28467,N_28989);
nor UO_760 (O_760,N_28664,N_29898);
xnor UO_761 (O_761,N_28008,N_28640);
or UO_762 (O_762,N_28851,N_29587);
nor UO_763 (O_763,N_29197,N_29673);
or UO_764 (O_764,N_29706,N_29736);
or UO_765 (O_765,N_28383,N_29345);
and UO_766 (O_766,N_28089,N_29127);
and UO_767 (O_767,N_29055,N_29029);
nor UO_768 (O_768,N_28611,N_28517);
xnor UO_769 (O_769,N_29270,N_28729);
or UO_770 (O_770,N_28224,N_28427);
xnor UO_771 (O_771,N_28953,N_28638);
nand UO_772 (O_772,N_29461,N_28210);
nand UO_773 (O_773,N_28750,N_29568);
nor UO_774 (O_774,N_29495,N_28667);
nor UO_775 (O_775,N_29374,N_28331);
xnor UO_776 (O_776,N_28933,N_28704);
and UO_777 (O_777,N_28693,N_29408);
and UO_778 (O_778,N_28353,N_29168);
or UO_779 (O_779,N_29299,N_29724);
xnor UO_780 (O_780,N_29601,N_28087);
nand UO_781 (O_781,N_29866,N_29152);
and UO_782 (O_782,N_28511,N_28039);
or UO_783 (O_783,N_29521,N_29940);
or UO_784 (O_784,N_28492,N_29828);
nor UO_785 (O_785,N_29160,N_28432);
nand UO_786 (O_786,N_29730,N_29015);
xor UO_787 (O_787,N_28740,N_28196);
or UO_788 (O_788,N_29632,N_29683);
nand UO_789 (O_789,N_28617,N_28747);
xor UO_790 (O_790,N_29141,N_29988);
nand UO_791 (O_791,N_29284,N_29022);
nor UO_792 (O_792,N_29873,N_29336);
nor UO_793 (O_793,N_29268,N_28359);
nand UO_794 (O_794,N_28677,N_29860);
nor UO_795 (O_795,N_29103,N_28285);
xnor UO_796 (O_796,N_29355,N_28560);
or UO_797 (O_797,N_29464,N_28732);
nand UO_798 (O_798,N_28535,N_28086);
or UO_799 (O_799,N_28931,N_29349);
nand UO_800 (O_800,N_28273,N_29375);
xor UO_801 (O_801,N_28994,N_29433);
nand UO_802 (O_802,N_29784,N_28538);
or UO_803 (O_803,N_29748,N_29490);
nand UO_804 (O_804,N_28266,N_29207);
xor UO_805 (O_805,N_29895,N_29305);
or UO_806 (O_806,N_29494,N_28892);
and UO_807 (O_807,N_29599,N_29646);
and UO_808 (O_808,N_29861,N_29049);
nor UO_809 (O_809,N_29755,N_29167);
nand UO_810 (O_810,N_28875,N_29107);
xor UO_811 (O_811,N_28622,N_28091);
or UO_812 (O_812,N_28584,N_29189);
or UO_813 (O_813,N_28853,N_29927);
xnor UO_814 (O_814,N_28395,N_28609);
nand UO_815 (O_815,N_29053,N_29824);
or UO_816 (O_816,N_28177,N_28771);
xnor UO_817 (O_817,N_29091,N_28624);
xnor UO_818 (O_818,N_28505,N_29157);
nor UO_819 (O_819,N_28984,N_29499);
or UO_820 (O_820,N_29522,N_28239);
xor UO_821 (O_821,N_29787,N_28924);
nor UO_822 (O_822,N_28533,N_29251);
or UO_823 (O_823,N_28435,N_28493);
nand UO_824 (O_824,N_29371,N_29400);
or UO_825 (O_825,N_29949,N_28400);
or UO_826 (O_826,N_29424,N_29108);
or UO_827 (O_827,N_28246,N_29894);
nand UO_828 (O_828,N_29304,N_28967);
or UO_829 (O_829,N_29631,N_28131);
and UO_830 (O_830,N_29020,N_28053);
or UO_831 (O_831,N_29737,N_29845);
or UO_832 (O_832,N_29295,N_29886);
or UO_833 (O_833,N_29783,N_28093);
nor UO_834 (O_834,N_28675,N_29801);
nor UO_835 (O_835,N_29021,N_28570);
or UO_836 (O_836,N_29950,N_28108);
nand UO_837 (O_837,N_29121,N_29822);
or UO_838 (O_838,N_28150,N_29459);
xnor UO_839 (O_839,N_29960,N_28956);
and UO_840 (O_840,N_29856,N_28752);
or UO_841 (O_841,N_29193,N_28896);
and UO_842 (O_842,N_28341,N_29799);
xnor UO_843 (O_843,N_28647,N_28318);
nand UO_844 (O_844,N_29602,N_29218);
nor UO_845 (O_845,N_28765,N_29670);
or UO_846 (O_846,N_29775,N_29515);
or UO_847 (O_847,N_28737,N_29425);
nand UO_848 (O_848,N_29234,N_29715);
nor UO_849 (O_849,N_29214,N_28159);
and UO_850 (O_850,N_28329,N_29904);
nand UO_851 (O_851,N_28366,N_28067);
xnor UO_852 (O_852,N_28661,N_28655);
nand UO_853 (O_853,N_28817,N_28860);
xnor UO_854 (O_854,N_28642,N_28174);
and UO_855 (O_855,N_28157,N_29146);
xor UO_856 (O_856,N_29518,N_29835);
xnor UO_857 (O_857,N_28848,N_28208);
xor UO_858 (O_858,N_29201,N_29340);
or UO_859 (O_859,N_29423,N_28184);
nor UO_860 (O_860,N_29929,N_29899);
and UO_861 (O_861,N_28092,N_29080);
xnor UO_862 (O_862,N_28475,N_28599);
or UO_863 (O_863,N_29181,N_28884);
and UO_864 (O_864,N_29654,N_29794);
xnor UO_865 (O_865,N_29987,N_29456);
nand UO_866 (O_866,N_28251,N_28520);
or UO_867 (O_867,N_29760,N_28378);
nand UO_868 (O_868,N_29458,N_29774);
and UO_869 (O_869,N_29863,N_28995);
nor UO_870 (O_870,N_28809,N_29347);
and UO_871 (O_871,N_28997,N_28725);
or UO_872 (O_872,N_29476,N_28534);
or UO_873 (O_873,N_29294,N_28448);
nor UO_874 (O_874,N_28576,N_28215);
or UO_875 (O_875,N_29976,N_29986);
or UO_876 (O_876,N_29008,N_28509);
nor UO_877 (O_877,N_29043,N_29980);
nor UO_878 (O_878,N_29592,N_28425);
nand UO_879 (O_879,N_29220,N_28874);
nand UO_880 (O_880,N_28216,N_28518);
and UO_881 (O_881,N_28821,N_28679);
nand UO_882 (O_882,N_28607,N_28214);
nor UO_883 (O_883,N_28223,N_28486);
nor UO_884 (O_884,N_28236,N_28985);
or UO_885 (O_885,N_29979,N_29586);
xor UO_886 (O_886,N_29283,N_29367);
xor UO_887 (O_887,N_28532,N_29329);
and UO_888 (O_888,N_29674,N_29954);
nor UO_889 (O_889,N_29050,N_29343);
and UO_890 (O_890,N_29219,N_28575);
nor UO_891 (O_891,N_28998,N_28623);
nor UO_892 (O_892,N_28774,N_28217);
nand UO_893 (O_893,N_29971,N_29913);
nor UO_894 (O_894,N_29767,N_29859);
xor UO_895 (O_895,N_29317,N_29396);
or UO_896 (O_896,N_28094,N_28085);
xor UO_897 (O_897,N_29178,N_28192);
and UO_898 (O_898,N_28601,N_28169);
or UO_899 (O_899,N_28656,N_29186);
xor UO_900 (O_900,N_29162,N_29063);
xnor UO_901 (O_901,N_29482,N_29113);
nand UO_902 (O_902,N_29791,N_28153);
and UO_903 (O_903,N_28939,N_29009);
and UO_904 (O_904,N_29908,N_28954);
xor UO_905 (O_905,N_29994,N_29637);
and UO_906 (O_906,N_28110,N_29447);
nor UO_907 (O_907,N_29993,N_29046);
nand UO_908 (O_908,N_29185,N_28580);
and UO_909 (O_909,N_28649,N_28502);
nand UO_910 (O_910,N_29194,N_28250);
nand UO_911 (O_911,N_29316,N_29457);
and UO_912 (O_912,N_28870,N_28970);
and UO_913 (O_913,N_29130,N_28349);
and UO_914 (O_914,N_28904,N_29286);
and UO_915 (O_915,N_29517,N_29565);
xor UO_916 (O_916,N_29663,N_28926);
and UO_917 (O_917,N_29763,N_29266);
xnor UO_918 (O_918,N_28260,N_28164);
nand UO_919 (O_919,N_28980,N_29723);
and UO_920 (O_920,N_29809,N_29384);
nand UO_921 (O_921,N_28959,N_29279);
xor UO_922 (O_922,N_29339,N_29924);
xor UO_923 (O_923,N_28240,N_29331);
nand UO_924 (O_924,N_29615,N_28673);
or UO_925 (O_925,N_28319,N_29546);
xnor UO_926 (O_926,N_28741,N_29768);
xnor UO_927 (O_927,N_29921,N_29678);
xnor UO_928 (O_928,N_29958,N_29922);
xor UO_929 (O_929,N_29451,N_28730);
xnor UO_930 (O_930,N_28258,N_28321);
xnor UO_931 (O_931,N_29604,N_29466);
nor UO_932 (O_932,N_28705,N_29001);
and UO_933 (O_933,N_29222,N_28457);
and UO_934 (O_934,N_28354,N_29584);
nor UO_935 (O_935,N_29780,N_29019);
nor UO_936 (O_936,N_29390,N_29981);
nor UO_937 (O_937,N_28859,N_29944);
xor UO_938 (O_938,N_29484,N_28237);
nor UO_939 (O_939,N_28600,N_29569);
nand UO_940 (O_940,N_29075,N_29241);
or UO_941 (O_941,N_28536,N_29702);
nand UO_942 (O_942,N_29373,N_28501);
or UO_943 (O_943,N_28429,N_28652);
nand UO_944 (O_944,N_29875,N_28293);
xor UO_945 (O_945,N_28806,N_28017);
and UO_946 (O_946,N_28695,N_28274);
and UO_947 (O_947,N_29563,N_28109);
nor UO_948 (O_948,N_28373,N_28392);
and UO_949 (O_949,N_29256,N_28172);
nor UO_950 (O_950,N_29691,N_29320);
nand UO_951 (O_951,N_28668,N_29445);
nor UO_952 (O_952,N_29440,N_29918);
xor UO_953 (O_953,N_29334,N_29136);
nor UO_954 (O_954,N_29038,N_29729);
and UO_955 (O_955,N_29368,N_29578);
and UO_956 (O_956,N_28676,N_28651);
nand UO_957 (O_957,N_29941,N_29874);
nor UO_958 (O_958,N_28564,N_28320);
and UO_959 (O_959,N_28785,N_29754);
nand UO_960 (O_960,N_29450,N_29313);
xor UO_961 (O_961,N_28339,N_29354);
or UO_962 (O_962,N_29557,N_29398);
xnor UO_963 (O_963,N_28744,N_29052);
or UO_964 (O_964,N_29068,N_29746);
nand UO_965 (O_965,N_29513,N_28006);
or UO_966 (O_966,N_28389,N_29379);
xnor UO_967 (O_967,N_29843,N_29756);
and UO_968 (O_968,N_29966,N_28688);
nand UO_969 (O_969,N_28311,N_28062);
or UO_970 (O_970,N_28000,N_28064);
nand UO_971 (O_971,N_29067,N_28381);
xor UO_972 (O_972,N_29635,N_29640);
xnor UO_973 (O_973,N_28451,N_28300);
xnor UO_974 (O_974,N_29849,N_28021);
xnor UO_975 (O_975,N_28431,N_29758);
or UO_976 (O_976,N_29428,N_28660);
xnor UO_977 (O_977,N_28061,N_29776);
or UO_978 (O_978,N_28865,N_28325);
xnor UO_979 (O_979,N_29489,N_28689);
and UO_980 (O_980,N_28621,N_28333);
xnor UO_981 (O_981,N_28423,N_29611);
xor UO_982 (O_982,N_28934,N_29115);
nand UO_983 (O_983,N_28795,N_28186);
xnor UO_984 (O_984,N_28134,N_29330);
xnor UO_985 (O_985,N_28297,N_28816);
nor UO_986 (O_986,N_28082,N_29070);
or UO_987 (O_987,N_29236,N_29182);
or UO_988 (O_988,N_28775,N_29056);
nand UO_989 (O_989,N_29817,N_28929);
nor UO_990 (O_990,N_28247,N_29486);
or UO_991 (O_991,N_29420,N_28588);
nand UO_992 (O_992,N_29888,N_29815);
or UO_993 (O_993,N_29007,N_29839);
and UO_994 (O_994,N_28384,N_29176);
xnor UO_995 (O_995,N_29677,N_29475);
nor UO_996 (O_996,N_29750,N_29128);
xor UO_997 (O_997,N_29077,N_28009);
and UO_998 (O_998,N_28367,N_28073);
nor UO_999 (O_999,N_28992,N_29171);
or UO_1000 (O_1000,N_29250,N_28316);
or UO_1001 (O_1001,N_28795,N_29716);
and UO_1002 (O_1002,N_28481,N_28999);
nor UO_1003 (O_1003,N_29694,N_28246);
nor UO_1004 (O_1004,N_28984,N_29152);
nor UO_1005 (O_1005,N_28264,N_28477);
and UO_1006 (O_1006,N_28761,N_29498);
and UO_1007 (O_1007,N_29714,N_28044);
nor UO_1008 (O_1008,N_28958,N_29319);
or UO_1009 (O_1009,N_29098,N_29176);
or UO_1010 (O_1010,N_28289,N_29658);
or UO_1011 (O_1011,N_28291,N_29393);
xnor UO_1012 (O_1012,N_29938,N_29984);
nand UO_1013 (O_1013,N_28300,N_28342);
and UO_1014 (O_1014,N_28813,N_28179);
xor UO_1015 (O_1015,N_28381,N_28821);
xnor UO_1016 (O_1016,N_28421,N_29420);
or UO_1017 (O_1017,N_28088,N_28349);
nor UO_1018 (O_1018,N_28903,N_29968);
or UO_1019 (O_1019,N_29228,N_28958);
nor UO_1020 (O_1020,N_29325,N_28708);
xor UO_1021 (O_1021,N_29615,N_28290);
nor UO_1022 (O_1022,N_29942,N_29037);
nand UO_1023 (O_1023,N_28062,N_28961);
nand UO_1024 (O_1024,N_28114,N_28120);
xnor UO_1025 (O_1025,N_28356,N_29194);
nor UO_1026 (O_1026,N_29340,N_29869);
nand UO_1027 (O_1027,N_28248,N_28373);
nor UO_1028 (O_1028,N_29300,N_28466);
nor UO_1029 (O_1029,N_29170,N_28496);
nand UO_1030 (O_1030,N_29532,N_28841);
or UO_1031 (O_1031,N_28580,N_29310);
xnor UO_1032 (O_1032,N_28291,N_28521);
nor UO_1033 (O_1033,N_29346,N_28593);
or UO_1034 (O_1034,N_28536,N_28363);
and UO_1035 (O_1035,N_28948,N_28768);
or UO_1036 (O_1036,N_28976,N_29027);
or UO_1037 (O_1037,N_28020,N_28169);
nor UO_1038 (O_1038,N_29158,N_29627);
nand UO_1039 (O_1039,N_28174,N_28295);
nor UO_1040 (O_1040,N_29586,N_28761);
nor UO_1041 (O_1041,N_28675,N_28927);
and UO_1042 (O_1042,N_29255,N_29172);
and UO_1043 (O_1043,N_28011,N_28867);
xnor UO_1044 (O_1044,N_29024,N_28270);
xor UO_1045 (O_1045,N_28713,N_28091);
nor UO_1046 (O_1046,N_29224,N_29226);
or UO_1047 (O_1047,N_29524,N_28568);
and UO_1048 (O_1048,N_28531,N_28415);
xnor UO_1049 (O_1049,N_29296,N_28387);
nand UO_1050 (O_1050,N_28012,N_29978);
and UO_1051 (O_1051,N_28510,N_29703);
nand UO_1052 (O_1052,N_29702,N_28122);
and UO_1053 (O_1053,N_29919,N_29320);
xnor UO_1054 (O_1054,N_29422,N_29028);
or UO_1055 (O_1055,N_28811,N_29388);
or UO_1056 (O_1056,N_28340,N_29955);
or UO_1057 (O_1057,N_28091,N_28522);
and UO_1058 (O_1058,N_29216,N_28300);
nor UO_1059 (O_1059,N_28992,N_28482);
xnor UO_1060 (O_1060,N_28852,N_28446);
or UO_1061 (O_1061,N_28886,N_29452);
nand UO_1062 (O_1062,N_29068,N_29898);
nand UO_1063 (O_1063,N_29870,N_29197);
or UO_1064 (O_1064,N_28707,N_29191);
xor UO_1065 (O_1065,N_28740,N_28616);
nor UO_1066 (O_1066,N_28460,N_29978);
nand UO_1067 (O_1067,N_28009,N_29124);
and UO_1068 (O_1068,N_29055,N_28772);
nand UO_1069 (O_1069,N_29314,N_29960);
xor UO_1070 (O_1070,N_29265,N_28037);
or UO_1071 (O_1071,N_29901,N_29956);
and UO_1072 (O_1072,N_28311,N_29709);
nand UO_1073 (O_1073,N_29404,N_29482);
or UO_1074 (O_1074,N_29102,N_28434);
or UO_1075 (O_1075,N_29712,N_28832);
nand UO_1076 (O_1076,N_28761,N_28035);
xor UO_1077 (O_1077,N_28814,N_29304);
xnor UO_1078 (O_1078,N_28605,N_29155);
xor UO_1079 (O_1079,N_28762,N_29226);
xor UO_1080 (O_1080,N_28421,N_29802);
nor UO_1081 (O_1081,N_29049,N_28046);
nor UO_1082 (O_1082,N_29378,N_29132);
nand UO_1083 (O_1083,N_29411,N_28272);
and UO_1084 (O_1084,N_28397,N_29079);
and UO_1085 (O_1085,N_29563,N_29038);
nor UO_1086 (O_1086,N_29595,N_28795);
and UO_1087 (O_1087,N_28896,N_28261);
nor UO_1088 (O_1088,N_28797,N_28559);
or UO_1089 (O_1089,N_28843,N_29722);
nor UO_1090 (O_1090,N_29721,N_28196);
nand UO_1091 (O_1091,N_29295,N_28707);
or UO_1092 (O_1092,N_29010,N_28283);
nand UO_1093 (O_1093,N_29202,N_28094);
xor UO_1094 (O_1094,N_28197,N_28705);
or UO_1095 (O_1095,N_29536,N_28099);
and UO_1096 (O_1096,N_28281,N_28974);
xnor UO_1097 (O_1097,N_28952,N_28466);
or UO_1098 (O_1098,N_28016,N_28062);
nand UO_1099 (O_1099,N_29644,N_28724);
nor UO_1100 (O_1100,N_28330,N_29296);
xnor UO_1101 (O_1101,N_29823,N_28589);
nor UO_1102 (O_1102,N_28705,N_28547);
or UO_1103 (O_1103,N_28994,N_28546);
or UO_1104 (O_1104,N_28820,N_29792);
nand UO_1105 (O_1105,N_28641,N_29942);
nor UO_1106 (O_1106,N_29045,N_29093);
xnor UO_1107 (O_1107,N_28323,N_28447);
or UO_1108 (O_1108,N_29238,N_29102);
or UO_1109 (O_1109,N_28489,N_29774);
xnor UO_1110 (O_1110,N_28618,N_29005);
nor UO_1111 (O_1111,N_28572,N_28323);
nand UO_1112 (O_1112,N_28451,N_28490);
or UO_1113 (O_1113,N_28291,N_28640);
and UO_1114 (O_1114,N_29831,N_29267);
nand UO_1115 (O_1115,N_28598,N_29682);
nand UO_1116 (O_1116,N_28196,N_28324);
xnor UO_1117 (O_1117,N_29497,N_28817);
nor UO_1118 (O_1118,N_29437,N_28142);
nor UO_1119 (O_1119,N_29926,N_28918);
and UO_1120 (O_1120,N_28061,N_29159);
xnor UO_1121 (O_1121,N_28950,N_28748);
nand UO_1122 (O_1122,N_29227,N_29281);
or UO_1123 (O_1123,N_28482,N_28688);
nor UO_1124 (O_1124,N_28437,N_29222);
xor UO_1125 (O_1125,N_28258,N_29124);
or UO_1126 (O_1126,N_28003,N_29486);
nand UO_1127 (O_1127,N_28033,N_29352);
nor UO_1128 (O_1128,N_28573,N_28423);
nand UO_1129 (O_1129,N_28975,N_29965);
or UO_1130 (O_1130,N_29982,N_28551);
or UO_1131 (O_1131,N_28780,N_28754);
nand UO_1132 (O_1132,N_29046,N_28988);
and UO_1133 (O_1133,N_28735,N_28822);
nor UO_1134 (O_1134,N_29963,N_28807);
xor UO_1135 (O_1135,N_29455,N_29031);
xnor UO_1136 (O_1136,N_28001,N_28911);
xnor UO_1137 (O_1137,N_28556,N_28760);
nor UO_1138 (O_1138,N_28969,N_29953);
nand UO_1139 (O_1139,N_28497,N_28994);
or UO_1140 (O_1140,N_29706,N_28595);
and UO_1141 (O_1141,N_28715,N_28049);
nand UO_1142 (O_1142,N_28269,N_28858);
or UO_1143 (O_1143,N_29585,N_29205);
xnor UO_1144 (O_1144,N_28710,N_28158);
or UO_1145 (O_1145,N_28038,N_28765);
nand UO_1146 (O_1146,N_29061,N_29440);
nand UO_1147 (O_1147,N_29525,N_29998);
xnor UO_1148 (O_1148,N_29427,N_28813);
nor UO_1149 (O_1149,N_29855,N_29783);
nand UO_1150 (O_1150,N_28669,N_28914);
xnor UO_1151 (O_1151,N_29736,N_28175);
and UO_1152 (O_1152,N_28604,N_29990);
and UO_1153 (O_1153,N_28952,N_29354);
nor UO_1154 (O_1154,N_28929,N_29539);
and UO_1155 (O_1155,N_29973,N_28789);
nand UO_1156 (O_1156,N_29864,N_28714);
or UO_1157 (O_1157,N_29366,N_28946);
nor UO_1158 (O_1158,N_28155,N_28756);
nor UO_1159 (O_1159,N_29942,N_28280);
or UO_1160 (O_1160,N_29484,N_29739);
or UO_1161 (O_1161,N_29450,N_28310);
nand UO_1162 (O_1162,N_29002,N_29264);
nand UO_1163 (O_1163,N_29649,N_28444);
xor UO_1164 (O_1164,N_29747,N_28256);
or UO_1165 (O_1165,N_29928,N_29023);
nor UO_1166 (O_1166,N_29301,N_29496);
nor UO_1167 (O_1167,N_29106,N_29224);
or UO_1168 (O_1168,N_28311,N_28167);
nor UO_1169 (O_1169,N_28973,N_29082);
nor UO_1170 (O_1170,N_28673,N_29870);
nand UO_1171 (O_1171,N_29034,N_29135);
nand UO_1172 (O_1172,N_29270,N_29729);
nand UO_1173 (O_1173,N_28348,N_29904);
xor UO_1174 (O_1174,N_28780,N_28729);
nor UO_1175 (O_1175,N_29906,N_29670);
nand UO_1176 (O_1176,N_28301,N_28642);
nand UO_1177 (O_1177,N_28616,N_29269);
and UO_1178 (O_1178,N_29316,N_29892);
xor UO_1179 (O_1179,N_28011,N_29674);
and UO_1180 (O_1180,N_29430,N_28981);
and UO_1181 (O_1181,N_28016,N_29403);
and UO_1182 (O_1182,N_29570,N_29836);
and UO_1183 (O_1183,N_29288,N_29553);
nand UO_1184 (O_1184,N_28287,N_28377);
nand UO_1185 (O_1185,N_29465,N_28888);
and UO_1186 (O_1186,N_29021,N_29303);
and UO_1187 (O_1187,N_28229,N_28512);
nand UO_1188 (O_1188,N_29155,N_29551);
or UO_1189 (O_1189,N_29231,N_29058);
and UO_1190 (O_1190,N_28697,N_28845);
xor UO_1191 (O_1191,N_28489,N_29736);
xnor UO_1192 (O_1192,N_29869,N_28413);
nor UO_1193 (O_1193,N_28863,N_29324);
nand UO_1194 (O_1194,N_28972,N_29795);
nand UO_1195 (O_1195,N_29208,N_28391);
xor UO_1196 (O_1196,N_28567,N_29466);
nor UO_1197 (O_1197,N_29080,N_28849);
and UO_1198 (O_1198,N_29232,N_29302);
nand UO_1199 (O_1199,N_29379,N_28674);
nor UO_1200 (O_1200,N_29061,N_28750);
xnor UO_1201 (O_1201,N_28722,N_29649);
or UO_1202 (O_1202,N_29701,N_28260);
xnor UO_1203 (O_1203,N_28865,N_28282);
xnor UO_1204 (O_1204,N_29308,N_29052);
nand UO_1205 (O_1205,N_29999,N_28225);
nor UO_1206 (O_1206,N_29858,N_29665);
nand UO_1207 (O_1207,N_28723,N_28559);
nand UO_1208 (O_1208,N_29236,N_28877);
xnor UO_1209 (O_1209,N_28921,N_29576);
nand UO_1210 (O_1210,N_28661,N_29452);
and UO_1211 (O_1211,N_29904,N_29348);
nor UO_1212 (O_1212,N_29474,N_28838);
nand UO_1213 (O_1213,N_28454,N_29151);
nor UO_1214 (O_1214,N_28472,N_29130);
xor UO_1215 (O_1215,N_28416,N_28983);
xor UO_1216 (O_1216,N_29553,N_28990);
and UO_1217 (O_1217,N_28419,N_29314);
or UO_1218 (O_1218,N_29620,N_29586);
xnor UO_1219 (O_1219,N_28135,N_28528);
or UO_1220 (O_1220,N_28183,N_28991);
or UO_1221 (O_1221,N_29094,N_28556);
nor UO_1222 (O_1222,N_28675,N_28670);
or UO_1223 (O_1223,N_29754,N_28718);
xor UO_1224 (O_1224,N_28902,N_29084);
or UO_1225 (O_1225,N_29713,N_29098);
nor UO_1226 (O_1226,N_29754,N_29473);
and UO_1227 (O_1227,N_29325,N_28069);
or UO_1228 (O_1228,N_28210,N_29884);
nor UO_1229 (O_1229,N_28991,N_28623);
and UO_1230 (O_1230,N_29173,N_28201);
nand UO_1231 (O_1231,N_29498,N_28058);
or UO_1232 (O_1232,N_28120,N_29129);
nand UO_1233 (O_1233,N_28974,N_29289);
nor UO_1234 (O_1234,N_28050,N_28641);
nand UO_1235 (O_1235,N_29123,N_29067);
xor UO_1236 (O_1236,N_28941,N_28947);
xor UO_1237 (O_1237,N_29014,N_28332);
and UO_1238 (O_1238,N_28445,N_28811);
and UO_1239 (O_1239,N_29573,N_29040);
nor UO_1240 (O_1240,N_29718,N_28576);
nor UO_1241 (O_1241,N_28527,N_28311);
xor UO_1242 (O_1242,N_28810,N_28612);
nand UO_1243 (O_1243,N_28655,N_29735);
nor UO_1244 (O_1244,N_29294,N_29157);
nand UO_1245 (O_1245,N_29479,N_28905);
nand UO_1246 (O_1246,N_28551,N_28631);
xor UO_1247 (O_1247,N_29415,N_28035);
nand UO_1248 (O_1248,N_29997,N_28796);
or UO_1249 (O_1249,N_29960,N_28504);
xor UO_1250 (O_1250,N_29896,N_28053);
nand UO_1251 (O_1251,N_29446,N_29406);
and UO_1252 (O_1252,N_28943,N_29145);
xor UO_1253 (O_1253,N_28186,N_28559);
or UO_1254 (O_1254,N_29696,N_28897);
nor UO_1255 (O_1255,N_29522,N_29107);
nor UO_1256 (O_1256,N_29405,N_28836);
nand UO_1257 (O_1257,N_28291,N_29426);
xnor UO_1258 (O_1258,N_29935,N_28919);
or UO_1259 (O_1259,N_28759,N_28798);
xnor UO_1260 (O_1260,N_29303,N_29467);
or UO_1261 (O_1261,N_28015,N_29035);
nand UO_1262 (O_1262,N_28378,N_29205);
or UO_1263 (O_1263,N_28256,N_28255);
xnor UO_1264 (O_1264,N_29555,N_28033);
nand UO_1265 (O_1265,N_28095,N_28079);
nor UO_1266 (O_1266,N_28400,N_28845);
and UO_1267 (O_1267,N_28992,N_29922);
nor UO_1268 (O_1268,N_28934,N_28776);
nor UO_1269 (O_1269,N_29595,N_29183);
or UO_1270 (O_1270,N_28482,N_29449);
or UO_1271 (O_1271,N_28634,N_29510);
or UO_1272 (O_1272,N_28553,N_29316);
nor UO_1273 (O_1273,N_28128,N_29225);
nand UO_1274 (O_1274,N_29726,N_29494);
or UO_1275 (O_1275,N_28828,N_28572);
nand UO_1276 (O_1276,N_29159,N_28325);
and UO_1277 (O_1277,N_28109,N_28305);
xnor UO_1278 (O_1278,N_28212,N_29033);
xnor UO_1279 (O_1279,N_29546,N_28500);
and UO_1280 (O_1280,N_28117,N_29412);
and UO_1281 (O_1281,N_29409,N_29225);
or UO_1282 (O_1282,N_28317,N_29878);
nor UO_1283 (O_1283,N_29088,N_28017);
nor UO_1284 (O_1284,N_29955,N_28844);
or UO_1285 (O_1285,N_28761,N_28899);
or UO_1286 (O_1286,N_29245,N_28448);
xnor UO_1287 (O_1287,N_29217,N_28168);
and UO_1288 (O_1288,N_29383,N_29322);
nor UO_1289 (O_1289,N_29211,N_29922);
xor UO_1290 (O_1290,N_28444,N_28379);
nand UO_1291 (O_1291,N_28586,N_28774);
and UO_1292 (O_1292,N_28491,N_28286);
nor UO_1293 (O_1293,N_29547,N_28777);
nor UO_1294 (O_1294,N_28307,N_29761);
or UO_1295 (O_1295,N_28300,N_29147);
and UO_1296 (O_1296,N_29334,N_29953);
or UO_1297 (O_1297,N_28491,N_29281);
or UO_1298 (O_1298,N_29509,N_28425);
or UO_1299 (O_1299,N_28838,N_28662);
nand UO_1300 (O_1300,N_28734,N_29402);
and UO_1301 (O_1301,N_29238,N_29661);
xnor UO_1302 (O_1302,N_28023,N_29054);
and UO_1303 (O_1303,N_29793,N_28916);
nor UO_1304 (O_1304,N_28386,N_29796);
and UO_1305 (O_1305,N_29175,N_28389);
or UO_1306 (O_1306,N_28982,N_29539);
nor UO_1307 (O_1307,N_29356,N_29959);
and UO_1308 (O_1308,N_29476,N_29992);
nor UO_1309 (O_1309,N_29972,N_29798);
and UO_1310 (O_1310,N_29035,N_29503);
nor UO_1311 (O_1311,N_29090,N_28974);
nand UO_1312 (O_1312,N_29586,N_29008);
and UO_1313 (O_1313,N_28418,N_28769);
and UO_1314 (O_1314,N_28394,N_29703);
nand UO_1315 (O_1315,N_28260,N_28327);
nor UO_1316 (O_1316,N_29478,N_29884);
nand UO_1317 (O_1317,N_28442,N_28709);
or UO_1318 (O_1318,N_28931,N_28316);
nand UO_1319 (O_1319,N_28236,N_29340);
and UO_1320 (O_1320,N_29472,N_29961);
nor UO_1321 (O_1321,N_29805,N_28106);
xnor UO_1322 (O_1322,N_28317,N_28659);
xor UO_1323 (O_1323,N_28904,N_28321);
or UO_1324 (O_1324,N_29507,N_28283);
xnor UO_1325 (O_1325,N_29448,N_28309);
nand UO_1326 (O_1326,N_29826,N_28177);
nor UO_1327 (O_1327,N_29307,N_28222);
and UO_1328 (O_1328,N_28552,N_29855);
or UO_1329 (O_1329,N_28926,N_29060);
xnor UO_1330 (O_1330,N_28439,N_28925);
xnor UO_1331 (O_1331,N_29240,N_28999);
nor UO_1332 (O_1332,N_29004,N_29199);
or UO_1333 (O_1333,N_29893,N_29710);
and UO_1334 (O_1334,N_29725,N_28374);
nand UO_1335 (O_1335,N_29623,N_28208);
nor UO_1336 (O_1336,N_28590,N_28720);
and UO_1337 (O_1337,N_29869,N_29077);
or UO_1338 (O_1338,N_29910,N_28255);
nor UO_1339 (O_1339,N_29856,N_29067);
nor UO_1340 (O_1340,N_28378,N_28556);
or UO_1341 (O_1341,N_29062,N_29752);
or UO_1342 (O_1342,N_28871,N_29021);
and UO_1343 (O_1343,N_28849,N_29565);
xnor UO_1344 (O_1344,N_28438,N_29993);
nand UO_1345 (O_1345,N_28408,N_29937);
and UO_1346 (O_1346,N_28592,N_29394);
or UO_1347 (O_1347,N_28996,N_28955);
xor UO_1348 (O_1348,N_29249,N_29817);
xnor UO_1349 (O_1349,N_29328,N_28753);
or UO_1350 (O_1350,N_28771,N_29501);
nand UO_1351 (O_1351,N_28336,N_29814);
and UO_1352 (O_1352,N_29221,N_29927);
xnor UO_1353 (O_1353,N_28776,N_28439);
nor UO_1354 (O_1354,N_29579,N_28134);
xnor UO_1355 (O_1355,N_28961,N_28259);
xor UO_1356 (O_1356,N_29909,N_29145);
nand UO_1357 (O_1357,N_28584,N_29857);
nand UO_1358 (O_1358,N_28808,N_29987);
nand UO_1359 (O_1359,N_29502,N_28317);
xnor UO_1360 (O_1360,N_28180,N_29008);
nand UO_1361 (O_1361,N_29601,N_29079);
nand UO_1362 (O_1362,N_28686,N_29100);
nand UO_1363 (O_1363,N_28664,N_29910);
nand UO_1364 (O_1364,N_29000,N_28335);
nor UO_1365 (O_1365,N_29726,N_29139);
or UO_1366 (O_1366,N_28528,N_28931);
nand UO_1367 (O_1367,N_28177,N_29700);
nand UO_1368 (O_1368,N_28230,N_29119);
nor UO_1369 (O_1369,N_29626,N_28408);
nor UO_1370 (O_1370,N_29765,N_28298);
nor UO_1371 (O_1371,N_29159,N_28158);
nand UO_1372 (O_1372,N_29292,N_29889);
and UO_1373 (O_1373,N_29589,N_28786);
and UO_1374 (O_1374,N_29339,N_28739);
or UO_1375 (O_1375,N_29258,N_29634);
nand UO_1376 (O_1376,N_29282,N_28512);
nand UO_1377 (O_1377,N_29744,N_29514);
nand UO_1378 (O_1378,N_28025,N_28377);
or UO_1379 (O_1379,N_28040,N_28297);
nor UO_1380 (O_1380,N_29852,N_29344);
nor UO_1381 (O_1381,N_29661,N_29105);
nand UO_1382 (O_1382,N_29093,N_28950);
and UO_1383 (O_1383,N_29314,N_29255);
and UO_1384 (O_1384,N_29132,N_28039);
xor UO_1385 (O_1385,N_28536,N_28023);
xnor UO_1386 (O_1386,N_29675,N_29397);
xor UO_1387 (O_1387,N_28001,N_29877);
and UO_1388 (O_1388,N_28676,N_28011);
nand UO_1389 (O_1389,N_29601,N_28347);
nand UO_1390 (O_1390,N_29174,N_28520);
and UO_1391 (O_1391,N_28889,N_29403);
nor UO_1392 (O_1392,N_28438,N_28392);
or UO_1393 (O_1393,N_28437,N_28281);
nand UO_1394 (O_1394,N_29642,N_29256);
nand UO_1395 (O_1395,N_29949,N_29507);
or UO_1396 (O_1396,N_28660,N_28547);
nand UO_1397 (O_1397,N_29120,N_28379);
nor UO_1398 (O_1398,N_29194,N_28691);
or UO_1399 (O_1399,N_29359,N_29533);
nand UO_1400 (O_1400,N_28856,N_28026);
nand UO_1401 (O_1401,N_29986,N_29622);
or UO_1402 (O_1402,N_28909,N_28106);
or UO_1403 (O_1403,N_29167,N_28744);
or UO_1404 (O_1404,N_28143,N_29581);
nor UO_1405 (O_1405,N_28795,N_28844);
nor UO_1406 (O_1406,N_28460,N_29879);
nor UO_1407 (O_1407,N_29627,N_29086);
xor UO_1408 (O_1408,N_28269,N_28070);
and UO_1409 (O_1409,N_28629,N_29740);
nand UO_1410 (O_1410,N_28171,N_28800);
nand UO_1411 (O_1411,N_29432,N_29649);
nor UO_1412 (O_1412,N_28403,N_28464);
xor UO_1413 (O_1413,N_28036,N_29011);
nand UO_1414 (O_1414,N_28750,N_29163);
or UO_1415 (O_1415,N_28035,N_29790);
or UO_1416 (O_1416,N_29561,N_29957);
nand UO_1417 (O_1417,N_29421,N_29971);
or UO_1418 (O_1418,N_28154,N_28365);
nand UO_1419 (O_1419,N_28719,N_28033);
xnor UO_1420 (O_1420,N_28957,N_28476);
nor UO_1421 (O_1421,N_28855,N_28474);
and UO_1422 (O_1422,N_29270,N_28342);
and UO_1423 (O_1423,N_28732,N_29258);
nor UO_1424 (O_1424,N_28773,N_29097);
nor UO_1425 (O_1425,N_28192,N_29620);
nand UO_1426 (O_1426,N_28803,N_29392);
or UO_1427 (O_1427,N_29498,N_29117);
nor UO_1428 (O_1428,N_29127,N_28799);
xor UO_1429 (O_1429,N_28316,N_28398);
xnor UO_1430 (O_1430,N_28835,N_29132);
nor UO_1431 (O_1431,N_29662,N_28612);
and UO_1432 (O_1432,N_28162,N_28237);
or UO_1433 (O_1433,N_29308,N_29069);
or UO_1434 (O_1434,N_28558,N_29249);
or UO_1435 (O_1435,N_29827,N_29629);
nor UO_1436 (O_1436,N_29995,N_28518);
or UO_1437 (O_1437,N_28116,N_29329);
or UO_1438 (O_1438,N_28577,N_29255);
nand UO_1439 (O_1439,N_29938,N_29339);
nand UO_1440 (O_1440,N_29918,N_28680);
nor UO_1441 (O_1441,N_29463,N_28299);
or UO_1442 (O_1442,N_28567,N_29186);
nor UO_1443 (O_1443,N_28291,N_29744);
nor UO_1444 (O_1444,N_28190,N_29964);
and UO_1445 (O_1445,N_28438,N_28002);
and UO_1446 (O_1446,N_28343,N_29843);
xor UO_1447 (O_1447,N_29264,N_29724);
xor UO_1448 (O_1448,N_28908,N_29745);
and UO_1449 (O_1449,N_29390,N_28677);
nand UO_1450 (O_1450,N_28894,N_28302);
xnor UO_1451 (O_1451,N_29393,N_28105);
or UO_1452 (O_1452,N_28327,N_28460);
xnor UO_1453 (O_1453,N_29419,N_28734);
xnor UO_1454 (O_1454,N_28844,N_28648);
nor UO_1455 (O_1455,N_29536,N_28845);
nand UO_1456 (O_1456,N_28854,N_29513);
and UO_1457 (O_1457,N_28720,N_28531);
nand UO_1458 (O_1458,N_28643,N_29100);
nor UO_1459 (O_1459,N_28826,N_29274);
nand UO_1460 (O_1460,N_28173,N_29100);
and UO_1461 (O_1461,N_28584,N_29698);
xnor UO_1462 (O_1462,N_28283,N_29366);
and UO_1463 (O_1463,N_28018,N_28014);
nor UO_1464 (O_1464,N_28611,N_28775);
nand UO_1465 (O_1465,N_29182,N_29188);
and UO_1466 (O_1466,N_29839,N_28210);
nor UO_1467 (O_1467,N_29158,N_29831);
nor UO_1468 (O_1468,N_29670,N_29458);
or UO_1469 (O_1469,N_29758,N_28315);
nor UO_1470 (O_1470,N_29969,N_29568);
xnor UO_1471 (O_1471,N_29073,N_29231);
nor UO_1472 (O_1472,N_28017,N_29414);
nor UO_1473 (O_1473,N_28581,N_28295);
xnor UO_1474 (O_1474,N_28214,N_29718);
or UO_1475 (O_1475,N_29362,N_28331);
xnor UO_1476 (O_1476,N_29884,N_28970);
nor UO_1477 (O_1477,N_28760,N_28995);
nor UO_1478 (O_1478,N_28122,N_29156);
and UO_1479 (O_1479,N_28532,N_29620);
nand UO_1480 (O_1480,N_29019,N_29633);
xnor UO_1481 (O_1481,N_29836,N_29760);
nor UO_1482 (O_1482,N_29660,N_29474);
nor UO_1483 (O_1483,N_29439,N_28167);
xor UO_1484 (O_1484,N_28366,N_28623);
and UO_1485 (O_1485,N_28844,N_29119);
nor UO_1486 (O_1486,N_28742,N_29323);
nor UO_1487 (O_1487,N_29782,N_29309);
and UO_1488 (O_1488,N_28679,N_29460);
nand UO_1489 (O_1489,N_29269,N_29827);
nor UO_1490 (O_1490,N_28029,N_29075);
xor UO_1491 (O_1491,N_28503,N_29236);
nor UO_1492 (O_1492,N_29692,N_28539);
nand UO_1493 (O_1493,N_28327,N_28206);
or UO_1494 (O_1494,N_29228,N_29391);
nand UO_1495 (O_1495,N_28624,N_29245);
nor UO_1496 (O_1496,N_29901,N_28888);
xor UO_1497 (O_1497,N_29820,N_29977);
xnor UO_1498 (O_1498,N_29977,N_28573);
and UO_1499 (O_1499,N_28969,N_29673);
nor UO_1500 (O_1500,N_29869,N_28411);
nand UO_1501 (O_1501,N_29477,N_29202);
xnor UO_1502 (O_1502,N_29988,N_28775);
and UO_1503 (O_1503,N_28136,N_29261);
or UO_1504 (O_1504,N_28369,N_28103);
and UO_1505 (O_1505,N_28815,N_28903);
xor UO_1506 (O_1506,N_29834,N_29564);
or UO_1507 (O_1507,N_28331,N_28138);
nand UO_1508 (O_1508,N_29643,N_28733);
nor UO_1509 (O_1509,N_29384,N_28030);
xnor UO_1510 (O_1510,N_29124,N_28420);
or UO_1511 (O_1511,N_28176,N_28340);
and UO_1512 (O_1512,N_28829,N_28543);
and UO_1513 (O_1513,N_28463,N_29361);
nor UO_1514 (O_1514,N_29806,N_29351);
nand UO_1515 (O_1515,N_29309,N_28382);
or UO_1516 (O_1516,N_29138,N_29337);
nor UO_1517 (O_1517,N_29434,N_29879);
xnor UO_1518 (O_1518,N_29516,N_29907);
xor UO_1519 (O_1519,N_28742,N_28496);
and UO_1520 (O_1520,N_29195,N_28810);
and UO_1521 (O_1521,N_29891,N_29501);
nand UO_1522 (O_1522,N_29932,N_29532);
or UO_1523 (O_1523,N_28896,N_29608);
nor UO_1524 (O_1524,N_28765,N_29071);
xor UO_1525 (O_1525,N_29174,N_29676);
nand UO_1526 (O_1526,N_28674,N_28829);
or UO_1527 (O_1527,N_28556,N_29388);
or UO_1528 (O_1528,N_29334,N_29658);
and UO_1529 (O_1529,N_28019,N_28664);
and UO_1530 (O_1530,N_28390,N_29738);
and UO_1531 (O_1531,N_28344,N_28270);
nor UO_1532 (O_1532,N_28618,N_28515);
nor UO_1533 (O_1533,N_28987,N_29971);
xnor UO_1534 (O_1534,N_28932,N_29615);
xor UO_1535 (O_1535,N_28049,N_29469);
or UO_1536 (O_1536,N_28407,N_29209);
nor UO_1537 (O_1537,N_29971,N_28532);
nor UO_1538 (O_1538,N_28730,N_28576);
nand UO_1539 (O_1539,N_28802,N_29857);
and UO_1540 (O_1540,N_28946,N_28128);
nand UO_1541 (O_1541,N_29568,N_29438);
nor UO_1542 (O_1542,N_28069,N_29032);
nand UO_1543 (O_1543,N_29033,N_29723);
nor UO_1544 (O_1544,N_29726,N_28435);
nand UO_1545 (O_1545,N_29159,N_29547);
nor UO_1546 (O_1546,N_28773,N_29944);
nand UO_1547 (O_1547,N_28242,N_28781);
nand UO_1548 (O_1548,N_29972,N_29187);
and UO_1549 (O_1549,N_28627,N_29633);
and UO_1550 (O_1550,N_28278,N_28130);
nand UO_1551 (O_1551,N_28094,N_29630);
nor UO_1552 (O_1552,N_28148,N_29428);
and UO_1553 (O_1553,N_28897,N_29005);
nand UO_1554 (O_1554,N_29402,N_28737);
xor UO_1555 (O_1555,N_28862,N_28955);
xnor UO_1556 (O_1556,N_28179,N_28802);
xor UO_1557 (O_1557,N_28334,N_28188);
xnor UO_1558 (O_1558,N_28498,N_29232);
and UO_1559 (O_1559,N_29454,N_28030);
nor UO_1560 (O_1560,N_29153,N_28588);
nand UO_1561 (O_1561,N_28259,N_29725);
nand UO_1562 (O_1562,N_28059,N_28286);
or UO_1563 (O_1563,N_28047,N_28034);
and UO_1564 (O_1564,N_29523,N_29446);
or UO_1565 (O_1565,N_28990,N_29046);
nor UO_1566 (O_1566,N_28550,N_28725);
nand UO_1567 (O_1567,N_29285,N_29411);
nand UO_1568 (O_1568,N_28997,N_28621);
or UO_1569 (O_1569,N_28518,N_29303);
nand UO_1570 (O_1570,N_29387,N_29606);
nor UO_1571 (O_1571,N_28830,N_29498);
nor UO_1572 (O_1572,N_29940,N_28077);
xor UO_1573 (O_1573,N_29731,N_29203);
or UO_1574 (O_1574,N_28267,N_28367);
and UO_1575 (O_1575,N_29334,N_29861);
or UO_1576 (O_1576,N_28662,N_28817);
nor UO_1577 (O_1577,N_28952,N_28423);
and UO_1578 (O_1578,N_29078,N_29568);
or UO_1579 (O_1579,N_29699,N_29922);
xor UO_1580 (O_1580,N_28570,N_29000);
nand UO_1581 (O_1581,N_28469,N_29284);
nand UO_1582 (O_1582,N_29931,N_28184);
nor UO_1583 (O_1583,N_28392,N_28214);
nor UO_1584 (O_1584,N_28475,N_29153);
xnor UO_1585 (O_1585,N_29739,N_29722);
and UO_1586 (O_1586,N_29173,N_28709);
xnor UO_1587 (O_1587,N_28175,N_29569);
nand UO_1588 (O_1588,N_29386,N_29328);
or UO_1589 (O_1589,N_28904,N_29939);
or UO_1590 (O_1590,N_28930,N_29871);
nand UO_1591 (O_1591,N_28777,N_29845);
xor UO_1592 (O_1592,N_28371,N_29024);
or UO_1593 (O_1593,N_29827,N_28053);
nand UO_1594 (O_1594,N_28223,N_29322);
nor UO_1595 (O_1595,N_29577,N_29218);
nor UO_1596 (O_1596,N_28855,N_29436);
nor UO_1597 (O_1597,N_29067,N_28064);
and UO_1598 (O_1598,N_28699,N_29596);
or UO_1599 (O_1599,N_28989,N_29451);
nand UO_1600 (O_1600,N_29262,N_28265);
nand UO_1601 (O_1601,N_29789,N_28810);
xnor UO_1602 (O_1602,N_28804,N_28471);
nand UO_1603 (O_1603,N_28408,N_28368);
nand UO_1604 (O_1604,N_29308,N_28136);
and UO_1605 (O_1605,N_29235,N_28643);
or UO_1606 (O_1606,N_29281,N_29674);
nor UO_1607 (O_1607,N_29055,N_28140);
xor UO_1608 (O_1608,N_29428,N_29902);
or UO_1609 (O_1609,N_28032,N_29432);
xor UO_1610 (O_1610,N_29888,N_29218);
nand UO_1611 (O_1611,N_28089,N_29273);
nand UO_1612 (O_1612,N_29681,N_28607);
nand UO_1613 (O_1613,N_29844,N_28121);
nand UO_1614 (O_1614,N_29625,N_29280);
xnor UO_1615 (O_1615,N_29022,N_29602);
nand UO_1616 (O_1616,N_29251,N_29932);
and UO_1617 (O_1617,N_28879,N_28573);
nor UO_1618 (O_1618,N_28169,N_28523);
or UO_1619 (O_1619,N_29632,N_29830);
and UO_1620 (O_1620,N_29259,N_28384);
xnor UO_1621 (O_1621,N_28256,N_29185);
nand UO_1622 (O_1622,N_28826,N_28368);
and UO_1623 (O_1623,N_28061,N_28845);
xor UO_1624 (O_1624,N_28980,N_28265);
and UO_1625 (O_1625,N_28446,N_29190);
nand UO_1626 (O_1626,N_28943,N_28197);
nand UO_1627 (O_1627,N_29347,N_29095);
xor UO_1628 (O_1628,N_28440,N_29825);
xor UO_1629 (O_1629,N_29160,N_28418);
nand UO_1630 (O_1630,N_29842,N_29457);
nor UO_1631 (O_1631,N_29203,N_28084);
or UO_1632 (O_1632,N_29654,N_29852);
or UO_1633 (O_1633,N_28466,N_28065);
xor UO_1634 (O_1634,N_28331,N_28776);
xnor UO_1635 (O_1635,N_29529,N_29057);
xnor UO_1636 (O_1636,N_28955,N_28303);
xnor UO_1637 (O_1637,N_29329,N_28936);
nand UO_1638 (O_1638,N_28316,N_29157);
nand UO_1639 (O_1639,N_29222,N_28627);
nand UO_1640 (O_1640,N_29457,N_29875);
or UO_1641 (O_1641,N_29108,N_29565);
xor UO_1642 (O_1642,N_29394,N_28317);
xor UO_1643 (O_1643,N_28607,N_28078);
or UO_1644 (O_1644,N_28542,N_29554);
and UO_1645 (O_1645,N_28195,N_28603);
xnor UO_1646 (O_1646,N_29870,N_29596);
xor UO_1647 (O_1647,N_28233,N_28097);
and UO_1648 (O_1648,N_29313,N_29098);
nand UO_1649 (O_1649,N_29422,N_28289);
xnor UO_1650 (O_1650,N_29188,N_29464);
nand UO_1651 (O_1651,N_28131,N_28503);
xnor UO_1652 (O_1652,N_29023,N_28805);
or UO_1653 (O_1653,N_29246,N_29387);
nor UO_1654 (O_1654,N_29557,N_28901);
and UO_1655 (O_1655,N_28061,N_29500);
nor UO_1656 (O_1656,N_29106,N_29362);
and UO_1657 (O_1657,N_28600,N_29726);
or UO_1658 (O_1658,N_29369,N_28318);
xnor UO_1659 (O_1659,N_28729,N_29691);
and UO_1660 (O_1660,N_29916,N_28052);
and UO_1661 (O_1661,N_29215,N_28358);
nor UO_1662 (O_1662,N_28943,N_29115);
or UO_1663 (O_1663,N_29676,N_29307);
and UO_1664 (O_1664,N_29186,N_28580);
nor UO_1665 (O_1665,N_28318,N_29845);
xnor UO_1666 (O_1666,N_29935,N_28463);
and UO_1667 (O_1667,N_28192,N_29830);
xnor UO_1668 (O_1668,N_29156,N_29144);
or UO_1669 (O_1669,N_29199,N_29423);
nor UO_1670 (O_1670,N_28327,N_28254);
nand UO_1671 (O_1671,N_29656,N_28067);
nand UO_1672 (O_1672,N_29041,N_28396);
or UO_1673 (O_1673,N_29121,N_29444);
xnor UO_1674 (O_1674,N_29012,N_29965);
and UO_1675 (O_1675,N_28001,N_28348);
xnor UO_1676 (O_1676,N_29846,N_29324);
xnor UO_1677 (O_1677,N_29367,N_29617);
nand UO_1678 (O_1678,N_29745,N_28929);
or UO_1679 (O_1679,N_28366,N_29929);
nand UO_1680 (O_1680,N_28469,N_28063);
nor UO_1681 (O_1681,N_28466,N_29793);
or UO_1682 (O_1682,N_29013,N_29315);
xnor UO_1683 (O_1683,N_29660,N_29624);
and UO_1684 (O_1684,N_28756,N_29197);
or UO_1685 (O_1685,N_29233,N_28057);
nand UO_1686 (O_1686,N_29801,N_28634);
and UO_1687 (O_1687,N_28048,N_29960);
or UO_1688 (O_1688,N_29166,N_28656);
nand UO_1689 (O_1689,N_28453,N_28009);
nor UO_1690 (O_1690,N_28901,N_28302);
xnor UO_1691 (O_1691,N_29816,N_29804);
and UO_1692 (O_1692,N_29892,N_29289);
nor UO_1693 (O_1693,N_28273,N_29636);
and UO_1694 (O_1694,N_28160,N_28939);
nor UO_1695 (O_1695,N_28586,N_28922);
xor UO_1696 (O_1696,N_29761,N_29317);
and UO_1697 (O_1697,N_29941,N_29593);
xnor UO_1698 (O_1698,N_29875,N_29453);
nand UO_1699 (O_1699,N_29202,N_28119);
nand UO_1700 (O_1700,N_28500,N_28035);
nor UO_1701 (O_1701,N_28934,N_28239);
or UO_1702 (O_1702,N_29655,N_28530);
nor UO_1703 (O_1703,N_28818,N_28418);
and UO_1704 (O_1704,N_28685,N_28325);
and UO_1705 (O_1705,N_28184,N_28254);
or UO_1706 (O_1706,N_28221,N_28714);
and UO_1707 (O_1707,N_28001,N_28610);
or UO_1708 (O_1708,N_28470,N_28135);
xnor UO_1709 (O_1709,N_28706,N_29265);
and UO_1710 (O_1710,N_28830,N_28216);
xor UO_1711 (O_1711,N_29111,N_29778);
nor UO_1712 (O_1712,N_29351,N_29133);
and UO_1713 (O_1713,N_28167,N_28922);
nor UO_1714 (O_1714,N_29285,N_29933);
xor UO_1715 (O_1715,N_29650,N_28489);
xnor UO_1716 (O_1716,N_28465,N_29493);
nand UO_1717 (O_1717,N_28041,N_29563);
nor UO_1718 (O_1718,N_29593,N_29838);
or UO_1719 (O_1719,N_29077,N_29717);
or UO_1720 (O_1720,N_29038,N_29814);
or UO_1721 (O_1721,N_29600,N_28748);
nor UO_1722 (O_1722,N_29128,N_29204);
nor UO_1723 (O_1723,N_29317,N_29415);
or UO_1724 (O_1724,N_29804,N_28163);
nor UO_1725 (O_1725,N_28052,N_29341);
and UO_1726 (O_1726,N_29189,N_29500);
xor UO_1727 (O_1727,N_28258,N_29669);
and UO_1728 (O_1728,N_29637,N_29932);
or UO_1729 (O_1729,N_29695,N_28202);
nor UO_1730 (O_1730,N_28443,N_28695);
and UO_1731 (O_1731,N_29767,N_28274);
nor UO_1732 (O_1732,N_28173,N_29022);
and UO_1733 (O_1733,N_29586,N_29843);
or UO_1734 (O_1734,N_29353,N_29792);
nand UO_1735 (O_1735,N_28681,N_29998);
or UO_1736 (O_1736,N_28748,N_29807);
nor UO_1737 (O_1737,N_29439,N_28513);
nor UO_1738 (O_1738,N_29688,N_28042);
nand UO_1739 (O_1739,N_29321,N_29052);
nand UO_1740 (O_1740,N_29916,N_28028);
and UO_1741 (O_1741,N_28487,N_29052);
nand UO_1742 (O_1742,N_29685,N_29668);
xnor UO_1743 (O_1743,N_28766,N_29624);
xor UO_1744 (O_1744,N_28275,N_29975);
nor UO_1745 (O_1745,N_28925,N_29608);
xor UO_1746 (O_1746,N_28033,N_28595);
nor UO_1747 (O_1747,N_28615,N_29930);
nor UO_1748 (O_1748,N_28239,N_28893);
nand UO_1749 (O_1749,N_29322,N_29041);
and UO_1750 (O_1750,N_29638,N_29922);
nor UO_1751 (O_1751,N_29648,N_29838);
and UO_1752 (O_1752,N_28275,N_28304);
or UO_1753 (O_1753,N_28782,N_28155);
and UO_1754 (O_1754,N_29064,N_29494);
xor UO_1755 (O_1755,N_28902,N_29393);
nor UO_1756 (O_1756,N_29530,N_28629);
nand UO_1757 (O_1757,N_29448,N_28044);
nand UO_1758 (O_1758,N_28222,N_28036);
nor UO_1759 (O_1759,N_28774,N_28132);
or UO_1760 (O_1760,N_29430,N_29294);
nor UO_1761 (O_1761,N_29524,N_29995);
nand UO_1762 (O_1762,N_29442,N_29672);
nand UO_1763 (O_1763,N_28371,N_29799);
nand UO_1764 (O_1764,N_29596,N_29180);
and UO_1765 (O_1765,N_28979,N_28233);
and UO_1766 (O_1766,N_28471,N_29888);
nand UO_1767 (O_1767,N_29367,N_29105);
or UO_1768 (O_1768,N_29917,N_28953);
or UO_1769 (O_1769,N_29123,N_28202);
nand UO_1770 (O_1770,N_28426,N_28148);
and UO_1771 (O_1771,N_28259,N_29945);
nor UO_1772 (O_1772,N_29915,N_28898);
xnor UO_1773 (O_1773,N_29803,N_28250);
nor UO_1774 (O_1774,N_29611,N_29746);
and UO_1775 (O_1775,N_29307,N_28603);
and UO_1776 (O_1776,N_29974,N_28984);
nand UO_1777 (O_1777,N_29068,N_29962);
xor UO_1778 (O_1778,N_29362,N_29814);
nor UO_1779 (O_1779,N_28520,N_29076);
nand UO_1780 (O_1780,N_28544,N_28374);
nor UO_1781 (O_1781,N_28994,N_28278);
xor UO_1782 (O_1782,N_28574,N_29344);
xor UO_1783 (O_1783,N_28103,N_28568);
xnor UO_1784 (O_1784,N_28958,N_29311);
or UO_1785 (O_1785,N_28888,N_29541);
nor UO_1786 (O_1786,N_28247,N_29128);
and UO_1787 (O_1787,N_28090,N_28244);
or UO_1788 (O_1788,N_28219,N_28238);
xnor UO_1789 (O_1789,N_29924,N_28985);
xnor UO_1790 (O_1790,N_29416,N_28285);
xor UO_1791 (O_1791,N_28633,N_28614);
xnor UO_1792 (O_1792,N_29294,N_28176);
or UO_1793 (O_1793,N_28162,N_28108);
or UO_1794 (O_1794,N_29533,N_29304);
nand UO_1795 (O_1795,N_29458,N_28876);
and UO_1796 (O_1796,N_29975,N_28610);
or UO_1797 (O_1797,N_29402,N_29932);
xor UO_1798 (O_1798,N_28727,N_29410);
and UO_1799 (O_1799,N_29222,N_29410);
nor UO_1800 (O_1800,N_29875,N_29300);
nor UO_1801 (O_1801,N_29681,N_29402);
and UO_1802 (O_1802,N_29847,N_29514);
xor UO_1803 (O_1803,N_28712,N_29754);
or UO_1804 (O_1804,N_28931,N_28231);
nor UO_1805 (O_1805,N_28246,N_28902);
xnor UO_1806 (O_1806,N_29018,N_28517);
or UO_1807 (O_1807,N_29437,N_28857);
nor UO_1808 (O_1808,N_28988,N_28320);
xnor UO_1809 (O_1809,N_28118,N_28935);
or UO_1810 (O_1810,N_28029,N_29035);
and UO_1811 (O_1811,N_28322,N_28284);
or UO_1812 (O_1812,N_28095,N_29233);
and UO_1813 (O_1813,N_28339,N_28074);
nand UO_1814 (O_1814,N_28933,N_28983);
nor UO_1815 (O_1815,N_28223,N_29156);
nor UO_1816 (O_1816,N_29953,N_28083);
nor UO_1817 (O_1817,N_28190,N_28067);
xor UO_1818 (O_1818,N_28299,N_29016);
xor UO_1819 (O_1819,N_28470,N_28633);
nor UO_1820 (O_1820,N_28058,N_29343);
nor UO_1821 (O_1821,N_29125,N_28985);
nor UO_1822 (O_1822,N_29138,N_29633);
xor UO_1823 (O_1823,N_28005,N_29789);
nand UO_1824 (O_1824,N_29630,N_28724);
and UO_1825 (O_1825,N_28717,N_28188);
or UO_1826 (O_1826,N_28301,N_28490);
nand UO_1827 (O_1827,N_28692,N_28555);
xor UO_1828 (O_1828,N_28849,N_29467);
nor UO_1829 (O_1829,N_28859,N_28269);
nand UO_1830 (O_1830,N_28320,N_29888);
or UO_1831 (O_1831,N_28774,N_29575);
nand UO_1832 (O_1832,N_28580,N_29620);
and UO_1833 (O_1833,N_29629,N_28333);
or UO_1834 (O_1834,N_28180,N_29247);
nor UO_1835 (O_1835,N_28558,N_29890);
and UO_1836 (O_1836,N_29354,N_29884);
nor UO_1837 (O_1837,N_28499,N_29172);
nor UO_1838 (O_1838,N_28809,N_29339);
or UO_1839 (O_1839,N_29323,N_28973);
or UO_1840 (O_1840,N_28395,N_29161);
and UO_1841 (O_1841,N_28385,N_28010);
xnor UO_1842 (O_1842,N_28303,N_28062);
nor UO_1843 (O_1843,N_28906,N_29672);
or UO_1844 (O_1844,N_28188,N_29394);
nand UO_1845 (O_1845,N_29083,N_29379);
and UO_1846 (O_1846,N_28633,N_29486);
nor UO_1847 (O_1847,N_28190,N_29342);
xor UO_1848 (O_1848,N_28689,N_29285);
and UO_1849 (O_1849,N_28560,N_28768);
or UO_1850 (O_1850,N_29378,N_29561);
and UO_1851 (O_1851,N_29298,N_29753);
or UO_1852 (O_1852,N_29860,N_29448);
and UO_1853 (O_1853,N_28064,N_29670);
and UO_1854 (O_1854,N_29979,N_29571);
or UO_1855 (O_1855,N_28992,N_28350);
and UO_1856 (O_1856,N_28939,N_28349);
xnor UO_1857 (O_1857,N_28636,N_29580);
or UO_1858 (O_1858,N_28539,N_28030);
nand UO_1859 (O_1859,N_28119,N_29701);
or UO_1860 (O_1860,N_29269,N_29099);
or UO_1861 (O_1861,N_28878,N_28390);
nor UO_1862 (O_1862,N_29774,N_28359);
or UO_1863 (O_1863,N_29299,N_28938);
and UO_1864 (O_1864,N_29518,N_28987);
nor UO_1865 (O_1865,N_29856,N_29413);
and UO_1866 (O_1866,N_28353,N_29455);
xnor UO_1867 (O_1867,N_29899,N_29762);
and UO_1868 (O_1868,N_29876,N_29589);
or UO_1869 (O_1869,N_28353,N_28779);
or UO_1870 (O_1870,N_28509,N_28577);
nand UO_1871 (O_1871,N_29799,N_29182);
nand UO_1872 (O_1872,N_29208,N_28574);
xor UO_1873 (O_1873,N_29334,N_29464);
xnor UO_1874 (O_1874,N_28428,N_28052);
xnor UO_1875 (O_1875,N_28667,N_29671);
xor UO_1876 (O_1876,N_28640,N_29872);
nand UO_1877 (O_1877,N_29222,N_28880);
nand UO_1878 (O_1878,N_29265,N_28194);
or UO_1879 (O_1879,N_29067,N_28183);
xnor UO_1880 (O_1880,N_29633,N_28054);
and UO_1881 (O_1881,N_28831,N_29859);
nand UO_1882 (O_1882,N_29555,N_29508);
xnor UO_1883 (O_1883,N_28724,N_28013);
or UO_1884 (O_1884,N_28075,N_28341);
and UO_1885 (O_1885,N_28182,N_29084);
nand UO_1886 (O_1886,N_28630,N_28575);
nor UO_1887 (O_1887,N_29102,N_28579);
nand UO_1888 (O_1888,N_29017,N_29824);
and UO_1889 (O_1889,N_28887,N_28827);
nand UO_1890 (O_1890,N_28271,N_28353);
and UO_1891 (O_1891,N_28344,N_28196);
nor UO_1892 (O_1892,N_28624,N_28400);
xor UO_1893 (O_1893,N_29164,N_28672);
nand UO_1894 (O_1894,N_28614,N_28748);
nand UO_1895 (O_1895,N_28524,N_29772);
nand UO_1896 (O_1896,N_29319,N_28666);
nand UO_1897 (O_1897,N_29801,N_28886);
xnor UO_1898 (O_1898,N_28261,N_29010);
nand UO_1899 (O_1899,N_28920,N_29282);
and UO_1900 (O_1900,N_28215,N_28134);
xor UO_1901 (O_1901,N_29923,N_28054);
xor UO_1902 (O_1902,N_28161,N_28519);
or UO_1903 (O_1903,N_28176,N_29347);
nand UO_1904 (O_1904,N_28557,N_28498);
or UO_1905 (O_1905,N_29049,N_29829);
nand UO_1906 (O_1906,N_29113,N_28100);
nor UO_1907 (O_1907,N_28867,N_29285);
nor UO_1908 (O_1908,N_28459,N_29658);
nor UO_1909 (O_1909,N_29562,N_28672);
nor UO_1910 (O_1910,N_29221,N_29822);
and UO_1911 (O_1911,N_28928,N_28001);
and UO_1912 (O_1912,N_29281,N_28431);
nand UO_1913 (O_1913,N_28081,N_29429);
or UO_1914 (O_1914,N_28391,N_29710);
or UO_1915 (O_1915,N_29815,N_28146);
xor UO_1916 (O_1916,N_29915,N_29693);
nand UO_1917 (O_1917,N_29668,N_29265);
xor UO_1918 (O_1918,N_28600,N_29570);
nor UO_1919 (O_1919,N_29931,N_28824);
nor UO_1920 (O_1920,N_28071,N_28275);
and UO_1921 (O_1921,N_29854,N_28450);
xnor UO_1922 (O_1922,N_29149,N_28937);
xnor UO_1923 (O_1923,N_28060,N_29836);
nand UO_1924 (O_1924,N_29212,N_28746);
nor UO_1925 (O_1925,N_28173,N_28283);
nor UO_1926 (O_1926,N_28534,N_28329);
nor UO_1927 (O_1927,N_28237,N_28873);
xor UO_1928 (O_1928,N_29316,N_28411);
and UO_1929 (O_1929,N_28725,N_28315);
nor UO_1930 (O_1930,N_29832,N_28779);
and UO_1931 (O_1931,N_28316,N_29411);
nor UO_1932 (O_1932,N_28393,N_29956);
or UO_1933 (O_1933,N_28133,N_28134);
nor UO_1934 (O_1934,N_29980,N_29886);
or UO_1935 (O_1935,N_29067,N_29352);
nand UO_1936 (O_1936,N_28077,N_28369);
and UO_1937 (O_1937,N_28503,N_28321);
or UO_1938 (O_1938,N_28376,N_28664);
and UO_1939 (O_1939,N_29916,N_29804);
and UO_1940 (O_1940,N_28760,N_29221);
xnor UO_1941 (O_1941,N_28223,N_28258);
xnor UO_1942 (O_1942,N_28610,N_28467);
nand UO_1943 (O_1943,N_28265,N_28098);
nor UO_1944 (O_1944,N_28399,N_28516);
nor UO_1945 (O_1945,N_28529,N_29314);
xnor UO_1946 (O_1946,N_29742,N_29546);
nor UO_1947 (O_1947,N_29537,N_29006);
xor UO_1948 (O_1948,N_28447,N_29579);
xor UO_1949 (O_1949,N_29328,N_28774);
or UO_1950 (O_1950,N_29988,N_29018);
or UO_1951 (O_1951,N_28887,N_29156);
xnor UO_1952 (O_1952,N_28877,N_29375);
nand UO_1953 (O_1953,N_29951,N_29921);
xnor UO_1954 (O_1954,N_29287,N_29759);
nor UO_1955 (O_1955,N_29599,N_29918);
xor UO_1956 (O_1956,N_29898,N_28558);
xor UO_1957 (O_1957,N_29547,N_28130);
nor UO_1958 (O_1958,N_29258,N_29661);
or UO_1959 (O_1959,N_29250,N_29288);
xnor UO_1960 (O_1960,N_28334,N_29455);
and UO_1961 (O_1961,N_29429,N_29390);
and UO_1962 (O_1962,N_29878,N_29327);
xnor UO_1963 (O_1963,N_29568,N_28072);
and UO_1964 (O_1964,N_29293,N_29865);
nor UO_1965 (O_1965,N_29262,N_29834);
nand UO_1966 (O_1966,N_28003,N_29337);
nand UO_1967 (O_1967,N_29824,N_28593);
and UO_1968 (O_1968,N_29367,N_28519);
or UO_1969 (O_1969,N_29948,N_28924);
nor UO_1970 (O_1970,N_28282,N_29715);
nor UO_1971 (O_1971,N_29612,N_28820);
xnor UO_1972 (O_1972,N_29690,N_28562);
and UO_1973 (O_1973,N_29276,N_29809);
nand UO_1974 (O_1974,N_28915,N_29965);
nand UO_1975 (O_1975,N_28460,N_28635);
nand UO_1976 (O_1976,N_29185,N_28069);
nand UO_1977 (O_1977,N_28433,N_28243);
and UO_1978 (O_1978,N_29319,N_29863);
nor UO_1979 (O_1979,N_28392,N_28633);
or UO_1980 (O_1980,N_29486,N_28671);
nor UO_1981 (O_1981,N_28147,N_29083);
and UO_1982 (O_1982,N_28497,N_28105);
xor UO_1983 (O_1983,N_28313,N_29420);
nand UO_1984 (O_1984,N_29607,N_29377);
and UO_1985 (O_1985,N_29339,N_28518);
and UO_1986 (O_1986,N_29964,N_28894);
and UO_1987 (O_1987,N_28522,N_29937);
and UO_1988 (O_1988,N_28966,N_28985);
xnor UO_1989 (O_1989,N_28696,N_28848);
or UO_1990 (O_1990,N_29566,N_28111);
and UO_1991 (O_1991,N_28515,N_29434);
xor UO_1992 (O_1992,N_28687,N_28319);
xnor UO_1993 (O_1993,N_29007,N_29450);
and UO_1994 (O_1994,N_28624,N_29111);
and UO_1995 (O_1995,N_29285,N_28787);
or UO_1996 (O_1996,N_29143,N_29217);
xor UO_1997 (O_1997,N_29049,N_28417);
and UO_1998 (O_1998,N_29134,N_29881);
xnor UO_1999 (O_1999,N_29105,N_29581);
nor UO_2000 (O_2000,N_29223,N_29862);
nand UO_2001 (O_2001,N_29515,N_28774);
nor UO_2002 (O_2002,N_28681,N_28165);
nor UO_2003 (O_2003,N_29192,N_29323);
xnor UO_2004 (O_2004,N_29547,N_28226);
nand UO_2005 (O_2005,N_29496,N_28087);
nand UO_2006 (O_2006,N_28520,N_29793);
or UO_2007 (O_2007,N_29367,N_29038);
nand UO_2008 (O_2008,N_28811,N_29680);
nor UO_2009 (O_2009,N_28306,N_28772);
nor UO_2010 (O_2010,N_28310,N_28627);
or UO_2011 (O_2011,N_29854,N_28026);
xor UO_2012 (O_2012,N_28870,N_29257);
or UO_2013 (O_2013,N_28208,N_29794);
and UO_2014 (O_2014,N_28745,N_29025);
nor UO_2015 (O_2015,N_28583,N_29613);
nand UO_2016 (O_2016,N_29225,N_29377);
nor UO_2017 (O_2017,N_28288,N_28836);
or UO_2018 (O_2018,N_29077,N_28194);
nor UO_2019 (O_2019,N_28995,N_28392);
nand UO_2020 (O_2020,N_28185,N_29489);
nor UO_2021 (O_2021,N_28638,N_28139);
and UO_2022 (O_2022,N_28714,N_29600);
and UO_2023 (O_2023,N_29804,N_29609);
nand UO_2024 (O_2024,N_29849,N_28824);
xnor UO_2025 (O_2025,N_28173,N_28233);
xnor UO_2026 (O_2026,N_28739,N_28622);
nand UO_2027 (O_2027,N_29597,N_29307);
or UO_2028 (O_2028,N_28780,N_28948);
and UO_2029 (O_2029,N_29169,N_28174);
nand UO_2030 (O_2030,N_29064,N_29635);
and UO_2031 (O_2031,N_29887,N_29967);
xnor UO_2032 (O_2032,N_28399,N_29806);
nor UO_2033 (O_2033,N_29702,N_28181);
or UO_2034 (O_2034,N_28350,N_29178);
xor UO_2035 (O_2035,N_29619,N_28507);
or UO_2036 (O_2036,N_28524,N_29412);
and UO_2037 (O_2037,N_29252,N_29477);
or UO_2038 (O_2038,N_28184,N_29936);
xor UO_2039 (O_2039,N_29648,N_29626);
or UO_2040 (O_2040,N_29428,N_28019);
and UO_2041 (O_2041,N_29204,N_28545);
nor UO_2042 (O_2042,N_28060,N_29448);
or UO_2043 (O_2043,N_29781,N_29010);
nand UO_2044 (O_2044,N_28864,N_28812);
xor UO_2045 (O_2045,N_29605,N_29257);
xnor UO_2046 (O_2046,N_28770,N_29780);
and UO_2047 (O_2047,N_29568,N_29385);
nand UO_2048 (O_2048,N_29573,N_28898);
nand UO_2049 (O_2049,N_28317,N_28084);
xnor UO_2050 (O_2050,N_28289,N_29405);
xor UO_2051 (O_2051,N_29731,N_28291);
nor UO_2052 (O_2052,N_29126,N_29195);
or UO_2053 (O_2053,N_28390,N_28836);
nor UO_2054 (O_2054,N_29979,N_28046);
nand UO_2055 (O_2055,N_29706,N_29430);
xor UO_2056 (O_2056,N_28711,N_29387);
xor UO_2057 (O_2057,N_28281,N_29263);
and UO_2058 (O_2058,N_29169,N_28859);
and UO_2059 (O_2059,N_28394,N_29718);
xnor UO_2060 (O_2060,N_28660,N_28919);
xnor UO_2061 (O_2061,N_29539,N_29788);
nand UO_2062 (O_2062,N_28839,N_29297);
nor UO_2063 (O_2063,N_29397,N_28457);
xnor UO_2064 (O_2064,N_28250,N_29514);
nand UO_2065 (O_2065,N_29152,N_28111);
or UO_2066 (O_2066,N_29713,N_29347);
or UO_2067 (O_2067,N_28253,N_29963);
and UO_2068 (O_2068,N_28280,N_28737);
xor UO_2069 (O_2069,N_29455,N_28317);
and UO_2070 (O_2070,N_29419,N_29334);
and UO_2071 (O_2071,N_29758,N_28600);
or UO_2072 (O_2072,N_28990,N_28943);
nor UO_2073 (O_2073,N_29220,N_28598);
and UO_2074 (O_2074,N_28550,N_29000);
and UO_2075 (O_2075,N_29784,N_29177);
xnor UO_2076 (O_2076,N_29894,N_28134);
and UO_2077 (O_2077,N_28468,N_28893);
nand UO_2078 (O_2078,N_28400,N_29905);
nor UO_2079 (O_2079,N_28433,N_28291);
or UO_2080 (O_2080,N_29587,N_28870);
nor UO_2081 (O_2081,N_28052,N_28230);
or UO_2082 (O_2082,N_29061,N_29374);
and UO_2083 (O_2083,N_29946,N_29277);
nor UO_2084 (O_2084,N_29399,N_29539);
or UO_2085 (O_2085,N_29760,N_28427);
nor UO_2086 (O_2086,N_28592,N_28702);
nand UO_2087 (O_2087,N_29775,N_29924);
nand UO_2088 (O_2088,N_28820,N_28849);
or UO_2089 (O_2089,N_28238,N_28798);
or UO_2090 (O_2090,N_29836,N_28863);
nand UO_2091 (O_2091,N_29884,N_28994);
or UO_2092 (O_2092,N_28253,N_28923);
xor UO_2093 (O_2093,N_28874,N_29823);
or UO_2094 (O_2094,N_29793,N_29529);
or UO_2095 (O_2095,N_29212,N_28491);
xor UO_2096 (O_2096,N_28731,N_29980);
and UO_2097 (O_2097,N_29481,N_29173);
and UO_2098 (O_2098,N_28972,N_29836);
nand UO_2099 (O_2099,N_29417,N_29271);
and UO_2100 (O_2100,N_28716,N_29948);
xnor UO_2101 (O_2101,N_28586,N_28460);
or UO_2102 (O_2102,N_29606,N_28258);
nand UO_2103 (O_2103,N_28821,N_28757);
and UO_2104 (O_2104,N_29309,N_29678);
nor UO_2105 (O_2105,N_28584,N_28155);
or UO_2106 (O_2106,N_29074,N_28877);
or UO_2107 (O_2107,N_29109,N_28474);
and UO_2108 (O_2108,N_29195,N_29617);
nand UO_2109 (O_2109,N_29658,N_28259);
and UO_2110 (O_2110,N_28802,N_29597);
nor UO_2111 (O_2111,N_28982,N_29279);
nand UO_2112 (O_2112,N_29187,N_29539);
nor UO_2113 (O_2113,N_28690,N_29905);
xor UO_2114 (O_2114,N_29130,N_29587);
xor UO_2115 (O_2115,N_28828,N_29485);
xnor UO_2116 (O_2116,N_28670,N_29949);
xnor UO_2117 (O_2117,N_29756,N_29729);
and UO_2118 (O_2118,N_29188,N_28445);
or UO_2119 (O_2119,N_28677,N_29543);
xor UO_2120 (O_2120,N_29612,N_28817);
nand UO_2121 (O_2121,N_28817,N_28984);
and UO_2122 (O_2122,N_29830,N_28755);
or UO_2123 (O_2123,N_29329,N_28719);
nand UO_2124 (O_2124,N_29249,N_29786);
or UO_2125 (O_2125,N_29887,N_28701);
nand UO_2126 (O_2126,N_29240,N_29538);
nand UO_2127 (O_2127,N_29446,N_29350);
or UO_2128 (O_2128,N_28922,N_28874);
and UO_2129 (O_2129,N_28732,N_29201);
and UO_2130 (O_2130,N_28089,N_29533);
xnor UO_2131 (O_2131,N_28980,N_28565);
or UO_2132 (O_2132,N_29975,N_29259);
nor UO_2133 (O_2133,N_29189,N_28411);
and UO_2134 (O_2134,N_29897,N_28341);
and UO_2135 (O_2135,N_29508,N_28418);
and UO_2136 (O_2136,N_29448,N_29036);
nand UO_2137 (O_2137,N_28479,N_28085);
xnor UO_2138 (O_2138,N_28826,N_28659);
nand UO_2139 (O_2139,N_29751,N_28211);
or UO_2140 (O_2140,N_29008,N_28296);
xor UO_2141 (O_2141,N_29744,N_29028);
nor UO_2142 (O_2142,N_28327,N_29009);
xnor UO_2143 (O_2143,N_28259,N_29501);
nor UO_2144 (O_2144,N_28018,N_29103);
nor UO_2145 (O_2145,N_28239,N_28548);
nor UO_2146 (O_2146,N_28365,N_29046);
or UO_2147 (O_2147,N_28958,N_28154);
or UO_2148 (O_2148,N_28438,N_28449);
and UO_2149 (O_2149,N_28915,N_29041);
nand UO_2150 (O_2150,N_29832,N_29288);
or UO_2151 (O_2151,N_28137,N_28290);
or UO_2152 (O_2152,N_28420,N_29859);
xor UO_2153 (O_2153,N_28004,N_28417);
nor UO_2154 (O_2154,N_28495,N_28472);
nor UO_2155 (O_2155,N_28270,N_28213);
nand UO_2156 (O_2156,N_29240,N_29152);
or UO_2157 (O_2157,N_28164,N_28566);
xnor UO_2158 (O_2158,N_29492,N_29743);
xnor UO_2159 (O_2159,N_28231,N_28550);
nand UO_2160 (O_2160,N_28768,N_28710);
nor UO_2161 (O_2161,N_29226,N_29409);
xnor UO_2162 (O_2162,N_28273,N_29148);
xnor UO_2163 (O_2163,N_28613,N_29154);
and UO_2164 (O_2164,N_28748,N_28948);
nor UO_2165 (O_2165,N_28712,N_28581);
nor UO_2166 (O_2166,N_28909,N_29524);
and UO_2167 (O_2167,N_28855,N_29972);
or UO_2168 (O_2168,N_29717,N_28649);
xnor UO_2169 (O_2169,N_28861,N_29910);
or UO_2170 (O_2170,N_29577,N_28032);
nor UO_2171 (O_2171,N_28135,N_29545);
or UO_2172 (O_2172,N_29306,N_28568);
nand UO_2173 (O_2173,N_29021,N_28853);
nor UO_2174 (O_2174,N_28508,N_29879);
or UO_2175 (O_2175,N_28111,N_29326);
xnor UO_2176 (O_2176,N_29227,N_29684);
nand UO_2177 (O_2177,N_28826,N_28279);
nor UO_2178 (O_2178,N_29048,N_28367);
nand UO_2179 (O_2179,N_29047,N_29569);
nand UO_2180 (O_2180,N_29424,N_28830);
nor UO_2181 (O_2181,N_29871,N_29370);
xnor UO_2182 (O_2182,N_29221,N_29623);
or UO_2183 (O_2183,N_28987,N_28869);
nor UO_2184 (O_2184,N_29070,N_28182);
xnor UO_2185 (O_2185,N_28592,N_28042);
and UO_2186 (O_2186,N_28104,N_28357);
or UO_2187 (O_2187,N_29509,N_29307);
xor UO_2188 (O_2188,N_28434,N_28498);
nor UO_2189 (O_2189,N_28687,N_28712);
and UO_2190 (O_2190,N_29710,N_28350);
xnor UO_2191 (O_2191,N_29653,N_29374);
xor UO_2192 (O_2192,N_29635,N_28000);
nand UO_2193 (O_2193,N_28394,N_28797);
nand UO_2194 (O_2194,N_29595,N_29427);
nand UO_2195 (O_2195,N_29660,N_28585);
nand UO_2196 (O_2196,N_28666,N_28539);
nor UO_2197 (O_2197,N_29852,N_29372);
nand UO_2198 (O_2198,N_28014,N_29336);
xor UO_2199 (O_2199,N_28048,N_28580);
nor UO_2200 (O_2200,N_29202,N_28416);
and UO_2201 (O_2201,N_29116,N_28249);
xnor UO_2202 (O_2202,N_29832,N_28063);
or UO_2203 (O_2203,N_28474,N_28856);
and UO_2204 (O_2204,N_29582,N_28591);
and UO_2205 (O_2205,N_29283,N_28002);
or UO_2206 (O_2206,N_28770,N_29781);
nand UO_2207 (O_2207,N_29179,N_28724);
xnor UO_2208 (O_2208,N_29068,N_28282);
or UO_2209 (O_2209,N_29512,N_28080);
nand UO_2210 (O_2210,N_28833,N_29246);
and UO_2211 (O_2211,N_29781,N_29758);
xor UO_2212 (O_2212,N_29015,N_29820);
nand UO_2213 (O_2213,N_28837,N_28417);
or UO_2214 (O_2214,N_28421,N_29531);
nand UO_2215 (O_2215,N_29383,N_29484);
nand UO_2216 (O_2216,N_28966,N_29816);
nand UO_2217 (O_2217,N_28179,N_28533);
xnor UO_2218 (O_2218,N_29403,N_28181);
or UO_2219 (O_2219,N_28709,N_29268);
nor UO_2220 (O_2220,N_28024,N_28649);
nand UO_2221 (O_2221,N_29864,N_28525);
xnor UO_2222 (O_2222,N_29304,N_28736);
xnor UO_2223 (O_2223,N_29770,N_28373);
nor UO_2224 (O_2224,N_28628,N_29435);
nand UO_2225 (O_2225,N_28810,N_28716);
or UO_2226 (O_2226,N_29191,N_28414);
xnor UO_2227 (O_2227,N_29582,N_28611);
nor UO_2228 (O_2228,N_29531,N_28133);
nor UO_2229 (O_2229,N_28091,N_28807);
xor UO_2230 (O_2230,N_28252,N_29427);
nor UO_2231 (O_2231,N_28075,N_28181);
nor UO_2232 (O_2232,N_29037,N_28256);
nand UO_2233 (O_2233,N_29236,N_28586);
or UO_2234 (O_2234,N_29332,N_29809);
nor UO_2235 (O_2235,N_29690,N_28842);
or UO_2236 (O_2236,N_28475,N_28267);
xnor UO_2237 (O_2237,N_28695,N_29580);
xor UO_2238 (O_2238,N_29795,N_29961);
xor UO_2239 (O_2239,N_29715,N_29351);
xnor UO_2240 (O_2240,N_29068,N_29023);
nand UO_2241 (O_2241,N_29754,N_29319);
nor UO_2242 (O_2242,N_29255,N_28150);
xor UO_2243 (O_2243,N_28094,N_29455);
and UO_2244 (O_2244,N_28857,N_29326);
and UO_2245 (O_2245,N_28156,N_29689);
and UO_2246 (O_2246,N_28135,N_28517);
nand UO_2247 (O_2247,N_28911,N_29793);
and UO_2248 (O_2248,N_29267,N_29937);
or UO_2249 (O_2249,N_29159,N_28512);
xor UO_2250 (O_2250,N_29556,N_29237);
nand UO_2251 (O_2251,N_29432,N_29448);
xor UO_2252 (O_2252,N_28649,N_29487);
and UO_2253 (O_2253,N_29342,N_28202);
nand UO_2254 (O_2254,N_29066,N_29241);
nand UO_2255 (O_2255,N_29045,N_29745);
or UO_2256 (O_2256,N_28438,N_28474);
or UO_2257 (O_2257,N_28328,N_29996);
nor UO_2258 (O_2258,N_28958,N_29829);
nor UO_2259 (O_2259,N_29461,N_29657);
nor UO_2260 (O_2260,N_28156,N_28760);
xnor UO_2261 (O_2261,N_29949,N_28772);
and UO_2262 (O_2262,N_29474,N_29627);
nor UO_2263 (O_2263,N_28217,N_29601);
nand UO_2264 (O_2264,N_29706,N_29316);
nand UO_2265 (O_2265,N_29674,N_28087);
nand UO_2266 (O_2266,N_28874,N_29995);
and UO_2267 (O_2267,N_29271,N_28550);
nor UO_2268 (O_2268,N_28907,N_29126);
nor UO_2269 (O_2269,N_29360,N_29634);
nand UO_2270 (O_2270,N_29711,N_29142);
or UO_2271 (O_2271,N_28493,N_28387);
or UO_2272 (O_2272,N_29020,N_28065);
xnor UO_2273 (O_2273,N_29471,N_28228);
nor UO_2274 (O_2274,N_29535,N_29267);
or UO_2275 (O_2275,N_28281,N_29783);
or UO_2276 (O_2276,N_29800,N_29083);
and UO_2277 (O_2277,N_28093,N_28256);
and UO_2278 (O_2278,N_28135,N_28217);
nor UO_2279 (O_2279,N_29174,N_28008);
nand UO_2280 (O_2280,N_28121,N_29283);
nand UO_2281 (O_2281,N_29354,N_28452);
and UO_2282 (O_2282,N_29507,N_29312);
and UO_2283 (O_2283,N_29707,N_28651);
nand UO_2284 (O_2284,N_29806,N_29818);
nand UO_2285 (O_2285,N_28784,N_28769);
xnor UO_2286 (O_2286,N_29293,N_28807);
and UO_2287 (O_2287,N_28202,N_28422);
nand UO_2288 (O_2288,N_29509,N_28307);
nor UO_2289 (O_2289,N_29237,N_28963);
xor UO_2290 (O_2290,N_28611,N_28579);
and UO_2291 (O_2291,N_28623,N_29156);
or UO_2292 (O_2292,N_28496,N_28337);
nor UO_2293 (O_2293,N_29819,N_29982);
and UO_2294 (O_2294,N_28946,N_28325);
xor UO_2295 (O_2295,N_28997,N_28422);
nand UO_2296 (O_2296,N_29954,N_28181);
nand UO_2297 (O_2297,N_29567,N_29894);
or UO_2298 (O_2298,N_28205,N_29849);
and UO_2299 (O_2299,N_28479,N_29273);
nand UO_2300 (O_2300,N_29381,N_29324);
nor UO_2301 (O_2301,N_29960,N_29877);
or UO_2302 (O_2302,N_28012,N_29764);
nand UO_2303 (O_2303,N_28857,N_29019);
xor UO_2304 (O_2304,N_29948,N_28667);
nor UO_2305 (O_2305,N_28930,N_28178);
nor UO_2306 (O_2306,N_28036,N_29076);
nor UO_2307 (O_2307,N_29125,N_28737);
nand UO_2308 (O_2308,N_28395,N_29394);
xnor UO_2309 (O_2309,N_28269,N_28322);
or UO_2310 (O_2310,N_28690,N_28240);
and UO_2311 (O_2311,N_28074,N_28909);
or UO_2312 (O_2312,N_28698,N_29843);
and UO_2313 (O_2313,N_29330,N_29853);
nor UO_2314 (O_2314,N_28941,N_29702);
or UO_2315 (O_2315,N_28970,N_28895);
nand UO_2316 (O_2316,N_29874,N_28433);
nor UO_2317 (O_2317,N_29644,N_29450);
xnor UO_2318 (O_2318,N_29462,N_28567);
nor UO_2319 (O_2319,N_28048,N_29038);
and UO_2320 (O_2320,N_28186,N_29553);
or UO_2321 (O_2321,N_29756,N_28767);
nor UO_2322 (O_2322,N_28368,N_29538);
nand UO_2323 (O_2323,N_28278,N_29589);
and UO_2324 (O_2324,N_29203,N_28145);
and UO_2325 (O_2325,N_29772,N_29196);
or UO_2326 (O_2326,N_28565,N_28524);
and UO_2327 (O_2327,N_29204,N_28006);
or UO_2328 (O_2328,N_28114,N_29212);
xnor UO_2329 (O_2329,N_28944,N_28950);
and UO_2330 (O_2330,N_28145,N_29335);
and UO_2331 (O_2331,N_28222,N_29156);
xnor UO_2332 (O_2332,N_28629,N_29220);
nor UO_2333 (O_2333,N_29991,N_28279);
and UO_2334 (O_2334,N_28015,N_29865);
nor UO_2335 (O_2335,N_28912,N_28884);
xor UO_2336 (O_2336,N_29191,N_29154);
nand UO_2337 (O_2337,N_29992,N_29827);
or UO_2338 (O_2338,N_28448,N_28293);
or UO_2339 (O_2339,N_28349,N_29617);
or UO_2340 (O_2340,N_29746,N_29706);
or UO_2341 (O_2341,N_29560,N_28726);
xor UO_2342 (O_2342,N_29409,N_29058);
xor UO_2343 (O_2343,N_28129,N_29681);
and UO_2344 (O_2344,N_29010,N_28444);
nand UO_2345 (O_2345,N_28930,N_29715);
nor UO_2346 (O_2346,N_29029,N_29653);
nand UO_2347 (O_2347,N_29126,N_28228);
xor UO_2348 (O_2348,N_28241,N_29009);
and UO_2349 (O_2349,N_29609,N_29115);
nor UO_2350 (O_2350,N_29826,N_29883);
and UO_2351 (O_2351,N_28944,N_28587);
nor UO_2352 (O_2352,N_29270,N_28624);
xnor UO_2353 (O_2353,N_29146,N_28413);
or UO_2354 (O_2354,N_28129,N_28203);
and UO_2355 (O_2355,N_28347,N_28413);
and UO_2356 (O_2356,N_28552,N_28444);
or UO_2357 (O_2357,N_29628,N_29085);
nand UO_2358 (O_2358,N_29625,N_29476);
nor UO_2359 (O_2359,N_29000,N_29256);
and UO_2360 (O_2360,N_28641,N_29920);
xor UO_2361 (O_2361,N_29657,N_28136);
nand UO_2362 (O_2362,N_29298,N_28778);
nor UO_2363 (O_2363,N_29068,N_28389);
xor UO_2364 (O_2364,N_28664,N_28096);
nand UO_2365 (O_2365,N_28127,N_28394);
or UO_2366 (O_2366,N_28362,N_28723);
or UO_2367 (O_2367,N_29296,N_28476);
and UO_2368 (O_2368,N_29603,N_28603);
and UO_2369 (O_2369,N_28804,N_29937);
and UO_2370 (O_2370,N_29999,N_28423);
and UO_2371 (O_2371,N_29273,N_28186);
and UO_2372 (O_2372,N_29504,N_29862);
or UO_2373 (O_2373,N_29947,N_29707);
or UO_2374 (O_2374,N_29498,N_28913);
or UO_2375 (O_2375,N_29765,N_29228);
nand UO_2376 (O_2376,N_29267,N_29495);
or UO_2377 (O_2377,N_28407,N_29694);
or UO_2378 (O_2378,N_28326,N_29151);
xor UO_2379 (O_2379,N_28702,N_28773);
nand UO_2380 (O_2380,N_29288,N_29530);
or UO_2381 (O_2381,N_29502,N_29578);
or UO_2382 (O_2382,N_29560,N_28917);
nor UO_2383 (O_2383,N_28275,N_29501);
or UO_2384 (O_2384,N_29579,N_29530);
or UO_2385 (O_2385,N_28522,N_29437);
nor UO_2386 (O_2386,N_29422,N_29433);
nor UO_2387 (O_2387,N_28282,N_28010);
or UO_2388 (O_2388,N_28190,N_28958);
nor UO_2389 (O_2389,N_28106,N_29057);
and UO_2390 (O_2390,N_29302,N_28632);
and UO_2391 (O_2391,N_28826,N_29204);
xor UO_2392 (O_2392,N_28338,N_29946);
or UO_2393 (O_2393,N_28541,N_29532);
and UO_2394 (O_2394,N_29544,N_28059);
or UO_2395 (O_2395,N_29620,N_28809);
and UO_2396 (O_2396,N_28453,N_28352);
nand UO_2397 (O_2397,N_28639,N_29878);
and UO_2398 (O_2398,N_29370,N_28512);
or UO_2399 (O_2399,N_29555,N_29340);
nor UO_2400 (O_2400,N_29323,N_29846);
and UO_2401 (O_2401,N_28677,N_28687);
nand UO_2402 (O_2402,N_28379,N_28629);
and UO_2403 (O_2403,N_28598,N_29902);
nor UO_2404 (O_2404,N_28108,N_29356);
or UO_2405 (O_2405,N_28115,N_29463);
and UO_2406 (O_2406,N_28016,N_29470);
xnor UO_2407 (O_2407,N_28921,N_29751);
and UO_2408 (O_2408,N_29770,N_28502);
nand UO_2409 (O_2409,N_28665,N_28590);
xor UO_2410 (O_2410,N_28651,N_28491);
nand UO_2411 (O_2411,N_28053,N_29911);
xor UO_2412 (O_2412,N_28778,N_28086);
nor UO_2413 (O_2413,N_28893,N_29212);
or UO_2414 (O_2414,N_29269,N_28744);
or UO_2415 (O_2415,N_29583,N_29072);
or UO_2416 (O_2416,N_29646,N_29689);
nand UO_2417 (O_2417,N_28653,N_29076);
nand UO_2418 (O_2418,N_29819,N_28668);
nor UO_2419 (O_2419,N_29307,N_29035);
or UO_2420 (O_2420,N_29067,N_28637);
nand UO_2421 (O_2421,N_28214,N_28255);
or UO_2422 (O_2422,N_29960,N_28964);
and UO_2423 (O_2423,N_29192,N_29864);
xor UO_2424 (O_2424,N_29875,N_28302);
nand UO_2425 (O_2425,N_28893,N_29588);
and UO_2426 (O_2426,N_29773,N_28069);
and UO_2427 (O_2427,N_29962,N_29108);
and UO_2428 (O_2428,N_28387,N_29530);
or UO_2429 (O_2429,N_29022,N_29397);
nand UO_2430 (O_2430,N_29995,N_28472);
nand UO_2431 (O_2431,N_29643,N_29588);
and UO_2432 (O_2432,N_29744,N_28062);
nand UO_2433 (O_2433,N_29710,N_29969);
and UO_2434 (O_2434,N_28878,N_29262);
and UO_2435 (O_2435,N_28402,N_29359);
or UO_2436 (O_2436,N_28018,N_29428);
or UO_2437 (O_2437,N_29410,N_28080);
xor UO_2438 (O_2438,N_28961,N_29292);
xor UO_2439 (O_2439,N_28025,N_29888);
nor UO_2440 (O_2440,N_28712,N_29172);
nand UO_2441 (O_2441,N_29845,N_28046);
or UO_2442 (O_2442,N_29752,N_28373);
xnor UO_2443 (O_2443,N_29847,N_29677);
xor UO_2444 (O_2444,N_29734,N_29850);
and UO_2445 (O_2445,N_29669,N_29459);
or UO_2446 (O_2446,N_29184,N_29745);
and UO_2447 (O_2447,N_28305,N_28895);
nor UO_2448 (O_2448,N_29781,N_29452);
nor UO_2449 (O_2449,N_29982,N_29814);
nand UO_2450 (O_2450,N_29292,N_29599);
nand UO_2451 (O_2451,N_29744,N_28481);
xor UO_2452 (O_2452,N_29721,N_28671);
or UO_2453 (O_2453,N_28205,N_28263);
nand UO_2454 (O_2454,N_28340,N_29737);
or UO_2455 (O_2455,N_28769,N_29871);
and UO_2456 (O_2456,N_29811,N_29773);
xnor UO_2457 (O_2457,N_29101,N_29924);
nor UO_2458 (O_2458,N_29253,N_29240);
xnor UO_2459 (O_2459,N_28978,N_28280);
nand UO_2460 (O_2460,N_28909,N_29240);
or UO_2461 (O_2461,N_28353,N_28504);
nor UO_2462 (O_2462,N_28692,N_29638);
xor UO_2463 (O_2463,N_29703,N_28479);
nand UO_2464 (O_2464,N_28982,N_28846);
xnor UO_2465 (O_2465,N_28521,N_28928);
xnor UO_2466 (O_2466,N_29517,N_28513);
or UO_2467 (O_2467,N_29639,N_28151);
xor UO_2468 (O_2468,N_29430,N_29261);
nand UO_2469 (O_2469,N_29258,N_28466);
or UO_2470 (O_2470,N_28614,N_29950);
or UO_2471 (O_2471,N_28748,N_29809);
or UO_2472 (O_2472,N_29648,N_29911);
nand UO_2473 (O_2473,N_29582,N_28891);
nor UO_2474 (O_2474,N_28512,N_28383);
nor UO_2475 (O_2475,N_29225,N_28146);
xnor UO_2476 (O_2476,N_28970,N_28502);
and UO_2477 (O_2477,N_29932,N_28858);
or UO_2478 (O_2478,N_29805,N_28833);
or UO_2479 (O_2479,N_28800,N_29346);
nand UO_2480 (O_2480,N_28024,N_29173);
or UO_2481 (O_2481,N_28680,N_29663);
or UO_2482 (O_2482,N_29967,N_29526);
nor UO_2483 (O_2483,N_29316,N_28627);
nand UO_2484 (O_2484,N_28371,N_28928);
nor UO_2485 (O_2485,N_28263,N_29768);
and UO_2486 (O_2486,N_28590,N_28580);
and UO_2487 (O_2487,N_28428,N_29635);
xnor UO_2488 (O_2488,N_28207,N_29929);
and UO_2489 (O_2489,N_29936,N_29645);
nor UO_2490 (O_2490,N_29009,N_28493);
and UO_2491 (O_2491,N_28488,N_29179);
or UO_2492 (O_2492,N_29345,N_28381);
nor UO_2493 (O_2493,N_28465,N_29948);
or UO_2494 (O_2494,N_28428,N_28972);
xor UO_2495 (O_2495,N_29897,N_29926);
nor UO_2496 (O_2496,N_28459,N_28056);
nand UO_2497 (O_2497,N_28167,N_29183);
xor UO_2498 (O_2498,N_29182,N_29981);
nand UO_2499 (O_2499,N_28431,N_28119);
nor UO_2500 (O_2500,N_29656,N_28751);
nand UO_2501 (O_2501,N_29429,N_29744);
nor UO_2502 (O_2502,N_29722,N_29483);
xnor UO_2503 (O_2503,N_29174,N_29190);
or UO_2504 (O_2504,N_28537,N_28043);
nor UO_2505 (O_2505,N_29065,N_28040);
nand UO_2506 (O_2506,N_29302,N_28257);
and UO_2507 (O_2507,N_28598,N_28499);
nand UO_2508 (O_2508,N_28557,N_28333);
and UO_2509 (O_2509,N_28413,N_28784);
and UO_2510 (O_2510,N_28181,N_29477);
or UO_2511 (O_2511,N_29532,N_28000);
nand UO_2512 (O_2512,N_28534,N_28221);
and UO_2513 (O_2513,N_29900,N_29258);
and UO_2514 (O_2514,N_29916,N_29244);
xor UO_2515 (O_2515,N_28256,N_28159);
nor UO_2516 (O_2516,N_29690,N_29883);
xor UO_2517 (O_2517,N_29334,N_28611);
nor UO_2518 (O_2518,N_28187,N_29127);
and UO_2519 (O_2519,N_29715,N_28400);
and UO_2520 (O_2520,N_28135,N_29956);
nor UO_2521 (O_2521,N_28416,N_28939);
xnor UO_2522 (O_2522,N_29766,N_29943);
nand UO_2523 (O_2523,N_28618,N_28788);
xor UO_2524 (O_2524,N_28438,N_29322);
xor UO_2525 (O_2525,N_29906,N_28194);
xnor UO_2526 (O_2526,N_29211,N_28216);
nand UO_2527 (O_2527,N_29159,N_28154);
xor UO_2528 (O_2528,N_28084,N_28301);
nor UO_2529 (O_2529,N_29607,N_28202);
or UO_2530 (O_2530,N_28926,N_29087);
and UO_2531 (O_2531,N_28040,N_29431);
xnor UO_2532 (O_2532,N_28028,N_28300);
nand UO_2533 (O_2533,N_28134,N_29455);
or UO_2534 (O_2534,N_28163,N_28753);
nand UO_2535 (O_2535,N_28217,N_29000);
nor UO_2536 (O_2536,N_28270,N_29503);
and UO_2537 (O_2537,N_28464,N_28430);
xor UO_2538 (O_2538,N_29352,N_28673);
or UO_2539 (O_2539,N_29005,N_29095);
nand UO_2540 (O_2540,N_28660,N_28069);
nor UO_2541 (O_2541,N_29393,N_28223);
nor UO_2542 (O_2542,N_29653,N_28842);
xnor UO_2543 (O_2543,N_28069,N_28394);
nand UO_2544 (O_2544,N_29451,N_28974);
or UO_2545 (O_2545,N_29216,N_29925);
and UO_2546 (O_2546,N_29490,N_28644);
xnor UO_2547 (O_2547,N_28858,N_29408);
xor UO_2548 (O_2548,N_28334,N_28435);
or UO_2549 (O_2549,N_28019,N_29056);
xnor UO_2550 (O_2550,N_29478,N_28085);
xnor UO_2551 (O_2551,N_29902,N_29393);
xor UO_2552 (O_2552,N_29687,N_29267);
xor UO_2553 (O_2553,N_29942,N_28569);
nor UO_2554 (O_2554,N_28332,N_29961);
or UO_2555 (O_2555,N_28447,N_29860);
xor UO_2556 (O_2556,N_28758,N_28904);
and UO_2557 (O_2557,N_29003,N_28130);
xor UO_2558 (O_2558,N_28853,N_28705);
xnor UO_2559 (O_2559,N_28830,N_29904);
nand UO_2560 (O_2560,N_29709,N_29161);
xnor UO_2561 (O_2561,N_28612,N_29805);
or UO_2562 (O_2562,N_28840,N_28313);
xor UO_2563 (O_2563,N_28399,N_28917);
xor UO_2564 (O_2564,N_28393,N_29480);
and UO_2565 (O_2565,N_29005,N_29628);
nor UO_2566 (O_2566,N_29446,N_28626);
nor UO_2567 (O_2567,N_28307,N_28479);
nand UO_2568 (O_2568,N_28196,N_28502);
and UO_2569 (O_2569,N_29135,N_28777);
or UO_2570 (O_2570,N_29074,N_29544);
nor UO_2571 (O_2571,N_28991,N_29987);
nor UO_2572 (O_2572,N_29035,N_28728);
nand UO_2573 (O_2573,N_28217,N_29024);
nand UO_2574 (O_2574,N_28926,N_28900);
xor UO_2575 (O_2575,N_29414,N_28228);
and UO_2576 (O_2576,N_28267,N_29949);
nand UO_2577 (O_2577,N_28164,N_29947);
or UO_2578 (O_2578,N_28506,N_28196);
xor UO_2579 (O_2579,N_28217,N_29029);
and UO_2580 (O_2580,N_28278,N_29676);
and UO_2581 (O_2581,N_29847,N_29175);
nand UO_2582 (O_2582,N_29411,N_28508);
nor UO_2583 (O_2583,N_28735,N_28798);
or UO_2584 (O_2584,N_29010,N_28533);
nor UO_2585 (O_2585,N_28166,N_28705);
and UO_2586 (O_2586,N_28635,N_29627);
nor UO_2587 (O_2587,N_29552,N_28470);
nor UO_2588 (O_2588,N_29471,N_28027);
xnor UO_2589 (O_2589,N_29178,N_29202);
nand UO_2590 (O_2590,N_28998,N_28233);
or UO_2591 (O_2591,N_29700,N_28045);
or UO_2592 (O_2592,N_28083,N_28223);
nor UO_2593 (O_2593,N_28232,N_28207);
nand UO_2594 (O_2594,N_29357,N_29403);
xor UO_2595 (O_2595,N_29016,N_28223);
nor UO_2596 (O_2596,N_28433,N_28416);
or UO_2597 (O_2597,N_29365,N_28204);
nand UO_2598 (O_2598,N_28000,N_29813);
xor UO_2599 (O_2599,N_29071,N_29856);
and UO_2600 (O_2600,N_29300,N_28425);
nor UO_2601 (O_2601,N_29153,N_29861);
nand UO_2602 (O_2602,N_29759,N_28843);
xor UO_2603 (O_2603,N_28910,N_29546);
nand UO_2604 (O_2604,N_28878,N_29120);
or UO_2605 (O_2605,N_28710,N_29834);
nand UO_2606 (O_2606,N_29939,N_29027);
and UO_2607 (O_2607,N_28884,N_29559);
nand UO_2608 (O_2608,N_29303,N_28846);
xnor UO_2609 (O_2609,N_28161,N_29189);
xnor UO_2610 (O_2610,N_29452,N_29643);
nor UO_2611 (O_2611,N_28981,N_29512);
nor UO_2612 (O_2612,N_28896,N_29741);
and UO_2613 (O_2613,N_28647,N_29687);
or UO_2614 (O_2614,N_28593,N_28058);
or UO_2615 (O_2615,N_28354,N_29742);
and UO_2616 (O_2616,N_28237,N_28371);
or UO_2617 (O_2617,N_29021,N_28925);
nor UO_2618 (O_2618,N_29735,N_28468);
and UO_2619 (O_2619,N_28770,N_28875);
or UO_2620 (O_2620,N_29145,N_29938);
nand UO_2621 (O_2621,N_29584,N_28815);
or UO_2622 (O_2622,N_28960,N_28710);
and UO_2623 (O_2623,N_29210,N_29799);
xnor UO_2624 (O_2624,N_29581,N_28950);
nor UO_2625 (O_2625,N_29267,N_29796);
or UO_2626 (O_2626,N_29636,N_29922);
nor UO_2627 (O_2627,N_29638,N_28771);
nand UO_2628 (O_2628,N_28920,N_28951);
nand UO_2629 (O_2629,N_28762,N_29806);
or UO_2630 (O_2630,N_28824,N_29319);
and UO_2631 (O_2631,N_28316,N_28086);
nand UO_2632 (O_2632,N_29574,N_29157);
and UO_2633 (O_2633,N_29461,N_29297);
nor UO_2634 (O_2634,N_28367,N_29886);
nand UO_2635 (O_2635,N_28097,N_29286);
and UO_2636 (O_2636,N_29742,N_29868);
or UO_2637 (O_2637,N_29677,N_29209);
or UO_2638 (O_2638,N_28655,N_29947);
and UO_2639 (O_2639,N_29808,N_29761);
nor UO_2640 (O_2640,N_29189,N_29018);
xor UO_2641 (O_2641,N_29049,N_29366);
nand UO_2642 (O_2642,N_28772,N_29451);
nor UO_2643 (O_2643,N_28869,N_28681);
or UO_2644 (O_2644,N_29029,N_28861);
xor UO_2645 (O_2645,N_28029,N_28482);
xor UO_2646 (O_2646,N_29494,N_28482);
nand UO_2647 (O_2647,N_29854,N_28879);
nor UO_2648 (O_2648,N_29425,N_28904);
xnor UO_2649 (O_2649,N_28495,N_29385);
xnor UO_2650 (O_2650,N_28065,N_29780);
or UO_2651 (O_2651,N_29818,N_29259);
and UO_2652 (O_2652,N_28786,N_28912);
or UO_2653 (O_2653,N_29537,N_29171);
or UO_2654 (O_2654,N_28332,N_28952);
nand UO_2655 (O_2655,N_28956,N_29734);
xor UO_2656 (O_2656,N_29456,N_28039);
or UO_2657 (O_2657,N_28669,N_28750);
nor UO_2658 (O_2658,N_29350,N_29341);
and UO_2659 (O_2659,N_28918,N_29505);
and UO_2660 (O_2660,N_28675,N_29780);
xor UO_2661 (O_2661,N_29359,N_28247);
xnor UO_2662 (O_2662,N_29105,N_28910);
nand UO_2663 (O_2663,N_29454,N_28860);
nor UO_2664 (O_2664,N_29176,N_29508);
or UO_2665 (O_2665,N_29125,N_28634);
or UO_2666 (O_2666,N_28997,N_28620);
or UO_2667 (O_2667,N_29351,N_29141);
and UO_2668 (O_2668,N_29733,N_28039);
or UO_2669 (O_2669,N_28733,N_29795);
nor UO_2670 (O_2670,N_29853,N_29902);
and UO_2671 (O_2671,N_28004,N_28436);
nand UO_2672 (O_2672,N_29493,N_28974);
nor UO_2673 (O_2673,N_28690,N_29862);
xnor UO_2674 (O_2674,N_28860,N_28612);
nor UO_2675 (O_2675,N_29056,N_29138);
xnor UO_2676 (O_2676,N_29121,N_29034);
nand UO_2677 (O_2677,N_28421,N_29490);
or UO_2678 (O_2678,N_29746,N_28312);
and UO_2679 (O_2679,N_28915,N_28299);
xnor UO_2680 (O_2680,N_29829,N_28047);
nor UO_2681 (O_2681,N_29573,N_28954);
or UO_2682 (O_2682,N_29151,N_29975);
or UO_2683 (O_2683,N_28332,N_29640);
and UO_2684 (O_2684,N_29762,N_29778);
or UO_2685 (O_2685,N_29475,N_29754);
xnor UO_2686 (O_2686,N_29976,N_28249);
nand UO_2687 (O_2687,N_29220,N_28987);
nand UO_2688 (O_2688,N_29678,N_29604);
or UO_2689 (O_2689,N_29539,N_28372);
nor UO_2690 (O_2690,N_28024,N_29198);
nor UO_2691 (O_2691,N_28633,N_28818);
nand UO_2692 (O_2692,N_29644,N_28617);
or UO_2693 (O_2693,N_29344,N_29376);
or UO_2694 (O_2694,N_29811,N_28079);
or UO_2695 (O_2695,N_28165,N_29991);
nand UO_2696 (O_2696,N_29514,N_29280);
nor UO_2697 (O_2697,N_29294,N_28540);
xor UO_2698 (O_2698,N_29397,N_28848);
and UO_2699 (O_2699,N_29263,N_28933);
xnor UO_2700 (O_2700,N_28327,N_28399);
nor UO_2701 (O_2701,N_28736,N_29124);
nand UO_2702 (O_2702,N_29686,N_28997);
nand UO_2703 (O_2703,N_29272,N_29637);
or UO_2704 (O_2704,N_28665,N_28700);
and UO_2705 (O_2705,N_28233,N_28961);
and UO_2706 (O_2706,N_28703,N_29446);
or UO_2707 (O_2707,N_29217,N_28047);
xnor UO_2708 (O_2708,N_29416,N_29659);
and UO_2709 (O_2709,N_28066,N_29002);
or UO_2710 (O_2710,N_29070,N_29489);
xor UO_2711 (O_2711,N_28534,N_28125);
or UO_2712 (O_2712,N_28071,N_28940);
xor UO_2713 (O_2713,N_28419,N_28210);
nor UO_2714 (O_2714,N_29033,N_29108);
xor UO_2715 (O_2715,N_28351,N_29257);
xnor UO_2716 (O_2716,N_28416,N_28461);
nand UO_2717 (O_2717,N_29244,N_28760);
or UO_2718 (O_2718,N_28847,N_28190);
nor UO_2719 (O_2719,N_29146,N_28030);
nand UO_2720 (O_2720,N_29913,N_28645);
nand UO_2721 (O_2721,N_29378,N_28394);
or UO_2722 (O_2722,N_29289,N_28108);
and UO_2723 (O_2723,N_28760,N_29492);
or UO_2724 (O_2724,N_28648,N_29640);
xor UO_2725 (O_2725,N_29955,N_28817);
nand UO_2726 (O_2726,N_28526,N_29348);
or UO_2727 (O_2727,N_28721,N_29219);
and UO_2728 (O_2728,N_29232,N_29753);
or UO_2729 (O_2729,N_28971,N_29485);
nand UO_2730 (O_2730,N_28163,N_29390);
nand UO_2731 (O_2731,N_29507,N_29284);
xnor UO_2732 (O_2732,N_28715,N_29202);
xnor UO_2733 (O_2733,N_28515,N_28658);
and UO_2734 (O_2734,N_29609,N_28711);
nand UO_2735 (O_2735,N_29080,N_28712);
or UO_2736 (O_2736,N_29527,N_29946);
nand UO_2737 (O_2737,N_29597,N_28134);
and UO_2738 (O_2738,N_28366,N_29496);
or UO_2739 (O_2739,N_28468,N_28276);
nand UO_2740 (O_2740,N_28831,N_29418);
and UO_2741 (O_2741,N_29470,N_29093);
and UO_2742 (O_2742,N_29820,N_28209);
nand UO_2743 (O_2743,N_29015,N_28504);
or UO_2744 (O_2744,N_28347,N_29501);
xor UO_2745 (O_2745,N_29976,N_29698);
nand UO_2746 (O_2746,N_28605,N_29478);
nor UO_2747 (O_2747,N_29138,N_29049);
nor UO_2748 (O_2748,N_28806,N_28657);
xor UO_2749 (O_2749,N_29540,N_29043);
or UO_2750 (O_2750,N_28673,N_29179);
nor UO_2751 (O_2751,N_28848,N_28181);
nor UO_2752 (O_2752,N_29758,N_28533);
and UO_2753 (O_2753,N_29348,N_28766);
or UO_2754 (O_2754,N_28388,N_29797);
nor UO_2755 (O_2755,N_29952,N_28380);
and UO_2756 (O_2756,N_29888,N_28586);
xnor UO_2757 (O_2757,N_29803,N_29714);
nor UO_2758 (O_2758,N_29930,N_28822);
nand UO_2759 (O_2759,N_29885,N_28556);
nor UO_2760 (O_2760,N_29411,N_28411);
xor UO_2761 (O_2761,N_29972,N_28302);
or UO_2762 (O_2762,N_28915,N_28728);
nand UO_2763 (O_2763,N_29787,N_29837);
nand UO_2764 (O_2764,N_29438,N_28220);
and UO_2765 (O_2765,N_28926,N_28265);
xor UO_2766 (O_2766,N_29440,N_29850);
nor UO_2767 (O_2767,N_28495,N_29783);
nor UO_2768 (O_2768,N_29957,N_28012);
nor UO_2769 (O_2769,N_28662,N_29794);
nor UO_2770 (O_2770,N_29104,N_29375);
nor UO_2771 (O_2771,N_28794,N_28633);
nor UO_2772 (O_2772,N_28928,N_28630);
xnor UO_2773 (O_2773,N_29328,N_28535);
nor UO_2774 (O_2774,N_28761,N_28124);
nor UO_2775 (O_2775,N_28986,N_28967);
and UO_2776 (O_2776,N_28581,N_28413);
xor UO_2777 (O_2777,N_28464,N_29487);
or UO_2778 (O_2778,N_29108,N_29935);
nand UO_2779 (O_2779,N_28814,N_29115);
xnor UO_2780 (O_2780,N_29196,N_29292);
xnor UO_2781 (O_2781,N_29768,N_29009);
or UO_2782 (O_2782,N_29193,N_28550);
xnor UO_2783 (O_2783,N_29356,N_29122);
or UO_2784 (O_2784,N_29286,N_28817);
and UO_2785 (O_2785,N_29017,N_28490);
and UO_2786 (O_2786,N_29699,N_29927);
or UO_2787 (O_2787,N_29647,N_29392);
nand UO_2788 (O_2788,N_29736,N_28926);
or UO_2789 (O_2789,N_29585,N_28693);
nand UO_2790 (O_2790,N_28040,N_29318);
and UO_2791 (O_2791,N_28875,N_28295);
nor UO_2792 (O_2792,N_29243,N_29411);
nand UO_2793 (O_2793,N_28413,N_28296);
or UO_2794 (O_2794,N_28743,N_28838);
xor UO_2795 (O_2795,N_29992,N_28458);
nand UO_2796 (O_2796,N_28490,N_28443);
xor UO_2797 (O_2797,N_29124,N_28229);
or UO_2798 (O_2798,N_28341,N_28928);
xor UO_2799 (O_2799,N_28093,N_29029);
nor UO_2800 (O_2800,N_28533,N_28548);
nand UO_2801 (O_2801,N_29772,N_28022);
and UO_2802 (O_2802,N_29838,N_28295);
and UO_2803 (O_2803,N_29291,N_28728);
and UO_2804 (O_2804,N_29800,N_28889);
xor UO_2805 (O_2805,N_28067,N_29790);
and UO_2806 (O_2806,N_29511,N_28698);
or UO_2807 (O_2807,N_28453,N_28723);
xnor UO_2808 (O_2808,N_28712,N_29962);
xnor UO_2809 (O_2809,N_28884,N_29995);
and UO_2810 (O_2810,N_29949,N_28747);
nor UO_2811 (O_2811,N_29229,N_28529);
xnor UO_2812 (O_2812,N_28761,N_28678);
and UO_2813 (O_2813,N_29878,N_29218);
and UO_2814 (O_2814,N_28270,N_28215);
xor UO_2815 (O_2815,N_28109,N_29017);
nor UO_2816 (O_2816,N_29851,N_28402);
nor UO_2817 (O_2817,N_29076,N_29032);
nand UO_2818 (O_2818,N_29347,N_29978);
nand UO_2819 (O_2819,N_28990,N_29478);
nand UO_2820 (O_2820,N_28355,N_29469);
nor UO_2821 (O_2821,N_29523,N_28276);
nand UO_2822 (O_2822,N_28422,N_29127);
or UO_2823 (O_2823,N_29835,N_29848);
and UO_2824 (O_2824,N_29477,N_29048);
and UO_2825 (O_2825,N_29443,N_29071);
xor UO_2826 (O_2826,N_28187,N_28178);
xor UO_2827 (O_2827,N_29972,N_29913);
xor UO_2828 (O_2828,N_29166,N_28000);
and UO_2829 (O_2829,N_29081,N_28834);
nor UO_2830 (O_2830,N_28402,N_29491);
nand UO_2831 (O_2831,N_29264,N_28565);
nand UO_2832 (O_2832,N_28136,N_29227);
and UO_2833 (O_2833,N_28881,N_28967);
nand UO_2834 (O_2834,N_28831,N_28349);
or UO_2835 (O_2835,N_29110,N_28132);
or UO_2836 (O_2836,N_28308,N_28188);
xor UO_2837 (O_2837,N_29625,N_29287);
xnor UO_2838 (O_2838,N_28804,N_28564);
xnor UO_2839 (O_2839,N_28544,N_28379);
and UO_2840 (O_2840,N_29694,N_29890);
nor UO_2841 (O_2841,N_28659,N_29502);
and UO_2842 (O_2842,N_28313,N_28177);
and UO_2843 (O_2843,N_28046,N_28759);
and UO_2844 (O_2844,N_29621,N_29311);
or UO_2845 (O_2845,N_29278,N_28009);
nor UO_2846 (O_2846,N_29687,N_28628);
nor UO_2847 (O_2847,N_28987,N_29359);
or UO_2848 (O_2848,N_29270,N_28531);
and UO_2849 (O_2849,N_28576,N_28591);
and UO_2850 (O_2850,N_29058,N_28065);
and UO_2851 (O_2851,N_29341,N_29575);
xnor UO_2852 (O_2852,N_28210,N_28966);
nand UO_2853 (O_2853,N_29839,N_29714);
or UO_2854 (O_2854,N_28013,N_28717);
or UO_2855 (O_2855,N_29930,N_28267);
or UO_2856 (O_2856,N_29829,N_29043);
nand UO_2857 (O_2857,N_28178,N_29829);
nand UO_2858 (O_2858,N_29682,N_29331);
nand UO_2859 (O_2859,N_28792,N_28187);
and UO_2860 (O_2860,N_29359,N_28146);
and UO_2861 (O_2861,N_28691,N_28936);
or UO_2862 (O_2862,N_29260,N_29369);
and UO_2863 (O_2863,N_28328,N_29052);
or UO_2864 (O_2864,N_29451,N_29750);
nand UO_2865 (O_2865,N_28152,N_29458);
or UO_2866 (O_2866,N_28681,N_28899);
and UO_2867 (O_2867,N_28533,N_29890);
or UO_2868 (O_2868,N_29584,N_28432);
or UO_2869 (O_2869,N_28235,N_28050);
nor UO_2870 (O_2870,N_29991,N_28536);
nand UO_2871 (O_2871,N_28389,N_29176);
or UO_2872 (O_2872,N_28515,N_28778);
nand UO_2873 (O_2873,N_29277,N_29775);
xor UO_2874 (O_2874,N_28026,N_28133);
xor UO_2875 (O_2875,N_28615,N_28507);
and UO_2876 (O_2876,N_29505,N_28781);
or UO_2877 (O_2877,N_29400,N_28477);
and UO_2878 (O_2878,N_28758,N_29080);
or UO_2879 (O_2879,N_29693,N_29461);
or UO_2880 (O_2880,N_29223,N_28547);
nand UO_2881 (O_2881,N_29291,N_28330);
or UO_2882 (O_2882,N_28659,N_28440);
xor UO_2883 (O_2883,N_28077,N_29958);
xnor UO_2884 (O_2884,N_29899,N_29039);
or UO_2885 (O_2885,N_29516,N_28429);
xor UO_2886 (O_2886,N_29630,N_28111);
nor UO_2887 (O_2887,N_29467,N_29372);
nor UO_2888 (O_2888,N_29406,N_28695);
nor UO_2889 (O_2889,N_29134,N_29428);
and UO_2890 (O_2890,N_29287,N_28366);
or UO_2891 (O_2891,N_29523,N_29567);
or UO_2892 (O_2892,N_29303,N_28338);
and UO_2893 (O_2893,N_28178,N_29231);
nor UO_2894 (O_2894,N_29021,N_28587);
nand UO_2895 (O_2895,N_29852,N_28478);
nor UO_2896 (O_2896,N_29237,N_29596);
and UO_2897 (O_2897,N_29411,N_28612);
or UO_2898 (O_2898,N_28838,N_29524);
nand UO_2899 (O_2899,N_28532,N_29345);
or UO_2900 (O_2900,N_28851,N_29086);
and UO_2901 (O_2901,N_28934,N_29364);
and UO_2902 (O_2902,N_29493,N_29509);
nand UO_2903 (O_2903,N_29648,N_28551);
and UO_2904 (O_2904,N_28511,N_28955);
nor UO_2905 (O_2905,N_29769,N_29352);
or UO_2906 (O_2906,N_29416,N_28817);
and UO_2907 (O_2907,N_29653,N_28228);
nor UO_2908 (O_2908,N_28183,N_29075);
nand UO_2909 (O_2909,N_28409,N_29607);
nor UO_2910 (O_2910,N_29888,N_28879);
and UO_2911 (O_2911,N_29055,N_28599);
nand UO_2912 (O_2912,N_29962,N_29275);
nor UO_2913 (O_2913,N_29557,N_28529);
and UO_2914 (O_2914,N_29123,N_29843);
or UO_2915 (O_2915,N_29007,N_29156);
or UO_2916 (O_2916,N_29762,N_28791);
xor UO_2917 (O_2917,N_28612,N_28893);
nor UO_2918 (O_2918,N_29541,N_28264);
or UO_2919 (O_2919,N_29313,N_28140);
and UO_2920 (O_2920,N_28224,N_29286);
nand UO_2921 (O_2921,N_29628,N_29186);
and UO_2922 (O_2922,N_28127,N_28600);
xnor UO_2923 (O_2923,N_29325,N_28651);
and UO_2924 (O_2924,N_29140,N_29751);
xor UO_2925 (O_2925,N_29690,N_29577);
nor UO_2926 (O_2926,N_28104,N_29749);
or UO_2927 (O_2927,N_28257,N_28519);
or UO_2928 (O_2928,N_28176,N_29785);
or UO_2929 (O_2929,N_29454,N_28466);
nor UO_2930 (O_2930,N_28890,N_29795);
or UO_2931 (O_2931,N_28886,N_28969);
nor UO_2932 (O_2932,N_28007,N_29432);
nand UO_2933 (O_2933,N_29333,N_29550);
xor UO_2934 (O_2934,N_29807,N_29196);
nor UO_2935 (O_2935,N_29376,N_29056);
nand UO_2936 (O_2936,N_29296,N_29378);
or UO_2937 (O_2937,N_29711,N_28841);
nor UO_2938 (O_2938,N_28867,N_28547);
or UO_2939 (O_2939,N_29745,N_28063);
and UO_2940 (O_2940,N_28924,N_29711);
nand UO_2941 (O_2941,N_29715,N_28806);
nor UO_2942 (O_2942,N_28903,N_28224);
nor UO_2943 (O_2943,N_29275,N_29203);
nand UO_2944 (O_2944,N_28925,N_29104);
nand UO_2945 (O_2945,N_28073,N_29541);
and UO_2946 (O_2946,N_29536,N_28648);
nand UO_2947 (O_2947,N_28348,N_29572);
and UO_2948 (O_2948,N_28955,N_29202);
nand UO_2949 (O_2949,N_28787,N_29229);
nor UO_2950 (O_2950,N_29740,N_28692);
or UO_2951 (O_2951,N_28395,N_29317);
xnor UO_2952 (O_2952,N_28929,N_28084);
or UO_2953 (O_2953,N_28803,N_28142);
or UO_2954 (O_2954,N_28222,N_28052);
xnor UO_2955 (O_2955,N_28782,N_28026);
or UO_2956 (O_2956,N_29192,N_29618);
nand UO_2957 (O_2957,N_29902,N_29290);
and UO_2958 (O_2958,N_29994,N_28794);
xnor UO_2959 (O_2959,N_29477,N_28011);
or UO_2960 (O_2960,N_29362,N_28271);
nand UO_2961 (O_2961,N_28332,N_29366);
xnor UO_2962 (O_2962,N_29134,N_29894);
xor UO_2963 (O_2963,N_29494,N_29103);
nor UO_2964 (O_2964,N_28769,N_29024);
and UO_2965 (O_2965,N_28741,N_28101);
nor UO_2966 (O_2966,N_29450,N_29444);
and UO_2967 (O_2967,N_29122,N_29223);
nand UO_2968 (O_2968,N_29675,N_29833);
nand UO_2969 (O_2969,N_29993,N_29048);
nand UO_2970 (O_2970,N_28349,N_28626);
xor UO_2971 (O_2971,N_28161,N_29164);
and UO_2972 (O_2972,N_28391,N_28114);
nor UO_2973 (O_2973,N_28033,N_28750);
and UO_2974 (O_2974,N_28143,N_29988);
xnor UO_2975 (O_2975,N_29415,N_29062);
or UO_2976 (O_2976,N_28912,N_29516);
or UO_2977 (O_2977,N_28277,N_29305);
nand UO_2978 (O_2978,N_28102,N_28276);
or UO_2979 (O_2979,N_29588,N_28103);
xor UO_2980 (O_2980,N_28452,N_28686);
nand UO_2981 (O_2981,N_29980,N_28093);
and UO_2982 (O_2982,N_29274,N_29322);
nor UO_2983 (O_2983,N_29186,N_28163);
xnor UO_2984 (O_2984,N_28724,N_29071);
nor UO_2985 (O_2985,N_28886,N_29730);
or UO_2986 (O_2986,N_29595,N_29513);
nor UO_2987 (O_2987,N_28346,N_28339);
nor UO_2988 (O_2988,N_28758,N_28938);
nand UO_2989 (O_2989,N_29305,N_29833);
and UO_2990 (O_2990,N_29789,N_29712);
nor UO_2991 (O_2991,N_28166,N_28939);
xor UO_2992 (O_2992,N_28510,N_29184);
or UO_2993 (O_2993,N_28667,N_28933);
xor UO_2994 (O_2994,N_28914,N_28211);
or UO_2995 (O_2995,N_29791,N_28147);
nand UO_2996 (O_2996,N_28190,N_28231);
and UO_2997 (O_2997,N_28595,N_29332);
or UO_2998 (O_2998,N_29400,N_28612);
or UO_2999 (O_2999,N_29475,N_29059);
or UO_3000 (O_3000,N_29292,N_28122);
nor UO_3001 (O_3001,N_29770,N_28059);
and UO_3002 (O_3002,N_29716,N_29731);
nor UO_3003 (O_3003,N_28745,N_29742);
xor UO_3004 (O_3004,N_28686,N_29291);
or UO_3005 (O_3005,N_28551,N_29207);
or UO_3006 (O_3006,N_29009,N_28332);
xnor UO_3007 (O_3007,N_28538,N_28661);
and UO_3008 (O_3008,N_28284,N_28842);
or UO_3009 (O_3009,N_29270,N_28455);
nor UO_3010 (O_3010,N_29195,N_28567);
or UO_3011 (O_3011,N_29077,N_29552);
xor UO_3012 (O_3012,N_28596,N_29770);
nor UO_3013 (O_3013,N_28978,N_28638);
xnor UO_3014 (O_3014,N_28434,N_28320);
and UO_3015 (O_3015,N_28255,N_29898);
nand UO_3016 (O_3016,N_28503,N_28149);
and UO_3017 (O_3017,N_28361,N_29449);
and UO_3018 (O_3018,N_28247,N_29192);
and UO_3019 (O_3019,N_28295,N_29268);
or UO_3020 (O_3020,N_29599,N_29012);
and UO_3021 (O_3021,N_28102,N_29282);
xnor UO_3022 (O_3022,N_29403,N_28400);
or UO_3023 (O_3023,N_28384,N_28086);
xnor UO_3024 (O_3024,N_29445,N_29046);
xor UO_3025 (O_3025,N_29143,N_28889);
xor UO_3026 (O_3026,N_29493,N_28461);
nand UO_3027 (O_3027,N_29365,N_28544);
and UO_3028 (O_3028,N_28278,N_28902);
or UO_3029 (O_3029,N_29282,N_28214);
nor UO_3030 (O_3030,N_29163,N_28771);
and UO_3031 (O_3031,N_28644,N_28381);
xor UO_3032 (O_3032,N_29875,N_28260);
and UO_3033 (O_3033,N_28983,N_28730);
and UO_3034 (O_3034,N_29653,N_28739);
xor UO_3035 (O_3035,N_29373,N_28976);
or UO_3036 (O_3036,N_29039,N_29555);
nor UO_3037 (O_3037,N_29595,N_29239);
or UO_3038 (O_3038,N_29040,N_29842);
and UO_3039 (O_3039,N_28157,N_28727);
or UO_3040 (O_3040,N_28122,N_29969);
and UO_3041 (O_3041,N_29603,N_28600);
and UO_3042 (O_3042,N_28245,N_29725);
or UO_3043 (O_3043,N_29128,N_29514);
nor UO_3044 (O_3044,N_28679,N_29856);
nand UO_3045 (O_3045,N_29045,N_29450);
nor UO_3046 (O_3046,N_29972,N_28905);
or UO_3047 (O_3047,N_29321,N_28206);
and UO_3048 (O_3048,N_28386,N_29863);
xor UO_3049 (O_3049,N_28664,N_28975);
nand UO_3050 (O_3050,N_29192,N_29750);
nand UO_3051 (O_3051,N_28265,N_29897);
and UO_3052 (O_3052,N_29250,N_28249);
and UO_3053 (O_3053,N_29869,N_28330);
nor UO_3054 (O_3054,N_29788,N_29168);
nor UO_3055 (O_3055,N_29345,N_28440);
xor UO_3056 (O_3056,N_29254,N_29772);
nand UO_3057 (O_3057,N_28964,N_29016);
xor UO_3058 (O_3058,N_29361,N_28006);
and UO_3059 (O_3059,N_29408,N_28817);
xnor UO_3060 (O_3060,N_28644,N_28572);
nor UO_3061 (O_3061,N_29187,N_28962);
and UO_3062 (O_3062,N_28612,N_29828);
nand UO_3063 (O_3063,N_29570,N_29828);
or UO_3064 (O_3064,N_29114,N_29760);
or UO_3065 (O_3065,N_29024,N_28783);
or UO_3066 (O_3066,N_29339,N_28612);
xnor UO_3067 (O_3067,N_29752,N_29248);
nor UO_3068 (O_3068,N_29064,N_28714);
nand UO_3069 (O_3069,N_29256,N_29910);
xor UO_3070 (O_3070,N_29250,N_29807);
nand UO_3071 (O_3071,N_29499,N_28339);
nor UO_3072 (O_3072,N_29155,N_28822);
and UO_3073 (O_3073,N_29337,N_28834);
or UO_3074 (O_3074,N_29236,N_28232);
nand UO_3075 (O_3075,N_28887,N_28520);
nor UO_3076 (O_3076,N_29474,N_29638);
nor UO_3077 (O_3077,N_28464,N_28022);
nand UO_3078 (O_3078,N_29259,N_28521);
nand UO_3079 (O_3079,N_28219,N_29462);
and UO_3080 (O_3080,N_29842,N_29749);
nand UO_3081 (O_3081,N_29919,N_28008);
xnor UO_3082 (O_3082,N_28910,N_28637);
or UO_3083 (O_3083,N_28445,N_28048);
nand UO_3084 (O_3084,N_28846,N_29662);
or UO_3085 (O_3085,N_28533,N_28003);
nor UO_3086 (O_3086,N_29092,N_29519);
and UO_3087 (O_3087,N_28169,N_28864);
nand UO_3088 (O_3088,N_28686,N_29766);
nand UO_3089 (O_3089,N_28977,N_29674);
nand UO_3090 (O_3090,N_28159,N_28719);
nand UO_3091 (O_3091,N_29774,N_28817);
or UO_3092 (O_3092,N_28806,N_29983);
and UO_3093 (O_3093,N_28237,N_28050);
or UO_3094 (O_3094,N_28712,N_29851);
nand UO_3095 (O_3095,N_29875,N_28193);
or UO_3096 (O_3096,N_28359,N_29780);
and UO_3097 (O_3097,N_29174,N_29025);
and UO_3098 (O_3098,N_29762,N_28079);
xnor UO_3099 (O_3099,N_28932,N_29219);
nor UO_3100 (O_3100,N_28378,N_29973);
nor UO_3101 (O_3101,N_28215,N_29467);
and UO_3102 (O_3102,N_29614,N_28360);
nor UO_3103 (O_3103,N_28367,N_29360);
nor UO_3104 (O_3104,N_29677,N_28133);
nand UO_3105 (O_3105,N_29769,N_29261);
nor UO_3106 (O_3106,N_28278,N_29346);
nor UO_3107 (O_3107,N_29929,N_29791);
nand UO_3108 (O_3108,N_29774,N_29478);
nand UO_3109 (O_3109,N_29594,N_28432);
nor UO_3110 (O_3110,N_29346,N_29993);
nand UO_3111 (O_3111,N_28605,N_28348);
nand UO_3112 (O_3112,N_28287,N_29473);
or UO_3113 (O_3113,N_29473,N_28375);
or UO_3114 (O_3114,N_28379,N_29411);
and UO_3115 (O_3115,N_29732,N_28200);
xor UO_3116 (O_3116,N_29610,N_28009);
nor UO_3117 (O_3117,N_28291,N_28988);
nor UO_3118 (O_3118,N_28772,N_29642);
xnor UO_3119 (O_3119,N_29025,N_28826);
or UO_3120 (O_3120,N_28538,N_28047);
nand UO_3121 (O_3121,N_28725,N_28473);
and UO_3122 (O_3122,N_29209,N_29287);
and UO_3123 (O_3123,N_29003,N_29568);
nand UO_3124 (O_3124,N_29812,N_29694);
nand UO_3125 (O_3125,N_29209,N_29741);
and UO_3126 (O_3126,N_28869,N_28606);
or UO_3127 (O_3127,N_28803,N_28931);
nand UO_3128 (O_3128,N_28931,N_29228);
or UO_3129 (O_3129,N_28519,N_28218);
nor UO_3130 (O_3130,N_28252,N_28627);
nand UO_3131 (O_3131,N_29575,N_28193);
nor UO_3132 (O_3132,N_29821,N_29963);
and UO_3133 (O_3133,N_28355,N_28670);
nand UO_3134 (O_3134,N_28980,N_28616);
and UO_3135 (O_3135,N_29361,N_28182);
nor UO_3136 (O_3136,N_28436,N_29862);
and UO_3137 (O_3137,N_29159,N_29964);
and UO_3138 (O_3138,N_28198,N_29890);
nor UO_3139 (O_3139,N_29250,N_28652);
xor UO_3140 (O_3140,N_28496,N_29951);
xnor UO_3141 (O_3141,N_28428,N_28011);
or UO_3142 (O_3142,N_29919,N_29035);
nor UO_3143 (O_3143,N_29801,N_28715);
or UO_3144 (O_3144,N_28475,N_28727);
and UO_3145 (O_3145,N_29853,N_29045);
nor UO_3146 (O_3146,N_29230,N_28219);
nor UO_3147 (O_3147,N_29119,N_29981);
xor UO_3148 (O_3148,N_29548,N_28520);
and UO_3149 (O_3149,N_28726,N_28227);
and UO_3150 (O_3150,N_28030,N_28081);
or UO_3151 (O_3151,N_28031,N_28024);
or UO_3152 (O_3152,N_28238,N_29773);
or UO_3153 (O_3153,N_28709,N_29088);
nand UO_3154 (O_3154,N_29361,N_29402);
or UO_3155 (O_3155,N_28148,N_29330);
or UO_3156 (O_3156,N_29688,N_29249);
or UO_3157 (O_3157,N_28394,N_28409);
and UO_3158 (O_3158,N_28424,N_28329);
and UO_3159 (O_3159,N_29945,N_28828);
nor UO_3160 (O_3160,N_28945,N_29307);
xor UO_3161 (O_3161,N_29018,N_28069);
xor UO_3162 (O_3162,N_29291,N_29648);
or UO_3163 (O_3163,N_28856,N_28011);
nand UO_3164 (O_3164,N_28880,N_29074);
or UO_3165 (O_3165,N_29354,N_29964);
and UO_3166 (O_3166,N_29659,N_28476);
xnor UO_3167 (O_3167,N_29777,N_29368);
nor UO_3168 (O_3168,N_29017,N_29448);
and UO_3169 (O_3169,N_28001,N_28079);
and UO_3170 (O_3170,N_28332,N_28759);
nor UO_3171 (O_3171,N_28773,N_28701);
xor UO_3172 (O_3172,N_28662,N_29086);
nand UO_3173 (O_3173,N_29075,N_29565);
or UO_3174 (O_3174,N_29564,N_29124);
or UO_3175 (O_3175,N_28916,N_29247);
nand UO_3176 (O_3176,N_28745,N_29414);
or UO_3177 (O_3177,N_29914,N_29608);
nand UO_3178 (O_3178,N_29401,N_29187);
or UO_3179 (O_3179,N_29267,N_28406);
nor UO_3180 (O_3180,N_29960,N_29948);
nor UO_3181 (O_3181,N_29874,N_28356);
nand UO_3182 (O_3182,N_28349,N_28192);
or UO_3183 (O_3183,N_29055,N_28980);
or UO_3184 (O_3184,N_28968,N_28917);
xor UO_3185 (O_3185,N_28548,N_29672);
and UO_3186 (O_3186,N_28823,N_28433);
nand UO_3187 (O_3187,N_29098,N_29644);
nand UO_3188 (O_3188,N_28820,N_29939);
and UO_3189 (O_3189,N_29142,N_29079);
nand UO_3190 (O_3190,N_28066,N_28877);
xnor UO_3191 (O_3191,N_28575,N_28673);
nor UO_3192 (O_3192,N_28067,N_28006);
or UO_3193 (O_3193,N_28169,N_29391);
nor UO_3194 (O_3194,N_28572,N_29974);
xnor UO_3195 (O_3195,N_28351,N_28272);
xor UO_3196 (O_3196,N_28597,N_28371);
nor UO_3197 (O_3197,N_28716,N_29163);
xor UO_3198 (O_3198,N_29998,N_29504);
nor UO_3199 (O_3199,N_29997,N_28065);
nor UO_3200 (O_3200,N_29719,N_28029);
and UO_3201 (O_3201,N_29151,N_29555);
xnor UO_3202 (O_3202,N_28136,N_28380);
nor UO_3203 (O_3203,N_28520,N_28016);
or UO_3204 (O_3204,N_29607,N_28996);
nand UO_3205 (O_3205,N_29538,N_28182);
xnor UO_3206 (O_3206,N_28087,N_29682);
nand UO_3207 (O_3207,N_29020,N_28333);
and UO_3208 (O_3208,N_29719,N_28470);
nor UO_3209 (O_3209,N_29036,N_29791);
nor UO_3210 (O_3210,N_29005,N_28888);
nand UO_3211 (O_3211,N_29420,N_29684);
xnor UO_3212 (O_3212,N_28768,N_28054);
nand UO_3213 (O_3213,N_28162,N_28158);
and UO_3214 (O_3214,N_29962,N_29226);
or UO_3215 (O_3215,N_29504,N_28488);
nand UO_3216 (O_3216,N_29297,N_28357);
xnor UO_3217 (O_3217,N_29854,N_28847);
or UO_3218 (O_3218,N_29964,N_28542);
and UO_3219 (O_3219,N_28023,N_29943);
or UO_3220 (O_3220,N_28199,N_29289);
or UO_3221 (O_3221,N_28136,N_28708);
xnor UO_3222 (O_3222,N_29524,N_28248);
or UO_3223 (O_3223,N_29691,N_28854);
nor UO_3224 (O_3224,N_29406,N_29912);
nor UO_3225 (O_3225,N_28169,N_29101);
nor UO_3226 (O_3226,N_29757,N_29704);
nor UO_3227 (O_3227,N_28192,N_29312);
nor UO_3228 (O_3228,N_28508,N_29506);
and UO_3229 (O_3229,N_28983,N_29068);
xnor UO_3230 (O_3230,N_29158,N_29147);
or UO_3231 (O_3231,N_28137,N_28837);
or UO_3232 (O_3232,N_29684,N_29568);
nand UO_3233 (O_3233,N_29017,N_29158);
xor UO_3234 (O_3234,N_28786,N_29132);
or UO_3235 (O_3235,N_28313,N_29121);
xnor UO_3236 (O_3236,N_28169,N_28847);
and UO_3237 (O_3237,N_28883,N_29980);
nor UO_3238 (O_3238,N_28782,N_29240);
nand UO_3239 (O_3239,N_29831,N_29704);
or UO_3240 (O_3240,N_28419,N_29689);
nand UO_3241 (O_3241,N_29297,N_29827);
nand UO_3242 (O_3242,N_28325,N_29976);
nand UO_3243 (O_3243,N_29869,N_28170);
xnor UO_3244 (O_3244,N_28385,N_29994);
xor UO_3245 (O_3245,N_29693,N_28635);
xor UO_3246 (O_3246,N_28773,N_29523);
or UO_3247 (O_3247,N_28158,N_28728);
or UO_3248 (O_3248,N_28581,N_28140);
and UO_3249 (O_3249,N_28366,N_29474);
nand UO_3250 (O_3250,N_29835,N_29126);
xnor UO_3251 (O_3251,N_29375,N_28417);
xnor UO_3252 (O_3252,N_29088,N_28326);
nor UO_3253 (O_3253,N_28923,N_28379);
nor UO_3254 (O_3254,N_29184,N_29298);
xor UO_3255 (O_3255,N_29548,N_29603);
and UO_3256 (O_3256,N_29900,N_28413);
nor UO_3257 (O_3257,N_29246,N_28888);
or UO_3258 (O_3258,N_29325,N_28003);
or UO_3259 (O_3259,N_29703,N_29751);
and UO_3260 (O_3260,N_29543,N_29124);
nand UO_3261 (O_3261,N_28095,N_28336);
xnor UO_3262 (O_3262,N_28889,N_29895);
and UO_3263 (O_3263,N_28471,N_29120);
or UO_3264 (O_3264,N_29249,N_28711);
xnor UO_3265 (O_3265,N_29758,N_29525);
and UO_3266 (O_3266,N_29932,N_29723);
nor UO_3267 (O_3267,N_28662,N_28056);
or UO_3268 (O_3268,N_28655,N_29842);
xor UO_3269 (O_3269,N_29533,N_29072);
xnor UO_3270 (O_3270,N_29912,N_28261);
nand UO_3271 (O_3271,N_29549,N_29604);
nand UO_3272 (O_3272,N_28152,N_29559);
or UO_3273 (O_3273,N_28585,N_28404);
or UO_3274 (O_3274,N_28853,N_29606);
nand UO_3275 (O_3275,N_29968,N_28335);
nand UO_3276 (O_3276,N_28225,N_28001);
and UO_3277 (O_3277,N_29801,N_29291);
or UO_3278 (O_3278,N_28744,N_28547);
or UO_3279 (O_3279,N_29047,N_28771);
nor UO_3280 (O_3280,N_29780,N_29059);
nor UO_3281 (O_3281,N_28107,N_28412);
nor UO_3282 (O_3282,N_28885,N_29048);
nor UO_3283 (O_3283,N_29557,N_29875);
nand UO_3284 (O_3284,N_29867,N_29806);
nand UO_3285 (O_3285,N_29458,N_28864);
xnor UO_3286 (O_3286,N_28171,N_28300);
nand UO_3287 (O_3287,N_28842,N_28157);
and UO_3288 (O_3288,N_29367,N_28192);
or UO_3289 (O_3289,N_28622,N_29094);
nand UO_3290 (O_3290,N_28507,N_28712);
nor UO_3291 (O_3291,N_28945,N_28999);
nand UO_3292 (O_3292,N_28949,N_28953);
and UO_3293 (O_3293,N_29538,N_28465);
nand UO_3294 (O_3294,N_28160,N_28082);
and UO_3295 (O_3295,N_28294,N_29933);
nand UO_3296 (O_3296,N_29657,N_28957);
or UO_3297 (O_3297,N_29558,N_29131);
xor UO_3298 (O_3298,N_28178,N_29557);
nor UO_3299 (O_3299,N_29923,N_29025);
nand UO_3300 (O_3300,N_28059,N_28223);
and UO_3301 (O_3301,N_28038,N_28209);
nand UO_3302 (O_3302,N_29888,N_28470);
nor UO_3303 (O_3303,N_29286,N_28630);
or UO_3304 (O_3304,N_28158,N_29547);
and UO_3305 (O_3305,N_28019,N_28677);
xnor UO_3306 (O_3306,N_29680,N_28345);
nand UO_3307 (O_3307,N_28112,N_29788);
or UO_3308 (O_3308,N_29628,N_28416);
nor UO_3309 (O_3309,N_28855,N_29386);
nor UO_3310 (O_3310,N_29222,N_29839);
nor UO_3311 (O_3311,N_28421,N_28723);
or UO_3312 (O_3312,N_28081,N_29301);
nor UO_3313 (O_3313,N_29768,N_28802);
nand UO_3314 (O_3314,N_29634,N_29183);
and UO_3315 (O_3315,N_28035,N_29652);
xnor UO_3316 (O_3316,N_29446,N_28426);
nor UO_3317 (O_3317,N_29144,N_28297);
xor UO_3318 (O_3318,N_28627,N_28965);
and UO_3319 (O_3319,N_28169,N_29528);
nand UO_3320 (O_3320,N_29193,N_29900);
nor UO_3321 (O_3321,N_29762,N_28164);
nand UO_3322 (O_3322,N_29266,N_28605);
or UO_3323 (O_3323,N_28782,N_28703);
or UO_3324 (O_3324,N_29112,N_29183);
nand UO_3325 (O_3325,N_29596,N_29613);
nand UO_3326 (O_3326,N_28176,N_28471);
or UO_3327 (O_3327,N_28573,N_28816);
and UO_3328 (O_3328,N_28286,N_28092);
nand UO_3329 (O_3329,N_29118,N_29894);
and UO_3330 (O_3330,N_28720,N_29185);
nand UO_3331 (O_3331,N_29493,N_28470);
and UO_3332 (O_3332,N_28324,N_28635);
and UO_3333 (O_3333,N_29549,N_28625);
nor UO_3334 (O_3334,N_29855,N_28436);
or UO_3335 (O_3335,N_29258,N_29762);
or UO_3336 (O_3336,N_29139,N_28533);
or UO_3337 (O_3337,N_29475,N_28668);
nand UO_3338 (O_3338,N_28413,N_29827);
xnor UO_3339 (O_3339,N_29001,N_29041);
xor UO_3340 (O_3340,N_29824,N_29332);
nand UO_3341 (O_3341,N_28394,N_28345);
and UO_3342 (O_3342,N_28645,N_29321);
and UO_3343 (O_3343,N_28710,N_28217);
or UO_3344 (O_3344,N_28317,N_29091);
xor UO_3345 (O_3345,N_28906,N_29868);
or UO_3346 (O_3346,N_29184,N_28559);
xnor UO_3347 (O_3347,N_29134,N_29496);
and UO_3348 (O_3348,N_29684,N_29411);
xor UO_3349 (O_3349,N_29136,N_29624);
and UO_3350 (O_3350,N_28959,N_28824);
nor UO_3351 (O_3351,N_28788,N_28616);
nand UO_3352 (O_3352,N_29931,N_28346);
xnor UO_3353 (O_3353,N_28469,N_29614);
nor UO_3354 (O_3354,N_29314,N_28958);
nor UO_3355 (O_3355,N_28294,N_28520);
xor UO_3356 (O_3356,N_28907,N_28347);
and UO_3357 (O_3357,N_28620,N_29666);
and UO_3358 (O_3358,N_29923,N_29566);
or UO_3359 (O_3359,N_29631,N_29997);
xnor UO_3360 (O_3360,N_28388,N_28154);
nor UO_3361 (O_3361,N_28344,N_29246);
nand UO_3362 (O_3362,N_29676,N_29142);
xnor UO_3363 (O_3363,N_29241,N_28417);
xor UO_3364 (O_3364,N_28870,N_28980);
nand UO_3365 (O_3365,N_29117,N_28047);
and UO_3366 (O_3366,N_28004,N_29788);
nor UO_3367 (O_3367,N_29155,N_28885);
nand UO_3368 (O_3368,N_28015,N_29967);
or UO_3369 (O_3369,N_29961,N_28807);
xor UO_3370 (O_3370,N_28799,N_29795);
and UO_3371 (O_3371,N_28792,N_28797);
and UO_3372 (O_3372,N_29454,N_28356);
and UO_3373 (O_3373,N_28704,N_28395);
and UO_3374 (O_3374,N_29831,N_29978);
and UO_3375 (O_3375,N_29367,N_28290);
and UO_3376 (O_3376,N_28080,N_28546);
nor UO_3377 (O_3377,N_29018,N_28813);
nor UO_3378 (O_3378,N_29323,N_29112);
or UO_3379 (O_3379,N_28221,N_29645);
or UO_3380 (O_3380,N_28842,N_28629);
and UO_3381 (O_3381,N_28724,N_29173);
xor UO_3382 (O_3382,N_28969,N_28192);
nor UO_3383 (O_3383,N_28622,N_28802);
xnor UO_3384 (O_3384,N_28397,N_29367);
and UO_3385 (O_3385,N_28669,N_28998);
nor UO_3386 (O_3386,N_29237,N_29187);
nor UO_3387 (O_3387,N_28729,N_28824);
xor UO_3388 (O_3388,N_29411,N_28244);
nor UO_3389 (O_3389,N_28342,N_29349);
and UO_3390 (O_3390,N_28582,N_29190);
xnor UO_3391 (O_3391,N_29850,N_29142);
and UO_3392 (O_3392,N_28836,N_29265);
xor UO_3393 (O_3393,N_28296,N_29297);
nor UO_3394 (O_3394,N_29413,N_28519);
and UO_3395 (O_3395,N_28839,N_29429);
xor UO_3396 (O_3396,N_29433,N_28267);
or UO_3397 (O_3397,N_29512,N_29451);
nor UO_3398 (O_3398,N_28762,N_29930);
nand UO_3399 (O_3399,N_29274,N_28109);
or UO_3400 (O_3400,N_28482,N_29560);
nor UO_3401 (O_3401,N_29160,N_29356);
and UO_3402 (O_3402,N_28009,N_28570);
or UO_3403 (O_3403,N_29691,N_29909);
xor UO_3404 (O_3404,N_29899,N_29657);
xor UO_3405 (O_3405,N_29722,N_29005);
and UO_3406 (O_3406,N_28674,N_28760);
nand UO_3407 (O_3407,N_29318,N_29615);
xnor UO_3408 (O_3408,N_28161,N_29316);
nand UO_3409 (O_3409,N_29575,N_28515);
xor UO_3410 (O_3410,N_28029,N_28481);
xor UO_3411 (O_3411,N_28294,N_29193);
nand UO_3412 (O_3412,N_29403,N_29854);
nand UO_3413 (O_3413,N_29180,N_29607);
xor UO_3414 (O_3414,N_28406,N_28123);
or UO_3415 (O_3415,N_28943,N_29388);
nor UO_3416 (O_3416,N_28654,N_28238);
nor UO_3417 (O_3417,N_28002,N_29602);
or UO_3418 (O_3418,N_29026,N_29928);
or UO_3419 (O_3419,N_28599,N_29879);
and UO_3420 (O_3420,N_28647,N_28937);
nand UO_3421 (O_3421,N_28734,N_28614);
xor UO_3422 (O_3422,N_29574,N_28355);
and UO_3423 (O_3423,N_29569,N_28687);
nor UO_3424 (O_3424,N_28403,N_29192);
xor UO_3425 (O_3425,N_28348,N_29268);
nand UO_3426 (O_3426,N_28008,N_28974);
and UO_3427 (O_3427,N_28608,N_29411);
nand UO_3428 (O_3428,N_29040,N_28675);
xor UO_3429 (O_3429,N_29926,N_28076);
or UO_3430 (O_3430,N_28941,N_29554);
nor UO_3431 (O_3431,N_28908,N_28112);
nor UO_3432 (O_3432,N_28021,N_28870);
or UO_3433 (O_3433,N_29470,N_28947);
and UO_3434 (O_3434,N_29933,N_28005);
xor UO_3435 (O_3435,N_28672,N_28913);
nor UO_3436 (O_3436,N_28396,N_29229);
xor UO_3437 (O_3437,N_28097,N_28936);
nor UO_3438 (O_3438,N_29582,N_29775);
and UO_3439 (O_3439,N_29696,N_28340);
and UO_3440 (O_3440,N_28160,N_28578);
nand UO_3441 (O_3441,N_29326,N_29120);
nand UO_3442 (O_3442,N_29474,N_29588);
nor UO_3443 (O_3443,N_28129,N_28084);
xnor UO_3444 (O_3444,N_28042,N_29367);
and UO_3445 (O_3445,N_28180,N_28750);
and UO_3446 (O_3446,N_28920,N_29603);
or UO_3447 (O_3447,N_29233,N_28016);
xor UO_3448 (O_3448,N_28128,N_28843);
xnor UO_3449 (O_3449,N_29825,N_29684);
nand UO_3450 (O_3450,N_29874,N_28715);
nor UO_3451 (O_3451,N_28688,N_29986);
or UO_3452 (O_3452,N_28113,N_29456);
nor UO_3453 (O_3453,N_29788,N_29078);
nand UO_3454 (O_3454,N_28371,N_28989);
or UO_3455 (O_3455,N_29325,N_29939);
and UO_3456 (O_3456,N_29574,N_28432);
nand UO_3457 (O_3457,N_29543,N_28394);
or UO_3458 (O_3458,N_29923,N_28862);
nor UO_3459 (O_3459,N_29052,N_29867);
nand UO_3460 (O_3460,N_29013,N_29470);
and UO_3461 (O_3461,N_29496,N_28345);
and UO_3462 (O_3462,N_29308,N_29329);
and UO_3463 (O_3463,N_29895,N_28464);
nand UO_3464 (O_3464,N_29414,N_29046);
nor UO_3465 (O_3465,N_28036,N_29166);
nor UO_3466 (O_3466,N_28780,N_28562);
xor UO_3467 (O_3467,N_29961,N_28155);
nor UO_3468 (O_3468,N_29474,N_28127);
nand UO_3469 (O_3469,N_28231,N_29801);
nor UO_3470 (O_3470,N_29511,N_29809);
or UO_3471 (O_3471,N_28591,N_28074);
xnor UO_3472 (O_3472,N_28978,N_28046);
nand UO_3473 (O_3473,N_28055,N_28698);
nand UO_3474 (O_3474,N_28650,N_28049);
xnor UO_3475 (O_3475,N_28793,N_28241);
or UO_3476 (O_3476,N_29147,N_29709);
nor UO_3477 (O_3477,N_29846,N_29575);
and UO_3478 (O_3478,N_28136,N_29513);
xnor UO_3479 (O_3479,N_29133,N_29062);
and UO_3480 (O_3480,N_28287,N_28324);
nor UO_3481 (O_3481,N_28353,N_29908);
nand UO_3482 (O_3482,N_29669,N_29446);
nand UO_3483 (O_3483,N_29279,N_28099);
xor UO_3484 (O_3484,N_28389,N_29882);
nand UO_3485 (O_3485,N_29580,N_29405);
and UO_3486 (O_3486,N_29936,N_28365);
nor UO_3487 (O_3487,N_28706,N_28420);
xnor UO_3488 (O_3488,N_29709,N_28697);
nor UO_3489 (O_3489,N_29189,N_28665);
xnor UO_3490 (O_3490,N_28041,N_29282);
nand UO_3491 (O_3491,N_29046,N_28875);
nand UO_3492 (O_3492,N_28817,N_28610);
nand UO_3493 (O_3493,N_28658,N_29070);
nand UO_3494 (O_3494,N_28750,N_29841);
xnor UO_3495 (O_3495,N_28555,N_28642);
xor UO_3496 (O_3496,N_29371,N_29147);
nor UO_3497 (O_3497,N_29393,N_29666);
xor UO_3498 (O_3498,N_29940,N_28202);
xor UO_3499 (O_3499,N_29465,N_29605);
endmodule