module basic_3000_30000_3500_15_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_1757,In_1972);
or U1 (N_1,In_1515,In_9);
nor U2 (N_2,In_422,In_579);
and U3 (N_3,In_1730,In_1268);
xor U4 (N_4,In_643,In_2744);
xnor U5 (N_5,In_2097,In_1829);
or U6 (N_6,In_2459,In_1255);
nor U7 (N_7,In_2855,In_2467);
nor U8 (N_8,In_2195,In_2548);
and U9 (N_9,In_2935,In_532);
nand U10 (N_10,In_1729,In_240);
or U11 (N_11,In_897,In_1622);
xnor U12 (N_12,In_1296,In_2342);
or U13 (N_13,In_1576,In_2835);
nor U14 (N_14,In_404,In_1173);
xor U15 (N_15,In_2767,In_233);
or U16 (N_16,In_2565,In_1837);
nor U17 (N_17,In_2185,In_2849);
nand U18 (N_18,In_1441,In_889);
and U19 (N_19,In_200,In_2899);
nor U20 (N_20,In_2211,In_392);
and U21 (N_21,In_1615,In_2666);
or U22 (N_22,In_2073,In_5);
and U23 (N_23,In_1625,In_2668);
nand U24 (N_24,In_1049,In_1984);
xnor U25 (N_25,In_309,In_2074);
xor U26 (N_26,In_1097,In_694);
nand U27 (N_27,In_1697,In_2594);
nand U28 (N_28,In_1880,In_1273);
xor U29 (N_29,In_1994,In_1955);
or U30 (N_30,In_2407,In_1485);
xnor U31 (N_31,In_2939,In_2660);
or U32 (N_32,In_2811,In_349);
and U33 (N_33,In_1127,In_443);
or U34 (N_34,In_2154,In_890);
and U35 (N_35,In_2403,In_1764);
nand U36 (N_36,In_102,In_1639);
or U37 (N_37,In_1967,In_2724);
and U38 (N_38,In_2485,In_1353);
or U39 (N_39,In_1520,In_263);
or U40 (N_40,In_1461,In_608);
nor U41 (N_41,In_2115,In_1487);
nor U42 (N_42,In_110,In_291);
and U43 (N_43,In_2947,In_1096);
nor U44 (N_44,In_2450,In_1653);
and U45 (N_45,In_1069,In_1936);
nand U46 (N_46,In_1449,In_356);
nand U47 (N_47,In_1166,In_2542);
nor U48 (N_48,In_256,In_316);
nand U49 (N_49,In_1411,In_2863);
xnor U50 (N_50,In_695,In_2901);
and U51 (N_51,In_1995,In_1738);
xnor U52 (N_52,In_963,In_375);
nor U53 (N_53,In_140,In_506);
xnor U54 (N_54,In_419,In_565);
xor U55 (N_55,In_2628,In_1116);
and U56 (N_56,In_846,In_2302);
nand U57 (N_57,In_571,In_2974);
or U58 (N_58,In_2694,In_1122);
nor U59 (N_59,In_207,In_2933);
nor U60 (N_60,In_1215,In_2975);
and U61 (N_61,In_2103,In_2556);
nor U62 (N_62,In_1529,In_1157);
nand U63 (N_63,In_1246,In_1134);
nand U64 (N_64,In_73,In_2189);
xor U65 (N_65,In_2824,In_71);
xnor U66 (N_66,In_642,In_59);
and U67 (N_67,In_307,In_1075);
and U68 (N_68,In_1964,In_1312);
xor U69 (N_69,In_231,In_330);
nand U70 (N_70,In_1684,In_1516);
nor U71 (N_71,In_1928,In_2969);
and U72 (N_72,In_2704,In_2807);
xor U73 (N_73,In_876,In_406);
and U74 (N_74,In_317,In_1045);
nor U75 (N_75,In_1490,In_798);
nand U76 (N_76,In_1798,In_1720);
xor U77 (N_77,In_2150,In_1915);
or U78 (N_78,In_235,In_1715);
or U79 (N_79,In_2310,In_1250);
and U80 (N_80,In_2952,In_2294);
or U81 (N_81,In_282,In_790);
and U82 (N_82,In_629,In_2845);
xnor U83 (N_83,In_1094,In_2481);
or U84 (N_84,In_97,In_1556);
nor U85 (N_85,In_2327,In_2651);
or U86 (N_86,In_2573,In_1130);
nor U87 (N_87,In_2910,In_638);
or U88 (N_88,In_938,In_2924);
and U89 (N_89,In_1547,In_450);
xor U90 (N_90,In_2945,In_2402);
and U91 (N_91,In_1532,In_2198);
xor U92 (N_92,In_2854,In_2546);
xor U93 (N_93,In_89,In_1396);
xnor U94 (N_94,In_1554,In_1488);
and U95 (N_95,In_2775,In_700);
xnor U96 (N_96,In_2822,In_816);
or U97 (N_97,In_388,In_1092);
or U98 (N_98,In_734,In_1227);
nand U99 (N_99,In_1111,In_1119);
or U100 (N_100,In_2898,In_430);
nor U101 (N_101,In_594,In_1793);
nand U102 (N_102,In_2196,In_2003);
and U103 (N_103,In_1899,In_1063);
nor U104 (N_104,In_2606,In_2426);
nand U105 (N_105,In_1950,In_2337);
xnor U106 (N_106,In_1983,In_2142);
nor U107 (N_107,In_2048,In_301);
nand U108 (N_108,In_2042,In_2858);
nor U109 (N_109,In_237,In_1067);
or U110 (N_110,In_1229,In_2970);
xnor U111 (N_111,In_2068,In_394);
nand U112 (N_112,In_280,In_504);
nand U113 (N_113,In_755,In_1608);
xnor U114 (N_114,In_150,In_2569);
nor U115 (N_115,In_455,In_198);
and U116 (N_116,In_1402,In_1618);
nand U117 (N_117,In_515,In_1714);
xnor U118 (N_118,In_1536,In_645);
nor U119 (N_119,In_473,In_1679);
nand U120 (N_120,In_329,In_261);
nand U121 (N_121,In_739,In_1176);
nor U122 (N_122,In_332,In_2997);
xor U123 (N_123,In_2033,In_2754);
nand U124 (N_124,In_1013,In_635);
nand U125 (N_125,In_2750,In_2380);
nand U126 (N_126,In_128,In_1648);
nor U127 (N_127,In_533,In_1438);
and U128 (N_128,In_2543,In_2298);
and U129 (N_129,In_1235,In_1373);
nand U130 (N_130,In_1976,In_1628);
nand U131 (N_131,In_1104,In_715);
xor U132 (N_132,In_221,In_2108);
nand U133 (N_133,In_2953,In_618);
and U134 (N_134,In_397,In_2813);
and U135 (N_135,In_1315,In_2167);
or U136 (N_136,In_2535,In_2549);
nand U137 (N_137,In_1643,In_575);
xor U138 (N_138,In_988,In_1454);
nand U139 (N_139,In_1718,In_2504);
nor U140 (N_140,In_475,In_288);
xor U141 (N_141,In_1511,In_478);
xor U142 (N_142,In_2879,In_2741);
or U143 (N_143,In_401,In_2261);
and U144 (N_144,In_713,In_2165);
or U145 (N_145,In_292,In_1813);
xnor U146 (N_146,In_797,In_610);
nand U147 (N_147,In_2179,In_290);
xor U148 (N_148,In_869,In_2597);
or U149 (N_149,In_820,In_2494);
nand U150 (N_150,In_66,In_1699);
nand U151 (N_151,In_636,In_1541);
nand U152 (N_152,In_2954,In_60);
xnor U153 (N_153,In_343,In_2508);
or U154 (N_154,In_298,In_666);
nor U155 (N_155,In_2739,In_452);
or U156 (N_156,In_314,In_108);
nor U157 (N_157,In_2518,In_1420);
nand U158 (N_158,In_1783,In_612);
nor U159 (N_159,In_593,In_2471);
nor U160 (N_160,In_2759,In_348);
or U161 (N_161,In_94,In_402);
nand U162 (N_162,In_2453,In_2787);
nand U163 (N_163,In_832,In_400);
nor U164 (N_164,In_2695,In_250);
nand U165 (N_165,In_468,In_481);
and U166 (N_166,In_1614,In_720);
or U167 (N_167,In_2778,In_2237);
and U168 (N_168,In_2032,In_2647);
nor U169 (N_169,In_948,In_2979);
nor U170 (N_170,In_1430,In_1211);
xnor U171 (N_171,In_366,In_1878);
and U172 (N_172,In_1076,In_1642);
or U173 (N_173,In_2591,In_2506);
nand U174 (N_174,In_95,In_1961);
xnor U175 (N_175,In_2434,In_433);
nor U176 (N_176,In_852,In_2877);
nand U177 (N_177,In_538,In_998);
xor U178 (N_178,In_2644,In_2375);
nor U179 (N_179,In_802,In_2861);
xor U180 (N_180,In_737,In_751);
and U181 (N_181,In_791,In_1392);
nand U182 (N_182,In_34,In_717);
or U183 (N_183,In_177,In_973);
nor U184 (N_184,In_1299,In_2214);
xor U185 (N_185,In_777,In_31);
nand U186 (N_186,In_1681,In_1318);
nor U187 (N_187,In_2550,In_1985);
nand U188 (N_188,In_1065,In_892);
or U189 (N_189,In_1968,In_1589);
xor U190 (N_190,In_2273,In_1140);
or U191 (N_191,In_2137,In_2119);
nand U192 (N_192,In_1393,In_1136);
or U193 (N_193,In_2981,In_1897);
nor U194 (N_194,In_752,In_2987);
or U195 (N_195,In_943,In_1858);
or U196 (N_196,In_1031,In_2101);
and U197 (N_197,In_238,In_1560);
nor U198 (N_198,In_2100,In_2642);
nor U199 (N_199,In_1760,In_1182);
and U200 (N_200,In_223,In_42);
nor U201 (N_201,In_2886,In_479);
or U202 (N_202,In_1371,In_2492);
nand U203 (N_203,In_1241,In_1727);
and U204 (N_204,In_2713,In_2392);
or U205 (N_205,In_1361,In_813);
xnor U206 (N_206,In_113,In_1933);
or U207 (N_207,In_2014,In_2900);
and U208 (N_208,In_2932,In_1394);
and U209 (N_209,In_1131,In_2571);
xor U210 (N_210,In_849,In_1501);
and U211 (N_211,In_1350,In_1991);
or U212 (N_212,In_1342,In_1217);
nand U213 (N_213,In_74,In_2602);
nor U214 (N_214,In_1053,In_1307);
nor U215 (N_215,In_1794,In_1975);
nor U216 (N_216,In_2430,In_28);
xnor U217 (N_217,In_143,In_2574);
nor U218 (N_218,In_2911,In_2373);
nand U219 (N_219,In_1708,In_744);
xor U220 (N_220,In_1455,In_2605);
nand U221 (N_221,In_531,In_1113);
or U222 (N_222,In_347,In_2645);
xor U223 (N_223,In_2278,In_1051);
or U224 (N_224,In_2120,In_2816);
or U225 (N_225,In_1934,In_365);
or U226 (N_226,In_139,In_1030);
or U227 (N_227,In_270,In_2624);
or U228 (N_228,In_771,In_1978);
nand U229 (N_229,In_2451,In_2307);
nand U230 (N_230,In_1670,In_85);
and U231 (N_231,In_20,In_2468);
or U232 (N_232,In_969,In_2993);
nand U233 (N_233,In_1374,In_1322);
nand U234 (N_234,In_1460,In_2285);
or U235 (N_235,In_2919,In_2681);
nor U236 (N_236,In_2288,In_2245);
nand U237 (N_237,In_2643,In_1224);
nand U238 (N_238,In_1190,In_1663);
xnor U239 (N_239,In_2149,In_663);
xnor U240 (N_240,In_1707,In_1973);
or U241 (N_241,In_1337,In_1918);
and U242 (N_242,In_1081,In_1925);
nand U243 (N_243,In_2332,In_2331);
or U244 (N_244,In_2062,In_1930);
nor U245 (N_245,In_2821,In_451);
nand U246 (N_246,In_2809,In_1220);
nor U247 (N_247,In_159,In_1167);
or U248 (N_248,In_1291,In_617);
and U249 (N_249,In_134,In_384);
xnor U250 (N_250,In_287,In_1204);
and U251 (N_251,In_1805,In_16);
xnor U252 (N_252,In_606,In_1476);
xor U253 (N_253,In_2353,In_1249);
xor U254 (N_254,In_976,In_583);
xor U255 (N_255,In_1875,In_1877);
or U256 (N_256,In_227,In_1348);
and U257 (N_257,In_417,In_1555);
xor U258 (N_258,In_1201,In_1789);
and U259 (N_259,In_1772,In_913);
nand U260 (N_260,In_427,In_1752);
nor U261 (N_261,In_500,In_1905);
and U262 (N_262,In_2072,In_996);
and U263 (N_263,In_1719,In_619);
or U264 (N_264,In_2841,In_1710);
nand U265 (N_265,In_589,In_1470);
or U266 (N_266,In_1381,In_493);
nor U267 (N_267,In_800,In_632);
and U268 (N_268,In_2792,In_118);
or U269 (N_269,In_2143,In_462);
xor U270 (N_270,In_242,In_949);
or U271 (N_271,In_197,In_2473);
nor U272 (N_272,In_144,In_1468);
nand U273 (N_273,In_1050,In_1629);
nand U274 (N_274,In_2665,In_2210);
xnor U275 (N_275,In_2613,In_115);
nand U276 (N_276,In_1799,In_665);
nor U277 (N_277,In_2520,In_2366);
and U278 (N_278,In_600,In_2322);
or U279 (N_279,In_2415,In_1557);
xor U280 (N_280,In_681,In_580);
or U281 (N_281,In_1304,In_1288);
xnor U282 (N_282,In_1916,In_458);
xor U283 (N_283,In_1329,In_1620);
xor U284 (N_284,In_385,In_631);
and U285 (N_285,In_2561,In_1607);
nand U286 (N_286,In_1538,In_2908);
nor U287 (N_287,In_2880,In_219);
nand U288 (N_288,In_1351,In_382);
and U289 (N_289,In_459,In_810);
nor U290 (N_290,In_561,In_2140);
nand U291 (N_291,In_1982,In_560);
or U292 (N_292,In_2055,In_611);
nand U293 (N_293,In_1635,In_1324);
xnor U294 (N_294,In_2918,In_1769);
nand U295 (N_295,In_1844,In_1827);
nand U296 (N_296,In_878,In_1841);
and U297 (N_297,In_2277,In_1997);
nand U298 (N_298,In_376,In_2840);
or U299 (N_299,In_1510,In_1347);
xor U300 (N_300,In_2823,In_2669);
and U301 (N_301,In_1726,In_2495);
xnor U302 (N_302,In_379,In_1832);
and U303 (N_303,In_1222,In_1514);
nor U304 (N_304,In_2354,In_360);
nand U305 (N_305,In_350,In_2563);
nand U306 (N_306,In_2769,In_2102);
nor U307 (N_307,In_2304,In_1019);
nand U308 (N_308,In_2007,In_858);
and U309 (N_309,In_2685,In_1723);
nand U310 (N_310,In_1422,In_2566);
or U311 (N_311,In_733,In_1571);
and U312 (N_312,In_906,In_123);
or U313 (N_313,In_1363,In_626);
nor U314 (N_314,In_1427,In_1894);
nor U315 (N_315,In_182,In_2675);
or U316 (N_316,In_1344,In_559);
nor U317 (N_317,In_1782,In_2343);
nand U318 (N_318,In_2967,In_648);
or U319 (N_319,In_2346,In_2552);
nand U320 (N_320,In_1044,In_2820);
xor U321 (N_321,In_770,In_2976);
nand U322 (N_322,In_604,In_1314);
or U323 (N_323,In_961,In_1284);
and U324 (N_324,In_758,In_12);
xor U325 (N_325,In_2173,In_1248);
nor U326 (N_326,In_148,In_1262);
nand U327 (N_327,In_1009,In_731);
nand U328 (N_328,In_1289,In_1587);
nand U329 (N_329,In_2251,In_1154);
nand U330 (N_330,In_1518,In_793);
and U331 (N_331,In_1179,In_2184);
nor U332 (N_332,In_1036,In_1156);
nand U333 (N_333,In_2096,In_336);
or U334 (N_334,In_225,In_705);
nand U335 (N_335,In_1594,In_2377);
nand U336 (N_336,In_1777,In_2087);
nand U337 (N_337,In_2972,In_2590);
xor U338 (N_338,In_2512,In_369);
or U339 (N_339,In_2837,In_2758);
or U340 (N_340,In_1264,In_2648);
and U341 (N_341,In_2162,In_2254);
or U342 (N_342,In_602,In_466);
nand U343 (N_343,In_480,In_1038);
nor U344 (N_344,In_726,In_1466);
or U345 (N_345,In_985,In_2742);
nor U346 (N_346,In_2784,In_2333);
or U347 (N_347,In_2361,In_1785);
xnor U348 (N_348,In_2051,In_2439);
or U349 (N_349,In_2397,In_2236);
nand U350 (N_350,In_2301,In_2045);
nand U351 (N_351,In_2844,In_625);
nand U352 (N_352,In_2351,In_264);
and U353 (N_353,In_2640,In_683);
and U354 (N_354,In_310,In_2313);
nor U355 (N_355,In_2129,In_1535);
xor U356 (N_356,In_2768,In_529);
and U357 (N_357,In_185,In_1048);
nand U358 (N_358,In_80,In_476);
and U359 (N_359,In_7,In_76);
nor U360 (N_360,In_2623,In_68);
nor U361 (N_361,In_2818,In_535);
and U362 (N_362,In_411,In_562);
xor U363 (N_363,In_135,In_1900);
nor U364 (N_364,In_2276,In_324);
and U365 (N_365,In_1502,In_1482);
and U366 (N_366,In_1701,In_1958);
nand U367 (N_367,In_886,In_2866);
nor U368 (N_368,In_1109,In_2282);
xor U369 (N_369,In_2169,In_2131);
nor U370 (N_370,In_173,In_2183);
nor U371 (N_371,In_860,In_1472);
or U372 (N_372,In_2308,In_1237);
and U373 (N_373,In_2336,In_1850);
and U374 (N_374,In_1064,In_2369);
nand U375 (N_375,In_35,In_1613);
or U376 (N_376,In_260,In_2796);
and U377 (N_377,In_1767,In_1566);
or U378 (N_378,In_2257,In_346);
nor U379 (N_379,In_1512,In_1114);
and U380 (N_380,In_2725,In_2622);
or U381 (N_381,In_2163,In_1459);
nand U382 (N_382,In_454,In_1093);
or U383 (N_383,In_2412,In_2729);
and U384 (N_384,In_1115,In_552);
and U385 (N_385,In_2540,In_440);
nand U386 (N_386,In_1839,In_161);
nor U387 (N_387,In_1882,In_370);
xnor U388 (N_388,In_2335,In_1671);
xor U389 (N_389,In_2255,In_2496);
and U390 (N_390,In_1887,In_1610);
nand U391 (N_391,In_1024,In_2612);
nand U392 (N_392,In_1243,In_2180);
or U393 (N_393,In_966,In_885);
or U394 (N_394,In_1469,In_274);
nand U395 (N_395,In_2509,In_101);
or U396 (N_396,In_2136,In_657);
nand U397 (N_397,In_2580,In_971);
or U398 (N_398,In_1879,In_2241);
nand U399 (N_399,In_1377,In_2851);
xnor U400 (N_400,In_2625,In_2719);
or U401 (N_401,In_2583,In_1216);
or U402 (N_402,In_2395,In_2526);
and U403 (N_403,In_226,In_447);
nand U404 (N_404,In_2105,In_1749);
or U405 (N_405,In_2349,In_1549);
nand U406 (N_406,In_2986,In_684);
or U407 (N_407,In_1517,In_1604);
xor U408 (N_408,In_2530,In_1132);
nor U409 (N_409,In_2368,In_1745);
xnor U410 (N_410,In_2128,In_434);
xor U411 (N_411,In_54,In_863);
xnor U412 (N_412,In_2921,In_2872);
nor U413 (N_413,In_916,In_2890);
or U414 (N_414,In_2348,In_2572);
or U415 (N_415,In_257,In_753);
nand U416 (N_416,In_1825,In_1807);
xnor U417 (N_417,In_2005,In_774);
nand U418 (N_418,In_2867,In_1254);
or U419 (N_419,In_120,In_549);
nand U420 (N_420,In_2607,In_105);
and U421 (N_421,In_1765,In_2035);
nor U422 (N_422,In_895,In_658);
nor U423 (N_423,In_748,In_659);
nand U424 (N_424,In_2040,In_2270);
xnor U425 (N_425,In_1090,In_1939);
or U426 (N_426,In_599,In_1695);
or U427 (N_427,In_546,In_2130);
nand U428 (N_428,In_912,In_127);
nand U429 (N_429,In_175,In_1509);
nor U430 (N_430,In_1321,In_2553);
xnor U431 (N_431,In_928,In_1378);
nand U432 (N_432,In_2079,In_2931);
nand U433 (N_433,In_934,In_429);
xnor U434 (N_434,In_1101,In_30);
nor U435 (N_435,In_1654,In_2155);
xor U436 (N_436,In_1100,In_1453);
xor U437 (N_437,In_2186,In_2983);
or U438 (N_438,In_980,In_2751);
nor U439 (N_439,In_1874,In_1492);
xor U440 (N_440,In_2021,In_2325);
nor U441 (N_441,In_843,In_2075);
nand U442 (N_442,In_1406,In_1369);
nor U443 (N_443,In_24,In_2896);
and U444 (N_444,In_1685,In_1938);
nor U445 (N_445,In_192,In_209);
and U446 (N_446,In_1595,In_1742);
nor U447 (N_447,In_981,In_1062);
nand U448 (N_448,In_1303,In_2959);
and U449 (N_449,In_2515,In_1848);
or U450 (N_450,In_2118,In_2437);
nand U451 (N_451,In_2047,In_799);
or U452 (N_452,In_1251,In_1521);
or U453 (N_453,In_2433,In_1739);
nand U454 (N_454,In_2001,In_1864);
and U455 (N_455,In_2996,In_2385);
nor U456 (N_456,In_2937,In_1669);
nand U457 (N_457,In_1448,In_352);
nor U458 (N_458,In_2199,In_2094);
nor U459 (N_459,In_891,In_413);
or U460 (N_460,In_1408,In_2568);
and U461 (N_461,In_968,In_2152);
and U462 (N_462,In_1687,In_2770);
and U463 (N_463,In_513,In_826);
nand U464 (N_464,In_106,In_569);
or U465 (N_465,In_2166,In_637);
xor U466 (N_466,In_1962,In_1506);
nand U467 (N_467,In_262,In_1853);
or U468 (N_468,In_902,In_2406);
and U469 (N_469,In_2803,In_241);
and U470 (N_470,In_760,In_555);
nand U471 (N_471,In_962,In_119);
nand U472 (N_472,In_1266,In_1418);
and U473 (N_473,In_2046,In_1568);
or U474 (N_474,In_1287,In_2610);
and U475 (N_475,In_725,In_1341);
and U476 (N_476,In_1898,In_2260);
and U477 (N_477,In_936,In_1705);
xor U478 (N_478,In_313,In_245);
and U479 (N_479,In_2206,In_2124);
xnor U480 (N_480,In_856,In_933);
and U481 (N_481,In_2708,In_1609);
nor U482 (N_482,In_2246,In_2239);
or U483 (N_483,In_2303,In_1680);
or U484 (N_484,In_2182,In_259);
or U485 (N_485,In_2955,In_1283);
nand U486 (N_486,In_1388,In_1770);
and U487 (N_487,In_1658,In_640);
or U488 (N_488,In_919,In_2773);
xor U489 (N_489,In_149,In_1138);
and U490 (N_490,In_829,In_1672);
nand U491 (N_491,In_2903,In_142);
nand U492 (N_492,In_1279,In_1980);
xnor U493 (N_493,In_2722,In_1728);
and U494 (N_494,In_1079,In_509);
or U495 (N_495,In_2193,In_2365);
xnor U496 (N_496,In_132,In_1451);
and U497 (N_497,In_2721,In_2043);
nor U498 (N_498,In_1689,In_2621);
or U499 (N_499,In_2295,In_764);
xnor U500 (N_500,In_1998,In_1796);
xnor U501 (N_501,In_1311,In_305);
nand U502 (N_502,In_1292,In_1932);
and U503 (N_503,In_901,In_1413);
and U504 (N_504,In_1158,In_1630);
nand U505 (N_505,In_2502,In_333);
or U506 (N_506,In_2799,In_2340);
nand U507 (N_507,In_364,In_2469);
xor U508 (N_508,In_780,In_378);
nor U509 (N_509,In_1137,In_37);
nand U510 (N_510,In_1498,In_1203);
or U511 (N_511,In_1564,In_1696);
nor U512 (N_512,In_2480,In_2629);
nor U513 (N_513,In_1446,In_1025);
or U514 (N_514,In_2203,In_2539);
nor U515 (N_515,In_86,In_265);
and U516 (N_516,In_1247,In_1776);
nor U517 (N_517,In_786,In_2444);
or U518 (N_518,In_2544,In_835);
and U519 (N_519,In_1285,In_2503);
and U520 (N_520,In_1073,In_1788);
or U521 (N_521,In_1724,In_2923);
nor U522 (N_522,In_2551,In_178);
or U523 (N_523,In_2106,In_582);
and U524 (N_524,In_104,In_993);
nand U525 (N_525,In_410,In_1198);
nor U526 (N_526,In_2363,In_1046);
nand U527 (N_527,In_2083,In_2902);
nor U528 (N_528,In_2168,In_2743);
nor U529 (N_529,In_222,In_39);
xnor U530 (N_530,In_1121,In_879);
nor U531 (N_531,In_1716,In_2151);
and U532 (N_532,In_2084,In_377);
and U533 (N_533,In_866,In_2593);
nor U534 (N_534,In_114,In_2541);
nand U535 (N_535,In_2882,In_1735);
nand U536 (N_536,In_2749,In_328);
or U537 (N_537,In_1457,In_577);
nand U538 (N_538,In_862,In_1412);
nor U539 (N_539,In_868,In_1231);
nor U540 (N_540,In_1209,In_1631);
and U541 (N_541,In_1035,In_1766);
or U542 (N_542,In_2922,In_2312);
or U543 (N_543,In_1087,In_1189);
xnor U544 (N_544,In_421,In_526);
nor U545 (N_545,In_2205,In_2692);
or U546 (N_546,In_776,In_2878);
nor U547 (N_547,In_1106,In_2012);
and U548 (N_548,In_1323,In_2232);
xnor U549 (N_549,In_294,In_279);
xor U550 (N_550,In_2009,In_296);
or U551 (N_551,In_1542,In_145);
nor U552 (N_552,In_44,In_1376);
or U553 (N_553,In_953,In_187);
xor U554 (N_554,In_1210,In_1494);
nor U555 (N_555,In_1744,In_2814);
nand U556 (N_556,In_2478,In_2227);
or U557 (N_557,In_572,In_395);
xor U558 (N_558,In_2740,In_2608);
nor U559 (N_559,In_474,In_1676);
and U560 (N_560,In_1043,In_79);
nor U561 (N_561,In_1824,In_2215);
nor U562 (N_562,In_63,In_2461);
and U563 (N_563,In_1496,In_2374);
and U564 (N_564,In_1395,In_539);
or U565 (N_565,In_1881,In_2705);
nor U566 (N_566,In_2104,In_2684);
nand U567 (N_567,In_121,In_1704);
nand U568 (N_568,In_2,In_954);
nor U569 (N_569,In_740,In_1462);
nand U570 (N_570,In_2875,In_534);
or U571 (N_571,In_1513,In_1503);
nor U572 (N_572,In_991,In_664);
or U573 (N_573,In_2059,In_2999);
and U574 (N_574,In_2576,In_1195);
xor U575 (N_575,In_1667,In_399);
nor U576 (N_576,In_109,In_2578);
and U577 (N_577,In_2345,In_1988);
nor U578 (N_578,In_438,In_183);
nand U579 (N_579,In_1095,In_2731);
and U580 (N_580,In_278,In_1354);
nor U581 (N_581,In_299,In_444);
nor U582 (N_582,In_850,In_1817);
xor U583 (N_583,In_2702,In_131);
or U584 (N_584,In_155,In_1085);
nor U585 (N_585,In_362,In_2533);
xor U586 (N_586,In_2292,In_2399);
and U587 (N_587,In_1456,In_373);
nand U588 (N_588,In_518,In_942);
nand U589 (N_589,In_372,In_2828);
xnor U590 (N_590,In_1372,In_1450);
xnor U591 (N_591,In_1971,In_2946);
or U592 (N_592,In_243,In_699);
or U593 (N_593,In_2982,In_1923);
nor U594 (N_594,In_1851,In_2693);
and U595 (N_595,In_2446,In_2943);
xor U596 (N_596,In_2213,In_2904);
or U597 (N_597,In_877,In_1661);
or U598 (N_598,In_1836,In_2977);
nand U599 (N_599,In_130,In_2280);
or U600 (N_600,In_590,In_1417);
nor U601 (N_601,In_1774,In_2829);
xnor U602 (N_602,In_55,In_2324);
or U603 (N_603,In_2626,In_2985);
xnor U604 (N_604,In_2575,In_188);
and U605 (N_605,In_2360,In_622);
nor U606 (N_606,In_170,In_983);
and U607 (N_607,In_1039,In_2715);
nand U608 (N_608,In_17,In_678);
nor U609 (N_609,In_2330,In_2326);
nor U610 (N_610,In_1903,In_483);
nor U611 (N_611,In_1585,In_1265);
nor U612 (N_612,In_2805,In_1274);
and U613 (N_613,In_2762,In_1349);
or U614 (N_614,In_1232,In_1191);
or U615 (N_615,In_160,In_2990);
xnor U616 (N_616,In_2170,In_1873);
and U617 (N_617,In_2786,In_323);
nand U618 (N_618,In_1996,In_841);
nor U619 (N_619,In_2887,In_1650);
and U620 (N_620,In_926,In_2030);
nor U621 (N_621,In_2058,In_542);
nor U622 (N_622,In_794,In_1345);
xnor U623 (N_623,In_940,In_831);
nor U624 (N_624,In_383,In_536);
nand U625 (N_625,In_1644,In_2222);
nor U626 (N_626,In_58,In_180);
or U627 (N_627,In_2928,In_520);
nand U628 (N_628,In_741,In_1177);
or U629 (N_629,In_677,In_662);
xnor U630 (N_630,In_2683,In_2601);
nor U631 (N_631,In_1768,In_2764);
nand U632 (N_632,In_1690,In_1447);
and U633 (N_633,In_1814,In_557);
and U634 (N_634,In_1702,In_2646);
nor U635 (N_635,In_2265,In_320);
nor U636 (N_636,In_1583,In_1077);
nor U637 (N_637,In_1202,In_2181);
and U638 (N_638,In_2275,In_293);
nand U639 (N_639,In_2416,In_2826);
xor U640 (N_640,In_2718,In_787);
nand U641 (N_641,In_2161,In_403);
nor U642 (N_642,In_1091,In_318);
or U643 (N_643,In_2405,In_2432);
and U644 (N_644,In_254,In_1647);
and U645 (N_645,In_2663,In_1306);
or U646 (N_646,In_2868,In_1543);
xor U647 (N_647,In_1992,In_566);
nor U648 (N_648,In_1548,In_1935);
and U649 (N_649,In_2798,In_1059);
or U650 (N_650,In_2984,In_2479);
nor U651 (N_651,In_2291,In_2714);
nand U652 (N_652,In_2893,In_53);
nor U653 (N_653,In_49,In_2266);
and U654 (N_654,In_1919,In_2268);
or U655 (N_655,In_355,In_2782);
xor U656 (N_656,In_2263,In_2655);
nand U657 (N_657,In_335,In_2121);
nand U658 (N_658,In_311,In_1298);
or U659 (N_659,In_903,In_647);
nand U660 (N_660,In_2790,In_1806);
or U661 (N_661,In_1149,In_2965);
or U662 (N_662,In_724,In_1740);
nor U663 (N_663,In_543,In_353);
nor U664 (N_664,In_1178,In_1965);
nand U665 (N_665,In_769,In_1142);
nand U666 (N_666,In_300,In_471);
xnor U667 (N_667,In_1596,In_2321);
xor U668 (N_668,In_972,In_331);
nand U669 (N_669,In_946,In_409);
xor U670 (N_670,In_2427,In_2204);
nand U671 (N_671,In_1828,In_432);
or U672 (N_672,In_2002,In_958);
nor U673 (N_673,In_2082,In_939);
xnor U674 (N_674,In_627,In_1599);
and U675 (N_675,In_117,In_1920);
nand U676 (N_676,In_653,In_482);
nor U677 (N_677,In_690,In_1660);
xor U678 (N_678,In_2585,In_93);
or U679 (N_679,In_1854,In_1436);
nor U680 (N_680,In_1056,In_1725);
xor U681 (N_681,In_1362,In_2435);
xnor U682 (N_682,In_1810,In_1924);
and U683 (N_683,In_1366,In_1908);
nand U684 (N_684,In_1921,In_232);
xnor U685 (N_685,In_2443,In_2086);
nor U686 (N_686,In_276,In_1474);
nand U687 (N_687,In_414,In_2971);
nand U688 (N_688,In_1588,In_2272);
or U689 (N_689,In_628,In_2909);
and U690 (N_690,In_986,In_2802);
nor U691 (N_691,In_1424,In_2973);
xnor U692 (N_692,In_179,In_2735);
and U693 (N_693,In_1277,In_1872);
and U694 (N_694,In_874,In_1301);
or U695 (N_695,In_2658,In_959);
or U696 (N_696,In_2966,In_437);
and U697 (N_697,In_295,In_1493);
and U698 (N_698,In_2486,In_1356);
nor U699 (N_699,In_698,In_1552);
and U700 (N_700,In_2733,In_2011);
and U701 (N_701,In_2554,In_2873);
xor U702 (N_702,In_2457,In_65);
nand U703 (N_703,In_2570,In_1055);
or U704 (N_704,In_2527,In_1790);
or U705 (N_705,In_545,In_327);
xnor U706 (N_706,In_308,In_408);
xor U707 (N_707,In_137,In_967);
and U708 (N_708,In_651,In_88);
or U709 (N_709,In_2008,In_1236);
or U710 (N_710,In_1904,In_2429);
and U711 (N_711,In_1172,In_1891);
nor U712 (N_712,In_199,In_167);
xor U713 (N_713,In_2493,In_827);
and U714 (N_714,In_2022,In_1275);
xor U715 (N_715,In_1592,In_964);
nand U716 (N_716,In_2689,In_2235);
xnor U717 (N_717,In_1159,In_165);
nand U718 (N_718,In_2906,In_1478);
xnor U719 (N_719,In_1259,In_1762);
nor U720 (N_720,In_2127,In_1748);
or U721 (N_721,In_441,In_22);
or U722 (N_722,In_1787,In_2053);
xnor U723 (N_723,In_729,In_523);
xor U724 (N_724,In_151,In_1781);
nor U725 (N_725,In_2560,In_1913);
xnor U726 (N_726,In_1483,In_911);
nand U727 (N_727,In_2187,In_2017);
nand U728 (N_728,In_2386,In_1193);
nor U729 (N_729,In_2487,In_1700);
and U730 (N_730,In_974,In_2484);
nor U731 (N_731,In_707,In_1037);
and U732 (N_732,In_1633,In_2727);
and U733 (N_733,In_1949,In_2995);
nor U734 (N_734,In_2224,In_814);
or U735 (N_735,In_46,In_2085);
or U736 (N_736,In_1437,In_880);
and U737 (N_737,In_613,In_91);
nand U738 (N_738,In_1270,In_2482);
nor U739 (N_739,In_100,In_1863);
or U740 (N_740,In_1066,In_1332);
xor U741 (N_741,In_1401,In_2419);
xnor U742 (N_742,In_2783,In_1712);
nand U743 (N_743,In_112,In_1601);
nor U744 (N_744,In_1333,In_1651);
xnor U745 (N_745,In_2315,In_193);
or U746 (N_746,In_2632,In_1623);
or U747 (N_747,In_2634,In_1086);
nand U748 (N_748,In_2800,In_896);
xnor U749 (N_749,In_1519,In_1228);
nor U750 (N_750,In_469,In_1577);
nor U751 (N_751,In_1367,In_1775);
nor U752 (N_752,In_540,In_2242);
and U753 (N_753,In_2159,In_92);
and U754 (N_754,In_803,In_2262);
and U755 (N_755,In_558,In_1545);
xor U756 (N_756,In_1755,In_2674);
xor U757 (N_757,In_2314,In_537);
xor U758 (N_758,In_2962,In_1162);
or U759 (N_759,In_1308,In_2233);
xnor U760 (N_760,In_2998,In_1107);
nor U761 (N_761,In_2942,In_1316);
xnor U762 (N_762,In_689,In_620);
nor U763 (N_763,In_1600,In_426);
nand U764 (N_764,In_1108,In_2226);
nor U765 (N_765,In_2637,In_909);
nor U766 (N_766,In_1442,In_214);
nand U767 (N_767,In_2825,In_2176);
or U768 (N_768,In_2905,In_1657);
nor U769 (N_769,In_405,In_359);
or U770 (N_770,In_2696,In_2631);
and U771 (N_771,In_1737,In_738);
nand U772 (N_772,In_2013,In_2667);
nand U773 (N_773,In_2144,In_484);
nor U774 (N_774,In_172,In_4);
nor U775 (N_775,In_2501,In_2116);
or U776 (N_776,In_1168,In_2620);
xnor U777 (N_777,In_1802,In_1859);
nand U778 (N_778,In_1835,In_807);
or U779 (N_779,In_1500,In_1171);
xor U780 (N_780,In_1857,In_920);
nor U781 (N_781,In_2113,In_1931);
xor U782 (N_782,In_2856,In_2545);
nand U783 (N_783,In_2038,In_2458);
and U784 (N_784,In_2209,In_2513);
nor U785 (N_785,In_2178,In_1885);
xor U786 (N_786,In_1815,In_1169);
xor U787 (N_787,In_714,In_788);
nor U788 (N_788,In_1758,In_2234);
xor U789 (N_789,In_2673,In_498);
xnor U790 (N_790,In_252,In_344);
or U791 (N_791,In_1186,In_2488);
nand U792 (N_792,In_2748,In_1071);
nor U793 (N_793,In_573,In_716);
nand U794 (N_794,In_1892,In_1890);
or U795 (N_795,In_1005,In_1884);
xnor U796 (N_796,In_485,In_675);
nand U797 (N_797,In_1688,In_2026);
or U798 (N_798,In_743,In_2491);
or U799 (N_799,In_2960,In_1914);
xnor U800 (N_800,In_1256,In_2247);
nor U801 (N_801,In_806,In_757);
nand U802 (N_802,In_1838,In_1305);
or U803 (N_803,In_1184,In_1736);
or U804 (N_804,In_203,In_682);
and U805 (N_805,In_2862,In_1397);
xor U806 (N_806,In_1591,In_1834);
or U807 (N_807,In_819,In_1602);
nor U808 (N_808,In_2389,In_285);
and U809 (N_809,In_578,In_2076);
xnor U810 (N_810,In_2148,In_1001);
xnor U811 (N_811,In_2664,In_1125);
nor U812 (N_812,In_2078,In_517);
or U813 (N_813,In_1867,In_2958);
and U814 (N_814,In_1358,In_146);
or U815 (N_815,In_839,In_1008);
and U816 (N_816,In_2250,In_1163);
or U817 (N_817,In_70,In_1993);
nor U818 (N_818,In_672,In_284);
and U819 (N_819,In_1732,In_1398);
xor U820 (N_820,In_2089,In_78);
xor U821 (N_821,In_1355,In_157);
nand U822 (N_822,In_1756,In_2004);
nor U823 (N_823,In_1429,In_2531);
nor U824 (N_824,In_2413,In_2789);
xnor U825 (N_825,In_1656,In_701);
nor U826 (N_826,In_2404,In_2428);
nor U827 (N_827,In_1105,In_1941);
xor U828 (N_828,In_1221,In_1328);
and U829 (N_829,In_2661,In_898);
or U830 (N_830,In_2992,In_1808);
or U831 (N_831,In_507,In_168);
nand U832 (N_832,In_2528,In_1664);
nor U833 (N_833,In_922,In_859);
nand U834 (N_834,In_2061,In_2586);
xnor U835 (N_835,In_587,In_2614);
xnor U836 (N_836,In_2316,In_64);
nor U837 (N_837,In_2926,In_1565);
or U838 (N_838,In_1860,In_1423);
or U839 (N_839,In_1310,In_646);
or U840 (N_840,In_217,In_2797);
and U841 (N_841,In_1733,In_1986);
nand U842 (N_842,In_1820,In_2016);
and U843 (N_843,In_1896,In_2028);
nor U844 (N_844,In_1539,In_2779);
nor U845 (N_845,In_2309,In_1070);
xnor U846 (N_846,In_2913,In_2132);
and U847 (N_847,In_2649,In_1868);
nand U848 (N_848,In_905,In_1909);
or U849 (N_849,In_1754,In_2256);
and U850 (N_850,In_2915,In_1145);
or U851 (N_851,In_1213,In_1068);
nand U852 (N_852,In_639,In_1886);
nor U853 (N_853,In_289,In_884);
nand U854 (N_854,In_1550,In_1057);
nor U855 (N_855,In_1020,In_1480);
nand U856 (N_856,In_875,In_194);
nand U857 (N_857,In_1528,In_1734);
nand U858 (N_858,In_2092,In_2448);
nand U859 (N_859,In_2732,In_730);
nor U860 (N_860,In_2391,In_576);
and U861 (N_861,In_607,In_2706);
or U862 (N_862,In_164,In_601);
xor U863 (N_863,In_1946,In_2794);
xnor U864 (N_864,In_522,In_415);
nand U865 (N_865,In_824,In_2188);
or U866 (N_866,In_2020,In_1467);
or U867 (N_867,In_2596,In_1942);
nand U868 (N_868,In_2044,In_1386);
nor U869 (N_869,In_661,In_857);
nor U870 (N_870,In_1999,In_2024);
nand U871 (N_871,In_1800,In_1444);
or U872 (N_872,In_1486,In_871);
nand U873 (N_873,In_2839,In_2852);
or U874 (N_874,In_306,In_2463);
nor U875 (N_875,In_955,In_2616);
or U876 (N_876,In_2452,In_1533);
nand U877 (N_877,In_525,In_2930);
nand U878 (N_878,In_2141,In_2460);
and U879 (N_879,In_84,In_2529);
or U880 (N_880,In_212,In_351);
or U881 (N_881,In_1578,In_927);
xnor U882 (N_882,In_277,In_326);
and U883 (N_883,In_719,In_2297);
or U884 (N_884,In_1691,In_2396);
xnor U885 (N_885,In_2650,In_1652);
nand U886 (N_886,In_2279,In_2847);
nor U887 (N_887,In_1319,In_2603);
nor U888 (N_888,In_1174,In_50);
and U889 (N_889,In_2698,In_2060);
and U890 (N_890,In_1260,In_766);
and U891 (N_891,In_975,In_1889);
xnor U892 (N_892,In_598,In_1317);
xor U893 (N_893,In_1979,In_472);
and U894 (N_894,In_2865,In_624);
nor U895 (N_895,In_169,In_1230);
and U896 (N_896,In_33,In_2347);
xnor U897 (N_897,In_1616,In_801);
nand U898 (N_898,In_45,In_1089);
or U899 (N_899,In_2356,In_1606);
nor U900 (N_900,In_1761,In_10);
nor U901 (N_901,In_2036,In_621);
nand U902 (N_902,In_271,In_997);
xor U903 (N_903,In_2929,In_2600);
xnor U904 (N_904,In_2988,In_873);
xnor U905 (N_905,In_490,In_381);
or U906 (N_906,In_1721,In_1847);
or U907 (N_907,In_2842,In_2598);
or U908 (N_908,In_1343,In_2883);
nand U909 (N_909,In_2804,In_1375);
or U910 (N_910,In_929,In_712);
nor U911 (N_911,In_679,In_1419);
nand U912 (N_912,In_2064,In_1893);
xor U913 (N_913,In_2534,In_947);
and U914 (N_914,In_2065,In_541);
xnor U915 (N_915,In_609,In_2371);
xor U916 (N_916,In_805,In_2860);
xor U917 (N_917,In_2107,In_1054);
or U918 (N_918,In_2766,In_528);
nand U919 (N_919,In_2212,In_2579);
nor U920 (N_920,In_1245,In_944);
or U921 (N_921,In_977,In_722);
and U922 (N_922,In_924,In_1148);
and U923 (N_923,In_138,In_1746);
nand U924 (N_924,In_872,In_1197);
or U925 (N_925,In_2027,In_796);
or U926 (N_926,In_2978,In_2088);
nor U927 (N_927,In_1294,In_2393);
xor U928 (N_928,In_1910,In_389);
nor U929 (N_929,In_211,In_1945);
or U930 (N_930,In_828,In_960);
nand U931 (N_931,In_1861,In_2511);
and U932 (N_932,In_1703,In_1646);
and U933 (N_933,In_1042,In_322);
nand U934 (N_934,In_830,In_1061);
nand U935 (N_935,In_25,In_1269);
xor U936 (N_936,In_708,In_2711);
nand U937 (N_937,In_1440,In_216);
and U938 (N_938,In_1225,In_2423);
nor U939 (N_939,In_41,In_1103);
or U940 (N_940,In_2135,In_62);
and U941 (N_941,In_742,In_2690);
and U942 (N_942,In_1300,In_1331);
xor U943 (N_943,In_2376,In_2510);
or U944 (N_944,In_1078,In_125);
and U945 (N_945,In_2582,In_1334);
xor U946 (N_946,In_1212,In_680);
and U947 (N_947,In_930,In_1579);
and U948 (N_948,In_1902,In_210);
xnor U949 (N_949,In_556,In_605);
nand U950 (N_950,In_1495,In_286);
nand U951 (N_951,In_2888,In_1843);
nor U952 (N_952,In_861,In_1033);
and U953 (N_953,In_319,In_524);
xor U954 (N_954,In_2726,In_2961);
and U955 (N_955,In_358,In_2652);
xor U956 (N_956,In_2093,In_2462);
nand U957 (N_957,In_436,In_2220);
and U958 (N_958,In_1403,In_688);
nor U959 (N_959,In_1432,In_570);
nor U960 (N_960,In_2831,In_2490);
nor U961 (N_961,In_2870,In_762);
or U962 (N_962,In_676,In_393);
or U963 (N_963,In_585,In_234);
nand U964 (N_964,In_0,In_1870);
and U965 (N_965,In_2000,In_1080);
nor U966 (N_966,In_2409,In_1026);
nor U967 (N_967,In_251,In_1387);
or U968 (N_968,In_1845,In_52);
and U969 (N_969,In_345,In_126);
nor U970 (N_970,In_90,In_2071);
and U971 (N_971,In_246,In_153);
nand U972 (N_972,In_2936,In_1389);
and U973 (N_973,In_649,In_914);
and U974 (N_974,In_1722,In_1574);
xor U975 (N_975,In_2387,In_1434);
nand U976 (N_976,In_2587,In_1384);
nand U977 (N_977,In_2745,In_1340);
nor U978 (N_978,In_567,In_1640);
and U979 (N_979,In_2871,In_48);
nand U980 (N_980,In_2207,In_1484);
nand U981 (N_981,In_2728,In_337);
xor U982 (N_982,In_1525,In_1041);
and U983 (N_983,In_1352,In_374);
and U984 (N_984,In_2109,In_2070);
or U985 (N_985,In_2676,In_1575);
nand U986 (N_986,In_275,In_2362);
or U987 (N_987,In_26,In_1821);
nor U988 (N_988,In_1951,In_2817);
nor U989 (N_989,In_1278,In_1206);
nand U990 (N_990,In_2208,In_1028);
xor U991 (N_991,In_865,In_883);
and U992 (N_992,In_822,In_1280);
nor U993 (N_993,In_1153,In_83);
or U994 (N_994,In_516,In_848);
and U995 (N_995,In_1146,In_213);
nand U996 (N_996,In_844,In_823);
or U997 (N_997,In_1795,In_881);
or U998 (N_998,In_1632,In_1597);
or U999 (N_999,In_368,In_746);
nor U1000 (N_1000,In_1218,In_1263);
xnor U1001 (N_1001,In_673,In_2838);
nand U1002 (N_1002,In_2846,In_122);
xnor U1003 (N_1003,In_789,In_548);
and U1004 (N_1004,In_1475,In_1869);
nor U1005 (N_1005,In_1023,In_2801);
nand U1006 (N_1006,In_1901,In_2379);
or U1007 (N_1007,In_1003,In_1849);
nor U1008 (N_1008,In_1404,In_1223);
nor U1009 (N_1009,In_1692,In_660);
or U1010 (N_1010,In_171,In_581);
xnor U1011 (N_1011,In_2394,In_2682);
and U1012 (N_1012,In_2589,In_2874);
xor U1013 (N_1013,In_1233,In_32);
nand U1014 (N_1014,In_965,In_2056);
nand U1015 (N_1015,In_2049,In_2716);
and U1016 (N_1016,In_1499,In_1662);
xor U1017 (N_1017,In_1219,In_2498);
nor U1018 (N_1018,In_363,In_2522);
nor U1019 (N_1019,In_1907,In_995);
nand U1020 (N_1020,In_1706,In_2177);
and U1021 (N_1021,In_494,In_1339);
or U1022 (N_1022,In_1649,In_312);
or U1023 (N_1023,In_181,In_2296);
and U1024 (N_1024,In_1751,In_1711);
nor U1025 (N_1025,In_1673,In_1809);
and U1026 (N_1026,In_496,In_1803);
and U1027 (N_1027,In_488,In_982);
and U1028 (N_1028,In_2917,In_2499);
and U1029 (N_1029,In_1855,In_837);
and U1030 (N_1030,In_1161,In_2067);
nor U1031 (N_1031,In_2638,In_1017);
xnor U1032 (N_1032,In_767,In_2099);
nor U1033 (N_1033,In_1391,In_1313);
xnor U1034 (N_1034,In_1581,In_1326);
nand U1035 (N_1035,In_1439,In_154);
and U1036 (N_1036,In_1842,In_1034);
or U1037 (N_1037,In_1012,In_1940);
xor U1038 (N_1038,In_1185,In_2876);
and U1039 (N_1039,In_2927,In_854);
nor U1040 (N_1040,In_2248,In_2243);
and U1041 (N_1041,In_2424,In_2039);
or U1042 (N_1042,In_2160,In_795);
nand U1043 (N_1043,In_825,In_1452);
nor U1044 (N_1044,In_1593,In_553);
or U1045 (N_1045,In_1431,In_1196);
nand U1046 (N_1046,In_2688,In_2662);
xor U1047 (N_1047,In_2581,In_1346);
xor U1048 (N_1048,In_1183,In_2476);
and U1049 (N_1049,In_1572,In_1937);
or U1050 (N_1050,In_2408,In_1636);
or U1051 (N_1051,In_2771,In_1947);
and U1052 (N_1052,In_2305,In_1508);
nand U1053 (N_1053,In_887,In_1698);
nand U1054 (N_1054,In_1379,In_923);
and U1055 (N_1055,In_2006,In_1252);
nand U1056 (N_1056,In_2925,In_1537);
nor U1057 (N_1057,In_2951,In_1523);
or U1058 (N_1058,In_2806,In_551);
and U1059 (N_1059,In_1006,In_1522);
nor U1060 (N_1060,In_2054,In_2611);
nand U1061 (N_1061,In_2761,In_1410);
or U1062 (N_1062,In_783,In_1207);
or U1063 (N_1063,In_2175,In_510);
nand U1064 (N_1064,In_487,In_3);
nand U1065 (N_1065,In_547,In_1040);
or U1066 (N_1066,In_1641,In_1253);
nand U1067 (N_1067,In_57,In_1731);
xnor U1068 (N_1068,In_761,In_2431);
and U1069 (N_1069,In_1926,In_792);
nand U1070 (N_1070,In_477,In_1621);
xor U1071 (N_1071,In_893,In_951);
nor U1072 (N_1072,In_1074,In_782);
nor U1073 (N_1073,In_407,In_2707);
nor U1074 (N_1074,In_354,In_2963);
nor U1075 (N_1075,In_195,In_1954);
xor U1076 (N_1076,In_2489,In_2382);
nand U1077 (N_1077,In_2194,In_2859);
xnor U1078 (N_1078,In_2281,In_2737);
or U1079 (N_1079,In_2401,In_1694);
nand U1080 (N_1080,In_2311,In_2240);
xnor U1081 (N_1081,In_1383,In_921);
nand U1082 (N_1082,In_244,In_564);
nand U1083 (N_1083,In_380,In_910);
and U1084 (N_1084,In_1082,In_2216);
nor U1085 (N_1085,In_1862,In_2843);
xor U1086 (N_1086,In_248,In_184);
nand U1087 (N_1087,In_2547,In_2980);
nor U1088 (N_1088,In_1141,In_396);
xor U1089 (N_1089,In_461,In_1281);
nand U1090 (N_1090,In_491,In_1481);
nor U1091 (N_1091,In_129,In_2505);
and U1092 (N_1092,In_2864,In_815);
and U1093 (N_1093,In_1977,In_1120);
xnor U1094 (N_1094,In_1027,In_107);
nor U1095 (N_1095,In_1876,In_1032);
and U1096 (N_1096,In_2521,In_845);
nor U1097 (N_1097,In_2025,In_704);
or U1098 (N_1098,In_2671,In_847);
or U1099 (N_1099,In_228,In_340);
nor U1100 (N_1100,In_303,In_918);
and U1101 (N_1101,In_670,In_1258);
xor U1102 (N_1102,In_2472,In_917);
nand U1103 (N_1103,In_2604,In_1407);
nor U1104 (N_1104,In_950,In_1990);
xnor U1105 (N_1105,In_2271,In_641);
and U1106 (N_1106,In_2869,In_1021);
nor U1107 (N_1107,In_990,In_1390);
xor U1108 (N_1108,In_667,In_2338);
nor U1109 (N_1109,In_2080,In_467);
xnor U1110 (N_1110,In_1152,In_2897);
nand U1111 (N_1111,In_2010,In_11);
xor U1112 (N_1112,In_1584,In_8);
nand U1113 (N_1113,In_1826,In_978);
xor U1114 (N_1114,In_2299,In_2223);
nor U1115 (N_1115,In_1368,In_2436);
or U1116 (N_1116,In_1072,In_644);
and U1117 (N_1117,In_1359,In_2289);
and U1118 (N_1118,In_1570,In_836);
and U1119 (N_1119,In_1959,In_1943);
or U1120 (N_1120,In_449,In_2018);
or U1121 (N_1121,In_781,In_1271);
xor U1122 (N_1122,In_2318,In_1558);
xor U1123 (N_1123,In_1385,In_14);
nor U1124 (N_1124,In_2122,In_1974);
nor U1125 (N_1125,In_1060,In_1922);
nor U1126 (N_1126,In_1123,In_82);
xor U1127 (N_1127,In_2050,In_1981);
xnor U1128 (N_1128,In_511,In_220);
and U1129 (N_1129,In_894,In_463);
nor U1130 (N_1130,In_984,In_702);
and U1131 (N_1131,In_2300,In_56);
or U1132 (N_1132,In_2133,In_1638);
xor U1133 (N_1133,In_2895,In_1617);
nand U1134 (N_1134,In_2599,In_808);
xor U1135 (N_1135,In_584,In_1987);
nand U1136 (N_1136,In_888,In_987);
or U1137 (N_1137,In_2781,In_999);
nand U1138 (N_1138,In_69,In_27);
and U1139 (N_1139,In_1970,In_2465);
nand U1140 (N_1140,In_266,In_2517);
xnor U1141 (N_1141,In_2383,In_957);
nand U1142 (N_1142,In_2584,In_1655);
and U1143 (N_1143,In_650,In_2264);
and U1144 (N_1144,In_502,In_156);
nor U1145 (N_1145,In_2023,In_696);
nand U1146 (N_1146,In_2153,In_633);
and U1147 (N_1147,In_711,In_1135);
or U1148 (N_1148,In_1261,In_51);
or U1149 (N_1149,In_1665,In_2615);
xnor U1150 (N_1150,In_1856,In_2090);
nor U1151 (N_1151,In_255,In_1192);
nand U1152 (N_1152,In_2218,In_745);
nor U1153 (N_1153,In_321,In_1823);
nand U1154 (N_1154,In_2795,In_544);
nor U1155 (N_1155,In_809,In_1416);
or U1156 (N_1156,In_15,In_1865);
nand U1157 (N_1157,In_2125,In_674);
or U1158 (N_1158,In_508,In_1058);
and U1159 (N_1159,In_1443,In_1473);
nor U1160 (N_1160,In_1002,In_842);
xor U1161 (N_1161,In_591,In_186);
and U1162 (N_1162,In_190,In_456);
nand U1163 (N_1163,In_1297,In_1409);
xnor U1164 (N_1164,In_900,In_2145);
and U1165 (N_1165,In_2788,In_2968);
and U1166 (N_1166,In_732,In_519);
nand U1167 (N_1167,In_249,In_1414);
nor U1168 (N_1168,In_2112,In_1463);
and U1169 (N_1169,In_281,In_834);
and U1170 (N_1170,In_2454,In_2077);
or U1171 (N_1171,In_1010,In_2827);
nor U1172 (N_1172,In_1445,In_1370);
nand U1173 (N_1173,In_2588,In_229);
nand U1174 (N_1174,In_2474,In_2483);
nor U1175 (N_1175,In_442,In_2680);
xor U1176 (N_1176,In_2949,In_2421);
nor U1177 (N_1177,In_29,In_652);
and U1178 (N_1178,In_596,In_391);
nand U1179 (N_1179,In_67,In_141);
and U1180 (N_1180,In_253,In_36);
xor U1181 (N_1181,In_1666,In_21);
nand U1182 (N_1182,In_1139,In_812);
nand U1183 (N_1183,In_1015,In_1779);
nor U1184 (N_1184,In_2425,In_778);
nand U1185 (N_1185,In_2378,In_2190);
xor U1186 (N_1186,In_1239,In_1563);
nand U1187 (N_1187,In_2191,In_2654);
or U1188 (N_1188,In_1458,In_390);
nor U1189 (N_1189,In_492,In_2710);
nand U1190 (N_1190,In_163,In_2329);
and U1191 (N_1191,In_334,In_1819);
nor U1192 (N_1192,In_1709,In_615);
xor U1193 (N_1193,In_2524,In_763);
and U1194 (N_1194,In_1717,In_386);
or U1195 (N_1195,In_1382,In_2500);
nand U1196 (N_1196,In_2941,In_189);
or U1197 (N_1197,In_2066,In_497);
nand U1198 (N_1198,In_2390,In_779);
and U1199 (N_1199,In_1743,In_937);
xnor U1200 (N_1200,In_2957,In_1759);
and U1201 (N_1201,In_206,In_2891);
nand U1202 (N_1202,In_2381,In_2138);
xnor U1203 (N_1203,In_2334,In_2730);
xnor U1204 (N_1204,In_592,In_1464);
and U1205 (N_1205,In_925,In_1302);
nand U1206 (N_1206,In_1561,In_2635);
nand U1207 (N_1207,In_1544,In_1428);
or U1208 (N_1208,In_77,In_302);
nand U1209 (N_1209,In_749,In_304);
xor U1210 (N_1210,In_2641,In_2497);
nand U1211 (N_1211,In_2146,In_692);
and U1212 (N_1212,In_2687,In_1018);
and U1213 (N_1213,In_514,In_1546);
or U1214 (N_1214,In_2738,In_979);
nor U1215 (N_1215,In_1433,In_597);
nand U1216 (N_1216,In_1110,In_668);
nand U1217 (N_1217,In_1605,In_2259);
nand U1218 (N_1218,In_1084,In_1686);
xor U1219 (N_1219,In_1426,In_445);
or U1220 (N_1220,In_2286,In_2158);
and U1221 (N_1221,In_1507,In_2139);
and U1222 (N_1222,In_709,In_1957);
nor U1223 (N_1223,In_1240,In_785);
xnor U1224 (N_1224,In_98,In_1360);
and U1225 (N_1225,In_2422,In_2780);
and U1226 (N_1226,In_1336,In_1155);
xor U1227 (N_1227,In_1812,In_162);
nand U1228 (N_1228,In_315,In_2627);
or U1229 (N_1229,In_703,In_2519);
and U1230 (N_1230,In_470,In_727);
nand U1231 (N_1231,In_2916,In_2657);
and U1232 (N_1232,In_2746,In_99);
nand U1233 (N_1233,In_1784,In_1399);
nand U1234 (N_1234,In_2755,In_338);
and U1235 (N_1235,In_2287,In_236);
or U1236 (N_1236,In_1582,In_623);
or U1237 (N_1237,In_595,In_1956);
nand U1238 (N_1238,In_2834,In_1801);
nand U1239 (N_1239,In_1267,In_1677);
and U1240 (N_1240,In_2449,In_1929);
or U1241 (N_1241,In_721,In_1208);
and U1242 (N_1242,In_1831,In_2595);
nor U1243 (N_1243,In_2940,In_1181);
or U1244 (N_1244,In_1400,In_2350);
nand U1245 (N_1245,In_1194,In_489);
xor U1246 (N_1246,In_1953,In_2934);
or U1247 (N_1247,In_2320,In_1952);
and U1248 (N_1248,In_1477,In_1117);
and U1249 (N_1249,In_124,In_1883);
and U1250 (N_1250,In_2833,In_1792);
nor U1251 (N_1251,In_1244,In_435);
nand U1252 (N_1252,In_833,In_2907);
and U1253 (N_1253,In_158,In_693);
xnor U1254 (N_1254,In_2052,In_1357);
and U1255 (N_1255,In_2410,In_1773);
and U1256 (N_1256,In_204,In_1047);
and U1257 (N_1257,In_1540,In_1645);
nor U1258 (N_1258,In_563,In_1948);
nand U1259 (N_1259,In_1471,In_811);
nor U1260 (N_1260,In_1804,In_2464);
or U1261 (N_1261,In_174,In_1771);
or U1262 (N_1262,In_2095,In_2274);
xnor U1263 (N_1263,In_2848,In_423);
xnor U1264 (N_1264,In_367,In_230);
nor U1265 (N_1265,In_2747,In_2201);
nor U1266 (N_1266,In_2920,In_817);
and U1267 (N_1267,In_1678,In_1200);
xor U1268 (N_1268,In_855,In_2231);
nand U1269 (N_1269,In_215,In_448);
nor U1270 (N_1270,In_686,In_756);
or U1271 (N_1271,In_1562,In_2339);
nor U1272 (N_1272,In_439,In_2639);
or U1273 (N_1273,In_1833,In_503);
or U1274 (N_1274,In_1559,In_687);
nor U1275 (N_1275,In_1611,In_935);
nand U1276 (N_1276,In_457,In_2244);
xnor U1277 (N_1277,In_932,In_2558);
or U1278 (N_1278,In_1415,In_2267);
nor U1279 (N_1279,In_460,In_2117);
nor U1280 (N_1280,In_2653,In_2656);
nor U1281 (N_1281,In_1619,In_297);
xnor U1282 (N_1282,In_2367,In_1282);
and U1283 (N_1283,In_2950,In_1126);
xnor U1284 (N_1284,In_1530,In_2466);
and U1285 (N_1285,In_2889,In_40);
nor U1286 (N_1286,In_2123,In_2703);
xor U1287 (N_1287,In_1906,In_2697);
nand U1288 (N_1288,In_1170,In_1118);
xnor U1289 (N_1289,In_1786,In_2857);
nand U1290 (N_1290,In_267,In_904);
nor U1291 (N_1291,In_1674,In_2284);
or U1292 (N_1292,In_669,In_2532);
and U1293 (N_1293,In_2525,In_754);
and U1294 (N_1294,In_1624,In_2670);
and U1295 (N_1295,In_2577,In_2359);
nor U1296 (N_1296,In_718,In_6);
nor U1297 (N_1297,In_2709,In_1421);
xor U1298 (N_1298,In_723,In_1960);
nand U1299 (N_1299,In_728,In_1797);
and U1300 (N_1300,In_864,In_2172);
or U1301 (N_1301,In_1822,In_2774);
nand U1302 (N_1302,In_804,In_1505);
xnor U1303 (N_1303,In_1226,In_2537);
or U1304 (N_1304,In_2701,In_2948);
nor U1305 (N_1305,In_2283,In_1405);
nand U1306 (N_1306,In_784,In_821);
or U1307 (N_1307,In_499,In_945);
or U1308 (N_1308,In_1830,In_908);
or U1309 (N_1309,In_2793,In_2516);
or U1310 (N_1310,In_1380,In_1052);
and U1311 (N_1311,In_505,In_1489);
or U1312 (N_1312,In_72,In_2029);
xnor U1313 (N_1313,In_2358,In_1272);
nand U1314 (N_1314,In_103,In_747);
nand U1315 (N_1315,In_2081,In_851);
or U1316 (N_1316,In_952,In_2219);
nand U1317 (N_1317,In_1165,In_2192);
nand U1318 (N_1318,In_1944,In_1214);
xnor U1319 (N_1319,In_706,In_111);
and U1320 (N_1320,In_2355,In_1320);
or U1321 (N_1321,In_371,In_941);
and U1322 (N_1322,In_2041,In_1164);
nand U1323 (N_1323,In_2760,In_1242);
or U1324 (N_1324,In_1022,In_1590);
and U1325 (N_1325,In_2853,In_2536);
or U1326 (N_1326,In_2514,In_61);
and U1327 (N_1327,In_1257,In_486);
nand U1328 (N_1328,In_2063,In_2812);
and U1329 (N_1329,In_773,In_2677);
nor U1330 (N_1330,In_554,In_1598);
or U1331 (N_1331,In_2659,In_2470);
and U1332 (N_1332,In_956,In_915);
and U1333 (N_1333,In_1016,In_2445);
nand U1334 (N_1334,In_1713,In_2567);
nor U1335 (N_1335,In_1763,In_574);
nand U1336 (N_1336,In_2678,In_2618);
nand U1337 (N_1337,In_750,In_1818);
xnor U1338 (N_1338,In_2752,In_416);
and U1339 (N_1339,In_1741,In_1465);
or U1340 (N_1340,In_2777,In_224);
or U1341 (N_1341,In_1112,In_1895);
xnor U1342 (N_1342,In_1083,In_2736);
and U1343 (N_1343,In_2019,In_899);
nand U1344 (N_1344,In_2850,In_2414);
nand U1345 (N_1345,In_2238,In_2034);
nor U1346 (N_1346,In_2200,In_568);
or U1347 (N_1347,In_38,In_2507);
or U1348 (N_1348,In_697,In_735);
and U1349 (N_1349,In_116,In_2564);
xor U1350 (N_1350,In_1205,In_1969);
or U1351 (N_1351,In_1811,In_671);
and U1352 (N_1352,In_2734,In_1626);
nor U1353 (N_1353,In_2617,In_630);
and U1354 (N_1354,In_1199,In_1238);
and U1355 (N_1355,In_2440,In_196);
nand U1356 (N_1356,In_2217,In_13);
nor U1357 (N_1357,In_428,In_136);
nor U1358 (N_1358,In_19,In_2609);
xnor U1359 (N_1359,In_1180,In_1780);
nand U1360 (N_1360,In_2111,In_1098);
nor U1361 (N_1361,In_772,In_2398);
xor U1362 (N_1362,In_2912,In_166);
xor U1363 (N_1363,In_2686,In_1524);
or U1364 (N_1364,In_269,In_1124);
nand U1365 (N_1365,In_1295,In_1364);
and U1366 (N_1366,In_1580,In_992);
and U1367 (N_1367,In_339,In_530);
and U1368 (N_1368,In_2633,In_1553);
nand U1369 (N_1369,In_425,In_768);
or U1370 (N_1370,In_1029,In_2370);
and U1371 (N_1371,In_1675,In_43);
nand U1372 (N_1372,In_1852,In_1286);
nand U1373 (N_1373,In_2344,In_1573);
nand U1374 (N_1374,In_1011,In_1840);
nand U1375 (N_1375,In_2438,In_656);
and U1376 (N_1376,In_2253,In_1088);
and U1377 (N_1377,In_418,In_1327);
xnor U1378 (N_1378,In_47,In_87);
and U1379 (N_1379,In_586,In_853);
and U1380 (N_1380,In_907,In_424);
xnor U1381 (N_1381,In_2197,In_273);
nor U1382 (N_1382,In_2555,In_2306);
nor U1383 (N_1383,In_2352,In_2114);
nand U1384 (N_1384,In_1966,In_147);
nor U1385 (N_1385,In_2258,In_2456);
xnor U1386 (N_1386,In_2763,In_18);
and U1387 (N_1387,In_1435,In_527);
xor U1388 (N_1388,In_2557,In_1627);
and U1389 (N_1389,In_765,In_634);
or U1390 (N_1390,In_2357,In_1014);
nand U1391 (N_1391,In_1963,In_2765);
xnor U1392 (N_1392,In_2411,In_2293);
xnor U1393 (N_1393,In_2229,In_654);
nor U1394 (N_1394,In_1531,In_2317);
nor U1395 (N_1395,In_1309,In_2384);
nand U1396 (N_1396,In_201,In_1846);
xor U1397 (N_1397,In_840,In_96);
and U1398 (N_1398,In_2723,In_512);
nand U1399 (N_1399,In_994,In_759);
or U1400 (N_1400,In_2720,In_1750);
nor U1401 (N_1401,In_2559,In_2174);
or U1402 (N_1402,In_1527,In_1747);
nand U1403 (N_1403,In_465,In_2538);
nor U1404 (N_1404,In_258,In_1151);
and U1405 (N_1405,In_1866,In_1504);
nor U1406 (N_1406,In_152,In_1682);
and U1407 (N_1407,In_2991,In_2776);
and U1408 (N_1408,In_838,In_2819);
or U1409 (N_1409,In_133,In_1491);
and U1410 (N_1410,In_2269,In_2126);
or U1411 (N_1411,In_1128,In_1634);
and U1412 (N_1412,In_1778,In_2037);
and U1413 (N_1413,In_2225,In_176);
and U1414 (N_1414,In_2810,In_81);
xnor U1415 (N_1415,In_691,In_2455);
nand U1416 (N_1416,In_588,In_2441);
or U1417 (N_1417,In_202,In_1150);
nor U1418 (N_1418,In_1917,In_2712);
and U1419 (N_1419,In_1497,In_616);
and U1420 (N_1420,In_501,In_2475);
nand U1421 (N_1421,In_453,In_387);
or U1422 (N_1422,In_2442,In_550);
nand U1423 (N_1423,In_341,In_2252);
nor U1424 (N_1424,In_1569,In_398);
xnor U1425 (N_1425,In_2753,In_446);
nand U1426 (N_1426,In_2938,In_1989);
or U1427 (N_1427,In_2323,In_2815);
nand U1428 (N_1428,In_1143,In_2892);
and U1429 (N_1429,In_1000,In_2400);
nor U1430 (N_1430,In_1330,In_2944);
nand U1431 (N_1431,In_2636,In_283);
and U1432 (N_1432,In_2832,In_1129);
or U1433 (N_1433,In_2228,In_2885);
or U1434 (N_1434,In_2290,In_1147);
nand U1435 (N_1435,In_2328,In_2785);
nand U1436 (N_1436,In_1175,In_2679);
and U1437 (N_1437,In_2341,In_1187);
or U1438 (N_1438,In_2069,In_2884);
or U1439 (N_1439,In_1612,In_1160);
or U1440 (N_1440,In_75,In_614);
nand U1441 (N_1441,In_931,In_710);
and U1442 (N_1442,In_1603,In_2757);
nor U1443 (N_1443,In_1791,In_2772);
nor U1444 (N_1444,In_495,In_239);
xor U1445 (N_1445,In_1102,In_1534);
xnor U1446 (N_1446,In_1099,In_342);
nor U1447 (N_1447,In_1753,In_1338);
xor U1448 (N_1448,In_1816,In_1133);
nand U1449 (N_1449,In_2700,In_2914);
nor U1450 (N_1450,In_2894,In_420);
nor U1451 (N_1451,In_870,In_2989);
or U1452 (N_1452,In_1479,In_2364);
or U1453 (N_1453,In_2672,In_655);
nand U1454 (N_1454,In_2836,In_1144);
nand U1455 (N_1455,In_2031,In_2249);
and U1456 (N_1456,In_1004,In_2388);
nor U1457 (N_1457,In_2091,In_2881);
nor U1458 (N_1458,In_2562,In_1335);
and U1459 (N_1459,In_1927,In_2447);
nor U1460 (N_1460,In_2477,In_1888);
and U1461 (N_1461,In_272,In_2372);
nor U1462 (N_1462,In_2319,In_2221);
and U1463 (N_1463,In_521,In_1586);
and U1464 (N_1464,In_2420,In_23);
and U1465 (N_1465,In_1325,In_2619);
xnor U1466 (N_1466,In_2808,In_1234);
xor U1467 (N_1467,In_736,In_1871);
and U1468 (N_1468,In_1912,In_1276);
xnor U1469 (N_1469,In_2691,In_2171);
nor U1470 (N_1470,In_2699,In_2057);
nor U1471 (N_1471,In_2134,In_2417);
nor U1472 (N_1472,In_989,In_2964);
nor U1473 (N_1473,In_2592,In_412);
xor U1474 (N_1474,In_2164,In_2523);
xor U1475 (N_1475,In_191,In_882);
nor U1476 (N_1476,In_208,In_1293);
xnor U1477 (N_1477,In_218,In_247);
or U1478 (N_1478,In_2756,In_2791);
nand U1479 (N_1479,In_1637,In_2230);
xnor U1480 (N_1480,In_357,In_431);
nand U1481 (N_1481,In_1567,In_1);
and U1482 (N_1482,In_325,In_361);
and U1483 (N_1483,In_2098,In_2156);
xnor U1484 (N_1484,In_1911,In_2630);
nor U1485 (N_1485,In_1668,In_1188);
or U1486 (N_1486,In_1693,In_464);
or U1487 (N_1487,In_2015,In_775);
nor U1488 (N_1488,In_2202,In_2147);
xnor U1489 (N_1489,In_2956,In_205);
nand U1490 (N_1490,In_1425,In_603);
or U1491 (N_1491,In_2418,In_2110);
and U1492 (N_1492,In_2157,In_818);
nand U1493 (N_1493,In_268,In_1365);
xnor U1494 (N_1494,In_1007,In_1526);
nor U1495 (N_1495,In_1290,In_867);
nand U1496 (N_1496,In_685,In_2830);
nand U1497 (N_1497,In_1551,In_2994);
xor U1498 (N_1498,In_1683,In_2717);
and U1499 (N_1499,In_1659,In_970);
nand U1500 (N_1500,In_1241,In_2701);
or U1501 (N_1501,In_795,In_2927);
and U1502 (N_1502,In_2030,In_2195);
xor U1503 (N_1503,In_1718,In_2482);
nor U1504 (N_1504,In_2674,In_1004);
xnor U1505 (N_1505,In_2877,In_1653);
xor U1506 (N_1506,In_1656,In_604);
nor U1507 (N_1507,In_837,In_2938);
nand U1508 (N_1508,In_625,In_125);
or U1509 (N_1509,In_2910,In_1475);
xor U1510 (N_1510,In_661,In_2732);
and U1511 (N_1511,In_1043,In_2663);
and U1512 (N_1512,In_1823,In_1588);
and U1513 (N_1513,In_2981,In_1576);
nor U1514 (N_1514,In_2566,In_1670);
nor U1515 (N_1515,In_205,In_2418);
xor U1516 (N_1516,In_2415,In_2381);
nor U1517 (N_1517,In_1338,In_2783);
nor U1518 (N_1518,In_1323,In_285);
xnor U1519 (N_1519,In_1532,In_2004);
and U1520 (N_1520,In_805,In_1728);
nor U1521 (N_1521,In_938,In_939);
nand U1522 (N_1522,In_1960,In_2332);
or U1523 (N_1523,In_870,In_1666);
and U1524 (N_1524,In_1120,In_2459);
nand U1525 (N_1525,In_601,In_2033);
nor U1526 (N_1526,In_937,In_2858);
and U1527 (N_1527,In_1222,In_2251);
and U1528 (N_1528,In_2513,In_2859);
and U1529 (N_1529,In_2783,In_1992);
and U1530 (N_1530,In_1871,In_1488);
nand U1531 (N_1531,In_2691,In_1980);
or U1532 (N_1532,In_388,In_230);
nor U1533 (N_1533,In_428,In_303);
xor U1534 (N_1534,In_563,In_2855);
nor U1535 (N_1535,In_1366,In_562);
nor U1536 (N_1536,In_1034,In_2714);
nand U1537 (N_1537,In_744,In_2280);
nand U1538 (N_1538,In_956,In_847);
nand U1539 (N_1539,In_1125,In_183);
and U1540 (N_1540,In_1704,In_2225);
nand U1541 (N_1541,In_745,In_654);
nand U1542 (N_1542,In_1088,In_114);
or U1543 (N_1543,In_1756,In_624);
nor U1544 (N_1544,In_1268,In_384);
nor U1545 (N_1545,In_2478,In_143);
or U1546 (N_1546,In_2803,In_891);
and U1547 (N_1547,In_2548,In_1981);
or U1548 (N_1548,In_2327,In_2009);
and U1549 (N_1549,In_1092,In_1387);
and U1550 (N_1550,In_1956,In_1518);
nor U1551 (N_1551,In_165,In_790);
nor U1552 (N_1552,In_1344,In_2065);
and U1553 (N_1553,In_2984,In_1050);
nor U1554 (N_1554,In_490,In_2514);
xnor U1555 (N_1555,In_1710,In_422);
and U1556 (N_1556,In_2088,In_1430);
and U1557 (N_1557,In_123,In_1198);
or U1558 (N_1558,In_2542,In_2692);
nor U1559 (N_1559,In_1690,In_2554);
nor U1560 (N_1560,In_2217,In_1478);
xor U1561 (N_1561,In_446,In_1742);
nand U1562 (N_1562,In_2967,In_1520);
and U1563 (N_1563,In_1652,In_1676);
and U1564 (N_1564,In_2430,In_1833);
or U1565 (N_1565,In_84,In_1911);
nand U1566 (N_1566,In_913,In_2877);
xor U1567 (N_1567,In_1239,In_2760);
nand U1568 (N_1568,In_2496,In_1126);
xor U1569 (N_1569,In_766,In_2168);
xnor U1570 (N_1570,In_1408,In_1285);
or U1571 (N_1571,In_2741,In_2986);
and U1572 (N_1572,In_1802,In_2246);
and U1573 (N_1573,In_2090,In_935);
or U1574 (N_1574,In_1423,In_924);
nor U1575 (N_1575,In_803,In_2287);
nand U1576 (N_1576,In_1030,In_2111);
nand U1577 (N_1577,In_2175,In_2605);
nor U1578 (N_1578,In_2664,In_1163);
nand U1579 (N_1579,In_778,In_1090);
nand U1580 (N_1580,In_2662,In_972);
and U1581 (N_1581,In_2518,In_205);
nand U1582 (N_1582,In_43,In_2465);
or U1583 (N_1583,In_1535,In_1514);
nor U1584 (N_1584,In_105,In_2498);
nor U1585 (N_1585,In_1915,In_498);
nand U1586 (N_1586,In_2132,In_232);
nand U1587 (N_1587,In_1436,In_1602);
and U1588 (N_1588,In_800,In_779);
and U1589 (N_1589,In_2230,In_592);
or U1590 (N_1590,In_734,In_75);
or U1591 (N_1591,In_217,In_2340);
and U1592 (N_1592,In_2697,In_2277);
nand U1593 (N_1593,In_2452,In_1311);
nand U1594 (N_1594,In_2938,In_1339);
or U1595 (N_1595,In_1183,In_2416);
nor U1596 (N_1596,In_1013,In_2873);
or U1597 (N_1597,In_2512,In_2338);
nand U1598 (N_1598,In_1386,In_1247);
and U1599 (N_1599,In_1626,In_2522);
nand U1600 (N_1600,In_2238,In_890);
nor U1601 (N_1601,In_9,In_251);
or U1602 (N_1602,In_1622,In_662);
xor U1603 (N_1603,In_2603,In_1627);
and U1604 (N_1604,In_2322,In_1881);
nand U1605 (N_1605,In_1766,In_2650);
nand U1606 (N_1606,In_629,In_268);
nand U1607 (N_1607,In_1669,In_1717);
and U1608 (N_1608,In_684,In_2304);
or U1609 (N_1609,In_1684,In_2120);
nor U1610 (N_1610,In_2743,In_1588);
or U1611 (N_1611,In_609,In_2081);
nand U1612 (N_1612,In_282,In_1500);
or U1613 (N_1613,In_1270,In_2283);
nor U1614 (N_1614,In_2019,In_1048);
or U1615 (N_1615,In_1380,In_2725);
and U1616 (N_1616,In_1,In_2204);
or U1617 (N_1617,In_2664,In_1230);
nand U1618 (N_1618,In_167,In_800);
nand U1619 (N_1619,In_1527,In_2532);
nor U1620 (N_1620,In_1549,In_1480);
nand U1621 (N_1621,In_1618,In_1805);
nor U1622 (N_1622,In_1951,In_87);
nand U1623 (N_1623,In_1229,In_2565);
or U1624 (N_1624,In_162,In_828);
xor U1625 (N_1625,In_2239,In_1341);
and U1626 (N_1626,In_2605,In_305);
and U1627 (N_1627,In_2967,In_2351);
xor U1628 (N_1628,In_2628,In_1120);
and U1629 (N_1629,In_1036,In_2396);
and U1630 (N_1630,In_1180,In_1596);
nand U1631 (N_1631,In_2078,In_2224);
xnor U1632 (N_1632,In_1860,In_716);
nor U1633 (N_1633,In_510,In_2734);
nor U1634 (N_1634,In_1293,In_32);
nand U1635 (N_1635,In_1458,In_316);
or U1636 (N_1636,In_573,In_754);
xor U1637 (N_1637,In_2008,In_1525);
xnor U1638 (N_1638,In_861,In_2000);
xnor U1639 (N_1639,In_1382,In_183);
and U1640 (N_1640,In_2164,In_383);
and U1641 (N_1641,In_365,In_2529);
or U1642 (N_1642,In_340,In_2059);
nand U1643 (N_1643,In_1578,In_2483);
or U1644 (N_1644,In_581,In_1797);
nor U1645 (N_1645,In_1086,In_1655);
nand U1646 (N_1646,In_430,In_1903);
or U1647 (N_1647,In_582,In_1316);
nand U1648 (N_1648,In_2273,In_794);
and U1649 (N_1649,In_814,In_1496);
xor U1650 (N_1650,In_653,In_2753);
xnor U1651 (N_1651,In_2935,In_1872);
nor U1652 (N_1652,In_1419,In_2030);
and U1653 (N_1653,In_1897,In_2295);
nor U1654 (N_1654,In_800,In_2105);
nand U1655 (N_1655,In_454,In_2837);
xnor U1656 (N_1656,In_2223,In_2365);
or U1657 (N_1657,In_1734,In_1217);
nand U1658 (N_1658,In_2204,In_1432);
and U1659 (N_1659,In_503,In_966);
nor U1660 (N_1660,In_872,In_1932);
or U1661 (N_1661,In_2622,In_2836);
nor U1662 (N_1662,In_363,In_2787);
nor U1663 (N_1663,In_2249,In_2849);
xnor U1664 (N_1664,In_1784,In_719);
xor U1665 (N_1665,In_1780,In_206);
nor U1666 (N_1666,In_1643,In_689);
or U1667 (N_1667,In_2672,In_188);
xnor U1668 (N_1668,In_1497,In_2742);
or U1669 (N_1669,In_1689,In_2021);
xor U1670 (N_1670,In_749,In_2459);
xnor U1671 (N_1671,In_207,In_1101);
xor U1672 (N_1672,In_1177,In_2127);
xor U1673 (N_1673,In_608,In_2069);
nand U1674 (N_1674,In_2046,In_2437);
nor U1675 (N_1675,In_2572,In_2819);
or U1676 (N_1676,In_421,In_1281);
nor U1677 (N_1677,In_2249,In_2382);
nor U1678 (N_1678,In_1659,In_679);
or U1679 (N_1679,In_97,In_2297);
nand U1680 (N_1680,In_1594,In_2594);
nand U1681 (N_1681,In_83,In_2314);
nor U1682 (N_1682,In_2732,In_2531);
or U1683 (N_1683,In_1010,In_2394);
xor U1684 (N_1684,In_2428,In_1658);
or U1685 (N_1685,In_2758,In_2733);
and U1686 (N_1686,In_928,In_1474);
xor U1687 (N_1687,In_2126,In_306);
nand U1688 (N_1688,In_2547,In_186);
nand U1689 (N_1689,In_1472,In_2221);
nor U1690 (N_1690,In_2301,In_2941);
nand U1691 (N_1691,In_1184,In_2623);
or U1692 (N_1692,In_1794,In_1098);
nand U1693 (N_1693,In_2697,In_2419);
xnor U1694 (N_1694,In_2859,In_2280);
nand U1695 (N_1695,In_2327,In_2155);
xor U1696 (N_1696,In_892,In_1583);
xnor U1697 (N_1697,In_2860,In_1975);
xor U1698 (N_1698,In_29,In_1950);
nor U1699 (N_1699,In_2897,In_721);
nor U1700 (N_1700,In_573,In_778);
and U1701 (N_1701,In_1422,In_2971);
and U1702 (N_1702,In_2465,In_2906);
nand U1703 (N_1703,In_2377,In_2959);
or U1704 (N_1704,In_2541,In_268);
nor U1705 (N_1705,In_1282,In_2376);
xor U1706 (N_1706,In_170,In_1756);
nand U1707 (N_1707,In_1081,In_2515);
or U1708 (N_1708,In_2805,In_2313);
nand U1709 (N_1709,In_1898,In_1343);
xnor U1710 (N_1710,In_618,In_721);
nor U1711 (N_1711,In_306,In_44);
xnor U1712 (N_1712,In_356,In_78);
and U1713 (N_1713,In_866,In_1315);
and U1714 (N_1714,In_1725,In_2171);
nand U1715 (N_1715,In_1605,In_1953);
xnor U1716 (N_1716,In_1386,In_1856);
and U1717 (N_1717,In_1379,In_871);
or U1718 (N_1718,In_2956,In_1148);
and U1719 (N_1719,In_1854,In_1870);
nand U1720 (N_1720,In_2213,In_1258);
xnor U1721 (N_1721,In_2371,In_2194);
or U1722 (N_1722,In_2964,In_2156);
or U1723 (N_1723,In_1550,In_933);
nor U1724 (N_1724,In_2004,In_2035);
or U1725 (N_1725,In_2746,In_22);
nand U1726 (N_1726,In_263,In_2450);
xnor U1727 (N_1727,In_1450,In_2010);
xnor U1728 (N_1728,In_2001,In_219);
nor U1729 (N_1729,In_2621,In_1466);
xor U1730 (N_1730,In_664,In_514);
or U1731 (N_1731,In_458,In_314);
nand U1732 (N_1732,In_2273,In_2767);
and U1733 (N_1733,In_1395,In_276);
nor U1734 (N_1734,In_8,In_1946);
or U1735 (N_1735,In_2235,In_662);
nand U1736 (N_1736,In_1723,In_2375);
nor U1737 (N_1737,In_776,In_579);
nor U1738 (N_1738,In_1943,In_959);
nor U1739 (N_1739,In_616,In_1189);
or U1740 (N_1740,In_2963,In_581);
and U1741 (N_1741,In_2155,In_1200);
xnor U1742 (N_1742,In_968,In_1107);
or U1743 (N_1743,In_2932,In_1128);
nand U1744 (N_1744,In_517,In_571);
and U1745 (N_1745,In_2973,In_2118);
and U1746 (N_1746,In_849,In_2282);
xnor U1747 (N_1747,In_2395,In_2070);
or U1748 (N_1748,In_703,In_1646);
and U1749 (N_1749,In_1886,In_587);
xnor U1750 (N_1750,In_987,In_1057);
or U1751 (N_1751,In_748,In_830);
or U1752 (N_1752,In_2602,In_531);
or U1753 (N_1753,In_227,In_97);
or U1754 (N_1754,In_659,In_1021);
and U1755 (N_1755,In_193,In_1272);
and U1756 (N_1756,In_1708,In_123);
nor U1757 (N_1757,In_394,In_960);
nand U1758 (N_1758,In_2731,In_1750);
and U1759 (N_1759,In_2992,In_116);
or U1760 (N_1760,In_460,In_1471);
nand U1761 (N_1761,In_10,In_470);
and U1762 (N_1762,In_848,In_1053);
nor U1763 (N_1763,In_2532,In_1031);
xor U1764 (N_1764,In_742,In_2342);
or U1765 (N_1765,In_2121,In_2504);
or U1766 (N_1766,In_1096,In_1905);
nor U1767 (N_1767,In_2891,In_816);
or U1768 (N_1768,In_383,In_625);
nand U1769 (N_1769,In_1333,In_1043);
nor U1770 (N_1770,In_1295,In_1562);
and U1771 (N_1771,In_1846,In_1193);
nand U1772 (N_1772,In_520,In_2452);
nor U1773 (N_1773,In_1372,In_2233);
xor U1774 (N_1774,In_2186,In_597);
or U1775 (N_1775,In_1477,In_538);
xor U1776 (N_1776,In_2090,In_1464);
xnor U1777 (N_1777,In_1214,In_497);
xnor U1778 (N_1778,In_1857,In_622);
nor U1779 (N_1779,In_1313,In_1007);
nor U1780 (N_1780,In_1985,In_66);
nor U1781 (N_1781,In_2545,In_2747);
xnor U1782 (N_1782,In_762,In_700);
xor U1783 (N_1783,In_2011,In_2586);
nand U1784 (N_1784,In_2771,In_1810);
nor U1785 (N_1785,In_2946,In_2677);
or U1786 (N_1786,In_483,In_2977);
or U1787 (N_1787,In_1348,In_2470);
and U1788 (N_1788,In_1312,In_1971);
xor U1789 (N_1789,In_1843,In_2867);
xnor U1790 (N_1790,In_1962,In_2649);
xnor U1791 (N_1791,In_1108,In_1190);
or U1792 (N_1792,In_2932,In_1571);
and U1793 (N_1793,In_1239,In_2323);
or U1794 (N_1794,In_201,In_2991);
xnor U1795 (N_1795,In_788,In_528);
nand U1796 (N_1796,In_1543,In_2946);
nand U1797 (N_1797,In_877,In_1643);
nand U1798 (N_1798,In_812,In_759);
and U1799 (N_1799,In_2914,In_178);
nand U1800 (N_1800,In_213,In_2761);
or U1801 (N_1801,In_385,In_1824);
nor U1802 (N_1802,In_2612,In_167);
and U1803 (N_1803,In_983,In_2577);
nor U1804 (N_1804,In_1070,In_2989);
or U1805 (N_1805,In_1520,In_1571);
and U1806 (N_1806,In_1209,In_520);
nand U1807 (N_1807,In_1194,In_579);
nand U1808 (N_1808,In_755,In_2645);
nand U1809 (N_1809,In_1821,In_2046);
and U1810 (N_1810,In_700,In_2575);
or U1811 (N_1811,In_374,In_15);
nor U1812 (N_1812,In_39,In_2698);
or U1813 (N_1813,In_2285,In_1772);
and U1814 (N_1814,In_2555,In_2512);
nand U1815 (N_1815,In_2108,In_436);
nand U1816 (N_1816,In_1152,In_2372);
nand U1817 (N_1817,In_1289,In_1790);
and U1818 (N_1818,In_323,In_1398);
nand U1819 (N_1819,In_2672,In_2013);
or U1820 (N_1820,In_889,In_1873);
nor U1821 (N_1821,In_2043,In_2245);
nand U1822 (N_1822,In_2776,In_2847);
xor U1823 (N_1823,In_2675,In_294);
nor U1824 (N_1824,In_2612,In_958);
nand U1825 (N_1825,In_2386,In_1488);
nor U1826 (N_1826,In_1068,In_2448);
nand U1827 (N_1827,In_1796,In_1739);
or U1828 (N_1828,In_2375,In_263);
and U1829 (N_1829,In_2462,In_185);
and U1830 (N_1830,In_1440,In_2514);
nor U1831 (N_1831,In_1564,In_449);
xor U1832 (N_1832,In_471,In_1345);
and U1833 (N_1833,In_1560,In_2256);
xnor U1834 (N_1834,In_1327,In_759);
and U1835 (N_1835,In_2951,In_2656);
nand U1836 (N_1836,In_45,In_1040);
xnor U1837 (N_1837,In_134,In_478);
xor U1838 (N_1838,In_2951,In_1516);
nand U1839 (N_1839,In_2671,In_1750);
or U1840 (N_1840,In_2749,In_2916);
xor U1841 (N_1841,In_288,In_2668);
and U1842 (N_1842,In_1201,In_2458);
and U1843 (N_1843,In_2080,In_753);
nand U1844 (N_1844,In_2734,In_1512);
xor U1845 (N_1845,In_1212,In_1071);
and U1846 (N_1846,In_2576,In_1637);
xnor U1847 (N_1847,In_1098,In_2115);
xor U1848 (N_1848,In_1196,In_1258);
nand U1849 (N_1849,In_1208,In_1721);
xnor U1850 (N_1850,In_2562,In_2060);
nand U1851 (N_1851,In_1966,In_2185);
nor U1852 (N_1852,In_1665,In_459);
or U1853 (N_1853,In_263,In_1796);
and U1854 (N_1854,In_289,In_322);
and U1855 (N_1855,In_2943,In_2310);
or U1856 (N_1856,In_1358,In_459);
or U1857 (N_1857,In_2571,In_491);
nor U1858 (N_1858,In_1081,In_46);
or U1859 (N_1859,In_2074,In_995);
xor U1860 (N_1860,In_891,In_152);
nand U1861 (N_1861,In_2226,In_2840);
xor U1862 (N_1862,In_51,In_695);
or U1863 (N_1863,In_1314,In_1151);
and U1864 (N_1864,In_1527,In_2149);
and U1865 (N_1865,In_64,In_2365);
nor U1866 (N_1866,In_1396,In_1452);
and U1867 (N_1867,In_2061,In_2839);
and U1868 (N_1868,In_1962,In_2002);
or U1869 (N_1869,In_1525,In_1359);
nand U1870 (N_1870,In_1450,In_181);
xnor U1871 (N_1871,In_210,In_917);
or U1872 (N_1872,In_2742,In_2026);
nor U1873 (N_1873,In_2286,In_1571);
or U1874 (N_1874,In_745,In_2888);
and U1875 (N_1875,In_1887,In_653);
and U1876 (N_1876,In_2323,In_121);
or U1877 (N_1877,In_2118,In_963);
nand U1878 (N_1878,In_2889,In_381);
nor U1879 (N_1879,In_2352,In_928);
xnor U1880 (N_1880,In_1820,In_1934);
xnor U1881 (N_1881,In_881,In_2027);
xor U1882 (N_1882,In_1838,In_842);
nor U1883 (N_1883,In_207,In_2876);
nor U1884 (N_1884,In_1305,In_2984);
xnor U1885 (N_1885,In_1962,In_689);
nor U1886 (N_1886,In_1476,In_930);
xnor U1887 (N_1887,In_1828,In_2968);
xnor U1888 (N_1888,In_1999,In_443);
and U1889 (N_1889,In_734,In_2569);
nand U1890 (N_1890,In_963,In_1660);
or U1891 (N_1891,In_2040,In_2024);
nand U1892 (N_1892,In_304,In_1715);
xnor U1893 (N_1893,In_2866,In_985);
or U1894 (N_1894,In_1540,In_2641);
xnor U1895 (N_1895,In_163,In_1276);
and U1896 (N_1896,In_1109,In_2615);
nand U1897 (N_1897,In_498,In_1315);
nor U1898 (N_1898,In_1853,In_1786);
nand U1899 (N_1899,In_901,In_1416);
and U1900 (N_1900,In_1181,In_1718);
xnor U1901 (N_1901,In_1785,In_1840);
and U1902 (N_1902,In_2422,In_386);
xor U1903 (N_1903,In_352,In_1669);
xor U1904 (N_1904,In_788,In_2310);
nand U1905 (N_1905,In_1501,In_492);
xnor U1906 (N_1906,In_185,In_233);
and U1907 (N_1907,In_20,In_1982);
nand U1908 (N_1908,In_746,In_621);
nand U1909 (N_1909,In_1679,In_1193);
xnor U1910 (N_1910,In_2630,In_2449);
nor U1911 (N_1911,In_1912,In_172);
xnor U1912 (N_1912,In_2269,In_2152);
and U1913 (N_1913,In_1723,In_184);
and U1914 (N_1914,In_19,In_524);
nor U1915 (N_1915,In_2291,In_2373);
or U1916 (N_1916,In_1172,In_2323);
nor U1917 (N_1917,In_104,In_2385);
or U1918 (N_1918,In_1457,In_966);
xor U1919 (N_1919,In_430,In_861);
or U1920 (N_1920,In_1299,In_951);
or U1921 (N_1921,In_313,In_2117);
or U1922 (N_1922,In_2364,In_1505);
nor U1923 (N_1923,In_2289,In_1388);
nand U1924 (N_1924,In_1568,In_2774);
and U1925 (N_1925,In_915,In_897);
or U1926 (N_1926,In_1498,In_1627);
or U1927 (N_1927,In_64,In_434);
and U1928 (N_1928,In_301,In_2155);
or U1929 (N_1929,In_2553,In_2361);
nor U1930 (N_1930,In_1838,In_810);
nand U1931 (N_1931,In_489,In_2634);
or U1932 (N_1932,In_63,In_367);
nand U1933 (N_1933,In_1068,In_2619);
or U1934 (N_1934,In_1279,In_1025);
xor U1935 (N_1935,In_1997,In_1350);
xnor U1936 (N_1936,In_1209,In_853);
and U1937 (N_1937,In_2251,In_192);
or U1938 (N_1938,In_688,In_2271);
or U1939 (N_1939,In_583,In_1157);
and U1940 (N_1940,In_1845,In_1654);
or U1941 (N_1941,In_866,In_2024);
nor U1942 (N_1942,In_1722,In_738);
nand U1943 (N_1943,In_2835,In_177);
or U1944 (N_1944,In_2792,In_816);
xnor U1945 (N_1945,In_2973,In_1558);
or U1946 (N_1946,In_1460,In_2897);
nor U1947 (N_1947,In_78,In_1894);
and U1948 (N_1948,In_1979,In_528);
nand U1949 (N_1949,In_1714,In_65);
nor U1950 (N_1950,In_618,In_550);
nor U1951 (N_1951,In_2891,In_885);
or U1952 (N_1952,In_2678,In_696);
nor U1953 (N_1953,In_1857,In_1441);
and U1954 (N_1954,In_1072,In_892);
nand U1955 (N_1955,In_1856,In_1720);
xor U1956 (N_1956,In_1176,In_2425);
and U1957 (N_1957,In_205,In_880);
xnor U1958 (N_1958,In_1351,In_2313);
xnor U1959 (N_1959,In_2107,In_2603);
or U1960 (N_1960,In_1656,In_2179);
and U1961 (N_1961,In_2690,In_534);
xor U1962 (N_1962,In_2521,In_187);
or U1963 (N_1963,In_1521,In_194);
or U1964 (N_1964,In_1600,In_2165);
or U1965 (N_1965,In_306,In_742);
and U1966 (N_1966,In_2725,In_279);
xor U1967 (N_1967,In_2477,In_774);
or U1968 (N_1968,In_2184,In_259);
nor U1969 (N_1969,In_1296,In_2797);
xnor U1970 (N_1970,In_745,In_2719);
nor U1971 (N_1971,In_172,In_2760);
and U1972 (N_1972,In_2330,In_71);
nor U1973 (N_1973,In_2194,In_1615);
and U1974 (N_1974,In_1145,In_824);
nor U1975 (N_1975,In_2155,In_1134);
xnor U1976 (N_1976,In_335,In_2497);
nor U1977 (N_1977,In_1580,In_1252);
or U1978 (N_1978,In_1291,In_121);
xor U1979 (N_1979,In_1030,In_1673);
or U1980 (N_1980,In_2593,In_2396);
xnor U1981 (N_1981,In_1685,In_2849);
or U1982 (N_1982,In_1161,In_2348);
or U1983 (N_1983,In_200,In_262);
xor U1984 (N_1984,In_193,In_2245);
and U1985 (N_1985,In_2489,In_1920);
nand U1986 (N_1986,In_1315,In_894);
and U1987 (N_1987,In_1231,In_1704);
nand U1988 (N_1988,In_2017,In_1143);
nor U1989 (N_1989,In_1031,In_2670);
nand U1990 (N_1990,In_1803,In_1684);
nand U1991 (N_1991,In_2637,In_1074);
nand U1992 (N_1992,In_1598,In_2197);
xor U1993 (N_1993,In_2387,In_1757);
or U1994 (N_1994,In_560,In_605);
xnor U1995 (N_1995,In_664,In_968);
and U1996 (N_1996,In_1195,In_1451);
or U1997 (N_1997,In_239,In_500);
xnor U1998 (N_1998,In_677,In_2583);
and U1999 (N_1999,In_2996,In_357);
nor U2000 (N_2000,N_1889,N_308);
and U2001 (N_2001,N_1246,N_1346);
or U2002 (N_2002,N_1549,N_1303);
or U2003 (N_2003,N_506,N_666);
nor U2004 (N_2004,N_1944,N_811);
nand U2005 (N_2005,N_1709,N_1379);
and U2006 (N_2006,N_1050,N_1197);
nor U2007 (N_2007,N_971,N_297);
nand U2008 (N_2008,N_658,N_252);
and U2009 (N_2009,N_1957,N_156);
and U2010 (N_2010,N_498,N_1684);
xnor U2011 (N_2011,N_647,N_1177);
and U2012 (N_2012,N_1567,N_448);
nand U2013 (N_2013,N_675,N_1774);
xnor U2014 (N_2014,N_19,N_1527);
nand U2015 (N_2015,N_578,N_492);
or U2016 (N_2016,N_1705,N_998);
nand U2017 (N_2017,N_1750,N_1471);
or U2018 (N_2018,N_1912,N_1490);
nand U2019 (N_2019,N_303,N_1109);
nand U2020 (N_2020,N_1036,N_1221);
and U2021 (N_2021,N_653,N_195);
or U2022 (N_2022,N_1649,N_97);
nor U2023 (N_2023,N_75,N_173);
and U2024 (N_2024,N_1333,N_287);
or U2025 (N_2025,N_322,N_103);
nand U2026 (N_2026,N_1207,N_1331);
or U2027 (N_2027,N_1658,N_275);
xnor U2028 (N_2028,N_736,N_662);
or U2029 (N_2029,N_990,N_1236);
nand U2030 (N_2030,N_1932,N_1640);
or U2031 (N_2031,N_686,N_503);
and U2032 (N_2032,N_1962,N_119);
and U2033 (N_2033,N_810,N_1343);
or U2034 (N_2034,N_70,N_1464);
and U2035 (N_2035,N_814,N_1964);
nor U2036 (N_2036,N_1818,N_1626);
or U2037 (N_2037,N_861,N_1310);
and U2038 (N_2038,N_419,N_1831);
and U2039 (N_2039,N_1934,N_1526);
nor U2040 (N_2040,N_299,N_237);
xor U2041 (N_2041,N_1542,N_1140);
or U2042 (N_2042,N_1332,N_1554);
or U2043 (N_2043,N_1399,N_1132);
nand U2044 (N_2044,N_1082,N_1564);
and U2045 (N_2045,N_1169,N_1397);
and U2046 (N_2046,N_842,N_1569);
and U2047 (N_2047,N_769,N_495);
nor U2048 (N_2048,N_777,N_228);
and U2049 (N_2049,N_1503,N_869);
and U2050 (N_2050,N_1773,N_460);
xnor U2051 (N_2051,N_1222,N_455);
or U2052 (N_2052,N_420,N_363);
nand U2053 (N_2053,N_1720,N_1173);
xnor U2054 (N_2054,N_440,N_213);
nand U2055 (N_2055,N_1297,N_1308);
or U2056 (N_2056,N_1877,N_596);
nand U2057 (N_2057,N_106,N_1941);
nand U2058 (N_2058,N_533,N_1698);
and U2059 (N_2059,N_1090,N_1585);
nor U2060 (N_2060,N_997,N_1270);
nor U2061 (N_2061,N_1563,N_25);
and U2062 (N_2062,N_1905,N_1063);
or U2063 (N_2063,N_1849,N_52);
or U2064 (N_2064,N_819,N_1095);
nor U2065 (N_2065,N_1494,N_1195);
and U2066 (N_2066,N_1410,N_940);
nor U2067 (N_2067,N_130,N_806);
nor U2068 (N_2068,N_1779,N_843);
and U2069 (N_2069,N_1495,N_1977);
and U2070 (N_2070,N_630,N_1047);
or U2071 (N_2071,N_1571,N_1361);
nand U2072 (N_2072,N_678,N_974);
xnor U2073 (N_2073,N_771,N_54);
xor U2074 (N_2074,N_1020,N_1989);
nand U2075 (N_2075,N_330,N_1428);
and U2076 (N_2076,N_1008,N_598);
nand U2077 (N_2077,N_668,N_165);
nand U2078 (N_2078,N_1943,N_946);
nor U2079 (N_2079,N_1443,N_1817);
or U2080 (N_2080,N_170,N_1556);
or U2081 (N_2081,N_501,N_584);
or U2082 (N_2082,N_1670,N_705);
nor U2083 (N_2083,N_952,N_133);
xnor U2084 (N_2084,N_1666,N_1856);
xor U2085 (N_2085,N_579,N_1199);
and U2086 (N_2086,N_1074,N_1775);
or U2087 (N_2087,N_527,N_1122);
and U2088 (N_2088,N_788,N_1088);
and U2089 (N_2089,N_982,N_374);
xor U2090 (N_2090,N_1159,N_1902);
and U2091 (N_2091,N_1472,N_354);
xor U2092 (N_2092,N_1129,N_111);
or U2093 (N_2093,N_1888,N_1809);
xnor U2094 (N_2094,N_922,N_1712);
nand U2095 (N_2095,N_1386,N_101);
and U2096 (N_2096,N_459,N_1694);
nand U2097 (N_2097,N_1198,N_1845);
nand U2098 (N_2098,N_548,N_1104);
or U2099 (N_2099,N_1053,N_1078);
xnor U2100 (N_2100,N_1741,N_642);
nand U2101 (N_2101,N_373,N_5);
xnor U2102 (N_2102,N_933,N_875);
or U2103 (N_2103,N_416,N_739);
or U2104 (N_2104,N_857,N_1073);
and U2105 (N_2105,N_1059,N_882);
nor U2106 (N_2106,N_1474,N_905);
xnor U2107 (N_2107,N_1422,N_337);
nand U2108 (N_2108,N_765,N_568);
or U2109 (N_2109,N_439,N_988);
xor U2110 (N_2110,N_123,N_1730);
or U2111 (N_2111,N_1016,N_741);
nor U2112 (N_2112,N_1478,N_1972);
and U2113 (N_2113,N_462,N_267);
xor U2114 (N_2114,N_1174,N_518);
nor U2115 (N_2115,N_1239,N_163);
nor U2116 (N_2116,N_1484,N_586);
or U2117 (N_2117,N_1430,N_1017);
nor U2118 (N_2118,N_384,N_1229);
or U2119 (N_2119,N_13,N_1249);
nand U2120 (N_2120,N_64,N_190);
xor U2121 (N_2121,N_394,N_189);
or U2122 (N_2122,N_733,N_1979);
and U2123 (N_2123,N_361,N_684);
nor U2124 (N_2124,N_1287,N_744);
and U2125 (N_2125,N_1228,N_1058);
nand U2126 (N_2126,N_632,N_604);
xor U2127 (N_2127,N_749,N_1141);
nor U2128 (N_2128,N_1444,N_104);
nor U2129 (N_2129,N_1445,N_834);
or U2130 (N_2130,N_754,N_281);
nor U2131 (N_2131,N_1955,N_1760);
and U2132 (N_2132,N_274,N_211);
and U2133 (N_2133,N_405,N_1810);
or U2134 (N_2134,N_1152,N_1096);
xor U2135 (N_2135,N_32,N_1544);
nand U2136 (N_2136,N_1392,N_468);
nor U2137 (N_2137,N_567,N_1057);
and U2138 (N_2138,N_561,N_196);
nand U2139 (N_2139,N_88,N_471);
xor U2140 (N_2140,N_402,N_1457);
nand U2141 (N_2141,N_1300,N_1196);
nand U2142 (N_2142,N_1796,N_1646);
xor U2143 (N_2143,N_1407,N_711);
xnor U2144 (N_2144,N_957,N_1751);
nor U2145 (N_2145,N_1041,N_1926);
xnor U2146 (N_2146,N_1248,N_396);
nand U2147 (N_2147,N_784,N_1841);
xor U2148 (N_2148,N_1328,N_535);
xnor U2149 (N_2149,N_450,N_531);
or U2150 (N_2150,N_1857,N_774);
and U2151 (N_2151,N_1752,N_981);
and U2152 (N_2152,N_1587,N_1986);
xnor U2153 (N_2153,N_232,N_43);
nor U2154 (N_2154,N_929,N_102);
nor U2155 (N_2155,N_86,N_142);
xor U2156 (N_2156,N_890,N_1367);
nand U2157 (N_2157,N_472,N_883);
or U2158 (N_2158,N_1903,N_3);
nor U2159 (N_2159,N_665,N_1434);
nand U2160 (N_2160,N_1825,N_1700);
nand U2161 (N_2161,N_209,N_1133);
nand U2162 (N_2162,N_1915,N_1015);
xor U2163 (N_2163,N_1225,N_1524);
nand U2164 (N_2164,N_277,N_1098);
xor U2165 (N_2165,N_1675,N_900);
and U2166 (N_2166,N_723,N_1769);
and U2167 (N_2167,N_783,N_1929);
nor U2168 (N_2168,N_781,N_114);
or U2169 (N_2169,N_184,N_848);
and U2170 (N_2170,N_790,N_1461);
nor U2171 (N_2171,N_689,N_706);
xor U2172 (N_2172,N_836,N_16);
nor U2173 (N_2173,N_227,N_325);
xnor U2174 (N_2174,N_704,N_1612);
xnor U2175 (N_2175,N_576,N_519);
nor U2176 (N_2176,N_71,N_934);
xnor U2177 (N_2177,N_1873,N_343);
nand U2178 (N_2178,N_26,N_1148);
nor U2179 (N_2179,N_1210,N_470);
nand U2180 (N_2180,N_1064,N_833);
xor U2181 (N_2181,N_1439,N_347);
and U2182 (N_2182,N_1488,N_1136);
or U2183 (N_2183,N_454,N_1548);
or U2184 (N_2184,N_1842,N_1650);
or U2185 (N_2185,N_1292,N_1353);
or U2186 (N_2186,N_641,N_832);
xor U2187 (N_2187,N_1493,N_1969);
nor U2188 (N_2188,N_558,N_1393);
or U2189 (N_2189,N_167,N_1628);
nor U2190 (N_2190,N_700,N_489);
and U2191 (N_2191,N_1150,N_1247);
or U2192 (N_2192,N_515,N_1261);
and U2193 (N_2193,N_1500,N_853);
or U2194 (N_2194,N_1010,N_961);
xnor U2195 (N_2195,N_1651,N_1718);
nor U2196 (N_2196,N_1324,N_1607);
nor U2197 (N_2197,N_939,N_1901);
nand U2198 (N_2198,N_796,N_1829);
nor U2199 (N_2199,N_913,N_1992);
nor U2200 (N_2200,N_1511,N_10);
and U2201 (N_2201,N_328,N_1865);
xnor U2202 (N_2202,N_645,N_614);
or U2203 (N_2203,N_15,N_1387);
nand U2204 (N_2204,N_608,N_96);
nand U2205 (N_2205,N_475,N_382);
nor U2206 (N_2206,N_538,N_1294);
or U2207 (N_2207,N_1509,N_594);
nand U2208 (N_2208,N_1258,N_135);
nor U2209 (N_2209,N_464,N_1147);
or U2210 (N_2210,N_1663,N_121);
and U2211 (N_2211,N_1031,N_1171);
nor U2212 (N_2212,N_1983,N_60);
xnor U2213 (N_2213,N_1999,N_1492);
nor U2214 (N_2214,N_391,N_1589);
nor U2215 (N_2215,N_1463,N_985);
nor U2216 (N_2216,N_422,N_1089);
nor U2217 (N_2217,N_1613,N_1762);
or U2218 (N_2218,N_891,N_992);
nand U2219 (N_2219,N_1719,N_1242);
xnor U2220 (N_2220,N_1798,N_873);
nor U2221 (N_2221,N_685,N_1723);
or U2222 (N_2222,N_17,N_1405);
xnor U2223 (N_2223,N_636,N_1925);
nor U2224 (N_2224,N_1900,N_480);
xnor U2225 (N_2225,N_461,N_1012);
and U2226 (N_2226,N_132,N_1470);
xor U2227 (N_2227,N_256,N_871);
nor U2228 (N_2228,N_1429,N_1037);
or U2229 (N_2229,N_523,N_755);
and U2230 (N_2230,N_1281,N_1562);
or U2231 (N_2231,N_807,N_0);
or U2232 (N_2232,N_65,N_1689);
and U2233 (N_2233,N_740,N_1459);
or U2234 (N_2234,N_158,N_1451);
xnor U2235 (N_2235,N_1413,N_964);
or U2236 (N_2236,N_399,N_1858);
nand U2237 (N_2237,N_1506,N_1203);
nor U2238 (N_2238,N_1508,N_888);
and U2239 (N_2239,N_839,N_1736);
nor U2240 (N_2240,N_1959,N_362);
xor U2241 (N_2241,N_591,N_1264);
nand U2242 (N_2242,N_296,N_1784);
and U2243 (N_2243,N_1610,N_1417);
or U2244 (N_2244,N_994,N_1114);
xnor U2245 (N_2245,N_1974,N_1603);
or U2246 (N_2246,N_1654,N_1418);
nor U2247 (N_2247,N_1921,N_366);
nor U2248 (N_2248,N_1595,N_657);
xor U2249 (N_2249,N_508,N_50);
and U2250 (N_2250,N_906,N_314);
nor U2251 (N_2251,N_878,N_1347);
and U2252 (N_2252,N_1906,N_400);
nor U2253 (N_2253,N_748,N_661);
and U2254 (N_2254,N_92,N_27);
and U2255 (N_2255,N_1642,N_1256);
xnor U2256 (N_2256,N_166,N_770);
or U2257 (N_2257,N_1739,N_1241);
or U2258 (N_2258,N_1803,N_1792);
nand U2259 (N_2259,N_476,N_85);
nand U2260 (N_2260,N_1048,N_682);
or U2261 (N_2261,N_681,N_247);
and U2262 (N_2262,N_1978,N_154);
nand U2263 (N_2263,N_203,N_432);
and U2264 (N_2264,N_1641,N_1458);
or U2265 (N_2265,N_1028,N_886);
nor U2266 (N_2266,N_1656,N_214);
nor U2267 (N_2267,N_1127,N_958);
and U2268 (N_2268,N_1269,N_491);
and U2269 (N_2269,N_1863,N_549);
xnor U2270 (N_2270,N_346,N_794);
nor U2271 (N_2271,N_1215,N_1910);
or U2272 (N_2272,N_1664,N_829);
or U2273 (N_2273,N_76,N_1312);
or U2274 (N_2274,N_1693,N_1100);
or U2275 (N_2275,N_671,N_947);
xor U2276 (N_2276,N_823,N_1305);
nand U2277 (N_2277,N_1625,N_1820);
or U2278 (N_2278,N_197,N_1446);
xor U2279 (N_2279,N_33,N_246);
and U2280 (N_2280,N_1685,N_1180);
nor U2281 (N_2281,N_1674,N_1273);
nor U2282 (N_2282,N_126,N_615);
nand U2283 (N_2283,N_644,N_320);
or U2284 (N_2284,N_1899,N_605);
xnor U2285 (N_2285,N_1194,N_626);
xor U2286 (N_2286,N_138,N_327);
nand U2287 (N_2287,N_1344,N_627);
nand U2288 (N_2288,N_802,N_124);
and U2289 (N_2289,N_772,N_932);
and U2290 (N_2290,N_667,N_659);
xor U2291 (N_2291,N_478,N_1348);
and U2292 (N_2292,N_1376,N_734);
or U2293 (N_2293,N_497,N_316);
nor U2294 (N_2294,N_437,N_1220);
nand U2295 (N_2295,N_1570,N_589);
nand U2296 (N_2296,N_1186,N_147);
xnor U2297 (N_2297,N_874,N_1620);
nor U2298 (N_2298,N_1091,N_1318);
nand U2299 (N_2299,N_1821,N_1178);
nor U2300 (N_2300,N_845,N_1237);
or U2301 (N_2301,N_1782,N_375);
nand U2302 (N_2302,N_118,N_1146);
nor U2303 (N_2303,N_1697,N_1802);
or U2304 (N_2304,N_481,N_731);
nand U2305 (N_2305,N_1665,N_1285);
nor U2306 (N_2306,N_1409,N_77);
xor U2307 (N_2307,N_1005,N_1815);
xnor U2308 (N_2308,N_973,N_1688);
xor U2309 (N_2309,N_306,N_1414);
xor U2310 (N_2310,N_1362,N_1812);
or U2311 (N_2311,N_1852,N_171);
or U2312 (N_2312,N_893,N_904);
and U2313 (N_2313,N_1371,N_1722);
nor U2314 (N_2314,N_813,N_707);
xor U2315 (N_2315,N_336,N_1584);
nor U2316 (N_2316,N_1531,N_1667);
and U2317 (N_2317,N_690,N_780);
or U2318 (N_2318,N_456,N_812);
xnor U2319 (N_2319,N_1891,N_1040);
nand U2320 (N_2320,N_804,N_380);
xor U2321 (N_2321,N_331,N_1853);
and U2322 (N_2322,N_1706,N_640);
nand U2323 (N_2323,N_553,N_1847);
nand U2324 (N_2324,N_1801,N_311);
xnor U2325 (N_2325,N_702,N_696);
nor U2326 (N_2326,N_1289,N_1864);
nand U2327 (N_2327,N_161,N_1381);
or U2328 (N_2328,N_240,N_999);
or U2329 (N_2329,N_332,N_1046);
or U2330 (N_2330,N_1499,N_513);
and U2331 (N_2331,N_127,N_1629);
nand U2332 (N_2332,N_715,N_951);
nand U2333 (N_2333,N_1257,N_319);
and U2334 (N_2334,N_151,N_1668);
or U2335 (N_2335,N_1102,N_517);
and U2336 (N_2336,N_1713,N_1271);
nand U2337 (N_2337,N_177,N_837);
nand U2338 (N_2338,N_1213,N_40);
or U2339 (N_2339,N_355,N_1763);
nor U2340 (N_2340,N_709,N_1093);
and U2341 (N_2341,N_944,N_1504);
or U2342 (N_2342,N_1683,N_1479);
nand U2343 (N_2343,N_773,N_1866);
xor U2344 (N_2344,N_881,N_372);
nand U2345 (N_2345,N_930,N_716);
and U2346 (N_2346,N_1183,N_729);
nand U2347 (N_2347,N_1475,N_1725);
nor U2348 (N_2348,N_387,N_344);
nand U2349 (N_2349,N_1936,N_187);
and U2350 (N_2350,N_863,N_620);
nand U2351 (N_2351,N_572,N_1816);
or U2352 (N_2352,N_750,N_443);
xnor U2353 (N_2353,N_1652,N_1365);
nor U2354 (N_2354,N_474,N_1505);
or U2355 (N_2355,N_699,N_1662);
and U2356 (N_2356,N_1609,N_188);
and U2357 (N_2357,N_1920,N_1594);
xnor U2358 (N_2358,N_1971,N_219);
xnor U2359 (N_2359,N_451,N_352);
or U2360 (N_2360,N_555,N_249);
nand U2361 (N_2361,N_182,N_1030);
or U2362 (N_2362,N_1937,N_270);
xnor U2363 (N_2363,N_1131,N_1756);
and U2364 (N_2364,N_683,N_1543);
and U2365 (N_2365,N_1070,N_1293);
nor U2366 (N_2366,N_1924,N_44);
and U2367 (N_2367,N_1582,N_1680);
nor U2368 (N_2368,N_1708,N_827);
or U2369 (N_2369,N_1276,N_1918);
xnor U2370 (N_2370,N_1072,N_315);
or U2371 (N_2371,N_1452,N_849);
and U2372 (N_2372,N_411,N_1184);
and U2373 (N_2373,N_1066,N_1994);
nand U2374 (N_2374,N_1118,N_864);
nor U2375 (N_2375,N_1370,N_1338);
xnor U2376 (N_2376,N_898,N_263);
xnor U2377 (N_2377,N_1211,N_1412);
and U2378 (N_2378,N_58,N_168);
and U2379 (N_2379,N_323,N_230);
nand U2380 (N_2380,N_1851,N_1309);
nand U2381 (N_2381,N_505,N_176);
xnor U2382 (N_2382,N_876,N_329);
xnor U2383 (N_2383,N_1356,N_424);
nand U2384 (N_2384,N_835,N_1797);
and U2385 (N_2385,N_1982,N_414);
and U2386 (N_2386,N_917,N_1254);
or U2387 (N_2387,N_49,N_1561);
and U2388 (N_2388,N_1454,N_634);
nor U2389 (N_2389,N_638,N_1787);
or U2390 (N_2390,N_1846,N_113);
nor U2391 (N_2391,N_1502,N_1243);
and U2392 (N_2392,N_390,N_376);
or U2393 (N_2393,N_1165,N_1075);
nor U2394 (N_2394,N_1111,N_674);
and U2395 (N_2395,N_1777,N_1436);
xnor U2396 (N_2396,N_703,N_1788);
nand U2397 (N_2397,N_826,N_108);
xor U2398 (N_2398,N_1726,N_1854);
xor U2399 (N_2399,N_63,N_95);
nand U2400 (N_2400,N_817,N_1876);
xor U2401 (N_2401,N_1768,N_321);
nand U2402 (N_2402,N_737,N_1168);
nand U2403 (N_2403,N_1704,N_157);
nand U2404 (N_2404,N_353,N_1345);
xnor U2405 (N_2405,N_379,N_1325);
or U2406 (N_2406,N_1933,N_1583);
and U2407 (N_2407,N_1185,N_570);
nor U2408 (N_2408,N_1151,N_447);
or U2409 (N_2409,N_1848,N_8);
xor U2410 (N_2410,N_1153,N_291);
nor U2411 (N_2411,N_1540,N_1014);
nor U2412 (N_2412,N_1251,N_1468);
or U2413 (N_2413,N_392,N_1621);
nor U2414 (N_2414,N_30,N_1604);
nor U2415 (N_2415,N_986,N_1106);
or U2416 (N_2416,N_824,N_365);
xnor U2417 (N_2417,N_1327,N_1678);
nand U2418 (N_2418,N_1080,N_1672);
nor U2419 (N_2419,N_356,N_1601);
and U2420 (N_2420,N_927,N_1882);
nor U2421 (N_2421,N_1702,N_766);
nor U2422 (N_2422,N_153,N_1455);
nor U2423 (N_2423,N_428,N_301);
and U2424 (N_2424,N_825,N_1602);
and U2425 (N_2425,N_1639,N_852);
xnor U2426 (N_2426,N_204,N_530);
nor U2427 (N_2427,N_1960,N_1340);
nor U2428 (N_2428,N_880,N_300);
and U2429 (N_2429,N_894,N_809);
or U2430 (N_2430,N_499,N_1135);
nor U2431 (N_2431,N_1265,N_960);
nand U2432 (N_2432,N_799,N_1988);
xor U2433 (N_2433,N_35,N_386);
nor U2434 (N_2434,N_1635,N_1330);
nand U2435 (N_2435,N_912,N_1872);
xnor U2436 (N_2436,N_1696,N_805);
and U2437 (N_2437,N_803,N_1512);
nand U2438 (N_2438,N_233,N_856);
nor U2439 (N_2439,N_742,N_250);
nor U2440 (N_2440,N_622,N_1052);
xnor U2441 (N_2441,N_87,N_672);
or U2442 (N_2442,N_200,N_159);
xnor U2443 (N_2443,N_225,N_324);
nor U2444 (N_2444,N_1002,N_925);
xor U2445 (N_2445,N_629,N_226);
nand U2446 (N_2446,N_68,N_692);
and U2447 (N_2447,N_643,N_1586);
or U2448 (N_2448,N_473,N_1482);
or U2449 (N_2449,N_1,N_1939);
nor U2450 (N_2450,N_1887,N_924);
nand U2451 (N_2451,N_1591,N_1208);
or U2452 (N_2452,N_406,N_1374);
or U2453 (N_2453,N_430,N_800);
or U2454 (N_2454,N_983,N_1749);
xnor U2455 (N_2455,N_1170,N_1204);
nor U2456 (N_2456,N_984,N_290);
and U2457 (N_2457,N_1322,N_820);
and U2458 (N_2458,N_1794,N_1808);
nand U2459 (N_2459,N_916,N_1137);
and U2460 (N_2460,N_1634,N_1023);
nor U2461 (N_2461,N_1401,N_1335);
and U2462 (N_2462,N_335,N_1703);
nor U2463 (N_2463,N_1867,N_1081);
and U2464 (N_2464,N_1862,N_131);
or U2465 (N_2465,N_646,N_1886);
nand U2466 (N_2466,N_409,N_1216);
nand U2467 (N_2467,N_1245,N_1715);
nor U2468 (N_2468,N_1307,N_341);
nand U2469 (N_2469,N_1800,N_1804);
nor U2470 (N_2470,N_1369,N_1441);
xor U2471 (N_2471,N_494,N_979);
and U2472 (N_2472,N_1973,N_312);
nor U2473 (N_2473,N_1290,N_996);
xnor U2474 (N_2474,N_1522,N_1230);
or U2475 (N_2475,N_479,N_1767);
or U2476 (N_2476,N_1315,N_1402);
nor U2477 (N_2477,N_1416,N_808);
xnor U2478 (N_2478,N_1596,N_921);
xnor U2479 (N_2479,N_66,N_500);
nand U2480 (N_2480,N_1227,N_738);
and U2481 (N_2481,N_1627,N_207);
xnor U2482 (N_2482,N_587,N_1489);
xnor U2483 (N_2483,N_1728,N_600);
or U2484 (N_2484,N_1298,N_1566);
nor U2485 (N_2485,N_956,N_791);
nor U2486 (N_2486,N_1590,N_1615);
nor U2487 (N_2487,N_968,N_1277);
or U2488 (N_2488,N_1415,N_1956);
or U2489 (N_2489,N_1477,N_655);
xor U2490 (N_2490,N_1669,N_23);
or U2491 (N_2491,N_1067,N_94);
nand U2492 (N_2492,N_1952,N_1234);
nand U2493 (N_2493,N_537,N_889);
xnor U2494 (N_2494,N_486,N_529);
or U2495 (N_2495,N_1027,N_278);
and U2496 (N_2496,N_434,N_417);
nand U2497 (N_2497,N_1286,N_745);
xnor U2498 (N_2498,N_569,N_1746);
nand U2499 (N_2499,N_69,N_1949);
nand U2500 (N_2500,N_1025,N_199);
and U2501 (N_2501,N_789,N_1717);
nor U2502 (N_2502,N_1976,N_1744);
nor U2503 (N_2503,N_1568,N_1007);
nor U2504 (N_2504,N_1737,N_453);
xnor U2505 (N_2505,N_1442,N_1167);
or U2506 (N_2506,N_1776,N_51);
nor U2507 (N_2507,N_144,N_611);
nand U2508 (N_2508,N_185,N_465);
nand U2509 (N_2509,N_1657,N_1288);
xor U2510 (N_2510,N_717,N_963);
nand U2511 (N_2511,N_284,N_1835);
or U2512 (N_2512,N_1212,N_78);
nor U2513 (N_2513,N_1618,N_962);
xor U2514 (N_2514,N_840,N_107);
nor U2515 (N_2515,N_574,N_1671);
nor U2516 (N_2516,N_1535,N_1130);
xor U2517 (N_2517,N_1143,N_937);
nor U2518 (N_2518,N_725,N_1144);
or U2519 (N_2519,N_902,N_1581);
nand U2520 (N_2520,N_46,N_268);
or U2521 (N_2521,N_1385,N_838);
nor U2522 (N_2522,N_1018,N_1614);
nand U2523 (N_2523,N_1447,N_1469);
nor U2524 (N_2524,N_191,N_273);
and U2525 (N_2525,N_1967,N_1633);
and U2526 (N_2526,N_1765,N_1101);
or U2527 (N_2527,N_467,N_493);
or U2528 (N_2528,N_433,N_1206);
nand U2529 (N_2529,N_452,N_318);
nand U2530 (N_2530,N_1467,N_1354);
or U2531 (N_2531,N_532,N_1968);
nor U2532 (N_2532,N_1121,N_1984);
and U2533 (N_2533,N_1259,N_1400);
nor U2534 (N_2534,N_413,N_1278);
or U2535 (N_2535,N_1466,N_56);
xor U2536 (N_2536,N_602,N_282);
nand U2537 (N_2537,N_1483,N_1079);
or U2538 (N_2538,N_1553,N_410);
nor U2539 (N_2539,N_79,N_1930);
and U2540 (N_2540,N_1546,N_911);
and U2541 (N_2541,N_1188,N_313);
nand U2542 (N_2542,N_1116,N_1826);
and U2543 (N_2543,N_1110,N_1735);
nand U2544 (N_2544,N_1911,N_1682);
nor U2545 (N_2545,N_116,N_955);
or U2546 (N_2546,N_1631,N_349);
nor U2547 (N_2547,N_20,N_757);
nand U2548 (N_2548,N_206,N_1084);
nand U2549 (N_2549,N_1313,N_1837);
nand U2550 (N_2550,N_1721,N_1420);
or U2551 (N_2551,N_792,N_285);
xor U2552 (N_2552,N_616,N_1557);
nor U2553 (N_2553,N_1827,N_1895);
nand U2554 (N_2554,N_220,N_248);
nor U2555 (N_2555,N_669,N_1062);
and U2556 (N_2556,N_82,N_431);
xnor U2557 (N_2557,N_348,N_762);
xor U2558 (N_2558,N_59,N_1380);
or U2559 (N_2559,N_1648,N_1859);
and U2560 (N_2560,N_1056,N_1179);
or U2561 (N_2561,N_977,N_698);
nor U2562 (N_2562,N_907,N_1883);
and U2563 (N_2563,N_1965,N_1339);
nand U2564 (N_2564,N_1908,N_1341);
nand U2565 (N_2565,N_160,N_469);
nor U2566 (N_2566,N_412,N_609);
nor U2567 (N_2567,N_1431,N_243);
and U2568 (N_2568,N_859,N_39);
and U2569 (N_2569,N_162,N_421);
and U2570 (N_2570,N_1395,N_1398);
nand U2571 (N_2571,N_989,N_1250);
nand U2572 (N_2572,N_1519,N_1574);
and U2573 (N_2573,N_1172,N_1537);
and U2574 (N_2574,N_1192,N_1742);
nand U2575 (N_2575,N_502,N_987);
xnor U2576 (N_2576,N_368,N_1753);
nor U2577 (N_2577,N_1359,N_1946);
xor U2578 (N_2578,N_1238,N_1731);
and U2579 (N_2579,N_67,N_202);
and U2580 (N_2580,N_242,N_143);
nor U2581 (N_2581,N_942,N_1071);
and U2582 (N_2582,N_266,N_855);
and U2583 (N_2583,N_993,N_1043);
xnor U2584 (N_2584,N_1793,N_631);
xnor U2585 (N_2585,N_45,N_520);
nor U2586 (N_2586,N_1755,N_1272);
nor U2587 (N_2587,N_1154,N_1606);
and U2588 (N_2588,N_235,N_1126);
nand U2589 (N_2589,N_1319,N_1991);
nand U2590 (N_2590,N_959,N_152);
or U2591 (N_2591,N_484,N_90);
xor U2592 (N_2592,N_1404,N_1822);
nor U2593 (N_2593,N_593,N_407);
or U2594 (N_2594,N_650,N_1868);
xor U2595 (N_2595,N_637,N_1611);
nand U2596 (N_2596,N_1103,N_726);
nand U2597 (N_2597,N_231,N_970);
xnor U2598 (N_2598,N_1433,N_1097);
and U2599 (N_2599,N_1954,N_721);
nand U2600 (N_2600,N_150,N_401);
xnor U2601 (N_2601,N_1661,N_241);
nor U2602 (N_2602,N_818,N_1790);
nand U2603 (N_2603,N_1382,N_1938);
or U2604 (N_2604,N_743,N_1843);
and U2605 (N_2605,N_169,N_1026);
xnor U2606 (N_2606,N_31,N_948);
and U2607 (N_2607,N_1985,N_1560);
and U2608 (N_2608,N_1855,N_487);
or U2609 (N_2609,N_1860,N_926);
nand U2610 (N_2610,N_1534,N_438);
or U2611 (N_2611,N_1187,N_1497);
or U2612 (N_2612,N_1158,N_81);
and U2613 (N_2613,N_403,N_128);
nand U2614 (N_2614,N_1734,N_560);
and U2615 (N_2615,N_680,N_1659);
xor U2616 (N_2616,N_1572,N_545);
or U2617 (N_2617,N_1958,N_80);
and U2618 (N_2618,N_1232,N_1350);
nand U2619 (N_2619,N_1280,N_1233);
and U2620 (N_2620,N_1510,N_710);
xnor U2621 (N_2621,N_155,N_1260);
xnor U2622 (N_2622,N_1372,N_601);
xnor U2623 (N_2623,N_728,N_1105);
nand U2624 (N_2624,N_109,N_1000);
or U2625 (N_2625,N_62,N_1149);
and U2626 (N_2626,N_1266,N_1120);
nor U2627 (N_2627,N_1083,N_844);
xor U2628 (N_2628,N_383,N_1283);
xnor U2629 (N_2629,N_795,N_931);
and U2630 (N_2630,N_1951,N_210);
xnor U2631 (N_2631,N_1757,N_514);
and U2632 (N_2632,N_691,N_1575);
nand U2633 (N_2633,N_1743,N_544);
xnor U2634 (N_2634,N_1833,N_1051);
and U2635 (N_2635,N_556,N_1157);
nor U2636 (N_2636,N_1360,N_1740);
and U2637 (N_2637,N_1299,N_975);
or U2638 (N_2638,N_1306,N_423);
nand U2639 (N_2639,N_1998,N_1772);
nand U2640 (N_2640,N_607,N_714);
or U2641 (N_2641,N_552,N_793);
xnor U2642 (N_2642,N_920,N_1966);
nor U2643 (N_2643,N_1301,N_449);
or U2644 (N_2644,N_1182,N_603);
nor U2645 (N_2645,N_903,N_540);
nor U2646 (N_2646,N_345,N_1637);
xor U2647 (N_2647,N_1128,N_1660);
and U2648 (N_2648,N_1437,N_1342);
or U2649 (N_2649,N_693,N_1677);
nand U2650 (N_2650,N_370,N_178);
xor U2651 (N_2651,N_897,N_628);
xor U2652 (N_2652,N_293,N_260);
nor U2653 (N_2653,N_1558,N_1275);
xnor U2654 (N_2654,N_488,N_1963);
nor U2655 (N_2655,N_1783,N_1928);
or U2656 (N_2656,N_1916,N_436);
nand U2657 (N_2657,N_181,N_180);
nor U2658 (N_2658,N_223,N_1547);
and U2659 (N_2659,N_1922,N_865);
or U2660 (N_2660,N_566,N_1013);
or U2661 (N_2661,N_1945,N_1496);
nor U2662 (N_2662,N_901,N_149);
nand U2663 (N_2663,N_1311,N_1164);
nand U2664 (N_2664,N_1644,N_1268);
nor U2665 (N_2665,N_1162,N_1781);
and U2666 (N_2666,N_1617,N_1068);
and U2667 (N_2667,N_1200,N_581);
or U2668 (N_2668,N_326,N_1541);
and U2669 (N_2669,N_1094,N_1806);
or U2670 (N_2670,N_229,N_854);
or U2671 (N_2671,N_679,N_1161);
nor U2672 (N_2672,N_1599,N_1861);
and U2673 (N_2673,N_1980,N_245);
nand U2674 (N_2674,N_198,N_541);
nand U2675 (N_2675,N_1223,N_1733);
nand U2676 (N_2676,N_1209,N_334);
and U2677 (N_2677,N_1065,N_923);
xor U2678 (N_2678,N_1533,N_444);
nand U2679 (N_2679,N_1219,N_1389);
xnor U2680 (N_2680,N_969,N_816);
or U2681 (N_2681,N_1727,N_292);
and U2682 (N_2682,N_619,N_831);
nor U2683 (N_2683,N_577,N_305);
nor U2684 (N_2684,N_1917,N_1758);
or U2685 (N_2685,N_381,N_28);
and U2686 (N_2686,N_1707,N_122);
xor U2687 (N_2687,N_1580,N_1545);
or U2688 (N_2688,N_1394,N_388);
nor U2689 (N_2689,N_1462,N_1745);
xor U2690 (N_2690,N_490,N_369);
nor U2691 (N_2691,N_1824,N_1732);
nor U2692 (N_2692,N_801,N_1579);
xnor U2693 (N_2693,N_1486,N_887);
nor U2694 (N_2694,N_1202,N_466);
nand U2695 (N_2695,N_1226,N_1565);
and U2696 (N_2696,N_1419,N_718);
and U2697 (N_2697,N_1729,N_877);
and U2698 (N_2698,N_1456,N_1898);
nor U2699 (N_2699,N_2,N_1160);
nor U2700 (N_2700,N_164,N_1576);
xor U2701 (N_2701,N_1119,N_1551);
xnor U2702 (N_2702,N_798,N_599);
nor U2703 (N_2703,N_846,N_953);
and U2704 (N_2704,N_208,N_730);
nor U2705 (N_2705,N_1766,N_768);
nand U2706 (N_2706,N_192,N_945);
and U2707 (N_2707,N_179,N_338);
nand U2708 (N_2708,N_575,N_307);
and U2709 (N_2709,N_512,N_976);
xor U2710 (N_2710,N_1780,N_105);
xor U2711 (N_2711,N_408,N_425);
nor U2712 (N_2712,N_652,N_870);
nand U2713 (N_2713,N_215,N_1244);
nor U2714 (N_2714,N_140,N_280);
and U2715 (N_2715,N_218,N_695);
and U2716 (N_2716,N_1525,N_309);
nor U2717 (N_2717,N_1701,N_760);
xnor U2718 (N_2718,N_1411,N_238);
nor U2719 (N_2719,N_509,N_1001);
nand U2720 (N_2720,N_610,N_1844);
xor U2721 (N_2721,N_1295,N_1336);
nor U2722 (N_2722,N_1189,N_1597);
and U2723 (N_2723,N_764,N_621);
nand U2724 (N_2724,N_1021,N_623);
nand U2725 (N_2725,N_914,N_193);
and U2726 (N_2726,N_1578,N_1099);
nand U2727 (N_2727,N_565,N_234);
nor U2728 (N_2728,N_1823,N_1435);
or U2729 (N_2729,N_1948,N_867);
xor U2730 (N_2730,N_1990,N_582);
or U2731 (N_2731,N_302,N_847);
and U2732 (N_2732,N_526,N_719);
nand U2733 (N_2733,N_9,N_648);
and U2734 (N_2734,N_186,N_1190);
nor U2735 (N_2735,N_89,N_651);
nor U2736 (N_2736,N_251,N_980);
and U2737 (N_2737,N_1909,N_995);
or U2738 (N_2738,N_860,N_289);
xnor U2739 (N_2739,N_1253,N_758);
and U2740 (N_2740,N_304,N_259);
or U2741 (N_2741,N_624,N_516);
or U2742 (N_2742,N_404,N_286);
and U2743 (N_2743,N_1042,N_1326);
or U2744 (N_2744,N_258,N_1296);
and U2745 (N_2745,N_1069,N_255);
and U2746 (N_2746,N_1880,N_221);
and U2747 (N_2747,N_1754,N_1029);
and U2748 (N_2748,N_539,N_427);
nor U2749 (N_2749,N_1592,N_253);
or U2750 (N_2750,N_1191,N_445);
nor U2751 (N_2751,N_1033,N_1940);
nor U2752 (N_2752,N_1274,N_649);
xor U2753 (N_2753,N_617,N_1323);
and U2754 (N_2754,N_1608,N_915);
and U2755 (N_2755,N_1600,N_1507);
and U2756 (N_2756,N_1913,N_1363);
and U2757 (N_2757,N_727,N_38);
or U2758 (N_2758,N_148,N_1791);
and U2759 (N_2759,N_967,N_521);
and U2760 (N_2760,N_895,N_446);
or U2761 (N_2761,N_1383,N_393);
xnor U2762 (N_2762,N_1517,N_174);
nor U2763 (N_2763,N_261,N_1830);
or U2764 (N_2764,N_1145,N_34);
nor U2765 (N_2765,N_358,N_892);
nor U2766 (N_2766,N_1947,N_1176);
xor U2767 (N_2767,N_554,N_14);
nor U2768 (N_2768,N_125,N_269);
or U2769 (N_2769,N_1676,N_1124);
xor U2770 (N_2770,N_1577,N_588);
and U2771 (N_2771,N_1515,N_279);
xnor U2772 (N_2772,N_919,N_1092);
and U2773 (N_2773,N_1019,N_112);
nand U2774 (N_2774,N_1423,N_776);
xor U2775 (N_2775,N_1764,N_1181);
or U2776 (N_2776,N_1539,N_1927);
xor U2777 (N_2777,N_288,N_625);
or U2778 (N_2778,N_534,N_585);
nor U2779 (N_2779,N_759,N_262);
or U2780 (N_2780,N_389,N_1559);
or U2781 (N_2781,N_763,N_1302);
or U2782 (N_2782,N_244,N_1624);
nor U2783 (N_2783,N_1373,N_767);
nor U2784 (N_2784,N_660,N_1573);
nand U2785 (N_2785,N_1291,N_1896);
or U2786 (N_2786,N_1390,N_74);
xor U2787 (N_2787,N_941,N_1337);
nor U2788 (N_2788,N_1117,N_1465);
and U2789 (N_2789,N_1355,N_1284);
or U2790 (N_2790,N_1997,N_1498);
nor U2791 (N_2791,N_224,N_1518);
and U2792 (N_2792,N_1653,N_1115);
and U2793 (N_2793,N_1163,N_1487);
or U2794 (N_2794,N_1473,N_546);
nor U2795 (N_2795,N_136,N_676);
nor U2796 (N_2796,N_1636,N_991);
or U2797 (N_2797,N_1352,N_426);
and U2798 (N_2798,N_1396,N_1786);
nor U2799 (N_2799,N_775,N_141);
xnor U2800 (N_2800,N_194,N_713);
xor U2801 (N_2801,N_732,N_1695);
nor U2802 (N_2802,N_1501,N_1440);
nor U2803 (N_2803,N_1425,N_1252);
and U2804 (N_2804,N_1645,N_73);
nor U2805 (N_2805,N_821,N_943);
nor U2806 (N_2806,N_339,N_639);
nand U2807 (N_2807,N_1819,N_360);
and U2808 (N_2808,N_841,N_949);
nor U2809 (N_2809,N_1142,N_656);
xor U2810 (N_2810,N_1426,N_1349);
xor U2811 (N_2811,N_1789,N_1799);
or U2812 (N_2812,N_367,N_850);
and U2813 (N_2813,N_1747,N_1970);
and U2814 (N_2814,N_257,N_1384);
nor U2815 (N_2815,N_688,N_201);
xnor U2816 (N_2816,N_1448,N_397);
and U2817 (N_2817,N_364,N_909);
or U2818 (N_2818,N_525,N_756);
nor U2819 (N_2819,N_673,N_1692);
or U2820 (N_2820,N_1134,N_1267);
nand U2821 (N_2821,N_559,N_18);
xnor U2822 (N_2822,N_635,N_1156);
xor U2823 (N_2823,N_1942,N_36);
or U2824 (N_2824,N_42,N_1836);
or U2825 (N_2825,N_654,N_222);
and U2826 (N_2826,N_1690,N_1491);
or U2827 (N_2827,N_1923,N_618);
and U2828 (N_2828,N_1598,N_24);
nand U2829 (N_2829,N_1552,N_722);
or U2830 (N_2830,N_47,N_1139);
nor U2831 (N_2831,N_697,N_1061);
nor U2832 (N_2832,N_1224,N_1453);
nand U2833 (N_2833,N_137,N_1795);
xor U2834 (N_2834,N_1262,N_1536);
or U2835 (N_2835,N_1304,N_595);
nor U2836 (N_2836,N_276,N_1314);
and U2837 (N_2837,N_1528,N_1112);
and U2838 (N_2838,N_1077,N_99);
nand U2839 (N_2839,N_48,N_1520);
xnor U2840 (N_2840,N_1450,N_1555);
and U2841 (N_2841,N_1421,N_1874);
nor U2842 (N_2842,N_1850,N_1605);
and U2843 (N_2843,N_938,N_1897);
or U2844 (N_2844,N_1060,N_1086);
xor U2845 (N_2845,N_1894,N_1366);
nor U2846 (N_2846,N_310,N_1530);
xor U2847 (N_2847,N_283,N_1885);
nor U2848 (N_2848,N_664,N_896);
nor U2849 (N_2849,N_510,N_1869);
nor U2850 (N_2850,N_1214,N_1687);
and U2851 (N_2851,N_378,N_1893);
and U2852 (N_2852,N_1588,N_1403);
nand U2853 (N_2853,N_1838,N_1316);
and U2854 (N_2854,N_435,N_830);
nand U2855 (N_2855,N_1714,N_966);
and U2856 (N_2856,N_1375,N_606);
nand U2857 (N_2857,N_477,N_1638);
nand U2858 (N_2858,N_1738,N_239);
nor U2859 (N_2859,N_1138,N_1813);
and U2860 (N_2860,N_751,N_1044);
and U2861 (N_2861,N_543,N_1240);
nor U2862 (N_2862,N_1805,N_183);
xnor U2863 (N_2863,N_1408,N_1391);
nand U2864 (N_2864,N_862,N_1006);
xnor U2865 (N_2865,N_217,N_398);
and U2866 (N_2866,N_371,N_1681);
or U2867 (N_2867,N_1778,N_1449);
nor U2868 (N_2868,N_918,N_1673);
or U2869 (N_2869,N_265,N_93);
nand U2870 (N_2870,N_1987,N_1364);
nor U2871 (N_2871,N_1513,N_1961);
nor U2872 (N_2872,N_1771,N_573);
nor U2873 (N_2873,N_1839,N_1358);
and U2874 (N_2874,N_1022,N_1871);
xnor U2875 (N_2875,N_340,N_41);
nor U2876 (N_2876,N_663,N_1904);
xnor U2877 (N_2877,N_442,N_1166);
and U2878 (N_2878,N_524,N_828);
nor U2879 (N_2879,N_720,N_562);
or U2880 (N_2880,N_866,N_1840);
or U2881 (N_2881,N_797,N_457);
xnor U2882 (N_2882,N_317,N_22);
and U2883 (N_2883,N_418,N_83);
nor U2884 (N_2884,N_1427,N_550);
nor U2885 (N_2885,N_708,N_1529);
xor U2886 (N_2886,N_1231,N_1785);
or U2887 (N_2887,N_1914,N_1175);
nand U2888 (N_2888,N_1034,N_129);
xnor U2889 (N_2889,N_458,N_1975);
xor U2890 (N_2890,N_295,N_212);
or U2891 (N_2891,N_1593,N_1623);
or U2892 (N_2892,N_175,N_1087);
or U2893 (N_2893,N_1485,N_1113);
nor U2894 (N_2894,N_885,N_1761);
nand U2895 (N_2895,N_1878,N_1832);
and U2896 (N_2896,N_753,N_1514);
or U2897 (N_2897,N_1811,N_1828);
xor U2898 (N_2898,N_511,N_1024);
xnor U2899 (N_2899,N_701,N_613);
or U2900 (N_2900,N_1351,N_1378);
nor U2901 (N_2901,N_55,N_272);
or U2902 (N_2902,N_1711,N_1432);
nor U2903 (N_2903,N_563,N_1691);
xor U2904 (N_2904,N_564,N_1996);
or U2905 (N_2905,N_746,N_1321);
nand U2906 (N_2906,N_1125,N_134);
nor U2907 (N_2907,N_1279,N_1724);
nand U2908 (N_2908,N_57,N_1320);
nand U2909 (N_2909,N_100,N_747);
xor U2910 (N_2910,N_29,N_1907);
nor U2911 (N_2911,N_1329,N_7);
and U2912 (N_2912,N_1388,N_37);
and U2913 (N_2913,N_4,N_712);
or U2914 (N_2914,N_1155,N_1950);
and U2915 (N_2915,N_633,N_1055);
nand U2916 (N_2916,N_117,N_1834);
or U2917 (N_2917,N_1881,N_687);
and U2918 (N_2918,N_1931,N_677);
nand U2919 (N_2919,N_1935,N_1981);
nand U2920 (N_2920,N_879,N_1193);
nor U2921 (N_2921,N_899,N_84);
nor U2922 (N_2922,N_11,N_359);
nand U2923 (N_2923,N_1699,N_1217);
nand U2924 (N_2924,N_858,N_120);
nor U2925 (N_2925,N_294,N_787);
and U2926 (N_2926,N_146,N_597);
and U2927 (N_2927,N_1054,N_236);
nand U2928 (N_2928,N_1045,N_884);
and U2929 (N_2929,N_954,N_350);
and U2930 (N_2930,N_98,N_528);
nand U2931 (N_2931,N_1255,N_583);
nand U2932 (N_2932,N_778,N_1870);
nor U2933 (N_2933,N_1480,N_592);
nor U2934 (N_2934,N_551,N_1521);
nor U2935 (N_2935,N_1647,N_872);
nand U2936 (N_2936,N_1770,N_694);
or U2937 (N_2937,N_547,N_1686);
nand U2938 (N_2938,N_1235,N_557);
or U2939 (N_2939,N_752,N_342);
or U2940 (N_2940,N_612,N_441);
and U2941 (N_2941,N_1679,N_205);
nor U2942 (N_2942,N_1550,N_1890);
xnor U2943 (N_2943,N_935,N_1995);
nand U2944 (N_2944,N_1108,N_1334);
nor U2945 (N_2945,N_785,N_936);
nand U2946 (N_2946,N_779,N_1201);
or U2947 (N_2947,N_298,N_1632);
or U2948 (N_2948,N_761,N_822);
or U2949 (N_2949,N_815,N_1205);
nor U2950 (N_2950,N_1035,N_1814);
nor U2951 (N_2951,N_12,N_115);
xor U2952 (N_2952,N_1038,N_1004);
xnor U2953 (N_2953,N_1011,N_724);
and U2954 (N_2954,N_72,N_1076);
or U2955 (N_2955,N_271,N_1317);
and U2956 (N_2956,N_61,N_463);
or U2957 (N_2957,N_1377,N_1368);
nor U2958 (N_2958,N_950,N_1919);
or U2959 (N_2959,N_536,N_972);
or U2960 (N_2960,N_395,N_910);
and U2961 (N_2961,N_482,N_1516);
nor U2962 (N_2962,N_429,N_1424);
or U2963 (N_2963,N_1049,N_978);
xor U2964 (N_2964,N_415,N_333);
or U2965 (N_2965,N_504,N_172);
and U2966 (N_2966,N_483,N_357);
and U2967 (N_2967,N_571,N_908);
and U2968 (N_2968,N_1622,N_139);
and U2969 (N_2969,N_1263,N_1875);
nand U2970 (N_2970,N_1107,N_1879);
nor U2971 (N_2971,N_542,N_928);
and U2972 (N_2972,N_1476,N_1748);
and U2973 (N_2973,N_1884,N_507);
nand U2974 (N_2974,N_782,N_496);
or U2975 (N_2975,N_735,N_145);
nand U2976 (N_2976,N_1123,N_1643);
nand U2977 (N_2977,N_377,N_1009);
xor U2978 (N_2978,N_851,N_53);
xor U2979 (N_2979,N_21,N_1003);
nand U2980 (N_2980,N_1406,N_385);
xor U2981 (N_2981,N_91,N_6);
nand U2982 (N_2982,N_965,N_1538);
or U2983 (N_2983,N_1993,N_216);
and U2984 (N_2984,N_868,N_580);
or U2985 (N_2985,N_670,N_1357);
nor U2986 (N_2986,N_1039,N_1807);
or U2987 (N_2987,N_110,N_1438);
or U2988 (N_2988,N_1892,N_1619);
nor U2989 (N_2989,N_1616,N_1460);
nor U2990 (N_2990,N_1218,N_1953);
nand U2991 (N_2991,N_485,N_254);
nor U2992 (N_2992,N_522,N_1085);
nand U2993 (N_2993,N_590,N_1481);
xor U2994 (N_2994,N_1532,N_1716);
or U2995 (N_2995,N_1032,N_1759);
nor U2996 (N_2996,N_1655,N_786);
nor U2997 (N_2997,N_1710,N_1282);
xnor U2998 (N_2998,N_1630,N_264);
xnor U2999 (N_2999,N_1523,N_351);
or U3000 (N_3000,N_593,N_1441);
or U3001 (N_3001,N_1668,N_1043);
or U3002 (N_3002,N_144,N_1617);
nand U3003 (N_3003,N_1360,N_665);
and U3004 (N_3004,N_1605,N_8);
or U3005 (N_3005,N_464,N_520);
nand U3006 (N_3006,N_1692,N_1622);
xnor U3007 (N_3007,N_1123,N_1010);
xnor U3008 (N_3008,N_1123,N_730);
and U3009 (N_3009,N_231,N_840);
or U3010 (N_3010,N_876,N_1690);
xnor U3011 (N_3011,N_1737,N_117);
or U3012 (N_3012,N_1595,N_1035);
xnor U3013 (N_3013,N_686,N_1751);
nand U3014 (N_3014,N_1763,N_610);
and U3015 (N_3015,N_916,N_200);
xnor U3016 (N_3016,N_1146,N_1625);
nor U3017 (N_3017,N_764,N_724);
and U3018 (N_3018,N_166,N_738);
nor U3019 (N_3019,N_1876,N_154);
nand U3020 (N_3020,N_454,N_305);
or U3021 (N_3021,N_660,N_964);
xnor U3022 (N_3022,N_1619,N_656);
and U3023 (N_3023,N_1262,N_1417);
nand U3024 (N_3024,N_1192,N_1567);
nor U3025 (N_3025,N_170,N_1395);
xor U3026 (N_3026,N_1,N_1794);
nor U3027 (N_3027,N_833,N_1495);
and U3028 (N_3028,N_489,N_1988);
and U3029 (N_3029,N_891,N_1104);
and U3030 (N_3030,N_322,N_1089);
xnor U3031 (N_3031,N_1548,N_1521);
nor U3032 (N_3032,N_69,N_1426);
or U3033 (N_3033,N_1366,N_1510);
or U3034 (N_3034,N_703,N_584);
nor U3035 (N_3035,N_1586,N_815);
or U3036 (N_3036,N_1772,N_101);
nor U3037 (N_3037,N_437,N_630);
nand U3038 (N_3038,N_1761,N_69);
or U3039 (N_3039,N_81,N_1924);
or U3040 (N_3040,N_1678,N_918);
and U3041 (N_3041,N_1222,N_1697);
nor U3042 (N_3042,N_1055,N_303);
and U3043 (N_3043,N_1060,N_300);
or U3044 (N_3044,N_249,N_370);
nor U3045 (N_3045,N_1875,N_354);
and U3046 (N_3046,N_878,N_1665);
and U3047 (N_3047,N_1092,N_1551);
nor U3048 (N_3048,N_896,N_1774);
nor U3049 (N_3049,N_1545,N_457);
or U3050 (N_3050,N_511,N_1185);
xor U3051 (N_3051,N_1064,N_362);
or U3052 (N_3052,N_7,N_339);
nor U3053 (N_3053,N_1527,N_1447);
xor U3054 (N_3054,N_1878,N_260);
xor U3055 (N_3055,N_836,N_1837);
or U3056 (N_3056,N_1609,N_398);
or U3057 (N_3057,N_217,N_662);
xnor U3058 (N_3058,N_1663,N_1005);
nand U3059 (N_3059,N_1172,N_799);
xnor U3060 (N_3060,N_1958,N_1325);
nor U3061 (N_3061,N_417,N_352);
xor U3062 (N_3062,N_967,N_1421);
and U3063 (N_3063,N_124,N_87);
and U3064 (N_3064,N_459,N_1796);
nor U3065 (N_3065,N_625,N_652);
nand U3066 (N_3066,N_953,N_1687);
nor U3067 (N_3067,N_1887,N_710);
or U3068 (N_3068,N_1184,N_288);
and U3069 (N_3069,N_1674,N_411);
and U3070 (N_3070,N_1522,N_302);
nand U3071 (N_3071,N_1630,N_750);
or U3072 (N_3072,N_1384,N_165);
and U3073 (N_3073,N_775,N_1571);
nand U3074 (N_3074,N_1840,N_1868);
nand U3075 (N_3075,N_1269,N_1437);
and U3076 (N_3076,N_1614,N_37);
nand U3077 (N_3077,N_679,N_1564);
xnor U3078 (N_3078,N_1726,N_1121);
and U3079 (N_3079,N_1551,N_1383);
and U3080 (N_3080,N_1936,N_82);
nand U3081 (N_3081,N_234,N_416);
nand U3082 (N_3082,N_1646,N_503);
xnor U3083 (N_3083,N_1696,N_312);
nand U3084 (N_3084,N_437,N_944);
nand U3085 (N_3085,N_137,N_1442);
or U3086 (N_3086,N_1676,N_1176);
and U3087 (N_3087,N_1795,N_1315);
or U3088 (N_3088,N_1529,N_964);
or U3089 (N_3089,N_549,N_604);
and U3090 (N_3090,N_839,N_114);
xnor U3091 (N_3091,N_1776,N_764);
and U3092 (N_3092,N_218,N_1688);
xnor U3093 (N_3093,N_1802,N_1481);
or U3094 (N_3094,N_1450,N_366);
xor U3095 (N_3095,N_926,N_868);
nor U3096 (N_3096,N_1293,N_604);
nand U3097 (N_3097,N_1041,N_830);
or U3098 (N_3098,N_1486,N_763);
nor U3099 (N_3099,N_977,N_1828);
nor U3100 (N_3100,N_1990,N_1227);
nand U3101 (N_3101,N_1038,N_1335);
xor U3102 (N_3102,N_1338,N_285);
or U3103 (N_3103,N_682,N_940);
or U3104 (N_3104,N_1173,N_588);
or U3105 (N_3105,N_802,N_1908);
and U3106 (N_3106,N_912,N_750);
nor U3107 (N_3107,N_1963,N_543);
nand U3108 (N_3108,N_1242,N_484);
or U3109 (N_3109,N_480,N_536);
xnor U3110 (N_3110,N_1518,N_1478);
nand U3111 (N_3111,N_292,N_605);
xor U3112 (N_3112,N_246,N_1614);
and U3113 (N_3113,N_950,N_1382);
nor U3114 (N_3114,N_161,N_1558);
and U3115 (N_3115,N_1811,N_1979);
nor U3116 (N_3116,N_1374,N_1213);
nand U3117 (N_3117,N_244,N_1530);
nand U3118 (N_3118,N_883,N_1505);
nand U3119 (N_3119,N_1451,N_1245);
and U3120 (N_3120,N_1394,N_266);
or U3121 (N_3121,N_1497,N_1685);
nor U3122 (N_3122,N_157,N_497);
and U3123 (N_3123,N_897,N_919);
and U3124 (N_3124,N_61,N_600);
or U3125 (N_3125,N_1420,N_1525);
nand U3126 (N_3126,N_1910,N_1781);
xnor U3127 (N_3127,N_1566,N_89);
or U3128 (N_3128,N_503,N_709);
and U3129 (N_3129,N_685,N_1970);
nor U3130 (N_3130,N_238,N_388);
nand U3131 (N_3131,N_616,N_623);
nand U3132 (N_3132,N_1582,N_818);
xnor U3133 (N_3133,N_378,N_1529);
nor U3134 (N_3134,N_398,N_450);
nand U3135 (N_3135,N_509,N_1266);
and U3136 (N_3136,N_1440,N_1438);
or U3137 (N_3137,N_1285,N_1614);
and U3138 (N_3138,N_1634,N_246);
nand U3139 (N_3139,N_424,N_604);
or U3140 (N_3140,N_870,N_1676);
xnor U3141 (N_3141,N_833,N_1549);
nor U3142 (N_3142,N_1642,N_1190);
or U3143 (N_3143,N_1790,N_1921);
or U3144 (N_3144,N_1159,N_1800);
nor U3145 (N_3145,N_632,N_1702);
and U3146 (N_3146,N_230,N_496);
nand U3147 (N_3147,N_422,N_234);
nor U3148 (N_3148,N_1066,N_578);
nor U3149 (N_3149,N_1987,N_1446);
nor U3150 (N_3150,N_1282,N_12);
xnor U3151 (N_3151,N_43,N_435);
nor U3152 (N_3152,N_891,N_1034);
and U3153 (N_3153,N_1119,N_68);
or U3154 (N_3154,N_1328,N_1837);
and U3155 (N_3155,N_1552,N_1104);
or U3156 (N_3156,N_78,N_1540);
nor U3157 (N_3157,N_548,N_296);
xor U3158 (N_3158,N_908,N_766);
and U3159 (N_3159,N_760,N_1650);
nand U3160 (N_3160,N_1020,N_1294);
nand U3161 (N_3161,N_475,N_1750);
nand U3162 (N_3162,N_1335,N_425);
nand U3163 (N_3163,N_904,N_278);
or U3164 (N_3164,N_1455,N_1833);
and U3165 (N_3165,N_1304,N_201);
and U3166 (N_3166,N_1749,N_660);
or U3167 (N_3167,N_460,N_211);
nor U3168 (N_3168,N_987,N_847);
nand U3169 (N_3169,N_1421,N_641);
and U3170 (N_3170,N_653,N_1880);
nand U3171 (N_3171,N_1142,N_1184);
or U3172 (N_3172,N_895,N_47);
or U3173 (N_3173,N_1331,N_1189);
or U3174 (N_3174,N_1957,N_419);
nand U3175 (N_3175,N_1648,N_1392);
and U3176 (N_3176,N_1840,N_800);
nor U3177 (N_3177,N_977,N_1824);
and U3178 (N_3178,N_530,N_1239);
nor U3179 (N_3179,N_196,N_1896);
nor U3180 (N_3180,N_1993,N_1598);
nand U3181 (N_3181,N_843,N_589);
nand U3182 (N_3182,N_389,N_1281);
nand U3183 (N_3183,N_218,N_572);
xor U3184 (N_3184,N_354,N_766);
xnor U3185 (N_3185,N_341,N_392);
and U3186 (N_3186,N_681,N_198);
and U3187 (N_3187,N_1592,N_1525);
nor U3188 (N_3188,N_1420,N_745);
nor U3189 (N_3189,N_1130,N_1151);
or U3190 (N_3190,N_1493,N_701);
nand U3191 (N_3191,N_1973,N_1126);
or U3192 (N_3192,N_1244,N_39);
and U3193 (N_3193,N_621,N_799);
nand U3194 (N_3194,N_455,N_507);
or U3195 (N_3195,N_450,N_768);
and U3196 (N_3196,N_957,N_1609);
or U3197 (N_3197,N_601,N_1255);
and U3198 (N_3198,N_532,N_1228);
and U3199 (N_3199,N_1578,N_279);
nand U3200 (N_3200,N_674,N_40);
xnor U3201 (N_3201,N_1547,N_1945);
and U3202 (N_3202,N_1499,N_436);
xnor U3203 (N_3203,N_985,N_1100);
or U3204 (N_3204,N_549,N_5);
and U3205 (N_3205,N_1278,N_1219);
or U3206 (N_3206,N_1092,N_1456);
and U3207 (N_3207,N_824,N_952);
and U3208 (N_3208,N_818,N_1061);
and U3209 (N_3209,N_1224,N_1084);
and U3210 (N_3210,N_771,N_1519);
xor U3211 (N_3211,N_703,N_913);
or U3212 (N_3212,N_1350,N_319);
or U3213 (N_3213,N_1188,N_1986);
or U3214 (N_3214,N_1712,N_744);
or U3215 (N_3215,N_1632,N_1676);
nand U3216 (N_3216,N_1067,N_226);
xor U3217 (N_3217,N_238,N_1501);
xor U3218 (N_3218,N_1386,N_179);
xor U3219 (N_3219,N_932,N_708);
nand U3220 (N_3220,N_1596,N_411);
nand U3221 (N_3221,N_1054,N_1416);
xor U3222 (N_3222,N_1352,N_555);
xnor U3223 (N_3223,N_185,N_319);
and U3224 (N_3224,N_875,N_1768);
and U3225 (N_3225,N_902,N_987);
nor U3226 (N_3226,N_284,N_422);
xor U3227 (N_3227,N_635,N_1722);
or U3228 (N_3228,N_1884,N_1545);
and U3229 (N_3229,N_1108,N_1222);
and U3230 (N_3230,N_1596,N_1515);
nand U3231 (N_3231,N_928,N_1812);
or U3232 (N_3232,N_1729,N_1394);
nand U3233 (N_3233,N_1221,N_461);
nor U3234 (N_3234,N_127,N_1668);
or U3235 (N_3235,N_675,N_603);
nor U3236 (N_3236,N_454,N_826);
nand U3237 (N_3237,N_942,N_1566);
and U3238 (N_3238,N_767,N_955);
xor U3239 (N_3239,N_1284,N_1739);
nor U3240 (N_3240,N_786,N_1545);
or U3241 (N_3241,N_1209,N_279);
or U3242 (N_3242,N_1438,N_1090);
xor U3243 (N_3243,N_1132,N_928);
nand U3244 (N_3244,N_1290,N_1492);
and U3245 (N_3245,N_608,N_1302);
or U3246 (N_3246,N_1698,N_694);
nor U3247 (N_3247,N_794,N_546);
xnor U3248 (N_3248,N_1533,N_104);
xor U3249 (N_3249,N_1852,N_71);
nand U3250 (N_3250,N_1461,N_1169);
xnor U3251 (N_3251,N_744,N_901);
nor U3252 (N_3252,N_1575,N_1930);
and U3253 (N_3253,N_1136,N_90);
nor U3254 (N_3254,N_1289,N_833);
or U3255 (N_3255,N_1711,N_314);
xor U3256 (N_3256,N_78,N_874);
nand U3257 (N_3257,N_435,N_805);
nor U3258 (N_3258,N_1485,N_947);
nor U3259 (N_3259,N_1189,N_1822);
nor U3260 (N_3260,N_1170,N_558);
or U3261 (N_3261,N_854,N_96);
or U3262 (N_3262,N_77,N_1016);
xnor U3263 (N_3263,N_1101,N_1655);
nor U3264 (N_3264,N_278,N_1213);
xor U3265 (N_3265,N_782,N_130);
xor U3266 (N_3266,N_287,N_830);
nor U3267 (N_3267,N_1570,N_1322);
or U3268 (N_3268,N_86,N_526);
xnor U3269 (N_3269,N_1450,N_1914);
nor U3270 (N_3270,N_1771,N_1346);
or U3271 (N_3271,N_666,N_502);
or U3272 (N_3272,N_1065,N_341);
nand U3273 (N_3273,N_1420,N_1806);
xor U3274 (N_3274,N_305,N_1856);
nand U3275 (N_3275,N_474,N_364);
nor U3276 (N_3276,N_232,N_443);
and U3277 (N_3277,N_1186,N_1338);
or U3278 (N_3278,N_1652,N_1093);
and U3279 (N_3279,N_587,N_338);
and U3280 (N_3280,N_335,N_1740);
or U3281 (N_3281,N_828,N_1238);
nor U3282 (N_3282,N_525,N_1653);
nor U3283 (N_3283,N_208,N_695);
nand U3284 (N_3284,N_776,N_160);
and U3285 (N_3285,N_1175,N_1164);
or U3286 (N_3286,N_281,N_1690);
or U3287 (N_3287,N_522,N_1540);
or U3288 (N_3288,N_1279,N_888);
and U3289 (N_3289,N_376,N_1810);
and U3290 (N_3290,N_267,N_738);
and U3291 (N_3291,N_388,N_1074);
xor U3292 (N_3292,N_730,N_1607);
and U3293 (N_3293,N_115,N_520);
nor U3294 (N_3294,N_1769,N_1866);
xor U3295 (N_3295,N_647,N_1529);
or U3296 (N_3296,N_52,N_886);
nand U3297 (N_3297,N_853,N_1975);
nor U3298 (N_3298,N_1320,N_1135);
or U3299 (N_3299,N_1384,N_1979);
and U3300 (N_3300,N_469,N_1651);
or U3301 (N_3301,N_1580,N_1142);
and U3302 (N_3302,N_1269,N_1163);
nor U3303 (N_3303,N_835,N_1012);
xor U3304 (N_3304,N_1479,N_1443);
or U3305 (N_3305,N_864,N_1246);
xnor U3306 (N_3306,N_653,N_526);
nand U3307 (N_3307,N_772,N_1416);
nor U3308 (N_3308,N_1750,N_746);
and U3309 (N_3309,N_1395,N_492);
nand U3310 (N_3310,N_1316,N_105);
xor U3311 (N_3311,N_1675,N_784);
nor U3312 (N_3312,N_1703,N_990);
and U3313 (N_3313,N_1770,N_1190);
nor U3314 (N_3314,N_1587,N_1074);
and U3315 (N_3315,N_904,N_921);
and U3316 (N_3316,N_978,N_1205);
nor U3317 (N_3317,N_1741,N_1083);
xnor U3318 (N_3318,N_1815,N_393);
xor U3319 (N_3319,N_1072,N_69);
xnor U3320 (N_3320,N_1376,N_552);
and U3321 (N_3321,N_294,N_1159);
nor U3322 (N_3322,N_863,N_175);
and U3323 (N_3323,N_723,N_1558);
nand U3324 (N_3324,N_1141,N_893);
or U3325 (N_3325,N_1988,N_338);
nand U3326 (N_3326,N_443,N_615);
and U3327 (N_3327,N_1746,N_433);
xnor U3328 (N_3328,N_904,N_977);
nor U3329 (N_3329,N_1381,N_946);
nand U3330 (N_3330,N_1675,N_133);
xnor U3331 (N_3331,N_1976,N_1645);
nor U3332 (N_3332,N_1255,N_1394);
nor U3333 (N_3333,N_377,N_1839);
nand U3334 (N_3334,N_1415,N_1073);
or U3335 (N_3335,N_1489,N_297);
nand U3336 (N_3336,N_965,N_737);
xor U3337 (N_3337,N_1467,N_1611);
or U3338 (N_3338,N_904,N_774);
nor U3339 (N_3339,N_297,N_248);
xnor U3340 (N_3340,N_1149,N_561);
nor U3341 (N_3341,N_657,N_514);
nand U3342 (N_3342,N_839,N_573);
xor U3343 (N_3343,N_1958,N_1588);
and U3344 (N_3344,N_1884,N_308);
and U3345 (N_3345,N_0,N_210);
or U3346 (N_3346,N_1034,N_140);
nor U3347 (N_3347,N_1783,N_1914);
and U3348 (N_3348,N_47,N_1647);
nor U3349 (N_3349,N_333,N_1514);
xnor U3350 (N_3350,N_1526,N_1991);
and U3351 (N_3351,N_1821,N_1735);
and U3352 (N_3352,N_1374,N_1405);
nand U3353 (N_3353,N_1782,N_881);
xor U3354 (N_3354,N_1337,N_1658);
nor U3355 (N_3355,N_1707,N_1425);
and U3356 (N_3356,N_728,N_1311);
or U3357 (N_3357,N_1929,N_484);
nand U3358 (N_3358,N_298,N_1328);
nor U3359 (N_3359,N_1206,N_1840);
or U3360 (N_3360,N_1317,N_1219);
and U3361 (N_3361,N_1898,N_843);
nor U3362 (N_3362,N_1913,N_1791);
nand U3363 (N_3363,N_1757,N_1347);
xnor U3364 (N_3364,N_648,N_681);
nor U3365 (N_3365,N_262,N_596);
or U3366 (N_3366,N_1760,N_720);
and U3367 (N_3367,N_977,N_1898);
xor U3368 (N_3368,N_359,N_1580);
or U3369 (N_3369,N_1126,N_1216);
or U3370 (N_3370,N_866,N_1493);
xnor U3371 (N_3371,N_240,N_1718);
xnor U3372 (N_3372,N_175,N_663);
nand U3373 (N_3373,N_51,N_1936);
and U3374 (N_3374,N_1561,N_937);
or U3375 (N_3375,N_238,N_593);
xnor U3376 (N_3376,N_1847,N_1766);
nand U3377 (N_3377,N_1920,N_663);
nand U3378 (N_3378,N_1101,N_1370);
or U3379 (N_3379,N_944,N_1131);
xnor U3380 (N_3380,N_555,N_1715);
nand U3381 (N_3381,N_1308,N_858);
nor U3382 (N_3382,N_1977,N_173);
and U3383 (N_3383,N_1243,N_1063);
nand U3384 (N_3384,N_732,N_1275);
xor U3385 (N_3385,N_1523,N_948);
nor U3386 (N_3386,N_1971,N_887);
xnor U3387 (N_3387,N_1323,N_278);
and U3388 (N_3388,N_461,N_1175);
nand U3389 (N_3389,N_11,N_22);
nor U3390 (N_3390,N_674,N_1830);
and U3391 (N_3391,N_1116,N_698);
xnor U3392 (N_3392,N_760,N_1165);
or U3393 (N_3393,N_1103,N_666);
xor U3394 (N_3394,N_619,N_153);
xor U3395 (N_3395,N_418,N_1748);
or U3396 (N_3396,N_281,N_808);
or U3397 (N_3397,N_1661,N_1950);
xor U3398 (N_3398,N_376,N_316);
nor U3399 (N_3399,N_1817,N_339);
nand U3400 (N_3400,N_1592,N_1197);
and U3401 (N_3401,N_284,N_1872);
and U3402 (N_3402,N_236,N_683);
xnor U3403 (N_3403,N_1618,N_1552);
xnor U3404 (N_3404,N_1582,N_1622);
nand U3405 (N_3405,N_234,N_87);
xnor U3406 (N_3406,N_1946,N_681);
nand U3407 (N_3407,N_296,N_363);
nand U3408 (N_3408,N_1413,N_312);
or U3409 (N_3409,N_1865,N_1875);
nand U3410 (N_3410,N_1470,N_643);
nor U3411 (N_3411,N_1315,N_1614);
xor U3412 (N_3412,N_849,N_1102);
xor U3413 (N_3413,N_1462,N_79);
nor U3414 (N_3414,N_80,N_1513);
and U3415 (N_3415,N_902,N_1131);
nor U3416 (N_3416,N_140,N_867);
nand U3417 (N_3417,N_796,N_301);
or U3418 (N_3418,N_972,N_1703);
nor U3419 (N_3419,N_1107,N_773);
and U3420 (N_3420,N_638,N_307);
or U3421 (N_3421,N_1096,N_91);
or U3422 (N_3422,N_1442,N_22);
nor U3423 (N_3423,N_1304,N_199);
xnor U3424 (N_3424,N_1778,N_1680);
and U3425 (N_3425,N_879,N_763);
nand U3426 (N_3426,N_1107,N_1521);
nand U3427 (N_3427,N_1287,N_807);
nor U3428 (N_3428,N_892,N_91);
or U3429 (N_3429,N_78,N_1803);
nand U3430 (N_3430,N_1958,N_343);
and U3431 (N_3431,N_845,N_1810);
nor U3432 (N_3432,N_1027,N_1553);
and U3433 (N_3433,N_259,N_1592);
nor U3434 (N_3434,N_1475,N_198);
nand U3435 (N_3435,N_1912,N_417);
nor U3436 (N_3436,N_659,N_1126);
xor U3437 (N_3437,N_231,N_73);
xor U3438 (N_3438,N_515,N_1228);
nor U3439 (N_3439,N_25,N_351);
nor U3440 (N_3440,N_185,N_1332);
nand U3441 (N_3441,N_1236,N_687);
xnor U3442 (N_3442,N_1362,N_1199);
xnor U3443 (N_3443,N_791,N_1815);
nor U3444 (N_3444,N_1831,N_1726);
and U3445 (N_3445,N_1892,N_1368);
or U3446 (N_3446,N_766,N_101);
and U3447 (N_3447,N_767,N_1229);
nor U3448 (N_3448,N_1097,N_947);
xnor U3449 (N_3449,N_1183,N_1096);
xnor U3450 (N_3450,N_1366,N_440);
nor U3451 (N_3451,N_1583,N_1574);
nand U3452 (N_3452,N_1250,N_27);
nor U3453 (N_3453,N_1802,N_478);
nor U3454 (N_3454,N_609,N_561);
and U3455 (N_3455,N_1070,N_1310);
xor U3456 (N_3456,N_291,N_1158);
xnor U3457 (N_3457,N_1506,N_1373);
or U3458 (N_3458,N_114,N_1812);
nor U3459 (N_3459,N_1706,N_1888);
and U3460 (N_3460,N_1880,N_702);
and U3461 (N_3461,N_708,N_220);
nor U3462 (N_3462,N_841,N_1749);
and U3463 (N_3463,N_108,N_142);
and U3464 (N_3464,N_1489,N_1169);
and U3465 (N_3465,N_640,N_1535);
or U3466 (N_3466,N_1301,N_1118);
or U3467 (N_3467,N_295,N_624);
and U3468 (N_3468,N_1714,N_481);
xnor U3469 (N_3469,N_351,N_1913);
and U3470 (N_3470,N_359,N_404);
xor U3471 (N_3471,N_1225,N_555);
and U3472 (N_3472,N_279,N_1850);
nor U3473 (N_3473,N_1640,N_845);
and U3474 (N_3474,N_146,N_1361);
or U3475 (N_3475,N_274,N_426);
nand U3476 (N_3476,N_1266,N_934);
and U3477 (N_3477,N_1845,N_358);
and U3478 (N_3478,N_1836,N_821);
and U3479 (N_3479,N_1339,N_1794);
or U3480 (N_3480,N_234,N_1705);
nand U3481 (N_3481,N_1363,N_1896);
nor U3482 (N_3482,N_1939,N_1037);
or U3483 (N_3483,N_728,N_512);
xor U3484 (N_3484,N_730,N_639);
nand U3485 (N_3485,N_1950,N_1028);
and U3486 (N_3486,N_722,N_959);
nor U3487 (N_3487,N_1149,N_1390);
xnor U3488 (N_3488,N_750,N_858);
nand U3489 (N_3489,N_1910,N_1867);
and U3490 (N_3490,N_1341,N_1286);
nor U3491 (N_3491,N_255,N_763);
and U3492 (N_3492,N_819,N_1305);
nand U3493 (N_3493,N_367,N_349);
and U3494 (N_3494,N_1787,N_1167);
xor U3495 (N_3495,N_616,N_600);
or U3496 (N_3496,N_471,N_133);
or U3497 (N_3497,N_1672,N_1064);
nor U3498 (N_3498,N_411,N_1944);
nand U3499 (N_3499,N_1084,N_1565);
nor U3500 (N_3500,N_245,N_1821);
nor U3501 (N_3501,N_172,N_377);
nor U3502 (N_3502,N_1708,N_97);
nand U3503 (N_3503,N_1470,N_1731);
or U3504 (N_3504,N_1870,N_1684);
xor U3505 (N_3505,N_1132,N_911);
nand U3506 (N_3506,N_837,N_1850);
nand U3507 (N_3507,N_324,N_76);
or U3508 (N_3508,N_1436,N_875);
or U3509 (N_3509,N_1161,N_466);
xnor U3510 (N_3510,N_137,N_1684);
nand U3511 (N_3511,N_1522,N_820);
or U3512 (N_3512,N_1318,N_1200);
xnor U3513 (N_3513,N_1259,N_1441);
and U3514 (N_3514,N_512,N_912);
or U3515 (N_3515,N_1964,N_1229);
or U3516 (N_3516,N_1519,N_1374);
or U3517 (N_3517,N_1273,N_1098);
xnor U3518 (N_3518,N_1878,N_543);
or U3519 (N_3519,N_841,N_1791);
and U3520 (N_3520,N_367,N_29);
nor U3521 (N_3521,N_1718,N_78);
xor U3522 (N_3522,N_1558,N_1070);
nor U3523 (N_3523,N_876,N_1138);
nand U3524 (N_3524,N_1550,N_729);
nand U3525 (N_3525,N_997,N_831);
xor U3526 (N_3526,N_1888,N_222);
or U3527 (N_3527,N_20,N_85);
nor U3528 (N_3528,N_127,N_381);
or U3529 (N_3529,N_860,N_790);
and U3530 (N_3530,N_87,N_16);
or U3531 (N_3531,N_1900,N_1196);
or U3532 (N_3532,N_761,N_1017);
and U3533 (N_3533,N_1728,N_1175);
and U3534 (N_3534,N_1523,N_1802);
nor U3535 (N_3535,N_1203,N_815);
and U3536 (N_3536,N_1709,N_1162);
nand U3537 (N_3537,N_1410,N_1917);
xnor U3538 (N_3538,N_180,N_1291);
nor U3539 (N_3539,N_5,N_1343);
nor U3540 (N_3540,N_397,N_176);
and U3541 (N_3541,N_516,N_261);
and U3542 (N_3542,N_679,N_136);
xor U3543 (N_3543,N_1188,N_590);
nor U3544 (N_3544,N_1203,N_832);
nor U3545 (N_3545,N_736,N_250);
or U3546 (N_3546,N_1421,N_1572);
and U3547 (N_3547,N_1925,N_1570);
nor U3548 (N_3548,N_725,N_627);
nor U3549 (N_3549,N_536,N_1345);
and U3550 (N_3550,N_85,N_1753);
nand U3551 (N_3551,N_298,N_766);
and U3552 (N_3552,N_134,N_1842);
xnor U3553 (N_3553,N_1814,N_131);
or U3554 (N_3554,N_973,N_1026);
nor U3555 (N_3555,N_258,N_1070);
and U3556 (N_3556,N_1600,N_1731);
or U3557 (N_3557,N_56,N_5);
and U3558 (N_3558,N_1047,N_383);
or U3559 (N_3559,N_1272,N_376);
or U3560 (N_3560,N_549,N_992);
xnor U3561 (N_3561,N_1729,N_1903);
xnor U3562 (N_3562,N_999,N_559);
xor U3563 (N_3563,N_1672,N_128);
nand U3564 (N_3564,N_1987,N_727);
and U3565 (N_3565,N_1606,N_1621);
and U3566 (N_3566,N_1605,N_176);
nand U3567 (N_3567,N_722,N_1340);
and U3568 (N_3568,N_1793,N_1210);
nand U3569 (N_3569,N_349,N_1422);
and U3570 (N_3570,N_1512,N_760);
nand U3571 (N_3571,N_1371,N_207);
xnor U3572 (N_3572,N_1450,N_207);
nand U3573 (N_3573,N_1145,N_1466);
xnor U3574 (N_3574,N_1283,N_815);
nor U3575 (N_3575,N_176,N_1745);
nor U3576 (N_3576,N_23,N_1872);
nand U3577 (N_3577,N_1364,N_1687);
and U3578 (N_3578,N_475,N_866);
xor U3579 (N_3579,N_267,N_882);
and U3580 (N_3580,N_856,N_467);
nand U3581 (N_3581,N_1204,N_443);
and U3582 (N_3582,N_1965,N_69);
nand U3583 (N_3583,N_1574,N_391);
nor U3584 (N_3584,N_557,N_1937);
nor U3585 (N_3585,N_1192,N_117);
nor U3586 (N_3586,N_1314,N_401);
nor U3587 (N_3587,N_81,N_1931);
xnor U3588 (N_3588,N_1356,N_231);
nor U3589 (N_3589,N_57,N_39);
and U3590 (N_3590,N_322,N_879);
xor U3591 (N_3591,N_1210,N_1524);
or U3592 (N_3592,N_545,N_1735);
or U3593 (N_3593,N_1499,N_1182);
or U3594 (N_3594,N_1621,N_562);
and U3595 (N_3595,N_907,N_339);
xor U3596 (N_3596,N_1600,N_1550);
xor U3597 (N_3597,N_1617,N_129);
nand U3598 (N_3598,N_1609,N_1111);
xnor U3599 (N_3599,N_1492,N_452);
and U3600 (N_3600,N_419,N_1246);
nor U3601 (N_3601,N_1192,N_1437);
or U3602 (N_3602,N_895,N_1461);
nand U3603 (N_3603,N_1841,N_899);
nand U3604 (N_3604,N_1220,N_1932);
nor U3605 (N_3605,N_910,N_645);
nor U3606 (N_3606,N_218,N_1882);
or U3607 (N_3607,N_210,N_1109);
or U3608 (N_3608,N_420,N_1014);
and U3609 (N_3609,N_1424,N_877);
xnor U3610 (N_3610,N_1276,N_1008);
nand U3611 (N_3611,N_722,N_1840);
or U3612 (N_3612,N_367,N_985);
or U3613 (N_3613,N_227,N_1283);
nand U3614 (N_3614,N_577,N_427);
xnor U3615 (N_3615,N_630,N_21);
or U3616 (N_3616,N_1408,N_1467);
nor U3617 (N_3617,N_138,N_949);
xnor U3618 (N_3618,N_326,N_1629);
or U3619 (N_3619,N_1131,N_823);
nor U3620 (N_3620,N_1976,N_295);
nor U3621 (N_3621,N_1782,N_486);
nor U3622 (N_3622,N_1512,N_14);
and U3623 (N_3623,N_885,N_1007);
or U3624 (N_3624,N_499,N_1296);
xor U3625 (N_3625,N_1640,N_1817);
and U3626 (N_3626,N_1031,N_1336);
xnor U3627 (N_3627,N_972,N_1953);
nand U3628 (N_3628,N_1487,N_1492);
or U3629 (N_3629,N_1017,N_1594);
nand U3630 (N_3630,N_927,N_1499);
and U3631 (N_3631,N_1226,N_1866);
nand U3632 (N_3632,N_957,N_1285);
or U3633 (N_3633,N_1164,N_701);
nor U3634 (N_3634,N_650,N_176);
xor U3635 (N_3635,N_1126,N_1944);
or U3636 (N_3636,N_676,N_1023);
nor U3637 (N_3637,N_1970,N_1907);
nand U3638 (N_3638,N_812,N_1309);
nor U3639 (N_3639,N_1267,N_1337);
nand U3640 (N_3640,N_669,N_1520);
nand U3641 (N_3641,N_313,N_1695);
xor U3642 (N_3642,N_699,N_995);
nand U3643 (N_3643,N_1679,N_1575);
xnor U3644 (N_3644,N_1854,N_1752);
xnor U3645 (N_3645,N_27,N_1071);
xor U3646 (N_3646,N_1489,N_1563);
nand U3647 (N_3647,N_863,N_1095);
xnor U3648 (N_3648,N_1548,N_1780);
nand U3649 (N_3649,N_698,N_350);
xnor U3650 (N_3650,N_1081,N_296);
xnor U3651 (N_3651,N_137,N_536);
or U3652 (N_3652,N_1499,N_53);
xnor U3653 (N_3653,N_1969,N_288);
xor U3654 (N_3654,N_1591,N_1517);
and U3655 (N_3655,N_177,N_238);
nor U3656 (N_3656,N_1718,N_587);
or U3657 (N_3657,N_1394,N_1364);
nor U3658 (N_3658,N_1921,N_1275);
nor U3659 (N_3659,N_236,N_1083);
or U3660 (N_3660,N_249,N_1712);
or U3661 (N_3661,N_464,N_925);
xnor U3662 (N_3662,N_460,N_1706);
nor U3663 (N_3663,N_802,N_1213);
and U3664 (N_3664,N_891,N_518);
nor U3665 (N_3665,N_1876,N_1358);
xnor U3666 (N_3666,N_977,N_1713);
xnor U3667 (N_3667,N_281,N_1846);
nor U3668 (N_3668,N_1299,N_1543);
nand U3669 (N_3669,N_1168,N_1245);
xor U3670 (N_3670,N_1858,N_472);
xnor U3671 (N_3671,N_1498,N_1410);
nand U3672 (N_3672,N_652,N_275);
or U3673 (N_3673,N_1038,N_1863);
nand U3674 (N_3674,N_65,N_939);
and U3675 (N_3675,N_1621,N_817);
and U3676 (N_3676,N_137,N_1476);
xnor U3677 (N_3677,N_752,N_1842);
nor U3678 (N_3678,N_1037,N_846);
xor U3679 (N_3679,N_901,N_949);
nor U3680 (N_3680,N_720,N_1796);
nor U3681 (N_3681,N_19,N_1943);
or U3682 (N_3682,N_949,N_1934);
or U3683 (N_3683,N_770,N_1991);
nand U3684 (N_3684,N_848,N_909);
and U3685 (N_3685,N_1674,N_250);
or U3686 (N_3686,N_965,N_571);
or U3687 (N_3687,N_1179,N_1247);
nand U3688 (N_3688,N_699,N_159);
or U3689 (N_3689,N_621,N_1386);
and U3690 (N_3690,N_28,N_1827);
or U3691 (N_3691,N_1449,N_1651);
xnor U3692 (N_3692,N_347,N_1967);
or U3693 (N_3693,N_1503,N_1734);
nand U3694 (N_3694,N_1256,N_1672);
and U3695 (N_3695,N_885,N_1383);
or U3696 (N_3696,N_1946,N_1538);
nand U3697 (N_3697,N_925,N_287);
nand U3698 (N_3698,N_1404,N_943);
and U3699 (N_3699,N_891,N_1782);
and U3700 (N_3700,N_726,N_39);
or U3701 (N_3701,N_240,N_110);
nand U3702 (N_3702,N_1731,N_861);
nand U3703 (N_3703,N_853,N_1530);
or U3704 (N_3704,N_525,N_394);
xnor U3705 (N_3705,N_296,N_211);
nand U3706 (N_3706,N_781,N_663);
nand U3707 (N_3707,N_1328,N_50);
nor U3708 (N_3708,N_433,N_1496);
and U3709 (N_3709,N_461,N_394);
nor U3710 (N_3710,N_1931,N_1443);
or U3711 (N_3711,N_772,N_1933);
and U3712 (N_3712,N_881,N_1256);
or U3713 (N_3713,N_1233,N_1513);
nor U3714 (N_3714,N_978,N_1067);
and U3715 (N_3715,N_1969,N_1991);
xor U3716 (N_3716,N_1289,N_1909);
nor U3717 (N_3717,N_1452,N_18);
or U3718 (N_3718,N_1474,N_958);
or U3719 (N_3719,N_1224,N_1788);
nand U3720 (N_3720,N_1443,N_1342);
or U3721 (N_3721,N_279,N_396);
or U3722 (N_3722,N_478,N_1657);
nor U3723 (N_3723,N_120,N_920);
nand U3724 (N_3724,N_755,N_1643);
nand U3725 (N_3725,N_1148,N_1258);
xor U3726 (N_3726,N_1972,N_163);
xnor U3727 (N_3727,N_664,N_1673);
and U3728 (N_3728,N_454,N_96);
nor U3729 (N_3729,N_1486,N_89);
nor U3730 (N_3730,N_541,N_791);
nand U3731 (N_3731,N_1444,N_388);
xor U3732 (N_3732,N_265,N_1798);
nor U3733 (N_3733,N_1469,N_1073);
and U3734 (N_3734,N_1723,N_1041);
and U3735 (N_3735,N_1968,N_164);
nor U3736 (N_3736,N_654,N_302);
xor U3737 (N_3737,N_419,N_1187);
and U3738 (N_3738,N_541,N_608);
nand U3739 (N_3739,N_793,N_1248);
xor U3740 (N_3740,N_993,N_1493);
nand U3741 (N_3741,N_1518,N_1861);
and U3742 (N_3742,N_764,N_1982);
and U3743 (N_3743,N_908,N_1495);
and U3744 (N_3744,N_1461,N_542);
nand U3745 (N_3745,N_832,N_1611);
xnor U3746 (N_3746,N_1975,N_42);
nand U3747 (N_3747,N_454,N_1235);
nor U3748 (N_3748,N_1409,N_385);
and U3749 (N_3749,N_943,N_1236);
or U3750 (N_3750,N_163,N_572);
nand U3751 (N_3751,N_490,N_1349);
and U3752 (N_3752,N_549,N_664);
nand U3753 (N_3753,N_1910,N_623);
nor U3754 (N_3754,N_1772,N_743);
or U3755 (N_3755,N_737,N_679);
nor U3756 (N_3756,N_151,N_1349);
and U3757 (N_3757,N_1899,N_979);
or U3758 (N_3758,N_580,N_1534);
nand U3759 (N_3759,N_593,N_768);
xor U3760 (N_3760,N_618,N_1603);
or U3761 (N_3761,N_857,N_277);
or U3762 (N_3762,N_406,N_1925);
xor U3763 (N_3763,N_1737,N_771);
xnor U3764 (N_3764,N_1661,N_1008);
nand U3765 (N_3765,N_1070,N_618);
xnor U3766 (N_3766,N_245,N_1837);
xor U3767 (N_3767,N_289,N_1354);
nor U3768 (N_3768,N_1201,N_1817);
or U3769 (N_3769,N_173,N_1575);
nand U3770 (N_3770,N_567,N_1610);
nor U3771 (N_3771,N_1595,N_1709);
xor U3772 (N_3772,N_867,N_1027);
xnor U3773 (N_3773,N_707,N_1420);
nor U3774 (N_3774,N_261,N_342);
and U3775 (N_3775,N_220,N_39);
nor U3776 (N_3776,N_1438,N_1994);
or U3777 (N_3777,N_476,N_118);
and U3778 (N_3778,N_5,N_1516);
and U3779 (N_3779,N_716,N_1675);
nor U3780 (N_3780,N_1162,N_1801);
xor U3781 (N_3781,N_1359,N_732);
xnor U3782 (N_3782,N_3,N_55);
nor U3783 (N_3783,N_306,N_1663);
and U3784 (N_3784,N_377,N_1933);
nor U3785 (N_3785,N_1926,N_1843);
nor U3786 (N_3786,N_1193,N_1289);
nand U3787 (N_3787,N_1963,N_1464);
xnor U3788 (N_3788,N_1630,N_1082);
xor U3789 (N_3789,N_824,N_816);
xnor U3790 (N_3790,N_530,N_456);
or U3791 (N_3791,N_1839,N_1060);
nor U3792 (N_3792,N_1612,N_245);
nand U3793 (N_3793,N_1508,N_1433);
and U3794 (N_3794,N_843,N_1571);
or U3795 (N_3795,N_877,N_671);
nand U3796 (N_3796,N_1264,N_882);
and U3797 (N_3797,N_1517,N_1014);
xor U3798 (N_3798,N_1436,N_564);
nand U3799 (N_3799,N_1325,N_1203);
nor U3800 (N_3800,N_910,N_624);
or U3801 (N_3801,N_1496,N_1897);
xor U3802 (N_3802,N_1214,N_1894);
nand U3803 (N_3803,N_1902,N_764);
nor U3804 (N_3804,N_861,N_1841);
xor U3805 (N_3805,N_1680,N_1278);
and U3806 (N_3806,N_1271,N_1892);
or U3807 (N_3807,N_1260,N_1903);
nand U3808 (N_3808,N_752,N_847);
or U3809 (N_3809,N_15,N_1765);
nor U3810 (N_3810,N_453,N_181);
or U3811 (N_3811,N_1843,N_917);
and U3812 (N_3812,N_1986,N_1947);
xor U3813 (N_3813,N_1488,N_1830);
or U3814 (N_3814,N_149,N_1562);
or U3815 (N_3815,N_1345,N_1773);
and U3816 (N_3816,N_830,N_1520);
or U3817 (N_3817,N_1273,N_997);
nor U3818 (N_3818,N_675,N_1180);
nor U3819 (N_3819,N_1001,N_661);
nor U3820 (N_3820,N_692,N_1892);
and U3821 (N_3821,N_276,N_1957);
xnor U3822 (N_3822,N_127,N_922);
or U3823 (N_3823,N_791,N_612);
and U3824 (N_3824,N_451,N_1138);
and U3825 (N_3825,N_1479,N_870);
xnor U3826 (N_3826,N_1223,N_1633);
and U3827 (N_3827,N_889,N_1545);
nand U3828 (N_3828,N_511,N_895);
or U3829 (N_3829,N_1491,N_1734);
and U3830 (N_3830,N_264,N_744);
nor U3831 (N_3831,N_1680,N_720);
or U3832 (N_3832,N_1503,N_285);
nand U3833 (N_3833,N_182,N_181);
xnor U3834 (N_3834,N_1353,N_169);
and U3835 (N_3835,N_1247,N_1595);
or U3836 (N_3836,N_621,N_1966);
nand U3837 (N_3837,N_1328,N_978);
nand U3838 (N_3838,N_178,N_1602);
nor U3839 (N_3839,N_771,N_1089);
nor U3840 (N_3840,N_322,N_571);
xnor U3841 (N_3841,N_1891,N_1654);
xnor U3842 (N_3842,N_1188,N_405);
and U3843 (N_3843,N_235,N_698);
nand U3844 (N_3844,N_1555,N_1361);
nor U3845 (N_3845,N_904,N_1834);
nor U3846 (N_3846,N_1441,N_1979);
xor U3847 (N_3847,N_1729,N_1917);
nor U3848 (N_3848,N_789,N_820);
nor U3849 (N_3849,N_79,N_416);
and U3850 (N_3850,N_1459,N_283);
or U3851 (N_3851,N_297,N_1801);
nand U3852 (N_3852,N_917,N_307);
xnor U3853 (N_3853,N_614,N_766);
or U3854 (N_3854,N_625,N_310);
or U3855 (N_3855,N_132,N_1344);
nand U3856 (N_3856,N_423,N_525);
or U3857 (N_3857,N_173,N_1318);
or U3858 (N_3858,N_171,N_63);
xor U3859 (N_3859,N_1909,N_1053);
and U3860 (N_3860,N_1154,N_1779);
nand U3861 (N_3861,N_1243,N_1206);
xnor U3862 (N_3862,N_1857,N_1307);
nor U3863 (N_3863,N_1084,N_1459);
or U3864 (N_3864,N_1953,N_1871);
or U3865 (N_3865,N_63,N_765);
or U3866 (N_3866,N_40,N_1564);
xor U3867 (N_3867,N_35,N_1876);
nor U3868 (N_3868,N_315,N_1307);
nor U3869 (N_3869,N_1745,N_1932);
xnor U3870 (N_3870,N_1156,N_296);
or U3871 (N_3871,N_1448,N_1571);
nand U3872 (N_3872,N_1449,N_292);
nand U3873 (N_3873,N_589,N_449);
nor U3874 (N_3874,N_677,N_794);
nand U3875 (N_3875,N_147,N_120);
and U3876 (N_3876,N_264,N_364);
or U3877 (N_3877,N_1554,N_175);
nand U3878 (N_3878,N_765,N_1940);
nor U3879 (N_3879,N_1239,N_582);
or U3880 (N_3880,N_115,N_124);
nand U3881 (N_3881,N_1558,N_1903);
nand U3882 (N_3882,N_591,N_1252);
xor U3883 (N_3883,N_1390,N_21);
nand U3884 (N_3884,N_1388,N_286);
or U3885 (N_3885,N_1340,N_1734);
nand U3886 (N_3886,N_305,N_608);
and U3887 (N_3887,N_171,N_1566);
and U3888 (N_3888,N_261,N_1945);
nand U3889 (N_3889,N_1516,N_1949);
or U3890 (N_3890,N_634,N_913);
nand U3891 (N_3891,N_741,N_61);
or U3892 (N_3892,N_1247,N_1787);
nand U3893 (N_3893,N_1261,N_1123);
or U3894 (N_3894,N_659,N_1192);
and U3895 (N_3895,N_357,N_1415);
or U3896 (N_3896,N_1700,N_52);
nand U3897 (N_3897,N_214,N_337);
or U3898 (N_3898,N_695,N_1273);
xor U3899 (N_3899,N_1486,N_1327);
or U3900 (N_3900,N_945,N_1908);
xor U3901 (N_3901,N_1228,N_24);
or U3902 (N_3902,N_1980,N_1323);
nor U3903 (N_3903,N_852,N_1880);
nand U3904 (N_3904,N_1090,N_1395);
or U3905 (N_3905,N_819,N_1680);
and U3906 (N_3906,N_941,N_1943);
nor U3907 (N_3907,N_255,N_1517);
nand U3908 (N_3908,N_699,N_183);
or U3909 (N_3909,N_1068,N_1041);
xnor U3910 (N_3910,N_1680,N_1068);
nor U3911 (N_3911,N_1414,N_1883);
xnor U3912 (N_3912,N_1425,N_90);
nand U3913 (N_3913,N_1579,N_634);
and U3914 (N_3914,N_1422,N_994);
or U3915 (N_3915,N_46,N_974);
or U3916 (N_3916,N_288,N_902);
or U3917 (N_3917,N_1009,N_1679);
or U3918 (N_3918,N_606,N_764);
and U3919 (N_3919,N_1956,N_747);
nor U3920 (N_3920,N_1676,N_936);
nor U3921 (N_3921,N_389,N_1620);
nand U3922 (N_3922,N_666,N_279);
and U3923 (N_3923,N_51,N_1385);
xor U3924 (N_3924,N_681,N_961);
or U3925 (N_3925,N_1440,N_850);
nor U3926 (N_3926,N_1563,N_1166);
nand U3927 (N_3927,N_360,N_1591);
or U3928 (N_3928,N_1707,N_172);
nand U3929 (N_3929,N_1494,N_278);
nand U3930 (N_3930,N_1236,N_67);
xnor U3931 (N_3931,N_189,N_385);
and U3932 (N_3932,N_274,N_678);
nand U3933 (N_3933,N_493,N_418);
xor U3934 (N_3934,N_104,N_1875);
nor U3935 (N_3935,N_1606,N_1674);
and U3936 (N_3936,N_1648,N_1263);
nor U3937 (N_3937,N_1149,N_1810);
xnor U3938 (N_3938,N_1403,N_1716);
or U3939 (N_3939,N_1021,N_1964);
xor U3940 (N_3940,N_344,N_1774);
xnor U3941 (N_3941,N_1349,N_359);
nand U3942 (N_3942,N_733,N_1955);
nor U3943 (N_3943,N_575,N_173);
or U3944 (N_3944,N_838,N_1235);
and U3945 (N_3945,N_214,N_1007);
or U3946 (N_3946,N_1049,N_1757);
and U3947 (N_3947,N_1586,N_1285);
and U3948 (N_3948,N_1839,N_1967);
nor U3949 (N_3949,N_1180,N_321);
or U3950 (N_3950,N_503,N_200);
nor U3951 (N_3951,N_631,N_405);
nor U3952 (N_3952,N_58,N_3);
and U3953 (N_3953,N_1602,N_711);
xor U3954 (N_3954,N_1645,N_922);
or U3955 (N_3955,N_938,N_564);
nor U3956 (N_3956,N_1264,N_1382);
and U3957 (N_3957,N_1622,N_562);
nand U3958 (N_3958,N_1686,N_196);
xor U3959 (N_3959,N_36,N_1389);
nand U3960 (N_3960,N_494,N_1812);
nor U3961 (N_3961,N_306,N_1998);
and U3962 (N_3962,N_190,N_50);
nor U3963 (N_3963,N_1173,N_1482);
nand U3964 (N_3964,N_465,N_413);
xnor U3965 (N_3965,N_1130,N_1490);
nor U3966 (N_3966,N_319,N_645);
nor U3967 (N_3967,N_751,N_583);
and U3968 (N_3968,N_611,N_1562);
nor U3969 (N_3969,N_561,N_849);
xnor U3970 (N_3970,N_130,N_265);
xnor U3971 (N_3971,N_657,N_317);
nand U3972 (N_3972,N_808,N_1527);
nand U3973 (N_3973,N_578,N_1087);
xnor U3974 (N_3974,N_523,N_474);
xor U3975 (N_3975,N_1808,N_1948);
xor U3976 (N_3976,N_1909,N_1528);
nor U3977 (N_3977,N_791,N_235);
xnor U3978 (N_3978,N_737,N_804);
nor U3979 (N_3979,N_1160,N_1986);
and U3980 (N_3980,N_1878,N_341);
xor U3981 (N_3981,N_1878,N_760);
nand U3982 (N_3982,N_810,N_1718);
nand U3983 (N_3983,N_446,N_950);
xor U3984 (N_3984,N_1328,N_1412);
nor U3985 (N_3985,N_924,N_948);
nand U3986 (N_3986,N_819,N_648);
or U3987 (N_3987,N_1134,N_231);
xor U3988 (N_3988,N_834,N_1273);
nand U3989 (N_3989,N_1877,N_832);
and U3990 (N_3990,N_1018,N_1839);
nor U3991 (N_3991,N_146,N_1281);
nand U3992 (N_3992,N_78,N_1971);
and U3993 (N_3993,N_387,N_1190);
and U3994 (N_3994,N_473,N_5);
nand U3995 (N_3995,N_1563,N_1142);
or U3996 (N_3996,N_1664,N_1858);
or U3997 (N_3997,N_858,N_1976);
nor U3998 (N_3998,N_1894,N_1770);
and U3999 (N_3999,N_465,N_519);
nor U4000 (N_4000,N_2464,N_3001);
xnor U4001 (N_4001,N_3411,N_3661);
and U4002 (N_4002,N_2296,N_3219);
xnor U4003 (N_4003,N_3009,N_3311);
xor U4004 (N_4004,N_3615,N_3913);
and U4005 (N_4005,N_2619,N_2831);
and U4006 (N_4006,N_3078,N_3731);
and U4007 (N_4007,N_3298,N_2964);
nand U4008 (N_4008,N_2309,N_3939);
and U4009 (N_4009,N_2771,N_2457);
and U4010 (N_4010,N_2555,N_2897);
or U4011 (N_4011,N_2682,N_3320);
or U4012 (N_4012,N_2183,N_3330);
nand U4013 (N_4013,N_2116,N_2124);
nor U4014 (N_4014,N_3186,N_2988);
nor U4015 (N_4015,N_2702,N_3758);
nand U4016 (N_4016,N_3395,N_3282);
xor U4017 (N_4017,N_2929,N_2516);
xor U4018 (N_4018,N_2668,N_2001);
and U4019 (N_4019,N_2291,N_3246);
or U4020 (N_4020,N_3930,N_2432);
nor U4021 (N_4021,N_2909,N_2152);
xnor U4022 (N_4022,N_2450,N_2692);
and U4023 (N_4023,N_3029,N_2382);
nand U4024 (N_4024,N_3610,N_2992);
xnor U4025 (N_4025,N_2572,N_2591);
nand U4026 (N_4026,N_3856,N_2347);
xnor U4027 (N_4027,N_2185,N_3477);
nor U4028 (N_4028,N_3710,N_3332);
or U4029 (N_4029,N_2958,N_3734);
xor U4030 (N_4030,N_3155,N_3592);
xor U4031 (N_4031,N_2114,N_2807);
nand U4032 (N_4032,N_2921,N_3805);
xor U4033 (N_4033,N_3464,N_3491);
and U4034 (N_4034,N_2491,N_2790);
and U4035 (N_4035,N_3069,N_3879);
nor U4036 (N_4036,N_3572,N_3110);
and U4037 (N_4037,N_2246,N_2028);
nand U4038 (N_4038,N_2214,N_3988);
nand U4039 (N_4039,N_3682,N_2280);
or U4040 (N_4040,N_2436,N_2804);
nor U4041 (N_4041,N_2313,N_2845);
or U4042 (N_4042,N_2784,N_2984);
xor U4043 (N_4043,N_3277,N_3142);
nor U4044 (N_4044,N_2446,N_3551);
nand U4045 (N_4045,N_3633,N_3989);
nor U4046 (N_4046,N_3972,N_2117);
or U4047 (N_4047,N_3354,N_3278);
nor U4048 (N_4048,N_3242,N_2602);
xnor U4049 (N_4049,N_3713,N_3562);
or U4050 (N_4050,N_3489,N_3567);
xnor U4051 (N_4051,N_3265,N_2365);
nand U4052 (N_4052,N_3653,N_2484);
nor U4053 (N_4053,N_2893,N_2403);
xnor U4054 (N_4054,N_3955,N_2725);
nor U4055 (N_4055,N_2521,N_3934);
nor U4056 (N_4056,N_3349,N_3138);
nor U4057 (N_4057,N_3150,N_3241);
nor U4058 (N_4058,N_3784,N_3201);
xnor U4059 (N_4059,N_3115,N_3695);
nor U4060 (N_4060,N_2690,N_2248);
or U4061 (N_4061,N_3649,N_2648);
and U4062 (N_4062,N_2107,N_3434);
and U4063 (N_4063,N_3835,N_2411);
nor U4064 (N_4064,N_3015,N_2581);
nand U4065 (N_4065,N_3670,N_3593);
and U4066 (N_4066,N_2137,N_2552);
and U4067 (N_4067,N_3403,N_3420);
nand U4068 (N_4068,N_2695,N_2273);
nor U4069 (N_4069,N_2935,N_2997);
and U4070 (N_4070,N_2612,N_3445);
nor U4071 (N_4071,N_3602,N_3747);
and U4072 (N_4072,N_3807,N_3970);
nand U4073 (N_4073,N_3995,N_3021);
xor U4074 (N_4074,N_2136,N_3373);
and U4075 (N_4075,N_2709,N_2086);
xnor U4076 (N_4076,N_2708,N_2064);
xnor U4077 (N_4077,N_3679,N_2119);
and U4078 (N_4078,N_3595,N_3739);
nor U4079 (N_4079,N_3941,N_3986);
and U4080 (N_4080,N_2355,N_2586);
xor U4081 (N_4081,N_2974,N_3270);
nor U4082 (N_4082,N_3753,N_3639);
xor U4083 (N_4083,N_2606,N_3351);
nor U4084 (N_4084,N_2386,N_2046);
or U4085 (N_4085,N_3478,N_2035);
nand U4086 (N_4086,N_2866,N_3427);
nand U4087 (N_4087,N_3568,N_3432);
xnor U4088 (N_4088,N_2179,N_2956);
xnor U4089 (N_4089,N_3273,N_3590);
or U4090 (N_4090,N_2818,N_2111);
nand U4091 (N_4091,N_2953,N_3218);
and U4092 (N_4092,N_3006,N_3124);
and U4093 (N_4093,N_3826,N_3512);
nand U4094 (N_4094,N_2765,N_2979);
nor U4095 (N_4095,N_2652,N_3974);
or U4096 (N_4096,N_3294,N_2821);
and U4097 (N_4097,N_2631,N_3863);
xor U4098 (N_4098,N_2167,N_2522);
or U4099 (N_4099,N_2898,N_2370);
and U4100 (N_4100,N_3908,N_2138);
nand U4101 (N_4101,N_3871,N_2633);
and U4102 (N_4102,N_2348,N_2081);
or U4103 (N_4103,N_3688,N_2775);
or U4104 (N_4104,N_3185,N_2384);
or U4105 (N_4105,N_2936,N_2683);
nand U4106 (N_4106,N_2196,N_3406);
nor U4107 (N_4107,N_2045,N_3724);
nand U4108 (N_4108,N_2677,N_2938);
or U4109 (N_4109,N_3093,N_2868);
nor U4110 (N_4110,N_3870,N_2063);
and U4111 (N_4111,N_3794,N_2846);
nand U4112 (N_4112,N_3869,N_2886);
nor U4113 (N_4113,N_3823,N_3013);
or U4114 (N_4114,N_2231,N_3254);
and U4115 (N_4115,N_2226,N_2377);
xnor U4116 (N_4116,N_3251,N_2959);
nand U4117 (N_4117,N_3914,N_2147);
xor U4118 (N_4118,N_2389,N_2926);
nor U4119 (N_4119,N_3224,N_2715);
xor U4120 (N_4120,N_2737,N_2778);
xor U4121 (N_4121,N_3574,N_2177);
and U4122 (N_4122,N_3090,N_3960);
nand U4123 (N_4123,N_2392,N_3719);
xor U4124 (N_4124,N_3180,N_2057);
nor U4125 (N_4125,N_2743,N_2582);
nor U4126 (N_4126,N_2139,N_2284);
xor U4127 (N_4127,N_3382,N_2029);
xor U4128 (N_4128,N_3165,N_2169);
and U4129 (N_4129,N_2325,N_3431);
nand U4130 (N_4130,N_2971,N_3943);
nor U4131 (N_4131,N_3517,N_2584);
xnor U4132 (N_4132,N_3617,N_2858);
nand U4133 (N_4133,N_2806,N_2085);
or U4134 (N_4134,N_2294,N_3644);
nor U4135 (N_4135,N_3120,N_2453);
and U4136 (N_4136,N_2299,N_3795);
xor U4137 (N_4137,N_3392,N_3746);
nor U4138 (N_4138,N_2131,N_3302);
nor U4139 (N_4139,N_2165,N_2551);
and U4140 (N_4140,N_2203,N_2418);
or U4141 (N_4141,N_3082,N_2258);
and U4142 (N_4142,N_2757,N_3689);
nor U4143 (N_4143,N_2388,N_3528);
nor U4144 (N_4144,N_3365,N_3369);
and U4145 (N_4145,N_3225,N_2078);
nand U4146 (N_4146,N_2895,N_3027);
xor U4147 (N_4147,N_3394,N_2053);
or U4148 (N_4148,N_2467,N_3969);
or U4149 (N_4149,N_3985,N_3628);
nor U4150 (N_4150,N_2130,N_2911);
nor U4151 (N_4151,N_3133,N_2217);
xnor U4152 (N_4152,N_2480,N_3907);
or U4153 (N_4153,N_3308,N_3741);
nand U4154 (N_4154,N_2982,N_2856);
xnor U4155 (N_4155,N_2040,N_2083);
nor U4156 (N_4156,N_2822,N_2470);
or U4157 (N_4157,N_3511,N_2622);
nor U4158 (N_4158,N_3089,N_2943);
and U4159 (N_4159,N_2242,N_2367);
xor U4160 (N_4160,N_2712,N_2786);
nand U4161 (N_4161,N_2884,N_2928);
xnor U4162 (N_4162,N_2329,N_2265);
and U4163 (N_4163,N_3591,N_3864);
and U4164 (N_4164,N_3164,N_2520);
xnor U4165 (N_4165,N_2642,N_3549);
xnor U4166 (N_4166,N_3999,N_3072);
and U4167 (N_4167,N_2674,N_2317);
xnor U4168 (N_4168,N_2571,N_2635);
nand U4169 (N_4169,N_2802,N_3978);
nand U4170 (N_4170,N_3624,N_3081);
or U4171 (N_4171,N_2832,N_3279);
and U4172 (N_4172,N_3813,N_3436);
or U4173 (N_4173,N_2463,N_2537);
nand U4174 (N_4174,N_2008,N_2404);
or U4175 (N_4175,N_2553,N_2202);
or U4176 (N_4176,N_2820,N_3229);
nand U4177 (N_4177,N_2980,N_2536);
or U4178 (N_4178,N_2198,N_2228);
nor U4179 (N_4179,N_3447,N_3776);
or U4180 (N_4180,N_2458,N_3402);
xnor U4181 (N_4181,N_3884,N_3367);
nor U4182 (N_4182,N_3240,N_3560);
xor U4183 (N_4183,N_2937,N_2590);
nor U4184 (N_4184,N_3126,N_3704);
nor U4185 (N_4185,N_3339,N_3195);
and U4186 (N_4186,N_3862,N_3696);
or U4187 (N_4187,N_2274,N_3428);
xnor U4188 (N_4188,N_3751,N_2047);
nand U4189 (N_4189,N_2499,N_2286);
xor U4190 (N_4190,N_2838,N_2208);
nand U4191 (N_4191,N_3505,N_2429);
xnor U4192 (N_4192,N_3071,N_3380);
or U4193 (N_4193,N_2426,N_3793);
or U4194 (N_4194,N_3641,N_3495);
xor U4195 (N_4195,N_3401,N_2961);
and U4196 (N_4196,N_2952,N_2339);
and U4197 (N_4197,N_3327,N_3346);
nor U4198 (N_4198,N_2252,N_2594);
nand U4199 (N_4199,N_3202,N_2297);
or U4200 (N_4200,N_2719,N_3711);
or U4201 (N_4201,N_3604,N_3375);
xnor U4202 (N_4202,N_2216,N_3391);
xor U4203 (N_4203,N_2283,N_2430);
nand U4204 (N_4204,N_3827,N_3386);
nor U4205 (N_4205,N_3141,N_2768);
or U4206 (N_4206,N_3233,N_3268);
nand U4207 (N_4207,N_3287,N_3601);
xnor U4208 (N_4208,N_2113,N_3681);
nor U4209 (N_4209,N_2335,N_2192);
nand U4210 (N_4210,N_3785,N_3291);
and U4211 (N_4211,N_3239,N_3822);
or U4212 (N_4212,N_2475,N_3662);
xor U4213 (N_4213,N_2155,N_2421);
or U4214 (N_4214,N_2570,N_3897);
xnor U4215 (N_4215,N_2595,N_2910);
or U4216 (N_4216,N_2565,N_2468);
nor U4217 (N_4217,N_3703,N_2874);
nand U4218 (N_4218,N_2995,N_3646);
or U4219 (N_4219,N_2496,N_2950);
nand U4220 (N_4220,N_2308,N_2190);
or U4221 (N_4221,N_3030,N_3285);
and U4222 (N_4222,N_3471,N_2067);
nor U4223 (N_4223,N_2412,N_3345);
xnor U4224 (N_4224,N_3638,N_3041);
or U4225 (N_4225,N_3714,N_3839);
nor U4226 (N_4226,N_3315,N_2942);
xnor U4227 (N_4227,N_3306,N_3749);
nand U4228 (N_4228,N_3461,N_3786);
nor U4229 (N_4229,N_2200,N_3850);
or U4230 (N_4230,N_2098,N_3422);
nor U4231 (N_4231,N_3026,N_2704);
and U4232 (N_4232,N_3190,N_3025);
xor U4233 (N_4233,N_2282,N_2160);
and U4234 (N_4234,N_3762,N_3396);
or U4235 (N_4235,N_3368,N_2454);
nand U4236 (N_4236,N_2905,N_2750);
or U4237 (N_4237,N_3815,N_2891);
nand U4238 (N_4238,N_2834,N_3852);
nor U4239 (N_4239,N_2962,N_3452);
nor U4240 (N_4240,N_3947,N_2172);
nor U4241 (N_4241,N_2506,N_3204);
nand U4242 (N_4242,N_3017,N_3114);
and U4243 (N_4243,N_2610,N_3607);
or U4244 (N_4244,N_3187,N_2121);
xor U4245 (N_4245,N_2292,N_3178);
nor U4246 (N_4246,N_2616,N_3555);
nor U4247 (N_4247,N_3656,N_3585);
nand U4248 (N_4248,N_3425,N_2842);
xor U4249 (N_4249,N_3458,N_3766);
xor U4250 (N_4250,N_3808,N_2833);
nor U4251 (N_4251,N_3665,N_3945);
or U4252 (N_4252,N_3954,N_2346);
nor U4253 (N_4253,N_3901,N_3159);
nor U4254 (N_4254,N_3650,N_3086);
nand U4255 (N_4255,N_2830,N_2176);
or U4256 (N_4256,N_3105,N_3235);
or U4257 (N_4257,N_2061,N_3987);
nor U4258 (N_4258,N_3821,N_2120);
xnor U4259 (N_4259,N_3557,N_3725);
and U4260 (N_4260,N_3258,N_3569);
or U4261 (N_4261,N_2498,N_3627);
or U4262 (N_4262,N_2321,N_2003);
xnor U4263 (N_4263,N_3586,N_3935);
or U4264 (N_4264,N_3408,N_3255);
xnor U4265 (N_4265,N_2788,N_2052);
nor U4266 (N_4266,N_2191,N_2628);
and U4267 (N_4267,N_3553,N_3232);
and U4268 (N_4268,N_2792,N_3664);
or U4269 (N_4269,N_2968,N_2032);
nand U4270 (N_4270,N_2826,N_3675);
nor U4271 (N_4271,N_2585,N_2759);
nand U4272 (N_4272,N_2206,N_2474);
and U4273 (N_4273,N_3767,N_2302);
nand U4274 (N_4274,N_2920,N_3630);
or U4275 (N_4275,N_3832,N_2976);
or U4276 (N_4276,N_3961,N_2043);
nor U4277 (N_4277,N_2890,N_2379);
nor U4278 (N_4278,N_3581,N_2075);
xnor U4279 (N_4279,N_3023,N_3117);
nand U4280 (N_4280,N_2157,N_3531);
nor U4281 (N_4281,N_2664,N_3454);
nor U4282 (N_4282,N_2481,N_3582);
nor U4283 (N_4283,N_3243,N_2713);
xnor U4284 (N_4284,N_3177,N_2438);
nand U4285 (N_4285,N_3274,N_2090);
xnor U4286 (N_4286,N_2564,N_2767);
or U4287 (N_4287,N_3635,N_2229);
nand U4288 (N_4288,N_2754,N_2727);
or U4289 (N_4289,N_2092,N_3867);
nor U4290 (N_4290,N_3062,N_3880);
or U4291 (N_4291,N_3981,N_2721);
and U4292 (N_4292,N_2326,N_2563);
or U4293 (N_4293,N_3004,N_2049);
xor U4294 (N_4294,N_2637,N_3775);
nor U4295 (N_4295,N_2666,N_3796);
nand U4296 (N_4296,N_2808,N_2828);
nor U4297 (N_4297,N_2009,N_2981);
or U4298 (N_4298,N_3777,N_2711);
and U4299 (N_4299,N_3353,N_3619);
and U4300 (N_4300,N_3504,N_3123);
and U4301 (N_4301,N_3313,N_3005);
nor U4302 (N_4302,N_2798,N_2401);
xor U4303 (N_4303,N_3651,N_2728);
or U4304 (N_4304,N_2235,N_2914);
nand U4305 (N_4305,N_3920,N_2882);
nor U4306 (N_4306,N_3119,N_2824);
and U4307 (N_4307,N_3686,N_3131);
xor U4308 (N_4308,N_3820,N_2796);
nand U4309 (N_4309,N_2048,N_3836);
and U4310 (N_4310,N_3338,N_2425);
nand U4311 (N_4311,N_3116,N_2378);
nor U4312 (N_4312,N_2253,N_3518);
xor U4313 (N_4313,N_2592,N_2060);
and U4314 (N_4314,N_3344,N_3659);
or U4315 (N_4315,N_2251,N_3660);
or U4316 (N_4316,N_2188,N_2904);
nand U4317 (N_4317,N_3618,N_2526);
xor U4318 (N_4318,N_2636,N_3498);
xor U4319 (N_4319,N_3781,N_3101);
nand U4320 (N_4320,N_3667,N_3446);
or U4321 (N_4321,N_3075,N_2673);
nand U4322 (N_4322,N_2689,N_2059);
nand U4323 (N_4323,N_2019,N_3390);
nand U4324 (N_4324,N_3448,N_3806);
xor U4325 (N_4325,N_2143,N_3033);
nor U4326 (N_4326,N_3830,N_2755);
and U4327 (N_4327,N_3673,N_3558);
nand U4328 (N_4328,N_3376,N_2529);
and U4329 (N_4329,N_3359,N_3429);
and U4330 (N_4330,N_3441,N_3991);
and U4331 (N_4331,N_2865,N_3797);
or U4332 (N_4332,N_2414,N_3109);
nor U4333 (N_4333,N_2773,N_2741);
nor U4334 (N_4334,N_3208,N_2675);
or U4335 (N_4335,N_3564,N_3065);
nand U4336 (N_4336,N_2505,N_2447);
or U4337 (N_4337,N_3666,N_2502);
nor U4338 (N_4338,N_2399,N_2605);
xor U4339 (N_4339,N_3860,N_3900);
xnor U4340 (N_4340,N_3457,N_3002);
xor U4341 (N_4341,N_2266,N_3486);
xor U4342 (N_4342,N_3616,N_3032);
or U4343 (N_4343,N_2512,N_3510);
xor U4344 (N_4344,N_2127,N_3061);
nor U4345 (N_4345,N_3305,N_3322);
nor U4346 (N_4346,N_3112,N_3397);
or U4347 (N_4347,N_2180,N_2779);
or U4348 (N_4348,N_3523,N_3014);
and U4349 (N_4349,N_2068,N_2716);
nand U4350 (N_4350,N_2860,N_2442);
or U4351 (N_4351,N_3140,N_3068);
xor U4352 (N_4352,N_2978,N_3791);
and U4353 (N_4353,N_2915,N_3297);
xnor U4354 (N_4354,N_3144,N_2030);
nand U4355 (N_4355,N_2247,N_3479);
and U4356 (N_4356,N_3275,N_3956);
and U4357 (N_4357,N_2527,N_2580);
nor U4358 (N_4358,N_2375,N_2410);
or U4359 (N_4359,N_3923,N_3054);
xor U4360 (N_4360,N_3137,N_3768);
or U4361 (N_4361,N_2237,N_3950);
and U4362 (N_4362,N_3709,N_3449);
or U4363 (N_4363,N_3887,N_2320);
nor U4364 (N_4364,N_2099,N_3642);
nand U4365 (N_4365,N_2991,N_3559);
or U4366 (N_4366,N_3070,N_3168);
xnor U4367 (N_4367,N_2366,N_3537);
and U4368 (N_4368,N_3631,N_3355);
and U4369 (N_4369,N_2659,N_3514);
xor U4370 (N_4370,N_2693,N_2658);
nand U4371 (N_4371,N_3566,N_3050);
and U4372 (N_4372,N_2070,N_2634);
or U4373 (N_4373,N_2678,N_3372);
nand U4374 (N_4374,N_2941,N_3818);
xor U4375 (N_4375,N_3608,N_2787);
xnor U4376 (N_4376,N_3056,N_2364);
nor U4377 (N_4377,N_3634,N_2118);
or U4378 (N_4378,N_2125,N_3938);
and U4379 (N_4379,N_2772,N_3470);
nor U4380 (N_4380,N_2360,N_2532);
or U4381 (N_4381,N_2531,N_2102);
and U4382 (N_4382,N_2620,N_2990);
nand U4383 (N_4383,N_3153,N_2256);
xnor U4384 (N_4384,N_2649,N_3861);
xor U4385 (N_4385,N_2327,N_2171);
and U4386 (N_4386,N_3962,N_2500);
nor U4387 (N_4387,N_3655,N_3356);
or U4388 (N_4388,N_2912,N_3430);
nand U4389 (N_4389,N_3910,N_2896);
or U4390 (N_4390,N_2069,N_3413);
nand U4391 (N_4391,N_2469,N_3894);
nand U4392 (N_4392,N_2900,N_2760);
and U4393 (N_4393,N_3847,N_3547);
or U4394 (N_4394,N_3252,N_3924);
or U4395 (N_4395,N_2331,N_2654);
nand U4396 (N_4396,N_2916,N_3883);
nand U4397 (N_4397,N_3903,N_2254);
nand U4398 (N_4398,N_2850,N_3335);
nor U4399 (N_4399,N_3842,N_2494);
nand U4400 (N_4400,N_2651,N_3216);
nand U4401 (N_4401,N_2660,N_3337);
nand U4402 (N_4402,N_3783,N_2431);
nor U4403 (N_4403,N_3417,N_3857);
or U4404 (N_4404,N_3473,N_3881);
nor U4405 (N_4405,N_2887,N_3849);
or U4406 (N_4406,N_2776,N_2084);
nor U4407 (N_4407,N_2372,N_2538);
nor U4408 (N_4408,N_3076,N_2394);
or U4409 (N_4409,N_2363,N_2645);
xnor U4410 (N_4410,N_3760,N_3721);
or U4411 (N_4411,N_3800,N_3088);
or U4412 (N_4412,N_2140,N_3223);
xor U4413 (N_4413,N_3096,N_3362);
nand U4414 (N_4414,N_3984,N_3248);
xnor U4415 (N_4415,N_2609,N_2764);
nand U4416 (N_4416,N_3175,N_2945);
nand U4417 (N_4417,N_3622,N_3173);
and U4418 (N_4418,N_2381,N_2794);
nor U4419 (N_4419,N_2174,N_3554);
nand U4420 (N_4420,N_2336,N_2220);
nor U4421 (N_4421,N_2753,N_2290);
and U4422 (N_4422,N_2097,N_2307);
xor U4423 (N_4423,N_2880,N_3439);
or U4424 (N_4424,N_2762,N_2777);
xor U4425 (N_4425,N_3176,N_3465);
nand U4426 (N_4426,N_2397,N_2782);
and U4427 (N_4427,N_2352,N_2879);
nor U4428 (N_4428,N_2688,N_3312);
or U4429 (N_4429,N_3043,N_3042);
or U4430 (N_4430,N_3637,N_2211);
nand U4431 (N_4431,N_2146,N_2669);
or U4432 (N_4432,N_2574,N_3927);
xor U4433 (N_4433,N_3750,N_2703);
and U4434 (N_4434,N_2262,N_3379);
and U4435 (N_4435,N_2402,N_2096);
nand U4436 (N_4436,N_2698,N_3718);
xnor U4437 (N_4437,N_2338,N_2508);
or U4438 (N_4438,N_3519,N_2298);
or U4439 (N_4439,N_2306,N_2983);
xnor U4440 (N_4440,N_3000,N_2295);
or U4441 (N_4441,N_3509,N_2607);
and U4442 (N_4442,N_2444,N_2110);
xnor U4443 (N_4443,N_3301,N_3276);
xnor U4444 (N_4444,N_2748,N_2015);
nor U4445 (N_4445,N_3334,N_3416);
or U4446 (N_4446,N_3500,N_2428);
nor U4447 (N_4447,N_3522,N_3544);
and U4448 (N_4448,N_3163,N_3036);
nor U4449 (N_4449,N_2437,N_3387);
nor U4450 (N_4450,N_3497,N_3503);
nor U4451 (N_4451,N_2545,N_3092);
nor U4452 (N_4452,N_2479,N_2733);
and U4453 (N_4453,N_2917,N_2744);
nor U4454 (N_4454,N_2800,N_3605);
or U4455 (N_4455,N_2857,N_3620);
nand U4456 (N_4456,N_2749,N_3583);
xor U4457 (N_4457,N_3019,N_3828);
or U4458 (N_4458,N_3959,N_3264);
nor U4459 (N_4459,N_3811,N_3524);
or U4460 (N_4460,N_2646,N_2026);
nand U4461 (N_4461,N_2161,N_2809);
nor U4462 (N_4462,N_2497,N_3371);
nor U4463 (N_4463,N_3426,N_3035);
xor U4464 (N_4464,N_2766,N_2473);
nand U4465 (N_4465,N_2623,N_2221);
or U4466 (N_4466,N_2908,N_3570);
xnor U4467 (N_4467,N_2051,N_3217);
nand U4468 (N_4468,N_2310,N_2903);
xor U4469 (N_4469,N_2626,N_2255);
and U4470 (N_4470,N_3802,N_2416);
and U4471 (N_4471,N_2279,N_3433);
nand U4472 (N_4472,N_2215,N_3121);
nor U4473 (N_4473,N_2686,N_3318);
nand U4474 (N_4474,N_2301,N_3091);
nor U4475 (N_4475,N_2907,N_2989);
nand U4476 (N_4476,N_2181,N_3290);
and U4477 (N_4477,N_3556,N_3694);
xnor U4478 (N_4478,N_3476,N_3462);
nor U4479 (N_4479,N_2345,N_3234);
nor U4480 (N_4480,N_3552,N_3657);
nand U4481 (N_4481,N_3674,N_3669);
nand U4482 (N_4482,N_2639,N_3643);
or U4483 (N_4483,N_2460,N_3496);
nor U4484 (N_4484,N_2333,N_3690);
and U4485 (N_4485,N_2621,N_3196);
and U4486 (N_4486,N_3381,N_3438);
or U4487 (N_4487,N_2549,N_2439);
nand U4488 (N_4488,N_2542,N_3323);
and U4489 (N_4489,N_2927,N_2476);
or U4490 (N_4490,N_3303,N_3325);
and U4491 (N_4491,N_2275,N_3937);
or U4492 (N_4492,N_2742,N_3911);
xor U4493 (N_4493,N_2705,N_3728);
or U4494 (N_4494,N_2449,N_2583);
and U4495 (N_4495,N_3525,N_2337);
xor U4496 (N_4496,N_2746,N_2629);
nor U4497 (N_4497,N_2354,N_2424);
and U4498 (N_4498,N_3717,N_2955);
or U4499 (N_4499,N_2488,N_2074);
and U4500 (N_4500,N_3506,N_2611);
xnor U4501 (N_4501,N_3933,N_2696);
and U4502 (N_4502,N_2932,N_3611);
xnor U4503 (N_4503,N_2079,N_3136);
or U4504 (N_4504,N_2644,N_2109);
xor U4505 (N_4505,N_3587,N_3412);
nand U4506 (N_4506,N_2287,N_2751);
and U4507 (N_4507,N_3157,N_3418);
and U4508 (N_4508,N_3085,N_3145);
nand U4509 (N_4509,N_3975,N_2257);
nand U4510 (N_4510,N_2135,N_2493);
or U4511 (N_4511,N_3629,N_3289);
nand U4512 (N_4512,N_2272,N_2947);
nor U4513 (N_4513,N_3834,N_3865);
nor U4514 (N_4514,N_3636,N_2815);
nand U4515 (N_4515,N_3490,N_2485);
nor U4516 (N_4516,N_2197,N_2260);
or U4517 (N_4517,N_2422,N_2546);
nor U4518 (N_4518,N_3460,N_3899);
nand U4519 (N_4519,N_3215,N_3329);
nor U4520 (N_4520,N_3450,N_2848);
and U4521 (N_4521,N_3771,N_3948);
or U4522 (N_4522,N_3726,N_2038);
xnor U4523 (N_4523,N_2350,N_3542);
xor U4524 (N_4524,N_3868,N_3370);
nand U4525 (N_4525,N_3296,N_2924);
nand U4526 (N_4526,N_3194,N_3102);
or U4527 (N_4527,N_3487,N_2745);
nand U4528 (N_4528,N_3118,N_3210);
nand U4529 (N_4529,N_3451,N_3108);
nand U4530 (N_4530,N_2840,N_3648);
xor U4531 (N_4531,N_3095,N_3310);
or U4532 (N_4532,N_2706,N_3996);
and U4533 (N_4533,N_2816,N_3754);
xor U4534 (N_4534,N_2902,N_3377);
xor U4535 (N_4535,N_3804,N_2173);
nor U4536 (N_4536,N_2625,N_3099);
nand U4537 (N_4537,N_3250,N_2729);
and U4538 (N_4538,N_3729,N_3389);
xnor U4539 (N_4539,N_2797,N_3409);
nor U4540 (N_4540,N_3423,N_2482);
nor U4541 (N_4541,N_3499,N_2986);
nor U4542 (N_4542,N_2371,N_3295);
xor U4543 (N_4543,N_2567,N_2811);
nand U4544 (N_4544,N_3189,N_2261);
nand U4545 (N_4545,N_2734,N_3331);
nand U4546 (N_4546,N_2044,N_3892);
and U4547 (N_4547,N_3925,N_2883);
nor U4548 (N_4548,N_3011,N_2210);
nand U4549 (N_4549,N_2685,N_2847);
and U4550 (N_4550,N_2730,N_3341);
or U4551 (N_4551,N_3501,N_3456);
and U4552 (N_4552,N_3854,N_3084);
xor U4553 (N_4553,N_3626,N_2182);
nand U4554 (N_4554,N_2836,N_3366);
and U4555 (N_4555,N_2018,N_2641);
nor U4556 (N_4556,N_2054,N_2667);
or U4557 (N_4557,N_2332,N_2509);
nor U4558 (N_4558,N_2672,N_2603);
or U4559 (N_4559,N_3982,N_3012);
and U4560 (N_4560,N_2653,N_2073);
and U4561 (N_4561,N_3442,N_2839);
or U4562 (N_4562,N_2328,N_3957);
nand U4563 (N_4563,N_3198,N_2710);
and U4564 (N_4564,N_2560,N_3336);
xor U4565 (N_4565,N_3513,N_2141);
nand U4566 (N_4566,N_3571,N_3779);
or U4567 (N_4567,N_3993,N_2888);
xor U4568 (N_4568,N_3735,N_3474);
nand U4569 (N_4569,N_3200,N_2525);
nand U4570 (N_4570,N_2691,N_2153);
and U4571 (N_4571,N_3563,N_3399);
nor U4572 (N_4572,N_2236,N_3761);
and U4573 (N_4573,N_2819,N_2738);
nor U4574 (N_4574,N_2000,N_2507);
nand U4575 (N_4575,N_2596,N_3106);
or U4576 (N_4576,N_3966,N_3931);
and U4577 (N_4577,N_2534,N_3221);
or U4578 (N_4578,N_2112,N_3541);
nor U4579 (N_4579,N_2873,N_2513);
nand U4580 (N_4580,N_3730,N_3702);
and U4581 (N_4581,N_3789,N_2376);
or U4582 (N_4582,N_3580,N_2101);
nand U4583 (N_4583,N_2087,N_2965);
or U4584 (N_4584,N_3594,N_2535);
or U4585 (N_4585,N_3024,N_2756);
nor U4586 (N_4586,N_3022,N_2071);
xor U4587 (N_4587,N_3663,N_3578);
xnor U4588 (N_4588,N_3918,N_3772);
and U4589 (N_4589,N_2913,N_2278);
or U4590 (N_4590,N_2150,N_3845);
nor U4591 (N_4591,N_2351,N_3833);
and U4592 (N_4592,N_3837,N_2960);
and U4593 (N_4593,N_2540,N_2814);
and U4594 (N_4594,N_2142,N_3171);
nand U4595 (N_4595,N_3316,N_2359);
xnor U4596 (N_4596,N_2230,N_2195);
and U4597 (N_4597,N_2993,N_3520);
or U4598 (N_4598,N_2556,N_3814);
and U4599 (N_4599,N_3151,N_3917);
nor U4600 (N_4600,N_3257,N_2440);
nand U4601 (N_4601,N_2277,N_2025);
or U4602 (N_4602,N_3016,N_2684);
nand U4603 (N_4603,N_3128,N_3886);
nor U4604 (N_4604,N_2657,N_3527);
nor U4605 (N_4605,N_3152,N_3819);
or U4606 (N_4606,N_3378,N_2362);
nand U4607 (N_4607,N_2881,N_2934);
nor U4608 (N_4608,N_3342,N_3148);
or U4609 (N_4609,N_3193,N_2168);
and U4610 (N_4610,N_2740,N_3851);
xnor U4611 (N_4611,N_3971,N_2036);
xnor U4612 (N_4612,N_3625,N_2383);
and U4613 (N_4613,N_3716,N_2722);
or U4614 (N_4614,N_2643,N_3983);
or U4615 (N_4615,N_3492,N_2514);
xnor U4616 (N_4616,N_2518,N_2853);
or U4617 (N_4617,N_2569,N_2393);
and U4618 (N_4618,N_3576,N_2353);
xor U4619 (N_4619,N_2205,N_2227);
or U4620 (N_4620,N_3535,N_3515);
or U4621 (N_4621,N_2483,N_2967);
nand U4622 (N_4622,N_3272,N_2922);
nor U4623 (N_4623,N_2793,N_3885);
xor U4624 (N_4624,N_3443,N_2323);
xnor U4625 (N_4625,N_3846,N_2162);
and U4626 (N_4626,N_2400,N_3684);
xor U4627 (N_4627,N_3994,N_2080);
or U4628 (N_4628,N_2864,N_2316);
nand U4629 (N_4629,N_2267,N_3130);
or U4630 (N_4630,N_3475,N_2234);
or U4631 (N_4631,N_2975,N_3953);
nor U4632 (N_4632,N_2419,N_3206);
and U4633 (N_4633,N_2213,N_2558);
nor U4634 (N_4634,N_3181,N_2547);
and U4635 (N_4635,N_2562,N_2471);
and U4636 (N_4636,N_3697,N_2655);
nand U4637 (N_4637,N_2184,N_2977);
and U4638 (N_4638,N_3536,N_2238);
and U4639 (N_4639,N_3949,N_2005);
nor U4640 (N_4640,N_2720,N_3074);
nand U4641 (N_4641,N_3748,N_3936);
and U4642 (N_4642,N_3598,N_2559);
or U4643 (N_4643,N_2761,N_2212);
or U4644 (N_4644,N_2533,N_2638);
or U4645 (N_4645,N_2770,N_2598);
nor U4646 (N_4646,N_2999,N_2923);
nor U4647 (N_4647,N_2024,N_2349);
and U4648 (N_4648,N_3149,N_3609);
nor U4649 (N_4649,N_2931,N_2434);
and U4650 (N_4650,N_3770,N_3468);
or U4651 (N_4651,N_3964,N_3192);
nor U4652 (N_4652,N_2058,N_3952);
or U4653 (N_4653,N_2561,N_2134);
and U4654 (N_4654,N_2700,N_2420);
nand U4655 (N_4655,N_2875,N_3902);
nand U4656 (N_4656,N_3079,N_2944);
xor U4657 (N_4657,N_3825,N_3266);
or U4658 (N_4658,N_2687,N_2245);
and U4659 (N_4659,N_2519,N_2825);
or U4660 (N_4660,N_3600,N_3259);
nor U4661 (N_4661,N_2813,N_2939);
xnor U4662 (N_4662,N_3533,N_2852);
and U4663 (N_4663,N_2361,N_2369);
nor U4664 (N_4664,N_3579,N_2726);
nor U4665 (N_4665,N_2163,N_3973);
or U4666 (N_4666,N_3671,N_2576);
and U4667 (N_4667,N_3191,N_2007);
nand U4668 (N_4668,N_3039,N_2614);
xor U4669 (N_4669,N_3053,N_3307);
nand U4670 (N_4670,N_2006,N_2731);
xor U4671 (N_4671,N_2014,N_3328);
nand U4672 (N_4672,N_2489,N_2341);
nor U4673 (N_4673,N_3589,N_3077);
xnor U4674 (N_4674,N_2827,N_2285);
nor U4675 (N_4675,N_3107,N_2854);
and U4676 (N_4676,N_2517,N_3502);
and U4677 (N_4677,N_3060,N_3699);
xor U4678 (N_4678,N_3172,N_2305);
or U4679 (N_4679,N_2264,N_3809);
nand U4680 (N_4680,N_3769,N_2849);
xnor U4681 (N_4681,N_2224,N_3098);
or U4682 (N_4682,N_3286,N_3018);
or U4683 (N_4683,N_3236,N_2630);
nor U4684 (N_4684,N_3787,N_2448);
nand U4685 (N_4685,N_3965,N_2878);
xor U4686 (N_4686,N_2544,N_2568);
nor U4687 (N_4687,N_2515,N_2501);
nand U4688 (N_4688,N_2785,N_2201);
nor U4689 (N_4689,N_2843,N_2918);
xnor U4690 (N_4690,N_2963,N_3031);
or U4691 (N_4691,N_3146,N_2694);
and U4692 (N_4692,N_3958,N_2933);
nand U4693 (N_4693,N_3799,N_2011);
or U4694 (N_4694,N_2413,N_3213);
or U4695 (N_4695,N_3599,N_3841);
nor U4696 (N_4696,N_2579,N_2799);
and U4697 (N_4697,N_3222,N_3757);
nand U4698 (N_4698,N_3358,N_3052);
xnor U4699 (N_4699,N_3540,N_2548);
nor U4700 (N_4700,N_3059,N_2342);
xnor U4701 (N_4701,N_3944,N_2010);
nor U4702 (N_4702,N_3737,N_3980);
xor U4703 (N_4703,N_3143,N_2632);
nand U4704 (N_4704,N_3040,N_3691);
and U4705 (N_4705,N_2618,N_2218);
nand U4706 (N_4706,N_2844,N_2670);
nor U4707 (N_4707,N_2543,N_2207);
nand U4708 (N_4708,N_2650,N_3237);
nor U4709 (N_4709,N_3742,N_2356);
and U4710 (N_4710,N_3238,N_3812);
or U4711 (N_4711,N_2503,N_2249);
and U4712 (N_4712,N_3467,N_2089);
and U4713 (N_4713,N_3113,N_3169);
or U4714 (N_4714,N_3269,N_3534);
and U4715 (N_4715,N_3603,N_3654);
and U4716 (N_4716,N_3979,N_3199);
or U4717 (N_4717,N_2012,N_3007);
nand U4718 (N_4718,N_3780,N_3227);
and U4719 (N_4719,N_2593,N_3384);
xnor U4720 (N_4720,N_3521,N_2919);
and U4721 (N_4721,N_2077,N_2578);
nand U4722 (N_4722,N_3680,N_2889);
nand U4723 (N_4723,N_2662,N_3493);
and U4724 (N_4724,N_3621,N_3293);
xnor U4725 (N_4725,N_3057,N_3708);
xnor U4726 (N_4726,N_2324,N_2042);
xor U4727 (N_4727,N_3840,N_2970);
nor U4728 (N_4728,N_3614,N_3921);
xor U4729 (N_4729,N_3508,N_3977);
and U4730 (N_4730,N_2504,N_3324);
nor U4731 (N_4731,N_3179,N_3890);
nand U4732 (N_4732,N_2647,N_3774);
nor U4733 (N_4733,N_2718,N_3055);
nand U4734 (N_4734,N_3584,N_3744);
or U4735 (N_4735,N_3701,N_2189);
or U4736 (N_4736,N_3104,N_2244);
nor U4737 (N_4737,N_3790,N_3488);
nor U4738 (N_4738,N_3385,N_3260);
nor U4739 (N_4739,N_2396,N_2066);
nor U4740 (N_4740,N_3135,N_3824);
nor U4741 (N_4741,N_2156,N_3008);
xnor U4742 (N_4742,N_3632,N_3577);
or U4743 (N_4743,N_3469,N_3759);
and U4744 (N_4744,N_2193,N_3707);
xor U4745 (N_4745,N_3565,N_3245);
nand U4746 (N_4746,N_3532,N_3909);
and U4747 (N_4747,N_3435,N_3051);
xor U4748 (N_4748,N_2405,N_2930);
xnor U4749 (N_4749,N_2835,N_2243);
or U4750 (N_4750,N_2149,N_3419);
nor U4751 (N_4751,N_2863,N_2587);
and U4752 (N_4752,N_3444,N_2062);
xnor U4753 (N_4753,N_3097,N_3882);
nor U4754 (N_4754,N_3606,N_3174);
nand U4755 (N_4755,N_2478,N_2222);
xnor U4756 (N_4756,N_2170,N_3896);
or U4757 (N_4757,N_3314,N_3546);
nand U4758 (N_4758,N_2311,N_2732);
nor U4759 (N_4759,N_2717,N_3732);
nor U4760 (N_4760,N_3858,N_3755);
nand U4761 (N_4761,N_2656,N_3915);
and U4762 (N_4762,N_2783,N_3727);
xnor U4763 (N_4763,N_2701,N_2186);
or U4764 (N_4764,N_3752,N_2957);
xnor U4765 (N_4765,N_2714,N_3678);
nor U4766 (N_4766,N_2966,N_3816);
nor U4767 (N_4767,N_2148,N_2608);
nor U4768 (N_4768,N_3951,N_3817);
and U4769 (N_4769,N_2510,N_3928);
and U4770 (N_4770,N_3067,N_3765);
nand U4771 (N_4771,N_3410,N_2225);
and U4772 (N_4772,N_3485,N_3158);
xnor U4773 (N_4773,N_2268,N_3877);
xor U4774 (N_4774,N_3612,N_2391);
nor U4775 (N_4775,N_3122,N_2472);
or U4776 (N_4776,N_3407,N_2315);
nor U4777 (N_4777,N_3687,N_3706);
or U4778 (N_4778,N_2837,N_2406);
nor U4779 (N_4779,N_2461,N_2859);
or U4780 (N_4780,N_3028,N_3782);
or U4781 (N_4781,N_2037,N_2407);
nand U4782 (N_4782,N_3209,N_2940);
or U4783 (N_4783,N_2899,N_3170);
nor U4784 (N_4784,N_3183,N_3919);
or U4785 (N_4785,N_3037,N_3803);
and U4786 (N_4786,N_3872,N_2219);
or U4787 (N_4787,N_3288,N_3677);
xnor U4788 (N_4788,N_2270,N_3575);
nand U4789 (N_4789,N_3244,N_2223);
xor U4790 (N_4790,N_3127,N_3685);
nor U4791 (N_4791,N_3182,N_3094);
nand U4792 (N_4792,N_3946,N_2577);
nor U4793 (N_4793,N_2303,N_2330);
xnor U4794 (N_4794,N_2041,N_3494);
and U4795 (N_4795,N_2758,N_3997);
xor U4796 (N_4796,N_3049,N_2663);
nand U4797 (N_4797,N_3350,N_3792);
nor U4798 (N_4798,N_2877,N_2697);
and U4799 (N_4799,N_2627,N_3773);
xnor U4800 (N_4800,N_2300,N_2435);
and U4801 (N_4801,N_3167,N_2823);
or U4802 (N_4802,N_2871,N_2707);
and U4803 (N_4803,N_3154,N_3374);
and U4804 (N_4804,N_2615,N_2948);
and U4805 (N_4805,N_2817,N_2573);
nand U4806 (N_4806,N_3249,N_3692);
nand U4807 (N_4807,N_2841,N_2679);
and U4808 (N_4808,N_2613,N_3672);
xor U4809 (N_4809,N_2949,N_2423);
xnor U4810 (N_4810,N_2604,N_2194);
xnor U4811 (N_4811,N_2312,N_3596);
nand U4812 (N_4812,N_3459,N_2803);
nor U4813 (N_4813,N_3893,N_2154);
and U4814 (N_4814,N_2829,N_3405);
xnor U4815 (N_4815,N_3976,N_3640);
and U4816 (N_4816,N_2699,N_3645);
or U4817 (N_4817,N_2343,N_3722);
nand U4818 (N_4818,N_3404,N_2851);
nor U4819 (N_4819,N_2017,N_3745);
and U4820 (N_4820,N_2151,N_2455);
nor U4821 (N_4821,N_2951,N_2892);
xor U4822 (N_4822,N_3211,N_2954);
xor U4823 (N_4823,N_3526,N_3848);
xor U4824 (N_4824,N_3214,N_3364);
and U4825 (N_4825,N_2665,N_2209);
and U4826 (N_4826,N_2998,N_2319);
xnor U4827 (N_4827,N_2969,N_2322);
nand U4828 (N_4828,N_2385,N_3888);
nand U4829 (N_4829,N_2002,N_3898);
nand U4830 (N_4830,N_2021,N_3588);
xnor U4831 (N_4831,N_3440,N_3271);
nand U4832 (N_4832,N_2946,N_3360);
nand U4833 (N_4833,N_2869,N_2289);
or U4834 (N_4834,N_3363,N_2133);
nand U4835 (N_4835,N_2723,N_3073);
and U4836 (N_4836,N_2390,N_2204);
nand U4837 (N_4837,N_3463,N_3788);
and U4838 (N_4838,N_3347,N_2250);
or U4839 (N_4839,N_3400,N_2056);
xnor U4840 (N_4840,N_2810,N_3889);
nor U4841 (N_4841,N_3317,N_3188);
or U4842 (N_4842,N_2128,N_2812);
and U4843 (N_4843,N_2082,N_2122);
nor U4844 (N_4844,N_3080,N_2158);
or U4845 (N_4845,N_3166,N_3044);
nand U4846 (N_4846,N_3147,N_3161);
and U4847 (N_4847,N_2022,N_2027);
nand U4848 (N_4848,N_3623,N_2259);
nand U4849 (N_4849,N_3348,N_3284);
and U4850 (N_4850,N_2736,N_3683);
xnor U4851 (N_4851,N_3453,N_2805);
nor U4852 (N_4852,N_3162,N_3658);
or U4853 (N_4853,N_3220,N_3020);
nor U4854 (N_4854,N_3160,N_2769);
or U4855 (N_4855,N_2088,N_2016);
nor U4856 (N_4856,N_3261,N_3134);
nor U4857 (N_4857,N_2452,N_2528);
and U4858 (N_4858,N_2395,N_3875);
nor U4859 (N_4859,N_3228,N_2492);
nor U4860 (N_4860,N_2987,N_3545);
or U4861 (N_4861,N_3756,N_2288);
or U4862 (N_4862,N_3963,N_3926);
and U4863 (N_4863,N_2380,N_3003);
or U4864 (N_4864,N_3357,N_2985);
nor U4865 (N_4865,N_2462,N_3083);
nand U4866 (N_4866,N_3992,N_2752);
nor U4867 (N_4867,N_3247,N_2076);
nor U4868 (N_4868,N_2539,N_2588);
nor U4869 (N_4869,N_2801,N_2676);
xor U4870 (N_4870,N_2013,N_2373);
and U4871 (N_4871,N_3668,N_3878);
or U4872 (N_4872,N_3652,N_2199);
nand U4873 (N_4873,N_2269,N_3466);
nor U4874 (N_4874,N_2304,N_2600);
nor U4875 (N_4875,N_3929,N_2735);
nand U4876 (N_4876,N_3529,N_2894);
or U4877 (N_4877,N_2640,N_2281);
nor U4878 (N_4878,N_2374,N_2340);
or U4879 (N_4879,N_2427,N_3844);
or U4880 (N_4880,N_2597,N_2318);
or U4881 (N_4881,N_2456,N_3740);
or U4882 (N_4882,N_2115,N_3916);
nor U4883 (N_4883,N_3763,N_3129);
xor U4884 (N_4884,N_3676,N_2123);
nor U4885 (N_4885,N_3415,N_3309);
xnor U4886 (N_4886,N_2867,N_2050);
or U4887 (N_4887,N_3383,N_3111);
xor U4888 (N_4888,N_2126,N_3398);
and U4889 (N_4889,N_2072,N_2415);
xnor U4890 (N_4890,N_2680,N_3904);
xnor U4891 (N_4891,N_2417,N_2566);
or U4892 (N_4892,N_2164,N_3810);
and U4893 (N_4893,N_3895,N_2144);
and U4894 (N_4894,N_3343,N_2906);
nand U4895 (N_4895,N_3738,N_2617);
nor U4896 (N_4896,N_3942,N_3340);
nor U4897 (N_4897,N_3231,N_2550);
nor U4898 (N_4898,N_2145,N_3698);
or U4899 (N_4899,N_2575,N_2240);
xor U4900 (N_4900,N_3715,N_2681);
nand U4901 (N_4901,N_3843,N_3139);
nand U4902 (N_4902,N_2232,N_3100);
and U4903 (N_4903,N_3829,N_2108);
xor U4904 (N_4904,N_3990,N_2443);
nor U4905 (N_4905,N_2523,N_2293);
or U4906 (N_4906,N_3263,N_3859);
xnor U4907 (N_4907,N_3855,N_3530);
and U4908 (N_4908,N_2105,N_3968);
nand U4909 (N_4909,N_2314,N_3253);
or U4910 (N_4910,N_3967,N_3733);
nand U4911 (N_4911,N_3472,N_2100);
nand U4912 (N_4912,N_3299,N_2885);
nand U4913 (N_4913,N_3778,N_2739);
nor U4914 (N_4914,N_3561,N_2132);
nor U4915 (N_4915,N_3321,N_2241);
nor U4916 (N_4916,N_2466,N_2486);
nor U4917 (N_4917,N_3801,N_3046);
nor U4918 (N_4918,N_3922,N_2409);
nand U4919 (N_4919,N_2004,N_2094);
nor U4920 (N_4920,N_3876,N_3212);
nor U4921 (N_4921,N_2724,N_3543);
xnor U4922 (N_4922,N_3712,N_3613);
nor U4923 (N_4923,N_3831,N_2387);
xnor U4924 (N_4924,N_2031,N_3230);
or U4925 (N_4925,N_3304,N_2747);
xnor U4926 (N_4926,N_3481,N_2530);
and U4927 (N_4927,N_2039,N_3048);
or U4928 (N_4928,N_3262,N_3421);
nor U4929 (N_4929,N_2093,N_2870);
or U4930 (N_4930,N_3292,N_2187);
and U4931 (N_4931,N_3538,N_2901);
nand U4932 (N_4932,N_2129,N_3038);
or U4933 (N_4933,N_3424,N_2490);
xnor U4934 (N_4934,N_3281,N_2239);
and U4935 (N_4935,N_3798,N_3184);
nand U4936 (N_4936,N_3932,N_3891);
nand U4937 (N_4937,N_2175,N_3010);
nor U4938 (N_4938,N_3507,N_2095);
and U4939 (N_4939,N_2973,N_2862);
nor U4940 (N_4940,N_3764,N_3693);
xor U4941 (N_4941,N_2445,N_2599);
or U4942 (N_4942,N_3197,N_3205);
nand U4943 (N_4943,N_3873,N_3414);
nand U4944 (N_4944,N_3480,N_3326);
nand U4945 (N_4945,N_2861,N_3103);
and U4946 (N_4946,N_2166,N_3548);
xor U4947 (N_4947,N_3573,N_2020);
nor U4948 (N_4948,N_2023,N_2601);
or U4949 (N_4949,N_2781,N_3207);
and U4950 (N_4950,N_3063,N_2358);
and U4951 (N_4951,N_3034,N_3125);
nand U4952 (N_4952,N_2524,N_2398);
nor U4953 (N_4953,N_3647,N_3482);
nor U4954 (N_4954,N_3906,N_2994);
nand U4955 (N_4955,N_3998,N_2795);
nor U4956 (N_4956,N_3940,N_3267);
nor U4957 (N_4957,N_3905,N_3736);
or U4958 (N_4958,N_2661,N_2065);
or U4959 (N_4959,N_3874,N_2033);
nand U4960 (N_4960,N_2178,N_2671);
nand U4961 (N_4961,N_3866,N_3064);
xor U4962 (N_4962,N_3087,N_3597);
and U4963 (N_4963,N_2451,N_2091);
or U4964 (N_4964,N_3066,N_2034);
nor U4965 (N_4965,N_3352,N_3720);
and U4966 (N_4966,N_3319,N_2487);
xnor U4967 (N_4967,N_3047,N_3393);
nand U4968 (N_4968,N_2276,N_2271);
nor U4969 (N_4969,N_2465,N_2511);
and U4970 (N_4970,N_2459,N_3388);
nand U4971 (N_4971,N_2554,N_2106);
xor U4972 (N_4972,N_2368,N_3045);
nand U4973 (N_4973,N_3705,N_2477);
or U4974 (N_4974,N_3743,N_3539);
nand U4975 (N_4975,N_2876,N_2408);
xor U4976 (N_4976,N_3300,N_2104);
nand U4977 (N_4977,N_3723,N_2780);
xnor U4978 (N_4978,N_2789,N_3333);
or U4979 (N_4979,N_3203,N_2495);
or U4980 (N_4980,N_3058,N_3838);
nand U4981 (N_4981,N_2972,N_3484);
xor U4982 (N_4982,N_3437,N_3156);
xnor U4983 (N_4983,N_3132,N_3283);
and U4984 (N_4984,N_3280,N_2344);
and U4985 (N_4985,N_3483,N_2855);
xnor U4986 (N_4986,N_2996,N_2433);
nor U4987 (N_4987,N_2441,N_3256);
xor U4988 (N_4988,N_2872,N_3226);
or U4989 (N_4989,N_2263,N_3361);
xnor U4990 (N_4990,N_2589,N_3700);
nor U4991 (N_4991,N_2624,N_3550);
and U4992 (N_4992,N_3516,N_2774);
nor U4993 (N_4993,N_2925,N_2159);
or U4994 (N_4994,N_2357,N_2103);
xnor U4995 (N_4995,N_3912,N_2763);
xnor U4996 (N_4996,N_2557,N_2334);
or U4997 (N_4997,N_2791,N_3853);
xor U4998 (N_4998,N_2055,N_2233);
or U4999 (N_4999,N_3455,N_2541);
or U5000 (N_5000,N_2588,N_2414);
and U5001 (N_5001,N_2803,N_2095);
nand U5002 (N_5002,N_3148,N_3548);
nor U5003 (N_5003,N_2240,N_2952);
nor U5004 (N_5004,N_2358,N_3505);
nand U5005 (N_5005,N_3226,N_2579);
nand U5006 (N_5006,N_2835,N_3831);
or U5007 (N_5007,N_2321,N_3168);
nand U5008 (N_5008,N_2800,N_3051);
and U5009 (N_5009,N_3792,N_2867);
nand U5010 (N_5010,N_2180,N_2888);
nor U5011 (N_5011,N_2340,N_3007);
nor U5012 (N_5012,N_2286,N_3547);
and U5013 (N_5013,N_2919,N_2978);
xor U5014 (N_5014,N_3809,N_2256);
xor U5015 (N_5015,N_3516,N_3902);
or U5016 (N_5016,N_3638,N_3904);
and U5017 (N_5017,N_2482,N_3240);
or U5018 (N_5018,N_3659,N_3680);
and U5019 (N_5019,N_3869,N_2124);
nand U5020 (N_5020,N_3324,N_3914);
or U5021 (N_5021,N_3331,N_2097);
xor U5022 (N_5022,N_2946,N_2735);
xor U5023 (N_5023,N_3062,N_3416);
xor U5024 (N_5024,N_3469,N_2341);
and U5025 (N_5025,N_3468,N_3472);
xor U5026 (N_5026,N_2698,N_3535);
nand U5027 (N_5027,N_3623,N_2245);
and U5028 (N_5028,N_3713,N_3506);
nor U5029 (N_5029,N_2461,N_3596);
or U5030 (N_5030,N_3948,N_3018);
xnor U5031 (N_5031,N_3743,N_3071);
xnor U5032 (N_5032,N_3349,N_3733);
nor U5033 (N_5033,N_3210,N_3933);
nand U5034 (N_5034,N_3930,N_3380);
nor U5035 (N_5035,N_2083,N_2697);
xor U5036 (N_5036,N_2465,N_3482);
xor U5037 (N_5037,N_3111,N_2744);
nand U5038 (N_5038,N_3842,N_2072);
nor U5039 (N_5039,N_2864,N_2973);
nand U5040 (N_5040,N_3636,N_3370);
xor U5041 (N_5041,N_2343,N_2468);
nand U5042 (N_5042,N_2904,N_3741);
nand U5043 (N_5043,N_2682,N_3906);
xor U5044 (N_5044,N_2187,N_2837);
nor U5045 (N_5045,N_3018,N_2658);
nand U5046 (N_5046,N_2049,N_2612);
nand U5047 (N_5047,N_3984,N_2256);
xnor U5048 (N_5048,N_3900,N_2729);
nor U5049 (N_5049,N_2775,N_3519);
and U5050 (N_5050,N_3466,N_2568);
and U5051 (N_5051,N_2122,N_2966);
or U5052 (N_5052,N_3781,N_3520);
and U5053 (N_5053,N_3386,N_2256);
nand U5054 (N_5054,N_3789,N_2229);
or U5055 (N_5055,N_2446,N_2578);
and U5056 (N_5056,N_2287,N_2663);
and U5057 (N_5057,N_2674,N_2110);
and U5058 (N_5058,N_2340,N_3947);
nand U5059 (N_5059,N_3695,N_2061);
xnor U5060 (N_5060,N_2186,N_2208);
xnor U5061 (N_5061,N_3933,N_2014);
xnor U5062 (N_5062,N_2500,N_3070);
and U5063 (N_5063,N_3553,N_2755);
nand U5064 (N_5064,N_3271,N_3269);
xnor U5065 (N_5065,N_3031,N_2451);
xnor U5066 (N_5066,N_2791,N_2212);
and U5067 (N_5067,N_2669,N_2163);
nand U5068 (N_5068,N_3800,N_2383);
xor U5069 (N_5069,N_2514,N_3865);
nand U5070 (N_5070,N_2725,N_2588);
xor U5071 (N_5071,N_3076,N_3025);
or U5072 (N_5072,N_3232,N_2093);
and U5073 (N_5073,N_2012,N_2276);
nor U5074 (N_5074,N_3002,N_3087);
nor U5075 (N_5075,N_2859,N_2424);
xor U5076 (N_5076,N_3677,N_3883);
nor U5077 (N_5077,N_2858,N_2476);
or U5078 (N_5078,N_2714,N_2383);
nand U5079 (N_5079,N_2488,N_3340);
nor U5080 (N_5080,N_3267,N_2037);
nor U5081 (N_5081,N_3548,N_3476);
and U5082 (N_5082,N_2327,N_3340);
or U5083 (N_5083,N_3690,N_2589);
and U5084 (N_5084,N_2561,N_3718);
and U5085 (N_5085,N_2627,N_3020);
xnor U5086 (N_5086,N_2213,N_3506);
or U5087 (N_5087,N_2777,N_2963);
nand U5088 (N_5088,N_2499,N_3343);
nand U5089 (N_5089,N_2468,N_3316);
and U5090 (N_5090,N_2773,N_3800);
nand U5091 (N_5091,N_2629,N_2575);
nor U5092 (N_5092,N_3771,N_3002);
nand U5093 (N_5093,N_2341,N_3312);
nor U5094 (N_5094,N_3170,N_3292);
nor U5095 (N_5095,N_2317,N_2749);
and U5096 (N_5096,N_2143,N_2930);
nor U5097 (N_5097,N_3850,N_2638);
xnor U5098 (N_5098,N_3613,N_2912);
nand U5099 (N_5099,N_3370,N_2920);
or U5100 (N_5100,N_2041,N_2557);
xor U5101 (N_5101,N_3795,N_3512);
nand U5102 (N_5102,N_2358,N_2573);
or U5103 (N_5103,N_2701,N_3777);
and U5104 (N_5104,N_3100,N_2920);
nand U5105 (N_5105,N_2791,N_2261);
and U5106 (N_5106,N_3469,N_3666);
and U5107 (N_5107,N_3963,N_2108);
or U5108 (N_5108,N_2709,N_2179);
and U5109 (N_5109,N_3312,N_3921);
nor U5110 (N_5110,N_2597,N_3369);
nor U5111 (N_5111,N_2519,N_2952);
or U5112 (N_5112,N_3127,N_2825);
or U5113 (N_5113,N_2515,N_3111);
xnor U5114 (N_5114,N_2490,N_3130);
xor U5115 (N_5115,N_3110,N_3350);
and U5116 (N_5116,N_2640,N_3408);
nor U5117 (N_5117,N_2473,N_2561);
nand U5118 (N_5118,N_3074,N_2676);
and U5119 (N_5119,N_3296,N_3494);
or U5120 (N_5120,N_3971,N_3573);
or U5121 (N_5121,N_2452,N_2931);
xor U5122 (N_5122,N_3106,N_3111);
xnor U5123 (N_5123,N_3334,N_3482);
and U5124 (N_5124,N_3168,N_3027);
nand U5125 (N_5125,N_2295,N_3253);
and U5126 (N_5126,N_3768,N_3267);
nand U5127 (N_5127,N_2816,N_2233);
or U5128 (N_5128,N_3498,N_2855);
or U5129 (N_5129,N_3891,N_2746);
or U5130 (N_5130,N_3931,N_3633);
nand U5131 (N_5131,N_3796,N_2554);
or U5132 (N_5132,N_3333,N_3198);
nor U5133 (N_5133,N_2384,N_3377);
or U5134 (N_5134,N_3500,N_2719);
and U5135 (N_5135,N_2072,N_3488);
or U5136 (N_5136,N_2937,N_3466);
nor U5137 (N_5137,N_3717,N_3798);
nor U5138 (N_5138,N_2061,N_3615);
or U5139 (N_5139,N_2304,N_3162);
and U5140 (N_5140,N_2953,N_3232);
xor U5141 (N_5141,N_2490,N_3126);
nor U5142 (N_5142,N_3924,N_2857);
and U5143 (N_5143,N_3108,N_3967);
xor U5144 (N_5144,N_2944,N_3934);
or U5145 (N_5145,N_2499,N_2219);
nand U5146 (N_5146,N_2513,N_3474);
nand U5147 (N_5147,N_2298,N_3649);
xnor U5148 (N_5148,N_3160,N_2272);
nand U5149 (N_5149,N_2203,N_2312);
xor U5150 (N_5150,N_2520,N_2322);
xor U5151 (N_5151,N_2868,N_3521);
nand U5152 (N_5152,N_3806,N_3026);
xnor U5153 (N_5153,N_2342,N_2374);
nand U5154 (N_5154,N_3651,N_2639);
nand U5155 (N_5155,N_2538,N_2297);
nand U5156 (N_5156,N_3220,N_2163);
or U5157 (N_5157,N_3629,N_3231);
xnor U5158 (N_5158,N_3551,N_2476);
and U5159 (N_5159,N_3268,N_3472);
nand U5160 (N_5160,N_2491,N_3556);
nand U5161 (N_5161,N_2714,N_2824);
and U5162 (N_5162,N_2356,N_3436);
or U5163 (N_5163,N_3442,N_2386);
and U5164 (N_5164,N_2323,N_2357);
xnor U5165 (N_5165,N_3006,N_2466);
and U5166 (N_5166,N_3720,N_3089);
or U5167 (N_5167,N_2763,N_2081);
nand U5168 (N_5168,N_3554,N_3092);
nand U5169 (N_5169,N_2181,N_2468);
xnor U5170 (N_5170,N_3195,N_2573);
or U5171 (N_5171,N_3826,N_3114);
and U5172 (N_5172,N_3056,N_2607);
xor U5173 (N_5173,N_3147,N_2028);
xor U5174 (N_5174,N_2327,N_2631);
nor U5175 (N_5175,N_3107,N_2419);
nand U5176 (N_5176,N_3389,N_2020);
or U5177 (N_5177,N_2713,N_2574);
nor U5178 (N_5178,N_2090,N_2876);
and U5179 (N_5179,N_2967,N_2889);
nor U5180 (N_5180,N_2354,N_3429);
or U5181 (N_5181,N_3885,N_2758);
nand U5182 (N_5182,N_3828,N_2668);
nor U5183 (N_5183,N_2940,N_3001);
and U5184 (N_5184,N_3621,N_3664);
nand U5185 (N_5185,N_2927,N_3520);
nor U5186 (N_5186,N_3020,N_2615);
xnor U5187 (N_5187,N_3676,N_2770);
nor U5188 (N_5188,N_3798,N_2736);
and U5189 (N_5189,N_2544,N_3327);
and U5190 (N_5190,N_2788,N_2700);
xnor U5191 (N_5191,N_3435,N_2913);
nor U5192 (N_5192,N_2884,N_3835);
nand U5193 (N_5193,N_2008,N_3470);
and U5194 (N_5194,N_3591,N_3691);
nand U5195 (N_5195,N_3661,N_3370);
nand U5196 (N_5196,N_2271,N_2280);
xnor U5197 (N_5197,N_2709,N_3922);
nor U5198 (N_5198,N_3667,N_2665);
and U5199 (N_5199,N_2471,N_3329);
and U5200 (N_5200,N_3542,N_3100);
and U5201 (N_5201,N_2670,N_2070);
or U5202 (N_5202,N_3694,N_3875);
nor U5203 (N_5203,N_2853,N_2697);
nor U5204 (N_5204,N_2275,N_2256);
xor U5205 (N_5205,N_3622,N_2110);
or U5206 (N_5206,N_3173,N_2862);
xor U5207 (N_5207,N_2611,N_2320);
nand U5208 (N_5208,N_2883,N_2478);
nor U5209 (N_5209,N_2860,N_2741);
nor U5210 (N_5210,N_2084,N_2850);
nor U5211 (N_5211,N_2523,N_3692);
and U5212 (N_5212,N_3560,N_2793);
nor U5213 (N_5213,N_2745,N_3096);
xor U5214 (N_5214,N_2555,N_3469);
or U5215 (N_5215,N_3356,N_2685);
or U5216 (N_5216,N_2099,N_2184);
and U5217 (N_5217,N_2480,N_3547);
nor U5218 (N_5218,N_2512,N_3727);
nor U5219 (N_5219,N_2709,N_3292);
nand U5220 (N_5220,N_3343,N_2540);
nor U5221 (N_5221,N_3748,N_2859);
or U5222 (N_5222,N_3159,N_3671);
xor U5223 (N_5223,N_2275,N_3464);
or U5224 (N_5224,N_2277,N_2069);
xnor U5225 (N_5225,N_2938,N_3858);
nor U5226 (N_5226,N_2021,N_3166);
xnor U5227 (N_5227,N_2911,N_2748);
and U5228 (N_5228,N_2073,N_3310);
nor U5229 (N_5229,N_2372,N_3183);
nor U5230 (N_5230,N_2072,N_2982);
and U5231 (N_5231,N_2989,N_2196);
xor U5232 (N_5232,N_3672,N_2484);
nand U5233 (N_5233,N_2532,N_3154);
nor U5234 (N_5234,N_3327,N_2880);
or U5235 (N_5235,N_3822,N_3161);
nor U5236 (N_5236,N_3292,N_3839);
or U5237 (N_5237,N_2402,N_3021);
or U5238 (N_5238,N_2439,N_2933);
xnor U5239 (N_5239,N_2135,N_3165);
xor U5240 (N_5240,N_2971,N_2932);
xor U5241 (N_5241,N_3047,N_3090);
or U5242 (N_5242,N_3558,N_3762);
nand U5243 (N_5243,N_3431,N_3382);
xnor U5244 (N_5244,N_2203,N_3466);
xor U5245 (N_5245,N_3182,N_3150);
nor U5246 (N_5246,N_3244,N_2287);
xnor U5247 (N_5247,N_3063,N_3245);
or U5248 (N_5248,N_2185,N_3280);
and U5249 (N_5249,N_3119,N_2158);
and U5250 (N_5250,N_2131,N_2591);
nor U5251 (N_5251,N_2661,N_3428);
nor U5252 (N_5252,N_3886,N_3058);
nor U5253 (N_5253,N_3259,N_2584);
and U5254 (N_5254,N_3066,N_3798);
nand U5255 (N_5255,N_2840,N_2758);
xor U5256 (N_5256,N_3167,N_3680);
xnor U5257 (N_5257,N_3146,N_3684);
nand U5258 (N_5258,N_3087,N_2046);
and U5259 (N_5259,N_2663,N_2598);
xnor U5260 (N_5260,N_2509,N_3988);
and U5261 (N_5261,N_3556,N_3771);
nor U5262 (N_5262,N_2690,N_2876);
and U5263 (N_5263,N_3941,N_3386);
and U5264 (N_5264,N_3496,N_2470);
nor U5265 (N_5265,N_2352,N_3861);
or U5266 (N_5266,N_2123,N_3160);
xnor U5267 (N_5267,N_3963,N_2208);
nor U5268 (N_5268,N_3981,N_2553);
xor U5269 (N_5269,N_2373,N_3824);
and U5270 (N_5270,N_3875,N_2190);
and U5271 (N_5271,N_3717,N_3593);
xnor U5272 (N_5272,N_2058,N_2401);
nor U5273 (N_5273,N_2940,N_2269);
nand U5274 (N_5274,N_2957,N_3980);
or U5275 (N_5275,N_2842,N_3835);
and U5276 (N_5276,N_2417,N_2829);
or U5277 (N_5277,N_2512,N_2409);
nand U5278 (N_5278,N_3644,N_3412);
nand U5279 (N_5279,N_2358,N_2697);
xor U5280 (N_5280,N_2280,N_2313);
nand U5281 (N_5281,N_2374,N_2545);
xnor U5282 (N_5282,N_2282,N_3007);
nor U5283 (N_5283,N_2601,N_3458);
and U5284 (N_5284,N_2175,N_3598);
nor U5285 (N_5285,N_3482,N_2586);
or U5286 (N_5286,N_2831,N_2779);
nand U5287 (N_5287,N_3515,N_2961);
xor U5288 (N_5288,N_3096,N_2062);
nand U5289 (N_5289,N_3178,N_3002);
nand U5290 (N_5290,N_3479,N_2931);
xor U5291 (N_5291,N_2117,N_2899);
or U5292 (N_5292,N_3266,N_3988);
nand U5293 (N_5293,N_3831,N_2628);
xor U5294 (N_5294,N_2573,N_3046);
and U5295 (N_5295,N_2563,N_2825);
nand U5296 (N_5296,N_3043,N_2415);
nor U5297 (N_5297,N_2010,N_3501);
nand U5298 (N_5298,N_2647,N_3924);
nor U5299 (N_5299,N_3281,N_2583);
nor U5300 (N_5300,N_3074,N_2973);
nor U5301 (N_5301,N_3385,N_3961);
or U5302 (N_5302,N_3731,N_2275);
and U5303 (N_5303,N_2451,N_3365);
nand U5304 (N_5304,N_3547,N_3457);
or U5305 (N_5305,N_2525,N_2106);
nor U5306 (N_5306,N_3576,N_3417);
and U5307 (N_5307,N_2149,N_3919);
or U5308 (N_5308,N_2521,N_3763);
nor U5309 (N_5309,N_2468,N_3665);
nor U5310 (N_5310,N_3753,N_3228);
or U5311 (N_5311,N_2659,N_2141);
nor U5312 (N_5312,N_2034,N_2220);
and U5313 (N_5313,N_3574,N_2345);
xor U5314 (N_5314,N_2215,N_2706);
xor U5315 (N_5315,N_2489,N_3726);
and U5316 (N_5316,N_2740,N_2573);
nand U5317 (N_5317,N_3218,N_3983);
nand U5318 (N_5318,N_2825,N_3362);
nand U5319 (N_5319,N_2494,N_3780);
nand U5320 (N_5320,N_2033,N_2380);
and U5321 (N_5321,N_2421,N_3626);
nand U5322 (N_5322,N_3347,N_2487);
nand U5323 (N_5323,N_3091,N_2673);
nor U5324 (N_5324,N_2680,N_3553);
and U5325 (N_5325,N_2397,N_3715);
nor U5326 (N_5326,N_3912,N_2959);
xor U5327 (N_5327,N_3026,N_2497);
or U5328 (N_5328,N_3907,N_3391);
nand U5329 (N_5329,N_3004,N_3425);
nand U5330 (N_5330,N_3487,N_2594);
or U5331 (N_5331,N_3496,N_3756);
and U5332 (N_5332,N_2846,N_2345);
nor U5333 (N_5333,N_2072,N_2280);
and U5334 (N_5334,N_2358,N_2891);
and U5335 (N_5335,N_3854,N_3964);
nand U5336 (N_5336,N_3179,N_3243);
xor U5337 (N_5337,N_3261,N_2540);
nand U5338 (N_5338,N_2445,N_2777);
and U5339 (N_5339,N_2862,N_3391);
nor U5340 (N_5340,N_3023,N_2906);
nand U5341 (N_5341,N_2478,N_3672);
nand U5342 (N_5342,N_2090,N_2916);
nand U5343 (N_5343,N_3414,N_3110);
or U5344 (N_5344,N_3683,N_3695);
nor U5345 (N_5345,N_3121,N_3059);
nor U5346 (N_5346,N_2040,N_2183);
nand U5347 (N_5347,N_2166,N_3379);
and U5348 (N_5348,N_3150,N_2722);
xnor U5349 (N_5349,N_3116,N_2747);
nor U5350 (N_5350,N_3160,N_2237);
xnor U5351 (N_5351,N_2774,N_3749);
nand U5352 (N_5352,N_3627,N_3891);
nor U5353 (N_5353,N_3821,N_3622);
or U5354 (N_5354,N_3538,N_2874);
and U5355 (N_5355,N_2484,N_3303);
xor U5356 (N_5356,N_2643,N_2508);
nand U5357 (N_5357,N_3746,N_3682);
nand U5358 (N_5358,N_2228,N_3790);
xnor U5359 (N_5359,N_2687,N_2047);
and U5360 (N_5360,N_3137,N_3984);
nor U5361 (N_5361,N_2165,N_2669);
nor U5362 (N_5362,N_3701,N_2009);
nand U5363 (N_5363,N_2837,N_3334);
nor U5364 (N_5364,N_2710,N_2298);
xor U5365 (N_5365,N_2709,N_3350);
or U5366 (N_5366,N_2186,N_2062);
nor U5367 (N_5367,N_3375,N_3681);
or U5368 (N_5368,N_2055,N_2056);
nor U5369 (N_5369,N_3349,N_3511);
and U5370 (N_5370,N_2250,N_3395);
nor U5371 (N_5371,N_3008,N_3195);
or U5372 (N_5372,N_3956,N_3352);
nand U5373 (N_5373,N_2149,N_3924);
xnor U5374 (N_5374,N_2689,N_3034);
xor U5375 (N_5375,N_2511,N_2417);
xnor U5376 (N_5376,N_3580,N_3099);
and U5377 (N_5377,N_3934,N_2334);
or U5378 (N_5378,N_2943,N_3752);
nor U5379 (N_5379,N_2805,N_3011);
and U5380 (N_5380,N_2482,N_3361);
nor U5381 (N_5381,N_3582,N_3633);
and U5382 (N_5382,N_3907,N_3142);
or U5383 (N_5383,N_3193,N_2032);
or U5384 (N_5384,N_3913,N_3944);
nor U5385 (N_5385,N_2085,N_2650);
xnor U5386 (N_5386,N_2802,N_3827);
xor U5387 (N_5387,N_2979,N_2947);
or U5388 (N_5388,N_2616,N_3892);
xnor U5389 (N_5389,N_3351,N_3211);
nor U5390 (N_5390,N_2045,N_2731);
nand U5391 (N_5391,N_3764,N_2841);
nand U5392 (N_5392,N_3070,N_2123);
or U5393 (N_5393,N_2158,N_2670);
nor U5394 (N_5394,N_3971,N_2760);
nor U5395 (N_5395,N_2103,N_2898);
nor U5396 (N_5396,N_2308,N_3594);
or U5397 (N_5397,N_2240,N_2940);
nand U5398 (N_5398,N_3289,N_2200);
nor U5399 (N_5399,N_2796,N_3542);
and U5400 (N_5400,N_2076,N_3985);
nor U5401 (N_5401,N_3903,N_2990);
xor U5402 (N_5402,N_2150,N_2208);
or U5403 (N_5403,N_3562,N_2161);
or U5404 (N_5404,N_3998,N_2892);
xor U5405 (N_5405,N_3948,N_3410);
and U5406 (N_5406,N_3717,N_2203);
or U5407 (N_5407,N_2082,N_3747);
nand U5408 (N_5408,N_3537,N_2137);
xnor U5409 (N_5409,N_2901,N_2131);
nand U5410 (N_5410,N_3906,N_2139);
or U5411 (N_5411,N_3364,N_3252);
xnor U5412 (N_5412,N_3044,N_2401);
nand U5413 (N_5413,N_2332,N_2971);
nand U5414 (N_5414,N_2622,N_2897);
or U5415 (N_5415,N_2797,N_3078);
nand U5416 (N_5416,N_3776,N_2262);
or U5417 (N_5417,N_2738,N_3855);
nor U5418 (N_5418,N_2529,N_2797);
or U5419 (N_5419,N_3107,N_3716);
xnor U5420 (N_5420,N_2869,N_3675);
or U5421 (N_5421,N_3898,N_3112);
nor U5422 (N_5422,N_3544,N_2345);
or U5423 (N_5423,N_2562,N_2718);
or U5424 (N_5424,N_2338,N_2156);
or U5425 (N_5425,N_2778,N_2394);
xor U5426 (N_5426,N_3643,N_3752);
and U5427 (N_5427,N_3260,N_2498);
nor U5428 (N_5428,N_2511,N_3166);
xnor U5429 (N_5429,N_2305,N_2989);
nand U5430 (N_5430,N_3999,N_2912);
or U5431 (N_5431,N_3098,N_2339);
or U5432 (N_5432,N_3053,N_3836);
nor U5433 (N_5433,N_2883,N_3713);
nor U5434 (N_5434,N_3541,N_2407);
nand U5435 (N_5435,N_3404,N_2948);
nor U5436 (N_5436,N_3720,N_2639);
or U5437 (N_5437,N_3715,N_3456);
and U5438 (N_5438,N_3425,N_2426);
xor U5439 (N_5439,N_2568,N_2324);
or U5440 (N_5440,N_2919,N_3885);
and U5441 (N_5441,N_3142,N_2666);
nand U5442 (N_5442,N_3424,N_2076);
nand U5443 (N_5443,N_2313,N_2896);
nand U5444 (N_5444,N_3335,N_3970);
nand U5445 (N_5445,N_2429,N_2419);
or U5446 (N_5446,N_3029,N_3754);
or U5447 (N_5447,N_2124,N_2211);
nand U5448 (N_5448,N_2542,N_3410);
nor U5449 (N_5449,N_2122,N_2032);
nor U5450 (N_5450,N_3713,N_3939);
xnor U5451 (N_5451,N_3770,N_3064);
xnor U5452 (N_5452,N_3706,N_3211);
nand U5453 (N_5453,N_2234,N_2263);
and U5454 (N_5454,N_3754,N_3219);
xor U5455 (N_5455,N_3324,N_2899);
xor U5456 (N_5456,N_3994,N_3185);
or U5457 (N_5457,N_2677,N_3642);
nor U5458 (N_5458,N_2446,N_2594);
or U5459 (N_5459,N_3082,N_3661);
nor U5460 (N_5460,N_2496,N_2629);
nor U5461 (N_5461,N_3548,N_3582);
nor U5462 (N_5462,N_3548,N_2867);
xnor U5463 (N_5463,N_2029,N_3551);
nand U5464 (N_5464,N_3879,N_3948);
xnor U5465 (N_5465,N_2743,N_3124);
or U5466 (N_5466,N_2585,N_3078);
nor U5467 (N_5467,N_2411,N_3146);
or U5468 (N_5468,N_3462,N_3508);
and U5469 (N_5469,N_2040,N_3597);
nor U5470 (N_5470,N_2916,N_3708);
nand U5471 (N_5471,N_2294,N_3128);
xnor U5472 (N_5472,N_3101,N_3203);
or U5473 (N_5473,N_3524,N_2570);
xnor U5474 (N_5474,N_2573,N_3079);
nand U5475 (N_5475,N_3189,N_3345);
xor U5476 (N_5476,N_3128,N_3634);
nand U5477 (N_5477,N_2749,N_3234);
xor U5478 (N_5478,N_3273,N_3312);
xnor U5479 (N_5479,N_2580,N_3398);
and U5480 (N_5480,N_3824,N_2317);
nand U5481 (N_5481,N_3541,N_3285);
nor U5482 (N_5482,N_2485,N_2972);
or U5483 (N_5483,N_2633,N_3631);
or U5484 (N_5484,N_2818,N_2908);
nor U5485 (N_5485,N_2468,N_2507);
nor U5486 (N_5486,N_2664,N_3311);
or U5487 (N_5487,N_3566,N_2361);
or U5488 (N_5488,N_2200,N_3215);
and U5489 (N_5489,N_3150,N_2486);
xnor U5490 (N_5490,N_2006,N_3550);
xnor U5491 (N_5491,N_3041,N_3544);
nor U5492 (N_5492,N_3728,N_3615);
nand U5493 (N_5493,N_2403,N_3791);
nor U5494 (N_5494,N_3944,N_3722);
xnor U5495 (N_5495,N_3441,N_2936);
and U5496 (N_5496,N_3700,N_2447);
xnor U5497 (N_5497,N_2501,N_3457);
or U5498 (N_5498,N_3862,N_2185);
and U5499 (N_5499,N_2538,N_3970);
and U5500 (N_5500,N_2786,N_3860);
nand U5501 (N_5501,N_3150,N_2074);
or U5502 (N_5502,N_3083,N_3380);
xor U5503 (N_5503,N_2144,N_3444);
nand U5504 (N_5504,N_2803,N_2823);
nor U5505 (N_5505,N_3787,N_3278);
nor U5506 (N_5506,N_2615,N_3678);
and U5507 (N_5507,N_3569,N_3105);
nand U5508 (N_5508,N_3558,N_2972);
xnor U5509 (N_5509,N_2309,N_3284);
or U5510 (N_5510,N_2614,N_3939);
xnor U5511 (N_5511,N_2210,N_2302);
nand U5512 (N_5512,N_3731,N_2878);
or U5513 (N_5513,N_2398,N_2270);
xnor U5514 (N_5514,N_2603,N_3251);
xnor U5515 (N_5515,N_2768,N_2002);
xnor U5516 (N_5516,N_3550,N_2123);
nor U5517 (N_5517,N_2834,N_3535);
nor U5518 (N_5518,N_3413,N_2954);
nand U5519 (N_5519,N_3925,N_2253);
nor U5520 (N_5520,N_2074,N_3503);
nor U5521 (N_5521,N_3132,N_3418);
nand U5522 (N_5522,N_2107,N_3155);
or U5523 (N_5523,N_3518,N_2739);
or U5524 (N_5524,N_3438,N_3004);
nor U5525 (N_5525,N_3933,N_3989);
nand U5526 (N_5526,N_3130,N_2327);
xor U5527 (N_5527,N_2566,N_2624);
or U5528 (N_5528,N_2677,N_2092);
or U5529 (N_5529,N_2501,N_3683);
and U5530 (N_5530,N_3445,N_2989);
nand U5531 (N_5531,N_2934,N_3345);
or U5532 (N_5532,N_2498,N_3090);
or U5533 (N_5533,N_2107,N_3415);
and U5534 (N_5534,N_3344,N_2131);
and U5535 (N_5535,N_3786,N_2674);
nor U5536 (N_5536,N_2364,N_2663);
nand U5537 (N_5537,N_3593,N_2168);
nand U5538 (N_5538,N_2462,N_2709);
or U5539 (N_5539,N_3051,N_3681);
xnor U5540 (N_5540,N_3080,N_3892);
nand U5541 (N_5541,N_2032,N_2587);
or U5542 (N_5542,N_3382,N_3702);
nor U5543 (N_5543,N_3164,N_3410);
nand U5544 (N_5544,N_3283,N_2444);
nor U5545 (N_5545,N_3182,N_2033);
nand U5546 (N_5546,N_3356,N_3465);
nor U5547 (N_5547,N_3588,N_2383);
or U5548 (N_5548,N_3963,N_2184);
or U5549 (N_5549,N_3074,N_2748);
nor U5550 (N_5550,N_3171,N_3801);
nor U5551 (N_5551,N_3614,N_3528);
and U5552 (N_5552,N_3866,N_3635);
and U5553 (N_5553,N_2017,N_2041);
nand U5554 (N_5554,N_2369,N_3674);
xor U5555 (N_5555,N_2426,N_3577);
nand U5556 (N_5556,N_3967,N_3177);
xor U5557 (N_5557,N_3842,N_2569);
nor U5558 (N_5558,N_2299,N_3944);
and U5559 (N_5559,N_2154,N_3064);
and U5560 (N_5560,N_2801,N_3063);
or U5561 (N_5561,N_2585,N_2270);
nand U5562 (N_5562,N_2245,N_2322);
and U5563 (N_5563,N_3947,N_3956);
and U5564 (N_5564,N_2175,N_2247);
nand U5565 (N_5565,N_2932,N_3807);
xor U5566 (N_5566,N_3309,N_3554);
nor U5567 (N_5567,N_3879,N_3286);
nor U5568 (N_5568,N_2594,N_2668);
or U5569 (N_5569,N_3099,N_2380);
or U5570 (N_5570,N_3474,N_3722);
nand U5571 (N_5571,N_3337,N_2931);
and U5572 (N_5572,N_2329,N_3584);
nor U5573 (N_5573,N_3817,N_3558);
or U5574 (N_5574,N_3397,N_3566);
xnor U5575 (N_5575,N_3989,N_2904);
xor U5576 (N_5576,N_3300,N_2536);
xnor U5577 (N_5577,N_2354,N_3421);
or U5578 (N_5578,N_2594,N_3927);
and U5579 (N_5579,N_3470,N_2180);
nand U5580 (N_5580,N_3108,N_2210);
or U5581 (N_5581,N_2329,N_2185);
and U5582 (N_5582,N_2327,N_2767);
or U5583 (N_5583,N_2636,N_3153);
xnor U5584 (N_5584,N_2484,N_2470);
nand U5585 (N_5585,N_2409,N_2625);
xnor U5586 (N_5586,N_3576,N_3481);
nand U5587 (N_5587,N_3751,N_3840);
and U5588 (N_5588,N_2225,N_2943);
or U5589 (N_5589,N_2441,N_2716);
and U5590 (N_5590,N_2348,N_2655);
and U5591 (N_5591,N_2435,N_2078);
nand U5592 (N_5592,N_2661,N_2421);
and U5593 (N_5593,N_2020,N_2885);
nand U5594 (N_5594,N_3133,N_3472);
and U5595 (N_5595,N_3109,N_3637);
nor U5596 (N_5596,N_3254,N_2651);
and U5597 (N_5597,N_3532,N_3597);
nand U5598 (N_5598,N_3065,N_3850);
nor U5599 (N_5599,N_3226,N_2900);
and U5600 (N_5600,N_2186,N_2762);
or U5601 (N_5601,N_3533,N_3516);
and U5602 (N_5602,N_3025,N_3515);
or U5603 (N_5603,N_2706,N_3927);
or U5604 (N_5604,N_3781,N_2761);
and U5605 (N_5605,N_3610,N_2169);
or U5606 (N_5606,N_2881,N_2176);
nor U5607 (N_5607,N_2529,N_2144);
nand U5608 (N_5608,N_3842,N_2842);
nor U5609 (N_5609,N_3321,N_3756);
xor U5610 (N_5610,N_2184,N_2837);
nor U5611 (N_5611,N_3148,N_3889);
xnor U5612 (N_5612,N_2469,N_2149);
and U5613 (N_5613,N_2498,N_2767);
nor U5614 (N_5614,N_2345,N_2479);
xor U5615 (N_5615,N_3810,N_3180);
or U5616 (N_5616,N_2410,N_2902);
nand U5617 (N_5617,N_3621,N_2958);
xnor U5618 (N_5618,N_3393,N_3334);
or U5619 (N_5619,N_2635,N_2700);
and U5620 (N_5620,N_2675,N_2930);
nand U5621 (N_5621,N_3687,N_2807);
and U5622 (N_5622,N_3549,N_3086);
nand U5623 (N_5623,N_3076,N_2620);
nand U5624 (N_5624,N_3612,N_2333);
nand U5625 (N_5625,N_3780,N_3919);
nor U5626 (N_5626,N_3001,N_2369);
nand U5627 (N_5627,N_2238,N_2942);
nand U5628 (N_5628,N_2232,N_3936);
nor U5629 (N_5629,N_3029,N_3450);
or U5630 (N_5630,N_3844,N_3319);
nor U5631 (N_5631,N_2797,N_2853);
xnor U5632 (N_5632,N_2887,N_3477);
nand U5633 (N_5633,N_2222,N_3379);
nand U5634 (N_5634,N_2841,N_3494);
nand U5635 (N_5635,N_2911,N_3179);
xnor U5636 (N_5636,N_3176,N_3984);
xor U5637 (N_5637,N_3645,N_2406);
nand U5638 (N_5638,N_2994,N_2423);
and U5639 (N_5639,N_2767,N_3299);
nor U5640 (N_5640,N_3360,N_2393);
or U5641 (N_5641,N_2879,N_3509);
and U5642 (N_5642,N_3611,N_2921);
and U5643 (N_5643,N_3094,N_2739);
nor U5644 (N_5644,N_3528,N_3405);
or U5645 (N_5645,N_3576,N_2778);
nor U5646 (N_5646,N_2737,N_3995);
or U5647 (N_5647,N_3344,N_2659);
nand U5648 (N_5648,N_2806,N_3809);
xor U5649 (N_5649,N_2942,N_3846);
nor U5650 (N_5650,N_2320,N_2268);
nor U5651 (N_5651,N_2597,N_3288);
and U5652 (N_5652,N_2904,N_2197);
xnor U5653 (N_5653,N_2615,N_3918);
or U5654 (N_5654,N_3652,N_3906);
and U5655 (N_5655,N_3341,N_2916);
or U5656 (N_5656,N_2443,N_3414);
nand U5657 (N_5657,N_3448,N_2077);
and U5658 (N_5658,N_3214,N_3272);
and U5659 (N_5659,N_3615,N_2933);
or U5660 (N_5660,N_2722,N_2190);
xor U5661 (N_5661,N_3333,N_2754);
xor U5662 (N_5662,N_3684,N_2584);
or U5663 (N_5663,N_2557,N_2046);
xor U5664 (N_5664,N_2410,N_2198);
nand U5665 (N_5665,N_2477,N_3130);
or U5666 (N_5666,N_3530,N_3148);
nor U5667 (N_5667,N_2685,N_2417);
nor U5668 (N_5668,N_2891,N_3252);
xnor U5669 (N_5669,N_3883,N_2098);
or U5670 (N_5670,N_2858,N_3482);
xor U5671 (N_5671,N_3741,N_2315);
xnor U5672 (N_5672,N_3629,N_3095);
nor U5673 (N_5673,N_3600,N_3027);
nor U5674 (N_5674,N_2196,N_2762);
and U5675 (N_5675,N_2686,N_3801);
and U5676 (N_5676,N_2902,N_3477);
and U5677 (N_5677,N_3137,N_2755);
or U5678 (N_5678,N_2969,N_3353);
and U5679 (N_5679,N_2616,N_3223);
nand U5680 (N_5680,N_2825,N_2166);
and U5681 (N_5681,N_3508,N_3700);
nor U5682 (N_5682,N_3954,N_2008);
nor U5683 (N_5683,N_2005,N_3904);
nor U5684 (N_5684,N_2544,N_3794);
or U5685 (N_5685,N_3407,N_3603);
xnor U5686 (N_5686,N_2097,N_2613);
and U5687 (N_5687,N_3108,N_3521);
nor U5688 (N_5688,N_2589,N_2988);
xnor U5689 (N_5689,N_3454,N_2560);
nand U5690 (N_5690,N_3379,N_3435);
nor U5691 (N_5691,N_3451,N_3706);
xor U5692 (N_5692,N_3028,N_3619);
and U5693 (N_5693,N_2958,N_3192);
and U5694 (N_5694,N_3015,N_2889);
or U5695 (N_5695,N_2133,N_3664);
or U5696 (N_5696,N_3366,N_3713);
xnor U5697 (N_5697,N_2650,N_2090);
nand U5698 (N_5698,N_2227,N_3481);
nor U5699 (N_5699,N_3697,N_2039);
and U5700 (N_5700,N_2586,N_3952);
nand U5701 (N_5701,N_2361,N_2613);
nand U5702 (N_5702,N_2381,N_3620);
or U5703 (N_5703,N_3423,N_3715);
nand U5704 (N_5704,N_2164,N_2175);
and U5705 (N_5705,N_3028,N_3636);
xor U5706 (N_5706,N_2142,N_3128);
and U5707 (N_5707,N_2289,N_3278);
xnor U5708 (N_5708,N_2403,N_3523);
xor U5709 (N_5709,N_3918,N_2741);
xor U5710 (N_5710,N_2389,N_3328);
xnor U5711 (N_5711,N_2134,N_3627);
xnor U5712 (N_5712,N_2261,N_2688);
nand U5713 (N_5713,N_3042,N_3254);
nor U5714 (N_5714,N_2711,N_2360);
or U5715 (N_5715,N_3211,N_2857);
xor U5716 (N_5716,N_2171,N_2712);
or U5717 (N_5717,N_2785,N_2272);
and U5718 (N_5718,N_3665,N_3207);
xnor U5719 (N_5719,N_3919,N_2333);
or U5720 (N_5720,N_3448,N_2673);
and U5721 (N_5721,N_2689,N_2719);
or U5722 (N_5722,N_2580,N_3295);
nor U5723 (N_5723,N_3611,N_2513);
nand U5724 (N_5724,N_3025,N_3065);
nand U5725 (N_5725,N_2994,N_3911);
nand U5726 (N_5726,N_2300,N_3763);
nand U5727 (N_5727,N_2633,N_3809);
and U5728 (N_5728,N_3916,N_3819);
nand U5729 (N_5729,N_3796,N_3042);
and U5730 (N_5730,N_2928,N_3605);
xnor U5731 (N_5731,N_2221,N_2842);
and U5732 (N_5732,N_2044,N_2157);
and U5733 (N_5733,N_3630,N_2721);
or U5734 (N_5734,N_2830,N_3295);
nor U5735 (N_5735,N_2173,N_3898);
xor U5736 (N_5736,N_2292,N_3938);
xor U5737 (N_5737,N_3479,N_3556);
and U5738 (N_5738,N_2520,N_3979);
xor U5739 (N_5739,N_2746,N_3469);
xnor U5740 (N_5740,N_3363,N_2179);
xor U5741 (N_5741,N_3645,N_3958);
xor U5742 (N_5742,N_3752,N_3626);
or U5743 (N_5743,N_2181,N_3040);
or U5744 (N_5744,N_3555,N_3678);
and U5745 (N_5745,N_2299,N_3436);
xnor U5746 (N_5746,N_3791,N_3122);
nand U5747 (N_5747,N_2962,N_3044);
and U5748 (N_5748,N_3878,N_2084);
nand U5749 (N_5749,N_2967,N_3903);
nand U5750 (N_5750,N_3506,N_2418);
nand U5751 (N_5751,N_3389,N_2688);
or U5752 (N_5752,N_2690,N_3460);
xor U5753 (N_5753,N_2900,N_2303);
nor U5754 (N_5754,N_3235,N_3075);
xnor U5755 (N_5755,N_2057,N_2930);
nand U5756 (N_5756,N_3626,N_2822);
and U5757 (N_5757,N_3745,N_2016);
nor U5758 (N_5758,N_3421,N_2216);
and U5759 (N_5759,N_3154,N_3169);
xnor U5760 (N_5760,N_3364,N_3082);
or U5761 (N_5761,N_2564,N_3315);
nand U5762 (N_5762,N_3977,N_3934);
nor U5763 (N_5763,N_3425,N_2304);
and U5764 (N_5764,N_3320,N_3415);
or U5765 (N_5765,N_3461,N_3133);
and U5766 (N_5766,N_3625,N_2173);
nand U5767 (N_5767,N_2388,N_3994);
xnor U5768 (N_5768,N_2074,N_3713);
or U5769 (N_5769,N_2780,N_3859);
or U5770 (N_5770,N_3276,N_2981);
nor U5771 (N_5771,N_2611,N_3795);
and U5772 (N_5772,N_2507,N_2945);
xor U5773 (N_5773,N_2953,N_3612);
and U5774 (N_5774,N_3637,N_3458);
nand U5775 (N_5775,N_2684,N_2029);
nor U5776 (N_5776,N_2062,N_3966);
nor U5777 (N_5777,N_3155,N_3010);
xnor U5778 (N_5778,N_3380,N_2995);
nor U5779 (N_5779,N_2741,N_3842);
xnor U5780 (N_5780,N_3915,N_2802);
nand U5781 (N_5781,N_2808,N_3399);
and U5782 (N_5782,N_3735,N_3370);
nor U5783 (N_5783,N_2603,N_3224);
nor U5784 (N_5784,N_3121,N_2651);
and U5785 (N_5785,N_3297,N_3246);
or U5786 (N_5786,N_2083,N_3026);
nor U5787 (N_5787,N_2821,N_3747);
nor U5788 (N_5788,N_2873,N_2338);
or U5789 (N_5789,N_2292,N_3950);
nand U5790 (N_5790,N_3307,N_3871);
or U5791 (N_5791,N_3122,N_2359);
xnor U5792 (N_5792,N_3898,N_3968);
and U5793 (N_5793,N_2241,N_3013);
nand U5794 (N_5794,N_2035,N_2429);
nand U5795 (N_5795,N_3611,N_2027);
xnor U5796 (N_5796,N_2144,N_2925);
nor U5797 (N_5797,N_3032,N_2363);
or U5798 (N_5798,N_3670,N_3874);
nor U5799 (N_5799,N_2870,N_2814);
and U5800 (N_5800,N_2504,N_3100);
nor U5801 (N_5801,N_2365,N_2138);
nand U5802 (N_5802,N_3788,N_3719);
and U5803 (N_5803,N_3243,N_2895);
and U5804 (N_5804,N_2264,N_2336);
xor U5805 (N_5805,N_3689,N_3365);
nand U5806 (N_5806,N_3517,N_2311);
nand U5807 (N_5807,N_2928,N_2657);
nor U5808 (N_5808,N_2787,N_3882);
xor U5809 (N_5809,N_2920,N_2959);
or U5810 (N_5810,N_3450,N_3832);
nor U5811 (N_5811,N_3979,N_3363);
and U5812 (N_5812,N_3175,N_3218);
xnor U5813 (N_5813,N_2543,N_2261);
nor U5814 (N_5814,N_3706,N_2762);
and U5815 (N_5815,N_3523,N_2755);
xor U5816 (N_5816,N_3860,N_3251);
nand U5817 (N_5817,N_2041,N_2087);
nand U5818 (N_5818,N_2944,N_3995);
xor U5819 (N_5819,N_2693,N_3792);
nand U5820 (N_5820,N_3101,N_2675);
or U5821 (N_5821,N_3503,N_2599);
nand U5822 (N_5822,N_2003,N_2805);
xnor U5823 (N_5823,N_3462,N_3306);
or U5824 (N_5824,N_3043,N_2296);
nor U5825 (N_5825,N_3538,N_2054);
and U5826 (N_5826,N_2562,N_3209);
nor U5827 (N_5827,N_2961,N_3055);
and U5828 (N_5828,N_2743,N_3167);
nand U5829 (N_5829,N_2953,N_2726);
and U5830 (N_5830,N_3835,N_3616);
and U5831 (N_5831,N_3215,N_3188);
nor U5832 (N_5832,N_2549,N_3893);
and U5833 (N_5833,N_3282,N_3956);
nand U5834 (N_5834,N_3317,N_2233);
nor U5835 (N_5835,N_3768,N_3037);
nor U5836 (N_5836,N_2645,N_3636);
xor U5837 (N_5837,N_3362,N_3288);
and U5838 (N_5838,N_3928,N_3866);
or U5839 (N_5839,N_3536,N_2406);
or U5840 (N_5840,N_3301,N_3350);
nor U5841 (N_5841,N_2113,N_3848);
nor U5842 (N_5842,N_3851,N_2878);
nor U5843 (N_5843,N_3853,N_2756);
xnor U5844 (N_5844,N_2863,N_2742);
and U5845 (N_5845,N_2471,N_2835);
xor U5846 (N_5846,N_3571,N_2327);
and U5847 (N_5847,N_3221,N_3977);
or U5848 (N_5848,N_2589,N_2362);
xor U5849 (N_5849,N_2659,N_3642);
nand U5850 (N_5850,N_3042,N_3318);
nand U5851 (N_5851,N_2634,N_2740);
or U5852 (N_5852,N_3354,N_3685);
and U5853 (N_5853,N_2984,N_3285);
nand U5854 (N_5854,N_3330,N_3149);
nor U5855 (N_5855,N_2307,N_2303);
nand U5856 (N_5856,N_3562,N_3153);
or U5857 (N_5857,N_3263,N_2321);
nor U5858 (N_5858,N_2439,N_3118);
xnor U5859 (N_5859,N_2522,N_3786);
nor U5860 (N_5860,N_3761,N_3601);
and U5861 (N_5861,N_2096,N_2178);
nor U5862 (N_5862,N_3096,N_3792);
nand U5863 (N_5863,N_3600,N_3246);
nor U5864 (N_5864,N_3601,N_2323);
nand U5865 (N_5865,N_3956,N_3303);
or U5866 (N_5866,N_2295,N_3264);
nand U5867 (N_5867,N_2940,N_2436);
and U5868 (N_5868,N_2050,N_2145);
nor U5869 (N_5869,N_3417,N_3541);
xor U5870 (N_5870,N_3909,N_3505);
xor U5871 (N_5871,N_2943,N_3831);
xnor U5872 (N_5872,N_3083,N_2631);
and U5873 (N_5873,N_3305,N_2306);
nor U5874 (N_5874,N_3035,N_2898);
xor U5875 (N_5875,N_2845,N_3361);
or U5876 (N_5876,N_2621,N_3614);
nand U5877 (N_5877,N_2721,N_2122);
nand U5878 (N_5878,N_3885,N_2914);
and U5879 (N_5879,N_2333,N_3666);
xor U5880 (N_5880,N_2563,N_3553);
nor U5881 (N_5881,N_2028,N_3307);
or U5882 (N_5882,N_3806,N_3006);
nand U5883 (N_5883,N_3560,N_3482);
and U5884 (N_5884,N_2941,N_3836);
xnor U5885 (N_5885,N_2792,N_3130);
nand U5886 (N_5886,N_2774,N_2642);
nor U5887 (N_5887,N_2388,N_3102);
nor U5888 (N_5888,N_2851,N_2324);
and U5889 (N_5889,N_2911,N_2437);
xnor U5890 (N_5890,N_3206,N_3123);
nor U5891 (N_5891,N_3656,N_3039);
or U5892 (N_5892,N_2308,N_2871);
and U5893 (N_5893,N_2266,N_2584);
and U5894 (N_5894,N_2518,N_2143);
xnor U5895 (N_5895,N_2000,N_3407);
nand U5896 (N_5896,N_3530,N_3791);
xnor U5897 (N_5897,N_2876,N_3410);
nand U5898 (N_5898,N_2382,N_3596);
or U5899 (N_5899,N_3306,N_3934);
xnor U5900 (N_5900,N_3652,N_2120);
nand U5901 (N_5901,N_2743,N_2434);
nand U5902 (N_5902,N_3429,N_2237);
nor U5903 (N_5903,N_3353,N_3143);
nand U5904 (N_5904,N_3617,N_2756);
nor U5905 (N_5905,N_3580,N_2488);
nand U5906 (N_5906,N_2366,N_2189);
nor U5907 (N_5907,N_3761,N_3176);
nand U5908 (N_5908,N_2329,N_3254);
or U5909 (N_5909,N_3966,N_2206);
nand U5910 (N_5910,N_3769,N_3007);
xor U5911 (N_5911,N_3879,N_3006);
nor U5912 (N_5912,N_2380,N_2268);
and U5913 (N_5913,N_3138,N_2974);
nand U5914 (N_5914,N_3338,N_3297);
or U5915 (N_5915,N_3079,N_3189);
nand U5916 (N_5916,N_2844,N_3052);
nand U5917 (N_5917,N_2594,N_2493);
xor U5918 (N_5918,N_3292,N_2099);
nor U5919 (N_5919,N_2624,N_3145);
nor U5920 (N_5920,N_3105,N_3593);
xnor U5921 (N_5921,N_2054,N_2779);
nor U5922 (N_5922,N_3928,N_2481);
and U5923 (N_5923,N_2657,N_3985);
xnor U5924 (N_5924,N_3190,N_3135);
nor U5925 (N_5925,N_2636,N_2905);
xnor U5926 (N_5926,N_3638,N_3368);
nor U5927 (N_5927,N_3245,N_2914);
or U5928 (N_5928,N_3429,N_2454);
or U5929 (N_5929,N_3863,N_3459);
nand U5930 (N_5930,N_2920,N_3580);
nand U5931 (N_5931,N_2383,N_2906);
and U5932 (N_5932,N_3875,N_3937);
or U5933 (N_5933,N_3447,N_2916);
nor U5934 (N_5934,N_3653,N_3904);
or U5935 (N_5935,N_3541,N_2158);
or U5936 (N_5936,N_3843,N_2386);
nand U5937 (N_5937,N_2858,N_3155);
xor U5938 (N_5938,N_2950,N_3113);
nor U5939 (N_5939,N_3959,N_2879);
and U5940 (N_5940,N_2349,N_3691);
xnor U5941 (N_5941,N_3598,N_2580);
xor U5942 (N_5942,N_2818,N_2815);
xor U5943 (N_5943,N_3556,N_3892);
xnor U5944 (N_5944,N_3518,N_3473);
nand U5945 (N_5945,N_3852,N_2930);
xnor U5946 (N_5946,N_3657,N_2847);
nand U5947 (N_5947,N_3697,N_2639);
nor U5948 (N_5948,N_3328,N_2444);
nand U5949 (N_5949,N_3931,N_2577);
nand U5950 (N_5950,N_2734,N_2021);
nor U5951 (N_5951,N_3814,N_3333);
nand U5952 (N_5952,N_2694,N_3153);
or U5953 (N_5953,N_2352,N_3172);
or U5954 (N_5954,N_3138,N_2349);
xor U5955 (N_5955,N_2993,N_2864);
nor U5956 (N_5956,N_2536,N_2644);
and U5957 (N_5957,N_3313,N_2978);
xnor U5958 (N_5958,N_2346,N_3118);
nand U5959 (N_5959,N_3956,N_2892);
and U5960 (N_5960,N_3670,N_3658);
nand U5961 (N_5961,N_3477,N_3280);
xnor U5962 (N_5962,N_3083,N_2269);
xnor U5963 (N_5963,N_3833,N_3696);
xnor U5964 (N_5964,N_3996,N_3491);
xor U5965 (N_5965,N_2481,N_3916);
xor U5966 (N_5966,N_2304,N_2932);
and U5967 (N_5967,N_2973,N_2786);
nor U5968 (N_5968,N_2374,N_3261);
nor U5969 (N_5969,N_3103,N_3861);
or U5970 (N_5970,N_3683,N_3506);
nand U5971 (N_5971,N_2474,N_3807);
nor U5972 (N_5972,N_3491,N_3898);
and U5973 (N_5973,N_3130,N_3257);
nor U5974 (N_5974,N_2045,N_2625);
and U5975 (N_5975,N_3558,N_3101);
nand U5976 (N_5976,N_2532,N_3589);
nor U5977 (N_5977,N_3909,N_3901);
and U5978 (N_5978,N_3745,N_2034);
nor U5979 (N_5979,N_2293,N_2171);
xnor U5980 (N_5980,N_2550,N_2320);
xor U5981 (N_5981,N_2352,N_3983);
or U5982 (N_5982,N_2052,N_3987);
nor U5983 (N_5983,N_3137,N_2502);
nand U5984 (N_5984,N_2367,N_2202);
nand U5985 (N_5985,N_3839,N_2789);
nand U5986 (N_5986,N_2380,N_3905);
or U5987 (N_5987,N_3621,N_3795);
or U5988 (N_5988,N_2393,N_2112);
xnor U5989 (N_5989,N_2494,N_2075);
nor U5990 (N_5990,N_3774,N_3068);
xnor U5991 (N_5991,N_3857,N_3138);
xnor U5992 (N_5992,N_3874,N_3927);
or U5993 (N_5993,N_2813,N_3683);
xnor U5994 (N_5994,N_2704,N_2111);
or U5995 (N_5995,N_3421,N_2614);
nor U5996 (N_5996,N_3157,N_2856);
nand U5997 (N_5997,N_2258,N_2780);
xor U5998 (N_5998,N_2713,N_3221);
and U5999 (N_5999,N_2771,N_3074);
nor U6000 (N_6000,N_4077,N_4714);
nand U6001 (N_6001,N_5750,N_4720);
or U6002 (N_6002,N_4243,N_5392);
nor U6003 (N_6003,N_5697,N_4986);
and U6004 (N_6004,N_5745,N_4215);
xor U6005 (N_6005,N_4245,N_5652);
nand U6006 (N_6006,N_5643,N_5889);
xnor U6007 (N_6007,N_5154,N_4414);
and U6008 (N_6008,N_5804,N_5007);
xnor U6009 (N_6009,N_5237,N_4502);
or U6010 (N_6010,N_5806,N_4405);
and U6011 (N_6011,N_4708,N_5972);
nand U6012 (N_6012,N_4059,N_5095);
or U6013 (N_6013,N_4134,N_5688);
xnor U6014 (N_6014,N_5408,N_5825);
or U6015 (N_6015,N_5908,N_5214);
and U6016 (N_6016,N_5228,N_5848);
and U6017 (N_6017,N_4854,N_5322);
or U6018 (N_6018,N_5348,N_5204);
xor U6019 (N_6019,N_5560,N_4571);
xnor U6020 (N_6020,N_5937,N_5633);
and U6021 (N_6021,N_4721,N_5160);
and U6022 (N_6022,N_4084,N_4892);
or U6023 (N_6023,N_5919,N_5630);
or U6024 (N_6024,N_4381,N_4881);
nand U6025 (N_6025,N_4840,N_4344);
nand U6026 (N_6026,N_5599,N_5024);
or U6027 (N_6027,N_5159,N_5991);
nand U6028 (N_6028,N_4993,N_4100);
nor U6029 (N_6029,N_4085,N_4334);
nor U6030 (N_6030,N_5453,N_5349);
or U6031 (N_6031,N_4285,N_5274);
xnor U6032 (N_6032,N_4821,N_4333);
nand U6033 (N_6033,N_5608,N_4609);
and U6034 (N_6034,N_5368,N_4107);
nor U6035 (N_6035,N_5865,N_5210);
or U6036 (N_6036,N_4770,N_4110);
or U6037 (N_6037,N_4646,N_4330);
nor U6038 (N_6038,N_5829,N_5696);
xnor U6039 (N_6039,N_5187,N_5715);
nor U6040 (N_6040,N_5665,N_4176);
nor U6041 (N_6041,N_5517,N_4384);
and U6042 (N_6042,N_5259,N_4070);
and U6043 (N_6043,N_5397,N_5583);
and U6044 (N_6044,N_5770,N_4751);
and U6045 (N_6045,N_4675,N_4196);
nand U6046 (N_6046,N_4411,N_5684);
nor U6047 (N_6047,N_4572,N_4471);
and U6048 (N_6048,N_5969,N_4064);
xor U6049 (N_6049,N_5957,N_4999);
and U6050 (N_6050,N_4580,N_5000);
nand U6051 (N_6051,N_4079,N_4331);
nand U6052 (N_6052,N_4387,N_5145);
nand U6053 (N_6053,N_4193,N_4119);
nor U6054 (N_6054,N_4737,N_4113);
nor U6055 (N_6055,N_5317,N_4259);
and U6056 (N_6056,N_5669,N_5768);
and U6057 (N_6057,N_5478,N_4308);
nor U6058 (N_6058,N_4250,N_5335);
nor U6059 (N_6059,N_4928,N_4154);
nand U6060 (N_6060,N_4857,N_4974);
xnor U6061 (N_6061,N_5577,N_4251);
nand U6062 (N_6062,N_5376,N_5078);
nor U6063 (N_6063,N_5915,N_4870);
nor U6064 (N_6064,N_4388,N_4997);
nand U6065 (N_6065,N_4915,N_4212);
nor U6066 (N_6066,N_5749,N_4000);
and U6067 (N_6067,N_4599,N_5133);
or U6068 (N_6068,N_5827,N_4191);
and U6069 (N_6069,N_5814,N_4712);
and U6070 (N_6070,N_4304,N_5138);
xor U6071 (N_6071,N_5288,N_5080);
nand U6072 (N_6072,N_4847,N_4539);
xnor U6073 (N_6073,N_5384,N_5420);
and U6074 (N_6074,N_5999,N_5815);
xnor U6075 (N_6075,N_5115,N_4981);
or U6076 (N_6076,N_4825,N_5977);
nand U6077 (N_6077,N_4172,N_4882);
nor U6078 (N_6078,N_5740,N_5019);
nor U6079 (N_6079,N_5315,N_5193);
xnor U6080 (N_6080,N_5216,N_5811);
nand U6081 (N_6081,N_4978,N_4739);
nand U6082 (N_6082,N_5037,N_4512);
or U6083 (N_6083,N_5600,N_5475);
xnor U6084 (N_6084,N_5620,N_5591);
and U6085 (N_6085,N_4188,N_4375);
xor U6086 (N_6086,N_5785,N_5904);
or U6087 (N_6087,N_4219,N_5757);
or U6088 (N_6088,N_4578,N_5933);
and U6089 (N_6089,N_5986,N_5332);
nand U6090 (N_6090,N_4274,N_5484);
nand U6091 (N_6091,N_4938,N_5916);
nor U6092 (N_6092,N_5661,N_5265);
nand U6093 (N_6093,N_5886,N_4783);
nand U6094 (N_6094,N_5361,N_4643);
nand U6095 (N_6095,N_4433,N_4908);
nor U6096 (N_6096,N_5711,N_4843);
xnor U6097 (N_6097,N_4062,N_4510);
xnor U6098 (N_6098,N_4587,N_4691);
or U6099 (N_6099,N_4164,N_4674);
and U6100 (N_6100,N_5358,N_5639);
or U6101 (N_6101,N_4715,N_5504);
xor U6102 (N_6102,N_4206,N_4836);
and U6103 (N_6103,N_4725,N_5981);
nand U6104 (N_6104,N_4702,N_4701);
xnor U6105 (N_6105,N_5497,N_5895);
nand U6106 (N_6106,N_5402,N_5020);
nand U6107 (N_6107,N_5248,N_5962);
or U6108 (N_6108,N_5920,N_4313);
nor U6109 (N_6109,N_5425,N_5858);
or U6110 (N_6110,N_4902,N_5334);
nor U6111 (N_6111,N_4924,N_4933);
or U6112 (N_6112,N_5628,N_5885);
xnor U6113 (N_6113,N_5911,N_5191);
xnor U6114 (N_6114,N_4228,N_5581);
or U6115 (N_6115,N_5224,N_5374);
nor U6116 (N_6116,N_5735,N_5050);
xor U6117 (N_6117,N_5952,N_4869);
nor U6118 (N_6118,N_5532,N_4929);
and U6119 (N_6119,N_5194,N_4896);
xor U6120 (N_6120,N_4416,N_5081);
xor U6121 (N_6121,N_4782,N_5738);
xnor U6122 (N_6122,N_5030,N_4383);
xnor U6123 (N_6123,N_5130,N_4368);
nor U6124 (N_6124,N_4460,N_5353);
or U6125 (N_6125,N_5968,N_5549);
xnor U6126 (N_6126,N_5192,N_4872);
and U6127 (N_6127,N_5752,N_5671);
or U6128 (N_6128,N_5898,N_4750);
or U6129 (N_6129,N_4067,N_4500);
nand U6130 (N_6130,N_4729,N_4366);
xor U6131 (N_6131,N_4781,N_4014);
or U6132 (N_6132,N_4099,N_4029);
and U6133 (N_6133,N_5277,N_5162);
or U6134 (N_6134,N_5439,N_5647);
nor U6135 (N_6135,N_4994,N_4307);
nand U6136 (N_6136,N_4832,N_5352);
nor U6137 (N_6137,N_4513,N_4830);
and U6138 (N_6138,N_5673,N_5562);
nand U6139 (N_6139,N_5239,N_5843);
or U6140 (N_6140,N_5813,N_5116);
nor U6141 (N_6141,N_4477,N_4867);
nand U6142 (N_6142,N_4422,N_4991);
and U6143 (N_6143,N_5817,N_4657);
xnor U6144 (N_6144,N_5987,N_4948);
xor U6145 (N_6145,N_4306,N_4864);
or U6146 (N_6146,N_5389,N_4287);
and U6147 (N_6147,N_5924,N_4229);
or U6148 (N_6148,N_4822,N_4341);
or U6149 (N_6149,N_4132,N_4158);
nand U6150 (N_6150,N_5294,N_5963);
and U6151 (N_6151,N_5896,N_4579);
and U6152 (N_6152,N_5153,N_5198);
and U6153 (N_6153,N_5642,N_5809);
xnor U6154 (N_6154,N_4470,N_5171);
nand U6155 (N_6155,N_4055,N_4973);
and U6156 (N_6156,N_5627,N_4240);
nand U6157 (N_6157,N_4793,N_5533);
or U6158 (N_6158,N_5270,N_5648);
nand U6159 (N_6159,N_4246,N_4412);
and U6160 (N_6160,N_5687,N_4216);
or U6161 (N_6161,N_4494,N_5452);
or U6162 (N_6162,N_5746,N_4036);
and U6163 (N_6163,N_5047,N_4258);
and U6164 (N_6164,N_4325,N_4849);
xnor U6165 (N_6165,N_4851,N_5939);
nand U6166 (N_6166,N_5728,N_4045);
or U6167 (N_6167,N_4071,N_5824);
or U6168 (N_6168,N_4226,N_5421);
and U6169 (N_6169,N_4311,N_5936);
xnor U6170 (N_6170,N_5427,N_5306);
or U6171 (N_6171,N_5678,N_5956);
nand U6172 (N_6172,N_5150,N_4147);
nand U6173 (N_6173,N_4761,N_4236);
nand U6174 (N_6174,N_5899,N_4249);
nand U6175 (N_6175,N_4338,N_4426);
xnor U6176 (N_6176,N_4631,N_5835);
nand U6177 (N_6177,N_4499,N_4063);
and U6178 (N_6178,N_4142,N_5996);
nand U6179 (N_6179,N_5503,N_4718);
nand U6180 (N_6180,N_4235,N_4069);
nand U6181 (N_6181,N_4976,N_4372);
xnor U6182 (N_6182,N_5207,N_4850);
xor U6183 (N_6183,N_4031,N_5959);
xnor U6184 (N_6184,N_5057,N_4361);
nor U6185 (N_6185,N_4440,N_4231);
and U6186 (N_6186,N_4597,N_4846);
nor U6187 (N_6187,N_4888,N_5670);
or U6188 (N_6188,N_4534,N_4032);
nand U6189 (N_6189,N_4696,N_4545);
or U6190 (N_6190,N_4364,N_5481);
or U6191 (N_6191,N_4875,N_4203);
or U6192 (N_6192,N_4054,N_5831);
xor U6193 (N_6193,N_5052,N_5313);
and U6194 (N_6194,N_5432,N_4151);
or U6195 (N_6195,N_5268,N_5656);
nor U6196 (N_6196,N_5840,N_5174);
xnor U6197 (N_6197,N_4816,N_4495);
or U6198 (N_6198,N_4261,N_5435);
and U6199 (N_6199,N_5685,N_5856);
xnor U6200 (N_6200,N_4607,N_5998);
xnor U6201 (N_6201,N_4509,N_5289);
xnor U6202 (N_6202,N_5531,N_4090);
xnor U6203 (N_6203,N_5488,N_5276);
or U6204 (N_6204,N_5949,N_4410);
and U6205 (N_6205,N_5461,N_4481);
nand U6206 (N_6206,N_4959,N_5424);
or U6207 (N_6207,N_5547,N_5788);
nand U6208 (N_6208,N_5753,N_5651);
nand U6209 (N_6209,N_4883,N_4838);
or U6210 (N_6210,N_5774,N_4027);
xor U6211 (N_6211,N_4967,N_4773);
and U6212 (N_6212,N_5383,N_5255);
nand U6213 (N_6213,N_4379,N_4706);
xor U6214 (N_6214,N_4417,N_5005);
nor U6215 (N_6215,N_4018,N_4536);
nand U6216 (N_6216,N_4957,N_4958);
and U6217 (N_6217,N_5377,N_5028);
xor U6218 (N_6218,N_4903,N_4615);
or U6219 (N_6219,N_4735,N_4394);
and U6220 (N_6220,N_4256,N_5305);
or U6221 (N_6221,N_5017,N_4709);
nor U6222 (N_6222,N_5499,N_4065);
and U6223 (N_6223,N_5181,N_4520);
or U6224 (N_6224,N_4004,N_4995);
nor U6225 (N_6225,N_5658,N_4019);
and U6226 (N_6226,N_4992,N_5645);
and U6227 (N_6227,N_4266,N_4421);
or U6228 (N_6228,N_4874,N_5942);
and U6229 (N_6229,N_4011,N_4068);
nand U6230 (N_6230,N_5786,N_4811);
or U6231 (N_6231,N_4698,N_5211);
xnor U6232 (N_6232,N_5931,N_4605);
nand U6233 (N_6233,N_5448,N_5233);
xnor U6234 (N_6234,N_4588,N_5852);
xor U6235 (N_6235,N_4886,N_4693);
nor U6236 (N_6236,N_4744,N_5505);
and U6237 (N_6237,N_4656,N_4819);
and U6238 (N_6238,N_4804,N_4877);
nor U6239 (N_6239,N_4655,N_4909);
xnor U6240 (N_6240,N_4209,N_5729);
xnor U6241 (N_6241,N_4526,N_4910);
xor U6242 (N_6242,N_4001,N_4893);
nand U6243 (N_6243,N_4121,N_4290);
nand U6244 (N_6244,N_5807,N_4747);
nor U6245 (N_6245,N_5590,N_5818);
nand U6246 (N_6246,N_4669,N_4895);
nand U6247 (N_6247,N_4323,N_5370);
nand U6248 (N_6248,N_5782,N_4469);
nor U6249 (N_6249,N_5482,N_5779);
nand U6250 (N_6250,N_5328,N_5554);
or U6251 (N_6251,N_4767,N_5837);
and U6252 (N_6252,N_5172,N_5287);
and U6253 (N_6253,N_5821,N_5457);
nand U6254 (N_6254,N_5002,N_4452);
nor U6255 (N_6255,N_5579,N_5681);
nand U6256 (N_6256,N_5300,N_5621);
and U6257 (N_6257,N_4522,N_4075);
nand U6258 (N_6258,N_5041,N_5777);
nand U6259 (N_6259,N_4367,N_4097);
nand U6260 (N_6260,N_5797,N_5411);
or U6261 (N_6261,N_4776,N_5367);
nor U6262 (N_6262,N_4941,N_4898);
xor U6263 (N_6263,N_5901,N_5561);
and U6264 (N_6264,N_4146,N_5350);
and U6265 (N_6265,N_5891,N_5597);
nor U6266 (N_6266,N_4982,N_4205);
or U6267 (N_6267,N_5780,N_4566);
xor U6268 (N_6268,N_5704,N_4723);
nor U6269 (N_6269,N_4859,N_4155);
xor U6270 (N_6270,N_5221,N_5739);
nor U6271 (N_6271,N_5379,N_4557);
or U6272 (N_6272,N_4345,N_5928);
or U6273 (N_6273,N_4899,N_4270);
and U6274 (N_6274,N_4565,N_5880);
nand U6275 (N_6275,N_5124,N_4663);
or U6276 (N_6276,N_5003,N_5567);
nand U6277 (N_6277,N_4091,N_4548);
xor U6278 (N_6278,N_4349,N_4803);
xor U6279 (N_6279,N_4006,N_5381);
nor U6280 (N_6280,N_5161,N_4668);
nand U6281 (N_6281,N_5209,N_4519);
and U6282 (N_6282,N_4913,N_4527);
and U6283 (N_6283,N_5553,N_4098);
nor U6284 (N_6284,N_5857,N_5229);
and U6285 (N_6285,N_5096,N_4204);
xnor U6286 (N_6286,N_5612,N_5245);
or U6287 (N_6287,N_5297,N_4862);
xor U6288 (N_6288,N_5853,N_4038);
xnor U6289 (N_6289,N_4983,N_4310);
nand U6290 (N_6290,N_5691,N_5631);
and U6291 (N_6291,N_5909,N_4809);
and U6292 (N_6292,N_5027,N_5613);
or U6293 (N_6293,N_5747,N_4213);
nor U6294 (N_6294,N_4165,N_4596);
nand U6295 (N_6295,N_4966,N_4476);
nand U6296 (N_6296,N_5605,N_5438);
nand U6297 (N_6297,N_5337,N_5065);
nand U6298 (N_6298,N_4074,N_4174);
xnor U6299 (N_6299,N_5012,N_4576);
xnor U6300 (N_6300,N_4745,N_4661);
and U6301 (N_6301,N_5218,N_4128);
nand U6302 (N_6302,N_4234,N_4719);
nand U6303 (N_6303,N_5431,N_4777);
and U6304 (N_6304,N_5066,N_4827);
or U6305 (N_6305,N_5601,N_4629);
xnor U6306 (N_6306,N_5165,N_4582);
xor U6307 (N_6307,N_5296,N_5575);
nand U6308 (N_6308,N_5527,N_5369);
and U6309 (N_6309,N_5925,N_4408);
nand U6310 (N_6310,N_4492,N_5450);
xor U6311 (N_6311,N_5801,N_5698);
and U6312 (N_6312,N_5934,N_4550);
nand U6313 (N_6313,N_4445,N_5536);
nor U6314 (N_6314,N_4732,N_4790);
nand U6315 (N_6315,N_5689,N_4563);
nand U6316 (N_6316,N_5359,N_5323);
or U6317 (N_6317,N_5357,N_5799);
nor U6318 (N_6318,N_4012,N_5246);
and U6319 (N_6319,N_5371,N_5914);
or U6320 (N_6320,N_4806,N_4778);
nor U6321 (N_6321,N_5451,N_5258);
xor U6322 (N_6322,N_4611,N_5314);
nand U6323 (N_6323,N_4736,N_5222);
nand U6324 (N_6324,N_5075,N_5775);
nor U6325 (N_6325,N_5646,N_4309);
nand U6326 (N_6326,N_4096,N_5466);
or U6327 (N_6327,N_5309,N_4278);
nor U6328 (N_6328,N_4224,N_5879);
and U6329 (N_6329,N_5347,N_5208);
or U6330 (N_6330,N_5197,N_5867);
nand U6331 (N_6331,N_5167,N_4552);
xnor U6332 (N_6332,N_4633,N_5176);
xor U6333 (N_6333,N_5113,N_5039);
or U6334 (N_6334,N_4961,N_5311);
nor U6335 (N_6335,N_5304,N_4700);
xor U6336 (N_6336,N_4116,N_5011);
nor U6337 (N_6337,N_5485,N_5913);
or U6338 (N_6338,N_5298,N_4301);
nor U6339 (N_6339,N_5655,N_4644);
and U6340 (N_6340,N_5624,N_4455);
and U6341 (N_6341,N_4123,N_5022);
xor U6342 (N_6342,N_4541,N_4490);
xnor U6343 (N_6343,N_5316,N_4659);
xor U6344 (N_6344,N_4363,N_4517);
nand U6345 (N_6345,N_5189,N_4628);
xor U6346 (N_6346,N_4717,N_4516);
nor U6347 (N_6347,N_5994,N_5773);
xor U6348 (N_6348,N_5226,N_5703);
nand U6349 (N_6349,N_4667,N_5792);
nor U6350 (N_6350,N_5566,N_5812);
and U6351 (N_6351,N_4507,N_4336);
or U6352 (N_6352,N_5892,N_5607);
or U6353 (N_6353,N_5206,N_5573);
nand U6354 (N_6354,N_4370,N_4762);
xor U6355 (N_6355,N_4124,N_4549);
nand U6356 (N_6356,N_5446,N_5091);
nor U6357 (N_6357,N_4501,N_4787);
nor U6358 (N_6358,N_4112,N_5490);
nand U6359 (N_6359,N_5751,N_4262);
xor U6360 (N_6360,N_4451,N_4227);
nand U6361 (N_6361,N_5064,N_5976);
nand U6362 (N_6362,N_4911,N_4662);
nand U6363 (N_6363,N_4242,N_4666);
nand U6364 (N_6364,N_5060,N_4694);
nand U6365 (N_6365,N_4956,N_5135);
and U6366 (N_6366,N_5958,N_4347);
nor U6367 (N_6367,N_5926,N_4211);
or U6368 (N_6368,N_5795,N_4923);
nand U6369 (N_6369,N_5238,N_5708);
and U6370 (N_6370,N_4918,N_5640);
xnor U6371 (N_6371,N_5122,N_5196);
xnor U6372 (N_6372,N_5604,N_5743);
xnor U6373 (N_6373,N_4463,N_4683);
nor U6374 (N_6374,N_4316,N_4194);
or U6375 (N_6375,N_4446,N_5378);
nor U6376 (N_6376,N_4880,N_4185);
nand U6377 (N_6377,N_4380,N_4044);
nand U6378 (N_6378,N_4947,N_4645);
xnor U6379 (N_6379,N_4152,N_5074);
or U6380 (N_6380,N_5049,N_5557);
or U6381 (N_6381,N_5592,N_4727);
or U6382 (N_6382,N_5727,N_4078);
nor U6383 (N_6383,N_5068,N_5111);
nor U6384 (N_6384,N_5516,N_5820);
and U6385 (N_6385,N_5653,N_5940);
xnor U6386 (N_6386,N_4459,N_4214);
nor U6387 (N_6387,N_5705,N_5980);
or U6388 (N_6388,N_5569,N_5292);
or U6389 (N_6389,N_4102,N_5282);
xor U6390 (N_6390,N_5512,N_4493);
or U6391 (N_6391,N_5731,N_5636);
nor U6392 (N_6392,N_5965,N_4855);
or U6393 (N_6393,N_4396,N_4884);
and U6394 (N_6394,N_4041,N_4756);
nor U6395 (N_6395,N_5866,N_4413);
or U6396 (N_6396,N_5458,N_5692);
or U6397 (N_6397,N_4868,N_5103);
nor U6398 (N_6398,N_5252,N_5638);
nand U6399 (N_6399,N_5372,N_5876);
nand U6400 (N_6400,N_5365,N_4429);
or U6401 (N_6401,N_5710,N_4275);
nand U6402 (N_6402,N_4786,N_5400);
xor U6403 (N_6403,N_4448,N_5186);
or U6404 (N_6404,N_4647,N_5834);
or U6405 (N_6405,N_4442,N_4949);
nor U6406 (N_6406,N_4390,N_4104);
and U6407 (N_6407,N_4449,N_5263);
nor U6408 (N_6408,N_4699,N_5230);
xnor U6409 (N_6409,N_5139,N_4178);
or U6410 (N_6410,N_4350,N_5326);
and U6411 (N_6411,N_4286,N_5051);
nor U6412 (N_6412,N_5616,N_4265);
or U6413 (N_6413,N_5542,N_4932);
nand U6414 (N_6414,N_4238,N_4603);
or U6415 (N_6415,N_5444,N_4473);
xor U6416 (N_6416,N_5736,N_5168);
nor U6417 (N_6417,N_4428,N_5870);
nor U6418 (N_6418,N_4374,N_4658);
nor U6419 (N_6419,N_4305,N_5240);
nand U6420 (N_6420,N_4837,N_4207);
xnor U6421 (N_6421,N_4639,N_4444);
or U6422 (N_6422,N_4860,N_5126);
or U6423 (N_6423,N_5844,N_4772);
nor U6424 (N_6424,N_5013,N_4082);
nor U6425 (N_6425,N_5953,N_4312);
or U6426 (N_6426,N_4060,N_4239);
xnor U6427 (N_6427,N_5423,N_5544);
nor U6428 (N_6428,N_5403,N_5734);
or U6429 (N_6429,N_5529,N_5173);
or U6430 (N_6430,N_4766,N_5416);
nand U6431 (N_6431,N_4392,N_5445);
and U6432 (N_6432,N_4889,N_5526);
xnor U6433 (N_6433,N_4759,N_4106);
nor U6434 (N_6434,N_5706,N_4263);
nor U6435 (N_6435,N_5059,N_4438);
nand U6436 (N_6436,N_4641,N_5073);
or U6437 (N_6437,N_5443,N_5395);
and U6438 (N_6438,N_4187,N_5971);
nor U6439 (N_6439,N_4876,N_4201);
or U6440 (N_6440,N_5570,N_4676);
nor U6441 (N_6441,N_5291,N_5278);
nor U6442 (N_6442,N_4020,N_4409);
xor U6443 (N_6443,N_5137,N_5618);
nor U6444 (N_6444,N_4337,N_5893);
or U6445 (N_6445,N_4220,N_5071);
xnor U6446 (N_6446,N_4535,N_4033);
nand U6447 (N_6447,N_5874,N_5143);
xnor U6448 (N_6448,N_4780,N_5872);
nor U6449 (N_6449,N_4475,N_4441);
and U6450 (N_6450,N_4362,N_4556);
nor U6451 (N_6451,N_5412,N_5267);
xnor U6452 (N_6452,N_4017,N_4705);
and U6453 (N_6453,N_4542,N_5295);
xor U6454 (N_6454,N_5548,N_4115);
nand U6455 (N_6455,N_5390,N_4692);
nand U6456 (N_6456,N_5083,N_4002);
xnor U6457 (N_6457,N_4504,N_5580);
nor U6458 (N_6458,N_5816,N_5520);
or U6459 (N_6459,N_4109,N_5941);
or U6460 (N_6460,N_4430,N_4192);
nor U6461 (N_6461,N_5227,N_5823);
xnor U6462 (N_6462,N_4665,N_4515);
xor U6463 (N_6463,N_5063,N_5511);
nand U6464 (N_6464,N_5910,N_4332);
xor U6465 (N_6465,N_4927,N_5978);
nand U6466 (N_6466,N_4007,N_5404);
or U6467 (N_6467,N_5680,N_4703);
or U6468 (N_6468,N_4197,N_5290);
and U6469 (N_6469,N_4671,N_5092);
nor U6470 (N_6470,N_5271,N_4985);
nor U6471 (N_6471,N_4039,N_5929);
or U6472 (N_6472,N_4133,N_5327);
or U6473 (N_6473,N_4606,N_5654);
nand U6474 (N_6474,N_4968,N_5748);
and U6475 (N_6475,N_4752,N_4955);
nor U6476 (N_6476,N_5995,N_5118);
or U6477 (N_6477,N_4291,N_5649);
and U6478 (N_6478,N_5031,N_5576);
xor U6479 (N_6479,N_5422,N_5758);
or U6480 (N_6480,N_4593,N_4105);
nand U6481 (N_6481,N_4839,N_4269);
and U6482 (N_6482,N_5860,N_5225);
or U6483 (N_6483,N_4354,N_5001);
or U6484 (N_6484,N_5521,N_5944);
and U6485 (N_6485,N_5447,N_4688);
and U6486 (N_6486,N_5360,N_4861);
nor U6487 (N_6487,N_5266,N_4389);
nor U6488 (N_6488,N_5563,N_4722);
xor U6489 (N_6489,N_4202,N_5702);
xor U6490 (N_6490,N_4799,N_5574);
nor U6491 (N_6491,N_4051,N_5254);
nand U6492 (N_6492,N_4279,N_4030);
xnor U6493 (N_6493,N_4462,N_5881);
xor U6494 (N_6494,N_4177,N_5720);
nand U6495 (N_6495,N_4126,N_5513);
nand U6496 (N_6496,N_4076,N_4163);
and U6497 (N_6497,N_5722,N_5890);
and U6498 (N_6498,N_4946,N_5343);
or U6499 (N_6499,N_5888,N_5851);
nand U6500 (N_6500,N_5112,N_5293);
nor U6501 (N_6501,N_5179,N_5067);
or U6502 (N_6502,N_5235,N_4061);
nand U6503 (N_6503,N_4586,N_4182);
xnor U6504 (N_6504,N_4798,N_4689);
and U6505 (N_6505,N_5869,N_4900);
nor U6506 (N_6506,N_4682,N_5663);
or U6507 (N_6507,N_4435,N_5528);
nand U6508 (N_6508,N_4025,N_5883);
or U6509 (N_6509,N_5522,N_5993);
xor U6510 (N_6510,N_4150,N_4594);
nor U6511 (N_6511,N_5862,N_5346);
xor U6512 (N_6512,N_4972,N_4088);
or U6513 (N_6513,N_5632,N_4619);
or U6514 (N_6514,N_4358,N_4208);
nor U6515 (N_6515,N_5213,N_4885);
and U6516 (N_6516,N_4942,N_4340);
xor U6517 (N_6517,N_5873,N_4613);
and U6518 (N_6518,N_4555,N_4057);
nor U6519 (N_6519,N_4087,N_5771);
or U6520 (N_6520,N_4289,N_5602);
nand U6521 (N_6521,N_5281,N_5088);
and U6522 (N_6522,N_5518,N_4636);
or U6523 (N_6523,N_5042,N_5543);
nor U6524 (N_6524,N_5641,N_4404);
nor U6525 (N_6525,N_4498,N_5146);
nand U6526 (N_6526,N_5501,N_4797);
or U6527 (N_6527,N_4111,N_4796);
nand U6528 (N_6528,N_4612,N_5107);
and U6529 (N_6529,N_5396,N_5086);
or U6530 (N_6530,N_4034,N_4618);
and U6531 (N_6531,N_4805,N_5810);
nand U6532 (N_6532,N_4093,N_4558);
nor U6533 (N_6533,N_5787,N_4528);
or U6534 (N_6534,N_4858,N_5056);
or U6535 (N_6535,N_4810,N_5912);
nor U6536 (N_6536,N_5538,N_4042);
xor U6537 (N_6537,N_4936,N_4468);
and U6538 (N_6538,N_4385,N_4685);
nand U6539 (N_6539,N_5463,N_4746);
xor U6540 (N_6540,N_5203,N_5690);
or U6541 (N_6541,N_5004,N_4382);
and U6542 (N_6542,N_5657,N_4791);
or U6543 (N_6543,N_5032,N_5033);
nand U6544 (N_6544,N_4268,N_5085);
or U6545 (N_6545,N_4648,N_5790);
nand U6546 (N_6546,N_4485,N_4021);
nor U6547 (N_6547,N_4866,N_4300);
xor U6548 (N_6548,N_5045,N_5307);
nand U6549 (N_6549,N_5125,N_5249);
xnor U6550 (N_6550,N_4232,N_5232);
or U6551 (N_6551,N_4785,N_4543);
nand U6552 (N_6552,N_4346,N_5954);
or U6553 (N_6553,N_5803,N_4189);
nand U6554 (N_6554,N_5855,N_4952);
nor U6555 (N_6555,N_4248,N_4166);
and U6556 (N_6556,N_5410,N_4436);
or U6557 (N_6557,N_4339,N_4028);
or U6558 (N_6558,N_4260,N_4407);
or U6559 (N_6559,N_5540,N_4853);
or U6560 (N_6560,N_4758,N_4393);
or U6561 (N_6561,N_4532,N_4406);
and U6562 (N_6562,N_4963,N_4120);
xnor U6563 (N_6563,N_4118,N_4604);
xnor U6564 (N_6564,N_5719,N_5302);
xnor U6565 (N_6565,N_4775,N_4351);
nor U6566 (N_6566,N_5635,N_5054);
or U6567 (N_6567,N_5283,N_5188);
and U6568 (N_6568,N_4454,N_4590);
nand U6569 (N_6569,N_4904,N_5364);
or U6570 (N_6570,N_4789,N_4939);
nor U6571 (N_6571,N_5426,N_4627);
and U6572 (N_6572,N_5683,N_5626);
or U6573 (N_6573,N_4564,N_5183);
nor U6574 (N_6574,N_5555,N_4420);
nor U6575 (N_6575,N_5498,N_4480);
nor U6576 (N_6576,N_4919,N_5712);
nor U6577 (N_6577,N_4686,N_5878);
or U6578 (N_6578,N_5467,N_4567);
nand U6579 (N_6579,N_5509,N_4733);
nor U6580 (N_6580,N_4402,N_4179);
or U6581 (N_6581,N_5637,N_5175);
nor U6582 (N_6582,N_5982,N_4478);
nand U6583 (N_6583,N_5048,N_4486);
or U6584 (N_6584,N_4769,N_4984);
nor U6585 (N_6585,N_4906,N_5742);
nand U6586 (N_6586,N_5151,N_4049);
nor U6587 (N_6587,N_5340,N_4833);
or U6588 (N_6588,N_4800,N_5725);
nand U6589 (N_6589,N_5955,N_4829);
xor U6590 (N_6590,N_4537,N_4324);
nand U6591 (N_6591,N_4056,N_5975);
or U6592 (N_6592,N_5662,N_5029);
nand U6593 (N_6593,N_4281,N_5262);
xor U6594 (N_6594,N_4386,N_5764);
or U6595 (N_6595,N_5760,N_5945);
nand U6596 (N_6596,N_4716,N_5355);
nand U6597 (N_6597,N_4373,N_5667);
and U6598 (N_6598,N_4755,N_5234);
nor U6599 (N_6599,N_5034,N_4820);
or U6600 (N_6600,N_4740,N_5716);
or U6601 (N_6601,N_5121,N_5483);
nor U6602 (N_6602,N_5487,N_4595);
xor U6603 (N_6603,N_4447,N_5339);
xnor U6604 (N_6604,N_5486,N_4953);
nor U6605 (N_6605,N_4734,N_5303);
or U6606 (N_6606,N_5442,N_4283);
nand U6607 (N_6607,N_5223,N_5784);
nand U6608 (N_6608,N_5260,N_5119);
xor U6609 (N_6609,N_5253,N_4640);
nor U6610 (N_6610,N_4879,N_5470);
nor U6611 (N_6611,N_5084,N_5380);
xor U6612 (N_6612,N_5611,N_5882);
and U6613 (N_6613,N_5756,N_5794);
and U6614 (N_6614,N_5140,N_4273);
and U6615 (N_6615,N_5158,N_4210);
or U6616 (N_6616,N_5109,N_4461);
xnor U6617 (N_6617,N_5619,N_5131);
nand U6618 (N_6618,N_4920,N_4742);
and U6619 (N_6619,N_4905,N_5164);
nor U6620 (N_6620,N_4378,N_5251);
xnor U6621 (N_6621,N_4148,N_5917);
xor U6622 (N_6622,N_4424,N_5184);
nor U6623 (N_6623,N_4602,N_4450);
or U6624 (N_6624,N_4288,N_5822);
nand U6625 (N_6625,N_5796,N_4267);
nor U6626 (N_6626,N_5464,N_5596);
or U6627 (N_6627,N_5104,N_5093);
or U6628 (N_6628,N_5471,N_4774);
nand U6629 (N_6629,N_4419,N_4637);
nand U6630 (N_6630,N_5550,N_4654);
and U6631 (N_6631,N_5247,N_5387);
xor U6632 (N_6632,N_4812,N_4488);
and U6633 (N_6633,N_4848,N_4704);
or U6634 (N_6634,N_4365,N_5718);
nand U6635 (N_6635,N_5850,N_5201);
nand U6636 (N_6636,N_4418,N_4137);
nand U6637 (N_6637,N_5582,N_5375);
and U6638 (N_6638,N_5868,N_4356);
or U6639 (N_6639,N_4546,N_5622);
and U6640 (N_6640,N_4127,N_5894);
nor U6641 (N_6641,N_5556,N_4670);
xor U6642 (N_6642,N_5449,N_5087);
nor U6643 (N_6643,N_5185,N_4951);
or U6644 (N_6644,N_4581,N_5036);
nand U6645 (N_6645,N_4763,N_4293);
or U6646 (N_6646,N_4934,N_4844);
and U6647 (N_6647,N_4022,N_4089);
xnor U6648 (N_6648,N_4965,N_4841);
or U6649 (N_6649,N_4095,N_4856);
nor U6650 (N_6650,N_4760,N_4653);
xor U6651 (N_6651,N_5769,N_5077);
nor U6652 (N_6652,N_5441,N_5391);
xnor U6653 (N_6653,N_4878,N_5331);
xor U6654 (N_6654,N_5589,N_5983);
nor U6655 (N_6655,N_4171,N_5406);
nand U6656 (N_6656,N_5524,N_5310);
nor U6657 (N_6657,N_5922,N_5385);
nor U6658 (N_6658,N_4784,N_4280);
or U6659 (N_6659,N_4253,N_5128);
or U6660 (N_6660,N_5010,N_5587);
and U6661 (N_6661,N_5847,N_5923);
or U6662 (N_6662,N_4523,N_5992);
or U6663 (N_6663,N_5496,N_4748);
xor U6664 (N_6664,N_5462,N_4757);
nor U6665 (N_6665,N_5275,N_4616);
nor U6666 (N_6666,N_5493,N_5166);
nor U6667 (N_6667,N_4035,N_5989);
and U6668 (N_6668,N_4989,N_4794);
nand U6669 (N_6669,N_4254,N_4474);
and U6670 (N_6670,N_4562,N_5826);
nand U6671 (N_6671,N_4945,N_4496);
or U6672 (N_6672,N_4971,N_5755);
nor U6673 (N_6673,N_4255,N_5440);
xnor U6674 (N_6674,N_4753,N_5625);
nand U6675 (N_6675,N_4817,N_4170);
or U6676 (N_6676,N_5997,N_5105);
nor U6677 (N_6677,N_4707,N_5428);
xor U6678 (N_6678,N_4591,N_5921);
or U6679 (N_6679,N_5805,N_5502);
and U6680 (N_6680,N_4970,N_5861);
or U6681 (N_6681,N_5887,N_4458);
and U6682 (N_6682,N_5677,N_4931);
xor U6683 (N_6683,N_5351,N_4195);
or U6684 (N_6684,N_4922,N_4092);
nand U6685 (N_6685,N_4114,N_5329);
or U6686 (N_6686,N_5394,N_4264);
nand U6687 (N_6687,N_4738,N_4353);
or U6688 (N_6688,N_4296,N_5182);
xnor U6689 (N_6689,N_5927,N_4944);
and U6690 (N_6690,N_4431,N_5155);
xnor U6691 (N_6691,N_5243,N_4801);
nand U6692 (N_6692,N_5950,N_4926);
and U6693 (N_6693,N_4013,N_5076);
and U6694 (N_6694,N_4479,N_5301);
nand U6695 (N_6695,N_4620,N_5819);
xor U6696 (N_6696,N_5906,N_4439);
or U6697 (N_6697,N_4538,N_4321);
xnor U6698 (N_6698,N_5800,N_5469);
or U6699 (N_6699,N_5018,N_5132);
nand U6700 (N_6700,N_5568,N_5699);
and U6701 (N_6701,N_5666,N_5284);
or U6702 (N_6702,N_4016,N_4397);
xnor U6703 (N_6703,N_5043,N_5058);
nand U6704 (N_6704,N_5539,N_4140);
or U6705 (N_6705,N_4598,N_5609);
and U6706 (N_6706,N_4108,N_5832);
xnor U6707 (N_6707,N_4181,N_5094);
or U6708 (N_6708,N_4575,N_4962);
xnor U6709 (N_6709,N_4048,N_5286);
nand U6710 (N_6710,N_4271,N_4754);
nor U6711 (N_6711,N_5098,N_5864);
nor U6712 (N_6712,N_4863,N_4401);
xor U6713 (N_6713,N_5798,N_5974);
xor U6714 (N_6714,N_5279,N_5675);
nand U6715 (N_6715,N_4651,N_5021);
nor U6716 (N_6716,N_5008,N_5772);
nand U6717 (N_6717,N_4257,N_4200);
nor U6718 (N_6718,N_5215,N_5717);
nor U6719 (N_6719,N_5016,N_5269);
xnor U6720 (N_6720,N_4135,N_4037);
nor U6721 (N_6721,N_5460,N_5783);
xor U6722 (N_6722,N_5617,N_5157);
and U6723 (N_6723,N_5127,N_5778);
or U6724 (N_6724,N_5754,N_4153);
xor U6725 (N_6725,N_4186,N_4570);
xor U6726 (N_6726,N_5430,N_5407);
xor U6727 (N_6727,N_5101,N_4871);
nor U6728 (N_6728,N_4072,N_5664);
xor U6729 (N_6729,N_5744,N_5897);
nor U6730 (N_6730,N_5090,N_5195);
xnor U6731 (N_6731,N_4680,N_4621);
xor U6732 (N_6732,N_5454,N_4466);
or U6733 (N_6733,N_4771,N_4937);
and U6734 (N_6734,N_5495,N_5551);
or U6735 (N_6735,N_5902,N_5436);
xor U6736 (N_6736,N_5659,N_5741);
and U6737 (N_6737,N_5110,N_5943);
and U6738 (N_6738,N_5836,N_4327);
xnor U6739 (N_6739,N_5615,N_5414);
and U6740 (N_6740,N_4980,N_4765);
xnor U6741 (N_6741,N_4489,N_5136);
nor U6742 (N_6742,N_4295,N_5985);
or U6743 (N_6743,N_4533,N_4518);
nor U6744 (N_6744,N_4907,N_5634);
or U6745 (N_6745,N_4834,N_5900);
or U6746 (N_6746,N_4073,N_5961);
nand U6747 (N_6747,N_5723,N_5776);
and U6748 (N_6748,N_5530,N_5242);
xor U6749 (N_6749,N_5951,N_4979);
or U6750 (N_6750,N_4890,N_4342);
nor U6751 (N_6751,N_4943,N_4823);
nor U6752 (N_6752,N_4162,N_5676);
xnor U6753 (N_6753,N_5948,N_4230);
xor U6754 (N_6754,N_4415,N_5219);
or U6755 (N_6755,N_5593,N_5062);
or U6756 (N_6756,N_5877,N_4503);
and U6757 (N_6757,N_4569,N_5767);
nand U6758 (N_6758,N_4282,N_4531);
nand U6759 (N_6759,N_5660,N_4672);
xor U6760 (N_6760,N_4139,N_4568);
nor U6761 (N_6761,N_5413,N_5356);
nand U6762 (N_6762,N_4617,N_4554);
nand U6763 (N_6763,N_5409,N_5578);
and U6764 (N_6764,N_5236,N_4852);
and U6765 (N_6765,N_5415,N_4247);
nand U6766 (N_6766,N_4094,N_4329);
or U6767 (N_6767,N_4768,N_5833);
nand U6768 (N_6768,N_4005,N_5713);
xor U6769 (N_6769,N_5838,N_5344);
or U6770 (N_6770,N_5319,N_4318);
xor U6771 (N_6771,N_4136,N_4749);
and U6772 (N_6772,N_5828,N_5546);
and U6773 (N_6773,N_4058,N_4403);
nand U6774 (N_6774,N_4925,N_5733);
nand U6775 (N_6775,N_5584,N_4547);
nor U6776 (N_6776,N_4015,N_5152);
and U6777 (N_6777,N_5644,N_4432);
xor U6778 (N_6778,N_5730,N_4614);
and U6779 (N_6779,N_5506,N_4277);
nand U6780 (N_6780,N_4818,N_5148);
nand U6781 (N_6781,N_4487,N_5695);
xor U6782 (N_6782,N_5134,N_4505);
and U6783 (N_6783,N_4726,N_4690);
xor U6784 (N_6784,N_5988,N_5875);
nor U6785 (N_6785,N_5545,N_5177);
and U6786 (N_6786,N_4315,N_5061);
and U6787 (N_6787,N_5973,N_5465);
nand U6788 (N_6788,N_4988,N_4660);
nand U6789 (N_6789,N_5672,N_5761);
and U6790 (N_6790,N_5565,N_4141);
and U6791 (N_6791,N_5217,N_4472);
xor U6792 (N_6792,N_5724,N_5342);
or U6793 (N_6793,N_4199,N_4464);
nor U6794 (N_6794,N_5594,N_5040);
nor U6795 (N_6795,N_5802,N_4710);
nand U6796 (N_6796,N_5079,N_5871);
xor U6797 (N_6797,N_5863,N_5534);
nor U6798 (N_6798,N_5362,N_4053);
and U6799 (N_6799,N_4156,N_5257);
nor U6800 (N_6800,N_4678,N_5363);
nand U6801 (N_6801,N_5964,N_4930);
nand U6802 (N_6802,N_5072,N_4457);
and U6803 (N_6803,N_4317,N_4608);
nor U6804 (N_6804,N_4623,N_4831);
nand U6805 (N_6805,N_5038,N_4292);
or U6806 (N_6806,N_5845,N_4921);
or U6807 (N_6807,N_4491,N_5070);
or U6808 (N_6808,N_4437,N_4456);
nand U6809 (N_6809,N_4551,N_5009);
xnor U6810 (N_6810,N_5984,N_4369);
nor U6811 (N_6811,N_4573,N_4625);
nor U6812 (N_6812,N_4023,N_5102);
xor U6813 (N_6813,N_5437,N_5726);
xnor U6814 (N_6814,N_4788,N_5682);
xor U6815 (N_6815,N_4497,N_5737);
and U6816 (N_6816,N_4086,N_4314);
and U6817 (N_6817,N_4183,N_5241);
nand U6818 (N_6818,N_5250,N_4009);
nand U6819 (N_6819,N_5333,N_4168);
nand U6820 (N_6820,N_5354,N_5603);
and U6821 (N_6821,N_5839,N_4894);
nand U6822 (N_6822,N_4996,N_5299);
nor U6823 (N_6823,N_4241,N_4008);
or U6824 (N_6824,N_5510,N_5679);
nand U6825 (N_6825,N_4355,N_4225);
or U6826 (N_6826,N_5433,N_4376);
xor U6827 (N_6827,N_5559,N_5564);
nor U6828 (N_6828,N_4521,N_5935);
or U6829 (N_6829,N_4377,N_5330);
and U6830 (N_6830,N_5830,N_5169);
and U6831 (N_6831,N_5552,N_4807);
xnor U6832 (N_6832,N_5123,N_4695);
nand U6833 (N_6833,N_4423,N_5586);
nand U6834 (N_6834,N_5614,N_4559);
nand U6835 (N_6835,N_4326,N_4328);
xor U6836 (N_6836,N_5100,N_4184);
or U6837 (N_6837,N_4352,N_4711);
nor U6838 (N_6838,N_4360,N_5523);
nor U6839 (N_6839,N_5500,N_5763);
xnor U6840 (N_6840,N_4730,N_4815);
xor U6841 (N_6841,N_5714,N_4540);
or U6842 (N_6842,N_4252,N_5459);
and U6843 (N_6843,N_5280,N_5244);
nor U6844 (N_6844,N_5709,N_4835);
and U6845 (N_6845,N_4465,N_5494);
xor U6846 (N_6846,N_4052,N_4960);
xnor U6847 (N_6847,N_4684,N_5338);
xor U6848 (N_6848,N_4222,N_5114);
nor U6849 (N_6849,N_4335,N_4322);
or U6850 (N_6850,N_5932,N_5854);
nor U6851 (N_6851,N_4160,N_4395);
and U6852 (N_6852,N_5907,N_4138);
nor U6853 (N_6853,N_5572,N_4359);
and U6854 (N_6854,N_5474,N_5595);
or U6855 (N_6855,N_4131,N_5382);
nand U6856 (N_6856,N_4357,N_4244);
or U6857 (N_6857,N_5859,N_4427);
and U6858 (N_6858,N_4897,N_5129);
xor U6859 (N_6859,N_4302,N_4144);
or U6860 (N_6860,N_4887,N_4294);
xnor U6861 (N_6861,N_5142,N_4975);
or U6862 (N_6862,N_4010,N_5492);
nand U6863 (N_6863,N_4802,N_4122);
and U6864 (N_6864,N_4145,N_4391);
or U6865 (N_6865,N_5508,N_5212);
nor U6866 (N_6866,N_4845,N_4987);
nor U6867 (N_6867,N_4650,N_5588);
and U6868 (N_6868,N_5884,N_5419);
and U6869 (N_6869,N_5418,N_4600);
xnor U6870 (N_6870,N_5650,N_5515);
xnor U6871 (N_6871,N_4741,N_4320);
nor U6872 (N_6872,N_4434,N_5960);
nand U6873 (N_6873,N_4198,N_4217);
xor U6874 (N_6874,N_5082,N_5674);
xnor U6875 (N_6875,N_5842,N_4814);
or U6876 (N_6876,N_4221,N_5366);
and U6877 (N_6877,N_4398,N_5220);
and U6878 (N_6878,N_5808,N_5434);
nor U6879 (N_6879,N_4977,N_4561);
nand U6880 (N_6880,N_4940,N_5200);
xnor U6881 (N_6881,N_5537,N_5015);
and U6882 (N_6882,N_5149,N_5399);
xnor U6883 (N_6883,N_5558,N_5629);
xnor U6884 (N_6884,N_4484,N_4681);
and U6885 (N_6885,N_5507,N_4634);
nand U6886 (N_6886,N_5905,N_4917);
nand U6887 (N_6887,N_5841,N_5272);
xnor U6888 (N_6888,N_4083,N_5312);
nand U6889 (N_6889,N_4525,N_4601);
and U6890 (N_6890,N_5035,N_4237);
nand U6891 (N_6891,N_5393,N_4592);
and U6892 (N_6892,N_5765,N_4964);
and U6893 (N_6893,N_4808,N_5261);
nor U6894 (N_6894,N_5525,N_4348);
and U6895 (N_6895,N_4129,N_5721);
nor U6896 (N_6896,N_5701,N_4443);
nand U6897 (N_6897,N_4159,N_4003);
xnor U6898 (N_6898,N_5489,N_4622);
xor U6899 (N_6899,N_5141,N_5006);
nand U6900 (N_6900,N_5325,N_4664);
or U6901 (N_6901,N_4585,N_4914);
or U6902 (N_6902,N_5762,N_4233);
xnor U6903 (N_6903,N_5069,N_4161);
or U6904 (N_6904,N_4916,N_4514);
xnor U6905 (N_6905,N_4792,N_5273);
nor U6906 (N_6906,N_4024,N_4284);
nor U6907 (N_6907,N_4117,N_5623);
xnor U6908 (N_6908,N_5264,N_4080);
or U6909 (N_6909,N_5585,N_5456);
xor U6910 (N_6910,N_5766,N_5256);
and U6911 (N_6911,N_4697,N_5781);
or U6912 (N_6912,N_5700,N_4276);
or U6913 (N_6913,N_5946,N_4299);
xor U6914 (N_6914,N_4584,N_5930);
xnor U6915 (N_6915,N_5535,N_5341);
xor U6916 (N_6916,N_4632,N_5791);
and U6917 (N_6917,N_5429,N_4954);
or U6918 (N_6918,N_4272,N_5202);
or U6919 (N_6919,N_4589,N_5903);
nor U6920 (N_6920,N_5732,N_5938);
and U6921 (N_6921,N_5401,N_4713);
and U6922 (N_6922,N_4677,N_4652);
nor U6923 (N_6923,N_5147,N_4130);
nor U6924 (N_6924,N_4046,N_5398);
or U6925 (N_6925,N_5231,N_4679);
and U6926 (N_6926,N_5308,N_4583);
nand U6927 (N_6927,N_5759,N_4143);
or U6928 (N_6928,N_4298,N_4731);
or U6929 (N_6929,N_4103,N_5846);
nand U6930 (N_6930,N_5044,N_5694);
nor U6931 (N_6931,N_5023,N_5966);
xor U6932 (N_6932,N_4673,N_5793);
xor U6933 (N_6933,N_4050,N_4218);
nand U6934 (N_6934,N_4610,N_4813);
and U6935 (N_6935,N_5707,N_4865);
and U6936 (N_6936,N_4649,N_4901);
xor U6937 (N_6937,N_4047,N_5089);
or U6938 (N_6938,N_5190,N_5373);
or U6939 (N_6939,N_5318,N_5668);
and U6940 (N_6940,N_5480,N_4912);
or U6941 (N_6941,N_5472,N_4467);
nor U6942 (N_6942,N_5686,N_4826);
or U6943 (N_6943,N_5099,N_5386);
or U6944 (N_6944,N_4998,N_4969);
or U6945 (N_6945,N_5117,N_5606);
and U6946 (N_6946,N_5026,N_4040);
xnor U6947 (N_6947,N_5345,N_5476);
or U6948 (N_6948,N_5170,N_4626);
and U6949 (N_6949,N_5947,N_5144);
nor U6950 (N_6950,N_5336,N_4425);
and U6951 (N_6951,N_5055,N_5320);
xor U6952 (N_6952,N_4190,N_4764);
or U6953 (N_6953,N_5046,N_5473);
nor U6954 (N_6954,N_5405,N_4453);
xor U6955 (N_6955,N_5967,N_4482);
and U6956 (N_6956,N_4223,N_4169);
xnor U6957 (N_6957,N_4950,N_5285);
or U6958 (N_6958,N_5468,N_4125);
or U6959 (N_6959,N_4935,N_5571);
xnor U6960 (N_6960,N_4624,N_4026);
xnor U6961 (N_6961,N_4180,N_5477);
or U6962 (N_6962,N_4297,N_4319);
xor U6963 (N_6963,N_4101,N_4399);
nand U6964 (N_6964,N_4066,N_5180);
and U6965 (N_6965,N_5163,N_4524);
nor U6966 (N_6966,N_4483,N_4157);
and U6967 (N_6967,N_4642,N_4724);
xor U6968 (N_6968,N_4687,N_5455);
nand U6969 (N_6969,N_4630,N_4828);
nor U6970 (N_6970,N_4173,N_5097);
nand U6971 (N_6971,N_4043,N_4167);
nand U6972 (N_6972,N_5178,N_5610);
and U6973 (N_6973,N_4149,N_5789);
and U6974 (N_6974,N_4728,N_5053);
xor U6975 (N_6975,N_4081,N_4303);
and U6976 (N_6976,N_5990,N_5514);
xnor U6977 (N_6977,N_5205,N_4574);
and U6978 (N_6978,N_5199,N_5979);
nand U6979 (N_6979,N_4508,N_4795);
xor U6980 (N_6980,N_4175,N_4544);
nor U6981 (N_6981,N_5014,N_4506);
or U6982 (N_6982,N_4891,N_4343);
or U6983 (N_6983,N_5120,N_5598);
xnor U6984 (N_6984,N_5108,N_4577);
and U6985 (N_6985,N_5324,N_4990);
nor U6986 (N_6986,N_4638,N_4824);
or U6987 (N_6987,N_5918,N_4842);
xnor U6988 (N_6988,N_4400,N_4635);
xnor U6989 (N_6989,N_4553,N_5479);
nand U6990 (N_6990,N_5388,N_5849);
nand U6991 (N_6991,N_5156,N_5519);
or U6992 (N_6992,N_4743,N_4779);
and U6993 (N_6993,N_4530,N_5025);
nor U6994 (N_6994,N_5970,N_4560);
xnor U6995 (N_6995,N_5106,N_5321);
and U6996 (N_6996,N_4371,N_5491);
nand U6997 (N_6997,N_4873,N_4511);
or U6998 (N_6998,N_4529,N_5417);
or U6999 (N_6999,N_5541,N_5693);
nand U7000 (N_7000,N_5262,N_4107);
nand U7001 (N_7001,N_5037,N_5267);
nor U7002 (N_7002,N_5248,N_5595);
nand U7003 (N_7003,N_5871,N_4608);
and U7004 (N_7004,N_5846,N_5713);
nand U7005 (N_7005,N_4648,N_4640);
nor U7006 (N_7006,N_5651,N_4671);
nand U7007 (N_7007,N_4000,N_4885);
and U7008 (N_7008,N_4220,N_4445);
xnor U7009 (N_7009,N_5785,N_4853);
and U7010 (N_7010,N_5808,N_4944);
and U7011 (N_7011,N_4836,N_4389);
or U7012 (N_7012,N_4452,N_4590);
nand U7013 (N_7013,N_5738,N_5796);
xnor U7014 (N_7014,N_4140,N_5826);
and U7015 (N_7015,N_4751,N_5576);
or U7016 (N_7016,N_4512,N_4042);
or U7017 (N_7017,N_5480,N_5504);
nor U7018 (N_7018,N_5185,N_5354);
nor U7019 (N_7019,N_4744,N_5460);
nand U7020 (N_7020,N_4555,N_4274);
or U7021 (N_7021,N_4983,N_5895);
xor U7022 (N_7022,N_4131,N_5338);
nand U7023 (N_7023,N_4308,N_4285);
or U7024 (N_7024,N_4151,N_5141);
or U7025 (N_7025,N_4817,N_4359);
nor U7026 (N_7026,N_4702,N_4450);
and U7027 (N_7027,N_4512,N_4889);
nor U7028 (N_7028,N_5216,N_4506);
nand U7029 (N_7029,N_5840,N_5695);
nand U7030 (N_7030,N_4340,N_4965);
xor U7031 (N_7031,N_5953,N_5653);
and U7032 (N_7032,N_4710,N_4725);
nand U7033 (N_7033,N_4788,N_4944);
nand U7034 (N_7034,N_4776,N_5109);
nand U7035 (N_7035,N_4303,N_4528);
or U7036 (N_7036,N_4703,N_4599);
nor U7037 (N_7037,N_4019,N_5725);
or U7038 (N_7038,N_5038,N_4791);
xnor U7039 (N_7039,N_4022,N_4736);
or U7040 (N_7040,N_5155,N_4280);
nor U7041 (N_7041,N_4078,N_4525);
xor U7042 (N_7042,N_4413,N_4116);
and U7043 (N_7043,N_4064,N_4867);
nand U7044 (N_7044,N_5358,N_4880);
and U7045 (N_7045,N_4293,N_4746);
xor U7046 (N_7046,N_4813,N_4258);
nor U7047 (N_7047,N_4367,N_5449);
xnor U7048 (N_7048,N_4725,N_4357);
nor U7049 (N_7049,N_5800,N_5528);
xnor U7050 (N_7050,N_4657,N_5458);
xnor U7051 (N_7051,N_5836,N_5191);
or U7052 (N_7052,N_5423,N_4882);
xnor U7053 (N_7053,N_5273,N_5119);
nor U7054 (N_7054,N_5278,N_4974);
or U7055 (N_7055,N_4870,N_5883);
xor U7056 (N_7056,N_4407,N_5848);
nor U7057 (N_7057,N_5788,N_5953);
nand U7058 (N_7058,N_5916,N_5047);
and U7059 (N_7059,N_4248,N_5477);
nand U7060 (N_7060,N_4345,N_4568);
or U7061 (N_7061,N_5102,N_4739);
nand U7062 (N_7062,N_4634,N_5776);
nand U7063 (N_7063,N_4530,N_4535);
nand U7064 (N_7064,N_5146,N_5427);
xnor U7065 (N_7065,N_5447,N_4101);
nand U7066 (N_7066,N_5974,N_4572);
nor U7067 (N_7067,N_5390,N_5985);
xor U7068 (N_7068,N_5957,N_5409);
or U7069 (N_7069,N_4767,N_5594);
xnor U7070 (N_7070,N_4049,N_4011);
nor U7071 (N_7071,N_5749,N_4010);
and U7072 (N_7072,N_4172,N_5900);
and U7073 (N_7073,N_4475,N_5177);
nor U7074 (N_7074,N_5343,N_4056);
nor U7075 (N_7075,N_4193,N_5463);
and U7076 (N_7076,N_4876,N_4828);
nand U7077 (N_7077,N_5725,N_4571);
nor U7078 (N_7078,N_4261,N_5911);
or U7079 (N_7079,N_5436,N_4004);
or U7080 (N_7080,N_4635,N_5892);
xnor U7081 (N_7081,N_5973,N_4662);
or U7082 (N_7082,N_5391,N_5687);
xnor U7083 (N_7083,N_5275,N_5496);
nor U7084 (N_7084,N_5464,N_5399);
xnor U7085 (N_7085,N_5688,N_4955);
xor U7086 (N_7086,N_4657,N_4194);
nand U7087 (N_7087,N_5237,N_5260);
and U7088 (N_7088,N_5194,N_5904);
nor U7089 (N_7089,N_5595,N_4447);
nand U7090 (N_7090,N_5223,N_4810);
xor U7091 (N_7091,N_5724,N_5463);
and U7092 (N_7092,N_4694,N_5336);
or U7093 (N_7093,N_5995,N_4588);
xnor U7094 (N_7094,N_5684,N_5780);
and U7095 (N_7095,N_4694,N_5644);
nor U7096 (N_7096,N_5221,N_4098);
or U7097 (N_7097,N_5386,N_5026);
and U7098 (N_7098,N_5841,N_5045);
xnor U7099 (N_7099,N_4724,N_4124);
nand U7100 (N_7100,N_4240,N_4718);
nor U7101 (N_7101,N_4298,N_5971);
nand U7102 (N_7102,N_5948,N_4852);
nand U7103 (N_7103,N_4328,N_5344);
nor U7104 (N_7104,N_4242,N_5167);
xor U7105 (N_7105,N_4774,N_4919);
or U7106 (N_7106,N_5467,N_5534);
and U7107 (N_7107,N_5604,N_5725);
and U7108 (N_7108,N_5211,N_5584);
xnor U7109 (N_7109,N_5849,N_4551);
nor U7110 (N_7110,N_4640,N_4761);
xnor U7111 (N_7111,N_4341,N_4896);
or U7112 (N_7112,N_4199,N_5580);
nand U7113 (N_7113,N_4297,N_4101);
and U7114 (N_7114,N_4168,N_5832);
xnor U7115 (N_7115,N_5564,N_5745);
nand U7116 (N_7116,N_5192,N_5128);
or U7117 (N_7117,N_5340,N_5647);
and U7118 (N_7118,N_4147,N_5923);
or U7119 (N_7119,N_4322,N_4553);
nand U7120 (N_7120,N_5840,N_4047);
xnor U7121 (N_7121,N_4444,N_4963);
nand U7122 (N_7122,N_4719,N_4429);
xor U7123 (N_7123,N_4572,N_5636);
and U7124 (N_7124,N_4259,N_5744);
xor U7125 (N_7125,N_5353,N_4922);
nor U7126 (N_7126,N_4503,N_4120);
or U7127 (N_7127,N_5209,N_5188);
and U7128 (N_7128,N_4849,N_5393);
nand U7129 (N_7129,N_4813,N_5522);
and U7130 (N_7130,N_5485,N_4925);
and U7131 (N_7131,N_4561,N_4754);
or U7132 (N_7132,N_5002,N_4165);
or U7133 (N_7133,N_4881,N_5647);
and U7134 (N_7134,N_5099,N_4511);
nor U7135 (N_7135,N_5962,N_5154);
and U7136 (N_7136,N_5391,N_4197);
nor U7137 (N_7137,N_4129,N_5882);
xor U7138 (N_7138,N_4596,N_4845);
nor U7139 (N_7139,N_4640,N_4823);
xnor U7140 (N_7140,N_4530,N_5821);
and U7141 (N_7141,N_4952,N_5281);
nor U7142 (N_7142,N_4693,N_4229);
nand U7143 (N_7143,N_4367,N_4160);
or U7144 (N_7144,N_4628,N_4895);
nor U7145 (N_7145,N_4472,N_5753);
nor U7146 (N_7146,N_5751,N_4188);
xnor U7147 (N_7147,N_4853,N_5816);
or U7148 (N_7148,N_4408,N_4150);
and U7149 (N_7149,N_4540,N_5734);
or U7150 (N_7150,N_4270,N_4108);
nor U7151 (N_7151,N_5316,N_4939);
or U7152 (N_7152,N_4718,N_5568);
nand U7153 (N_7153,N_5792,N_5513);
nor U7154 (N_7154,N_5334,N_4183);
nand U7155 (N_7155,N_4828,N_5412);
or U7156 (N_7156,N_4532,N_5630);
xnor U7157 (N_7157,N_5702,N_4852);
nand U7158 (N_7158,N_4295,N_4699);
xor U7159 (N_7159,N_5744,N_5005);
nand U7160 (N_7160,N_4231,N_4636);
or U7161 (N_7161,N_5037,N_5088);
xor U7162 (N_7162,N_4205,N_4921);
nor U7163 (N_7163,N_5661,N_5335);
and U7164 (N_7164,N_5773,N_5744);
or U7165 (N_7165,N_4979,N_4311);
nor U7166 (N_7166,N_5166,N_5045);
nand U7167 (N_7167,N_5628,N_4292);
nor U7168 (N_7168,N_5607,N_5380);
or U7169 (N_7169,N_4673,N_5788);
nor U7170 (N_7170,N_4377,N_4572);
xor U7171 (N_7171,N_4098,N_4564);
xnor U7172 (N_7172,N_5359,N_4230);
and U7173 (N_7173,N_5476,N_5378);
nor U7174 (N_7174,N_4382,N_5329);
xor U7175 (N_7175,N_5140,N_4952);
and U7176 (N_7176,N_5411,N_5739);
nor U7177 (N_7177,N_4394,N_5477);
xnor U7178 (N_7178,N_4249,N_5797);
nand U7179 (N_7179,N_4934,N_4564);
or U7180 (N_7180,N_5462,N_5537);
nand U7181 (N_7181,N_5428,N_4872);
xnor U7182 (N_7182,N_5074,N_5223);
xor U7183 (N_7183,N_4664,N_4465);
and U7184 (N_7184,N_5305,N_5479);
and U7185 (N_7185,N_5364,N_4562);
nand U7186 (N_7186,N_4887,N_4682);
or U7187 (N_7187,N_4724,N_4050);
or U7188 (N_7188,N_4635,N_5640);
nand U7189 (N_7189,N_4393,N_4859);
nand U7190 (N_7190,N_4428,N_5228);
nor U7191 (N_7191,N_5013,N_4904);
nor U7192 (N_7192,N_5231,N_5588);
xnor U7193 (N_7193,N_5883,N_5471);
nand U7194 (N_7194,N_5202,N_4760);
and U7195 (N_7195,N_4867,N_5426);
and U7196 (N_7196,N_4452,N_5261);
nand U7197 (N_7197,N_4492,N_5477);
xor U7198 (N_7198,N_4871,N_5079);
and U7199 (N_7199,N_4738,N_5542);
xor U7200 (N_7200,N_5659,N_5982);
nand U7201 (N_7201,N_5403,N_4290);
nand U7202 (N_7202,N_5175,N_4486);
or U7203 (N_7203,N_5662,N_5533);
and U7204 (N_7204,N_4351,N_4142);
nor U7205 (N_7205,N_5875,N_4901);
xor U7206 (N_7206,N_5793,N_5407);
and U7207 (N_7207,N_4541,N_4267);
xor U7208 (N_7208,N_5597,N_4969);
nor U7209 (N_7209,N_5037,N_4269);
and U7210 (N_7210,N_4351,N_5277);
and U7211 (N_7211,N_4741,N_4482);
and U7212 (N_7212,N_5184,N_4689);
and U7213 (N_7213,N_4618,N_5456);
and U7214 (N_7214,N_5489,N_5626);
and U7215 (N_7215,N_4018,N_4319);
xor U7216 (N_7216,N_5937,N_4033);
or U7217 (N_7217,N_5570,N_4034);
nor U7218 (N_7218,N_5030,N_4957);
xnor U7219 (N_7219,N_4981,N_5327);
and U7220 (N_7220,N_5234,N_4749);
xor U7221 (N_7221,N_5629,N_5006);
and U7222 (N_7222,N_4174,N_5275);
nand U7223 (N_7223,N_4192,N_5279);
or U7224 (N_7224,N_4629,N_4288);
or U7225 (N_7225,N_4427,N_5512);
nand U7226 (N_7226,N_4560,N_4697);
xnor U7227 (N_7227,N_4057,N_5998);
or U7228 (N_7228,N_4285,N_5343);
nand U7229 (N_7229,N_5564,N_5103);
nand U7230 (N_7230,N_5776,N_5811);
and U7231 (N_7231,N_4085,N_5691);
nor U7232 (N_7232,N_5742,N_4005);
or U7233 (N_7233,N_5486,N_4755);
xnor U7234 (N_7234,N_5730,N_4402);
nand U7235 (N_7235,N_5347,N_5979);
nor U7236 (N_7236,N_5902,N_4084);
and U7237 (N_7237,N_5265,N_5057);
and U7238 (N_7238,N_5766,N_5651);
nand U7239 (N_7239,N_4774,N_5566);
xnor U7240 (N_7240,N_5441,N_5108);
and U7241 (N_7241,N_4910,N_4882);
nor U7242 (N_7242,N_5111,N_4625);
nand U7243 (N_7243,N_5300,N_4816);
or U7244 (N_7244,N_5648,N_5362);
or U7245 (N_7245,N_5361,N_5375);
or U7246 (N_7246,N_5828,N_5371);
and U7247 (N_7247,N_5797,N_5912);
or U7248 (N_7248,N_4393,N_4582);
nor U7249 (N_7249,N_4562,N_4453);
xnor U7250 (N_7250,N_4095,N_5744);
nand U7251 (N_7251,N_4958,N_4808);
and U7252 (N_7252,N_4863,N_4335);
nor U7253 (N_7253,N_4424,N_5714);
or U7254 (N_7254,N_5299,N_4755);
or U7255 (N_7255,N_4821,N_4881);
and U7256 (N_7256,N_4329,N_4706);
nand U7257 (N_7257,N_4573,N_4714);
nand U7258 (N_7258,N_5140,N_5022);
xnor U7259 (N_7259,N_4460,N_4920);
or U7260 (N_7260,N_5088,N_5365);
nand U7261 (N_7261,N_5320,N_4723);
nor U7262 (N_7262,N_5455,N_5800);
nor U7263 (N_7263,N_5529,N_5878);
nand U7264 (N_7264,N_4215,N_4555);
and U7265 (N_7265,N_5703,N_4733);
xnor U7266 (N_7266,N_5083,N_4181);
xnor U7267 (N_7267,N_4538,N_4413);
or U7268 (N_7268,N_4916,N_5350);
or U7269 (N_7269,N_4943,N_4653);
nor U7270 (N_7270,N_5697,N_5876);
xor U7271 (N_7271,N_4309,N_5081);
xor U7272 (N_7272,N_4194,N_4779);
or U7273 (N_7273,N_5966,N_5381);
and U7274 (N_7274,N_4326,N_4338);
nor U7275 (N_7275,N_5977,N_4770);
xor U7276 (N_7276,N_4470,N_4852);
xor U7277 (N_7277,N_4086,N_4652);
or U7278 (N_7278,N_4572,N_5303);
xor U7279 (N_7279,N_5438,N_4768);
nand U7280 (N_7280,N_5615,N_4220);
and U7281 (N_7281,N_5969,N_4206);
and U7282 (N_7282,N_5460,N_5664);
and U7283 (N_7283,N_4230,N_5230);
nand U7284 (N_7284,N_5402,N_4420);
nand U7285 (N_7285,N_4593,N_5426);
nor U7286 (N_7286,N_5184,N_5350);
nand U7287 (N_7287,N_4072,N_5277);
or U7288 (N_7288,N_4533,N_5975);
nand U7289 (N_7289,N_4789,N_5938);
nor U7290 (N_7290,N_4970,N_5961);
nand U7291 (N_7291,N_4738,N_4344);
and U7292 (N_7292,N_5867,N_4885);
nand U7293 (N_7293,N_5551,N_5460);
and U7294 (N_7294,N_5506,N_5052);
nand U7295 (N_7295,N_5765,N_5282);
xor U7296 (N_7296,N_5776,N_5351);
and U7297 (N_7297,N_4920,N_5772);
xnor U7298 (N_7298,N_4943,N_4421);
nand U7299 (N_7299,N_5033,N_4416);
nor U7300 (N_7300,N_4243,N_4614);
or U7301 (N_7301,N_5430,N_4634);
nand U7302 (N_7302,N_5674,N_5353);
nand U7303 (N_7303,N_5927,N_4273);
and U7304 (N_7304,N_4361,N_5276);
nor U7305 (N_7305,N_5262,N_4284);
nor U7306 (N_7306,N_4631,N_4190);
xor U7307 (N_7307,N_4546,N_5769);
nand U7308 (N_7308,N_5897,N_4348);
nand U7309 (N_7309,N_5876,N_4349);
nand U7310 (N_7310,N_5873,N_4008);
and U7311 (N_7311,N_5371,N_5392);
nor U7312 (N_7312,N_4416,N_4504);
nand U7313 (N_7313,N_4678,N_5718);
and U7314 (N_7314,N_4616,N_5610);
nor U7315 (N_7315,N_4284,N_4191);
nor U7316 (N_7316,N_5470,N_5669);
xor U7317 (N_7317,N_4447,N_5282);
xnor U7318 (N_7318,N_4443,N_4554);
or U7319 (N_7319,N_5013,N_5405);
nor U7320 (N_7320,N_5130,N_5611);
or U7321 (N_7321,N_4630,N_4783);
and U7322 (N_7322,N_4635,N_5106);
nor U7323 (N_7323,N_4785,N_4674);
and U7324 (N_7324,N_4907,N_5751);
nand U7325 (N_7325,N_4194,N_4966);
and U7326 (N_7326,N_5435,N_4941);
or U7327 (N_7327,N_4742,N_4709);
xor U7328 (N_7328,N_4967,N_4972);
and U7329 (N_7329,N_5226,N_5068);
nor U7330 (N_7330,N_5038,N_5102);
or U7331 (N_7331,N_4484,N_4125);
xor U7332 (N_7332,N_4583,N_5187);
xor U7333 (N_7333,N_5226,N_4968);
xnor U7334 (N_7334,N_4874,N_4178);
nor U7335 (N_7335,N_4267,N_4657);
nor U7336 (N_7336,N_5881,N_5630);
nand U7337 (N_7337,N_4225,N_4223);
nor U7338 (N_7338,N_4107,N_5078);
or U7339 (N_7339,N_4686,N_5355);
xor U7340 (N_7340,N_4690,N_5351);
and U7341 (N_7341,N_5067,N_5352);
xor U7342 (N_7342,N_4440,N_5056);
and U7343 (N_7343,N_4783,N_4613);
and U7344 (N_7344,N_4955,N_4915);
and U7345 (N_7345,N_4716,N_5056);
nand U7346 (N_7346,N_4211,N_4119);
and U7347 (N_7347,N_4777,N_5700);
nand U7348 (N_7348,N_4132,N_5811);
or U7349 (N_7349,N_4807,N_4456);
and U7350 (N_7350,N_4000,N_4661);
nand U7351 (N_7351,N_5531,N_5661);
xnor U7352 (N_7352,N_5273,N_5070);
xnor U7353 (N_7353,N_4250,N_5634);
nand U7354 (N_7354,N_5890,N_5699);
nand U7355 (N_7355,N_4133,N_5642);
or U7356 (N_7356,N_4963,N_4111);
xor U7357 (N_7357,N_5059,N_4511);
nand U7358 (N_7358,N_4033,N_5123);
nand U7359 (N_7359,N_5933,N_5899);
nor U7360 (N_7360,N_4791,N_4532);
nand U7361 (N_7361,N_5902,N_5466);
and U7362 (N_7362,N_5259,N_5507);
nor U7363 (N_7363,N_5324,N_4815);
nand U7364 (N_7364,N_4243,N_5483);
and U7365 (N_7365,N_5274,N_5293);
nor U7366 (N_7366,N_5671,N_4620);
nor U7367 (N_7367,N_5351,N_5975);
and U7368 (N_7368,N_4506,N_4132);
xor U7369 (N_7369,N_5007,N_5129);
nor U7370 (N_7370,N_4906,N_5197);
or U7371 (N_7371,N_5477,N_5994);
nand U7372 (N_7372,N_4053,N_5170);
xor U7373 (N_7373,N_4275,N_5929);
and U7374 (N_7374,N_4117,N_4502);
nor U7375 (N_7375,N_5535,N_4298);
and U7376 (N_7376,N_4835,N_5924);
or U7377 (N_7377,N_5467,N_5506);
nor U7378 (N_7378,N_4274,N_5856);
xor U7379 (N_7379,N_4378,N_4054);
xnor U7380 (N_7380,N_5926,N_4974);
nand U7381 (N_7381,N_4091,N_5551);
or U7382 (N_7382,N_5023,N_4876);
and U7383 (N_7383,N_4741,N_4141);
or U7384 (N_7384,N_4073,N_4639);
or U7385 (N_7385,N_5484,N_5503);
nor U7386 (N_7386,N_4557,N_5824);
nor U7387 (N_7387,N_5036,N_4192);
and U7388 (N_7388,N_4326,N_5178);
nand U7389 (N_7389,N_5582,N_4199);
nor U7390 (N_7390,N_4023,N_5348);
or U7391 (N_7391,N_5612,N_5379);
nand U7392 (N_7392,N_5029,N_5138);
nor U7393 (N_7393,N_5042,N_4206);
nor U7394 (N_7394,N_4295,N_5106);
nor U7395 (N_7395,N_5847,N_5167);
nor U7396 (N_7396,N_4357,N_4159);
and U7397 (N_7397,N_4831,N_4441);
nor U7398 (N_7398,N_5209,N_5719);
nor U7399 (N_7399,N_4310,N_4997);
xnor U7400 (N_7400,N_4660,N_4356);
or U7401 (N_7401,N_4242,N_5959);
nand U7402 (N_7402,N_4406,N_5941);
or U7403 (N_7403,N_5986,N_4180);
xor U7404 (N_7404,N_5019,N_4842);
and U7405 (N_7405,N_5670,N_5146);
xnor U7406 (N_7406,N_5225,N_5589);
nand U7407 (N_7407,N_5846,N_4600);
nor U7408 (N_7408,N_4193,N_4843);
or U7409 (N_7409,N_4515,N_4305);
and U7410 (N_7410,N_5399,N_4659);
xnor U7411 (N_7411,N_4811,N_5780);
or U7412 (N_7412,N_5191,N_4427);
xor U7413 (N_7413,N_5514,N_5014);
nor U7414 (N_7414,N_4729,N_5154);
xnor U7415 (N_7415,N_4986,N_5916);
and U7416 (N_7416,N_5109,N_5384);
or U7417 (N_7417,N_4327,N_5240);
nor U7418 (N_7418,N_4846,N_5626);
xnor U7419 (N_7419,N_5866,N_4703);
xor U7420 (N_7420,N_5257,N_5600);
and U7421 (N_7421,N_5135,N_4403);
xnor U7422 (N_7422,N_5894,N_4850);
nand U7423 (N_7423,N_4863,N_4484);
nand U7424 (N_7424,N_5047,N_4145);
and U7425 (N_7425,N_4672,N_5268);
nor U7426 (N_7426,N_5621,N_5529);
and U7427 (N_7427,N_4806,N_4980);
xnor U7428 (N_7428,N_4016,N_4627);
and U7429 (N_7429,N_5930,N_5088);
and U7430 (N_7430,N_4028,N_4931);
xnor U7431 (N_7431,N_4736,N_4527);
or U7432 (N_7432,N_4681,N_5147);
and U7433 (N_7433,N_4763,N_4804);
nor U7434 (N_7434,N_5203,N_4037);
xnor U7435 (N_7435,N_4302,N_4127);
nand U7436 (N_7436,N_4865,N_4933);
and U7437 (N_7437,N_4602,N_4180);
and U7438 (N_7438,N_5874,N_5897);
nor U7439 (N_7439,N_4242,N_4913);
nand U7440 (N_7440,N_4106,N_5023);
or U7441 (N_7441,N_5219,N_4379);
xnor U7442 (N_7442,N_5963,N_5639);
or U7443 (N_7443,N_4522,N_4341);
and U7444 (N_7444,N_5644,N_5767);
xor U7445 (N_7445,N_5718,N_4732);
xor U7446 (N_7446,N_5030,N_4986);
and U7447 (N_7447,N_5516,N_4030);
nand U7448 (N_7448,N_5686,N_4636);
nand U7449 (N_7449,N_4264,N_4877);
nor U7450 (N_7450,N_5173,N_5596);
nor U7451 (N_7451,N_4554,N_5509);
nor U7452 (N_7452,N_4920,N_4975);
or U7453 (N_7453,N_4315,N_4265);
nand U7454 (N_7454,N_4624,N_4788);
nand U7455 (N_7455,N_5710,N_4633);
xnor U7456 (N_7456,N_4678,N_4993);
or U7457 (N_7457,N_4723,N_5286);
nand U7458 (N_7458,N_4551,N_4465);
or U7459 (N_7459,N_4118,N_5719);
xnor U7460 (N_7460,N_5730,N_4512);
and U7461 (N_7461,N_5599,N_5518);
nor U7462 (N_7462,N_4287,N_4696);
xor U7463 (N_7463,N_4015,N_4142);
xor U7464 (N_7464,N_4302,N_5446);
and U7465 (N_7465,N_4131,N_4340);
and U7466 (N_7466,N_5751,N_5738);
and U7467 (N_7467,N_4695,N_5016);
and U7468 (N_7468,N_5487,N_4518);
nand U7469 (N_7469,N_4528,N_4369);
or U7470 (N_7470,N_4969,N_4277);
nand U7471 (N_7471,N_5552,N_5848);
and U7472 (N_7472,N_4758,N_5964);
nand U7473 (N_7473,N_4744,N_4423);
xor U7474 (N_7474,N_5195,N_4766);
xor U7475 (N_7475,N_4648,N_4898);
xor U7476 (N_7476,N_4629,N_4611);
and U7477 (N_7477,N_4115,N_4890);
nand U7478 (N_7478,N_4824,N_5000);
xnor U7479 (N_7479,N_5116,N_4486);
nor U7480 (N_7480,N_5529,N_5535);
nor U7481 (N_7481,N_4766,N_5730);
or U7482 (N_7482,N_5804,N_5018);
nand U7483 (N_7483,N_4019,N_5260);
xnor U7484 (N_7484,N_4312,N_4849);
or U7485 (N_7485,N_4246,N_4865);
nand U7486 (N_7486,N_5110,N_4064);
and U7487 (N_7487,N_5483,N_4520);
xor U7488 (N_7488,N_4516,N_5301);
or U7489 (N_7489,N_5601,N_4093);
and U7490 (N_7490,N_4247,N_5786);
nand U7491 (N_7491,N_5795,N_4217);
nand U7492 (N_7492,N_4736,N_4490);
xnor U7493 (N_7493,N_4492,N_5200);
nand U7494 (N_7494,N_4074,N_4884);
nor U7495 (N_7495,N_5388,N_4545);
and U7496 (N_7496,N_5638,N_5173);
xnor U7497 (N_7497,N_4629,N_4107);
nor U7498 (N_7498,N_5378,N_4679);
or U7499 (N_7499,N_4308,N_5220);
and U7500 (N_7500,N_5381,N_5425);
and U7501 (N_7501,N_5215,N_4508);
nor U7502 (N_7502,N_5425,N_4316);
or U7503 (N_7503,N_5055,N_5340);
nand U7504 (N_7504,N_5083,N_5117);
nand U7505 (N_7505,N_4450,N_5779);
or U7506 (N_7506,N_4373,N_5786);
xor U7507 (N_7507,N_4762,N_5991);
or U7508 (N_7508,N_4474,N_5325);
and U7509 (N_7509,N_5350,N_5848);
nor U7510 (N_7510,N_5376,N_4931);
or U7511 (N_7511,N_4706,N_5872);
and U7512 (N_7512,N_5681,N_4314);
and U7513 (N_7513,N_4544,N_5249);
nand U7514 (N_7514,N_5875,N_5795);
or U7515 (N_7515,N_4074,N_4835);
or U7516 (N_7516,N_5523,N_5316);
and U7517 (N_7517,N_5903,N_4932);
xnor U7518 (N_7518,N_5980,N_4963);
or U7519 (N_7519,N_4424,N_4736);
xor U7520 (N_7520,N_5630,N_5615);
nor U7521 (N_7521,N_5186,N_4151);
nand U7522 (N_7522,N_4060,N_5053);
or U7523 (N_7523,N_5458,N_4269);
and U7524 (N_7524,N_5580,N_5451);
and U7525 (N_7525,N_4692,N_5750);
or U7526 (N_7526,N_4262,N_4604);
xor U7527 (N_7527,N_5237,N_5361);
or U7528 (N_7528,N_5938,N_4044);
xnor U7529 (N_7529,N_5434,N_4489);
xor U7530 (N_7530,N_5473,N_5581);
nor U7531 (N_7531,N_4110,N_4932);
nand U7532 (N_7532,N_5600,N_4467);
and U7533 (N_7533,N_5662,N_4276);
nor U7534 (N_7534,N_4723,N_5256);
xnor U7535 (N_7535,N_5886,N_5761);
or U7536 (N_7536,N_4208,N_5085);
and U7537 (N_7537,N_4845,N_5281);
or U7538 (N_7538,N_5198,N_5358);
xnor U7539 (N_7539,N_4536,N_4306);
xor U7540 (N_7540,N_5063,N_4245);
xnor U7541 (N_7541,N_4555,N_4353);
nor U7542 (N_7542,N_4817,N_4994);
and U7543 (N_7543,N_5318,N_4335);
and U7544 (N_7544,N_5823,N_5369);
nor U7545 (N_7545,N_5470,N_5787);
and U7546 (N_7546,N_5907,N_4715);
xor U7547 (N_7547,N_4162,N_4245);
or U7548 (N_7548,N_4001,N_5827);
nor U7549 (N_7549,N_4162,N_5338);
xor U7550 (N_7550,N_4968,N_4581);
xnor U7551 (N_7551,N_5548,N_5374);
xnor U7552 (N_7552,N_4778,N_4037);
or U7553 (N_7553,N_4197,N_4595);
nor U7554 (N_7554,N_5480,N_5718);
nor U7555 (N_7555,N_5462,N_4894);
and U7556 (N_7556,N_4389,N_5015);
nor U7557 (N_7557,N_5933,N_4142);
and U7558 (N_7558,N_4139,N_4465);
and U7559 (N_7559,N_5342,N_4071);
xnor U7560 (N_7560,N_5511,N_4238);
nor U7561 (N_7561,N_5945,N_5229);
or U7562 (N_7562,N_4612,N_4725);
or U7563 (N_7563,N_4411,N_4366);
nand U7564 (N_7564,N_5925,N_5514);
or U7565 (N_7565,N_4188,N_5074);
xor U7566 (N_7566,N_4076,N_5761);
and U7567 (N_7567,N_5189,N_5253);
xnor U7568 (N_7568,N_5640,N_4315);
or U7569 (N_7569,N_5084,N_4521);
xnor U7570 (N_7570,N_4959,N_4519);
nor U7571 (N_7571,N_5050,N_5570);
nand U7572 (N_7572,N_4720,N_5258);
nor U7573 (N_7573,N_4208,N_4113);
or U7574 (N_7574,N_4622,N_4439);
and U7575 (N_7575,N_4632,N_4495);
xor U7576 (N_7576,N_4012,N_5324);
nand U7577 (N_7577,N_4346,N_4157);
xnor U7578 (N_7578,N_4955,N_4125);
xor U7579 (N_7579,N_5242,N_4439);
or U7580 (N_7580,N_4244,N_4654);
or U7581 (N_7581,N_5696,N_5312);
xnor U7582 (N_7582,N_5912,N_5411);
nand U7583 (N_7583,N_4265,N_5063);
nand U7584 (N_7584,N_5145,N_4632);
and U7585 (N_7585,N_5206,N_5296);
and U7586 (N_7586,N_4910,N_4620);
and U7587 (N_7587,N_4190,N_4375);
nor U7588 (N_7588,N_4399,N_5961);
or U7589 (N_7589,N_4561,N_4687);
or U7590 (N_7590,N_5305,N_5044);
xor U7591 (N_7591,N_5706,N_4384);
xor U7592 (N_7592,N_4836,N_5653);
xnor U7593 (N_7593,N_5798,N_4336);
and U7594 (N_7594,N_5467,N_5083);
and U7595 (N_7595,N_4293,N_4902);
xor U7596 (N_7596,N_4429,N_5697);
nand U7597 (N_7597,N_4441,N_5526);
xnor U7598 (N_7598,N_4895,N_5681);
nor U7599 (N_7599,N_4837,N_4224);
nand U7600 (N_7600,N_4354,N_5194);
nand U7601 (N_7601,N_4849,N_4550);
and U7602 (N_7602,N_5342,N_5660);
and U7603 (N_7603,N_4730,N_5620);
or U7604 (N_7604,N_4795,N_4714);
nand U7605 (N_7605,N_5599,N_4965);
and U7606 (N_7606,N_4466,N_5182);
xor U7607 (N_7607,N_4967,N_4371);
nor U7608 (N_7608,N_5553,N_5675);
or U7609 (N_7609,N_5916,N_5029);
xnor U7610 (N_7610,N_5371,N_5083);
xnor U7611 (N_7611,N_5268,N_5183);
nor U7612 (N_7612,N_4707,N_5373);
or U7613 (N_7613,N_4163,N_5254);
nor U7614 (N_7614,N_4407,N_4908);
and U7615 (N_7615,N_5077,N_4102);
nor U7616 (N_7616,N_4973,N_5074);
nand U7617 (N_7617,N_5107,N_4279);
nor U7618 (N_7618,N_4706,N_4000);
and U7619 (N_7619,N_5630,N_5584);
nor U7620 (N_7620,N_5442,N_5229);
or U7621 (N_7621,N_4686,N_5175);
xnor U7622 (N_7622,N_4243,N_4712);
nor U7623 (N_7623,N_4222,N_5158);
xnor U7624 (N_7624,N_5603,N_4867);
or U7625 (N_7625,N_4848,N_4214);
and U7626 (N_7626,N_5431,N_4468);
or U7627 (N_7627,N_4400,N_4389);
or U7628 (N_7628,N_4407,N_5537);
or U7629 (N_7629,N_4061,N_4446);
or U7630 (N_7630,N_5860,N_5261);
or U7631 (N_7631,N_5228,N_5384);
or U7632 (N_7632,N_5110,N_4592);
xnor U7633 (N_7633,N_4451,N_5046);
or U7634 (N_7634,N_5598,N_5961);
nor U7635 (N_7635,N_5513,N_5223);
xnor U7636 (N_7636,N_5784,N_4783);
nor U7637 (N_7637,N_5358,N_5007);
or U7638 (N_7638,N_4376,N_5386);
nand U7639 (N_7639,N_4896,N_5524);
xor U7640 (N_7640,N_5810,N_4508);
and U7641 (N_7641,N_4551,N_5338);
xnor U7642 (N_7642,N_4458,N_4165);
nor U7643 (N_7643,N_4669,N_4784);
nor U7644 (N_7644,N_5356,N_4975);
and U7645 (N_7645,N_5258,N_5443);
nand U7646 (N_7646,N_5820,N_4329);
and U7647 (N_7647,N_5975,N_4103);
nor U7648 (N_7648,N_5894,N_5432);
or U7649 (N_7649,N_4691,N_4938);
or U7650 (N_7650,N_5006,N_4768);
nor U7651 (N_7651,N_4341,N_5789);
or U7652 (N_7652,N_5349,N_4548);
or U7653 (N_7653,N_4132,N_5568);
and U7654 (N_7654,N_4441,N_4616);
nand U7655 (N_7655,N_5287,N_4458);
or U7656 (N_7656,N_4022,N_5683);
or U7657 (N_7657,N_4031,N_4109);
xnor U7658 (N_7658,N_5631,N_4378);
xor U7659 (N_7659,N_5628,N_4384);
nand U7660 (N_7660,N_5929,N_5694);
nand U7661 (N_7661,N_4313,N_4400);
or U7662 (N_7662,N_5230,N_4843);
xnor U7663 (N_7663,N_5114,N_5253);
nor U7664 (N_7664,N_5597,N_4598);
nand U7665 (N_7665,N_5264,N_4372);
or U7666 (N_7666,N_4603,N_4322);
or U7667 (N_7667,N_5940,N_4978);
or U7668 (N_7668,N_4647,N_4382);
and U7669 (N_7669,N_4909,N_4721);
or U7670 (N_7670,N_4087,N_4960);
xor U7671 (N_7671,N_5035,N_5825);
nand U7672 (N_7672,N_5902,N_5673);
xor U7673 (N_7673,N_5655,N_4904);
nand U7674 (N_7674,N_5558,N_4965);
nor U7675 (N_7675,N_4421,N_5378);
xnor U7676 (N_7676,N_4565,N_5963);
nor U7677 (N_7677,N_4046,N_4209);
nor U7678 (N_7678,N_5179,N_5923);
nand U7679 (N_7679,N_5643,N_5740);
or U7680 (N_7680,N_4777,N_4072);
and U7681 (N_7681,N_5823,N_5421);
nor U7682 (N_7682,N_5617,N_4320);
or U7683 (N_7683,N_5679,N_4356);
xnor U7684 (N_7684,N_5027,N_5926);
nand U7685 (N_7685,N_4839,N_5535);
and U7686 (N_7686,N_4305,N_5425);
nor U7687 (N_7687,N_5270,N_4139);
nand U7688 (N_7688,N_5301,N_4831);
nand U7689 (N_7689,N_5763,N_5653);
xor U7690 (N_7690,N_4837,N_5559);
or U7691 (N_7691,N_5297,N_5214);
nor U7692 (N_7692,N_4490,N_5902);
or U7693 (N_7693,N_5851,N_4287);
nor U7694 (N_7694,N_4664,N_4730);
or U7695 (N_7695,N_5164,N_4246);
nand U7696 (N_7696,N_5219,N_4457);
and U7697 (N_7697,N_5529,N_4894);
nand U7698 (N_7698,N_4409,N_4399);
or U7699 (N_7699,N_5252,N_5789);
nand U7700 (N_7700,N_4417,N_4663);
nand U7701 (N_7701,N_5049,N_5903);
nor U7702 (N_7702,N_4431,N_5173);
and U7703 (N_7703,N_5789,N_5499);
xnor U7704 (N_7704,N_4215,N_4109);
nor U7705 (N_7705,N_5136,N_4231);
or U7706 (N_7706,N_5791,N_4295);
xnor U7707 (N_7707,N_4673,N_5372);
xor U7708 (N_7708,N_4288,N_4776);
xor U7709 (N_7709,N_4804,N_5671);
nand U7710 (N_7710,N_5056,N_5617);
and U7711 (N_7711,N_5080,N_5626);
xnor U7712 (N_7712,N_4513,N_4866);
nor U7713 (N_7713,N_5848,N_4204);
nor U7714 (N_7714,N_5533,N_4760);
nand U7715 (N_7715,N_5735,N_4950);
and U7716 (N_7716,N_4260,N_5580);
nor U7717 (N_7717,N_4838,N_4311);
nor U7718 (N_7718,N_4020,N_4563);
and U7719 (N_7719,N_4548,N_4781);
nor U7720 (N_7720,N_4357,N_4458);
nand U7721 (N_7721,N_4857,N_5802);
or U7722 (N_7722,N_4546,N_5112);
and U7723 (N_7723,N_5068,N_4383);
nor U7724 (N_7724,N_4112,N_5449);
and U7725 (N_7725,N_4647,N_4587);
or U7726 (N_7726,N_5856,N_4895);
nor U7727 (N_7727,N_4000,N_5972);
and U7728 (N_7728,N_4254,N_5164);
xor U7729 (N_7729,N_5393,N_4782);
or U7730 (N_7730,N_4354,N_5826);
and U7731 (N_7731,N_4852,N_4248);
nand U7732 (N_7732,N_4434,N_5503);
nor U7733 (N_7733,N_5620,N_5831);
xor U7734 (N_7734,N_5581,N_5559);
or U7735 (N_7735,N_5185,N_5047);
and U7736 (N_7736,N_5066,N_5515);
nor U7737 (N_7737,N_5874,N_5980);
xor U7738 (N_7738,N_5604,N_4804);
nand U7739 (N_7739,N_5346,N_4748);
nor U7740 (N_7740,N_5898,N_5675);
or U7741 (N_7741,N_4368,N_5662);
or U7742 (N_7742,N_4944,N_4443);
nor U7743 (N_7743,N_5179,N_5582);
and U7744 (N_7744,N_5794,N_5633);
xnor U7745 (N_7745,N_5711,N_4857);
xor U7746 (N_7746,N_5782,N_5891);
and U7747 (N_7747,N_5313,N_4408);
and U7748 (N_7748,N_4314,N_4115);
nor U7749 (N_7749,N_4494,N_4807);
nand U7750 (N_7750,N_5878,N_4883);
nand U7751 (N_7751,N_4217,N_5239);
nand U7752 (N_7752,N_4155,N_5666);
or U7753 (N_7753,N_4262,N_5418);
or U7754 (N_7754,N_5680,N_4192);
nor U7755 (N_7755,N_5382,N_4779);
nand U7756 (N_7756,N_5871,N_5907);
nor U7757 (N_7757,N_5343,N_4278);
xor U7758 (N_7758,N_5856,N_5248);
nor U7759 (N_7759,N_4688,N_5579);
nor U7760 (N_7760,N_5838,N_5282);
nand U7761 (N_7761,N_4019,N_4437);
nor U7762 (N_7762,N_4065,N_4871);
and U7763 (N_7763,N_5404,N_4285);
and U7764 (N_7764,N_4537,N_4337);
xor U7765 (N_7765,N_4973,N_5215);
and U7766 (N_7766,N_4610,N_5431);
nor U7767 (N_7767,N_4373,N_4125);
xor U7768 (N_7768,N_4579,N_5871);
and U7769 (N_7769,N_4489,N_4065);
and U7770 (N_7770,N_4292,N_4570);
and U7771 (N_7771,N_5463,N_4265);
nor U7772 (N_7772,N_4173,N_4600);
nand U7773 (N_7773,N_4975,N_5049);
or U7774 (N_7774,N_5993,N_5046);
and U7775 (N_7775,N_4284,N_4867);
nor U7776 (N_7776,N_5936,N_5578);
nand U7777 (N_7777,N_5665,N_4683);
and U7778 (N_7778,N_5915,N_4318);
nor U7779 (N_7779,N_5809,N_4675);
or U7780 (N_7780,N_5606,N_5721);
xor U7781 (N_7781,N_5568,N_5325);
nor U7782 (N_7782,N_5974,N_5465);
nor U7783 (N_7783,N_5311,N_5016);
nand U7784 (N_7784,N_4467,N_4424);
and U7785 (N_7785,N_5504,N_4163);
and U7786 (N_7786,N_4187,N_5521);
nand U7787 (N_7787,N_5072,N_5125);
xnor U7788 (N_7788,N_4701,N_4987);
xnor U7789 (N_7789,N_5724,N_5621);
or U7790 (N_7790,N_5019,N_5109);
xnor U7791 (N_7791,N_4605,N_5450);
nand U7792 (N_7792,N_4062,N_4189);
and U7793 (N_7793,N_5790,N_5849);
xnor U7794 (N_7794,N_4942,N_5906);
and U7795 (N_7795,N_4800,N_4725);
nand U7796 (N_7796,N_4875,N_5566);
xor U7797 (N_7797,N_4727,N_5729);
xor U7798 (N_7798,N_5756,N_4161);
nand U7799 (N_7799,N_4958,N_4066);
xor U7800 (N_7800,N_5709,N_4580);
or U7801 (N_7801,N_4630,N_4449);
and U7802 (N_7802,N_5345,N_5339);
and U7803 (N_7803,N_5912,N_4825);
xnor U7804 (N_7804,N_5831,N_4050);
xnor U7805 (N_7805,N_4109,N_4847);
and U7806 (N_7806,N_4712,N_4619);
nand U7807 (N_7807,N_4346,N_4328);
xor U7808 (N_7808,N_4666,N_5545);
nand U7809 (N_7809,N_5348,N_4559);
and U7810 (N_7810,N_4055,N_4924);
nor U7811 (N_7811,N_4041,N_4479);
nand U7812 (N_7812,N_4555,N_4436);
and U7813 (N_7813,N_4992,N_4672);
nand U7814 (N_7814,N_5235,N_4890);
nand U7815 (N_7815,N_5878,N_5369);
and U7816 (N_7816,N_5116,N_4948);
nand U7817 (N_7817,N_4949,N_5897);
nor U7818 (N_7818,N_5994,N_5719);
nand U7819 (N_7819,N_5632,N_5199);
nor U7820 (N_7820,N_4526,N_5521);
xnor U7821 (N_7821,N_5656,N_5672);
nand U7822 (N_7822,N_5190,N_4997);
nor U7823 (N_7823,N_4152,N_5596);
xor U7824 (N_7824,N_5059,N_5123);
or U7825 (N_7825,N_4832,N_5769);
nand U7826 (N_7826,N_4700,N_4358);
and U7827 (N_7827,N_4264,N_5574);
or U7828 (N_7828,N_5075,N_4013);
nor U7829 (N_7829,N_5943,N_5222);
and U7830 (N_7830,N_5317,N_4733);
nor U7831 (N_7831,N_4742,N_5391);
and U7832 (N_7832,N_5908,N_4769);
nor U7833 (N_7833,N_5124,N_5899);
xor U7834 (N_7834,N_4639,N_5954);
and U7835 (N_7835,N_5296,N_5541);
or U7836 (N_7836,N_4171,N_5069);
or U7837 (N_7837,N_4033,N_4187);
nor U7838 (N_7838,N_4020,N_4762);
nand U7839 (N_7839,N_5089,N_5010);
or U7840 (N_7840,N_4600,N_5849);
nor U7841 (N_7841,N_4423,N_5001);
nor U7842 (N_7842,N_4653,N_5181);
xnor U7843 (N_7843,N_5632,N_5438);
and U7844 (N_7844,N_4771,N_5833);
xor U7845 (N_7845,N_5671,N_4537);
or U7846 (N_7846,N_4729,N_5394);
xnor U7847 (N_7847,N_5529,N_5781);
nand U7848 (N_7848,N_4739,N_5169);
or U7849 (N_7849,N_4638,N_5666);
xnor U7850 (N_7850,N_4325,N_4183);
and U7851 (N_7851,N_5829,N_5597);
nor U7852 (N_7852,N_5860,N_4613);
and U7853 (N_7853,N_5520,N_4204);
or U7854 (N_7854,N_5339,N_5340);
or U7855 (N_7855,N_4683,N_4116);
nor U7856 (N_7856,N_4218,N_5778);
nor U7857 (N_7857,N_5494,N_4162);
nor U7858 (N_7858,N_4417,N_4520);
nor U7859 (N_7859,N_4530,N_5311);
nor U7860 (N_7860,N_4327,N_4285);
xor U7861 (N_7861,N_4753,N_5230);
and U7862 (N_7862,N_4251,N_5178);
or U7863 (N_7863,N_4522,N_4027);
xor U7864 (N_7864,N_4958,N_5826);
xor U7865 (N_7865,N_4551,N_5555);
nor U7866 (N_7866,N_5081,N_5017);
or U7867 (N_7867,N_4305,N_5136);
and U7868 (N_7868,N_4299,N_4336);
or U7869 (N_7869,N_5910,N_4113);
or U7870 (N_7870,N_4169,N_4452);
or U7871 (N_7871,N_4472,N_4520);
xor U7872 (N_7872,N_4966,N_5777);
nor U7873 (N_7873,N_4034,N_4002);
and U7874 (N_7874,N_5518,N_4275);
nand U7875 (N_7875,N_5802,N_4799);
nand U7876 (N_7876,N_4922,N_5842);
nor U7877 (N_7877,N_5994,N_5322);
nor U7878 (N_7878,N_4286,N_5005);
nand U7879 (N_7879,N_4606,N_4589);
nand U7880 (N_7880,N_5798,N_4440);
nor U7881 (N_7881,N_4986,N_5339);
nor U7882 (N_7882,N_4308,N_4206);
or U7883 (N_7883,N_4975,N_5564);
nor U7884 (N_7884,N_5627,N_5952);
nand U7885 (N_7885,N_5263,N_5630);
nand U7886 (N_7886,N_4441,N_5766);
or U7887 (N_7887,N_5705,N_5546);
nand U7888 (N_7888,N_5177,N_5487);
xor U7889 (N_7889,N_4057,N_5845);
or U7890 (N_7890,N_5195,N_5674);
nor U7891 (N_7891,N_4310,N_4190);
nor U7892 (N_7892,N_4371,N_4339);
or U7893 (N_7893,N_5649,N_5657);
nor U7894 (N_7894,N_5871,N_4542);
nand U7895 (N_7895,N_5033,N_5663);
and U7896 (N_7896,N_5984,N_4404);
nor U7897 (N_7897,N_4095,N_5595);
and U7898 (N_7898,N_4295,N_4102);
nand U7899 (N_7899,N_4656,N_4368);
nand U7900 (N_7900,N_4080,N_4090);
xor U7901 (N_7901,N_4545,N_4659);
or U7902 (N_7902,N_5283,N_4407);
or U7903 (N_7903,N_4395,N_4735);
or U7904 (N_7904,N_5376,N_4013);
xnor U7905 (N_7905,N_5645,N_5777);
nand U7906 (N_7906,N_5459,N_5947);
and U7907 (N_7907,N_4588,N_4015);
nor U7908 (N_7908,N_5203,N_5375);
nand U7909 (N_7909,N_4981,N_4055);
nand U7910 (N_7910,N_4591,N_4868);
nor U7911 (N_7911,N_4431,N_4056);
or U7912 (N_7912,N_5304,N_4306);
xnor U7913 (N_7913,N_4694,N_4266);
nor U7914 (N_7914,N_4709,N_5040);
nor U7915 (N_7915,N_5697,N_4985);
nand U7916 (N_7916,N_5888,N_4060);
and U7917 (N_7917,N_5051,N_4768);
nand U7918 (N_7918,N_4700,N_5180);
nand U7919 (N_7919,N_4827,N_4269);
xnor U7920 (N_7920,N_4484,N_5826);
xor U7921 (N_7921,N_4790,N_5324);
or U7922 (N_7922,N_4846,N_5592);
xor U7923 (N_7923,N_4462,N_4621);
and U7924 (N_7924,N_5313,N_4148);
nor U7925 (N_7925,N_4693,N_5382);
nor U7926 (N_7926,N_4489,N_4861);
and U7927 (N_7927,N_4803,N_5024);
xor U7928 (N_7928,N_4025,N_5574);
nor U7929 (N_7929,N_4061,N_5726);
or U7930 (N_7930,N_4391,N_4394);
nand U7931 (N_7931,N_4443,N_4791);
nor U7932 (N_7932,N_5209,N_4214);
and U7933 (N_7933,N_4355,N_4749);
nor U7934 (N_7934,N_5041,N_5548);
nand U7935 (N_7935,N_4162,N_5061);
or U7936 (N_7936,N_5921,N_4554);
nand U7937 (N_7937,N_4695,N_4126);
or U7938 (N_7938,N_4373,N_5949);
and U7939 (N_7939,N_4683,N_5225);
or U7940 (N_7940,N_5467,N_4931);
or U7941 (N_7941,N_4087,N_5441);
nand U7942 (N_7942,N_5251,N_4977);
and U7943 (N_7943,N_4567,N_5714);
and U7944 (N_7944,N_4737,N_4148);
nor U7945 (N_7945,N_5405,N_5356);
or U7946 (N_7946,N_4446,N_4090);
or U7947 (N_7947,N_4080,N_5352);
nor U7948 (N_7948,N_5532,N_4024);
or U7949 (N_7949,N_5204,N_4180);
nand U7950 (N_7950,N_4465,N_5403);
nor U7951 (N_7951,N_5577,N_4433);
nor U7952 (N_7952,N_5860,N_4728);
or U7953 (N_7953,N_5624,N_5207);
or U7954 (N_7954,N_4316,N_5507);
and U7955 (N_7955,N_4318,N_4093);
or U7956 (N_7956,N_4984,N_5102);
nand U7957 (N_7957,N_5495,N_5637);
nor U7958 (N_7958,N_5650,N_5706);
nor U7959 (N_7959,N_4516,N_4902);
or U7960 (N_7960,N_4042,N_5074);
nor U7961 (N_7961,N_5580,N_5381);
and U7962 (N_7962,N_4779,N_4636);
xor U7963 (N_7963,N_5734,N_5967);
xnor U7964 (N_7964,N_5394,N_4433);
and U7965 (N_7965,N_5164,N_4331);
nor U7966 (N_7966,N_4325,N_5300);
xor U7967 (N_7967,N_4574,N_4388);
nand U7968 (N_7968,N_4734,N_5856);
xnor U7969 (N_7969,N_4393,N_5676);
xnor U7970 (N_7970,N_5986,N_4217);
nor U7971 (N_7971,N_4364,N_5776);
nand U7972 (N_7972,N_4529,N_5495);
and U7973 (N_7973,N_5278,N_5748);
xnor U7974 (N_7974,N_5161,N_5637);
nand U7975 (N_7975,N_4773,N_5970);
nand U7976 (N_7976,N_4590,N_5384);
nor U7977 (N_7977,N_5625,N_4907);
and U7978 (N_7978,N_4391,N_5425);
nor U7979 (N_7979,N_4612,N_5407);
xnor U7980 (N_7980,N_4802,N_5682);
or U7981 (N_7981,N_5467,N_4971);
nor U7982 (N_7982,N_4853,N_5483);
nand U7983 (N_7983,N_5942,N_5528);
nand U7984 (N_7984,N_5283,N_4935);
and U7985 (N_7985,N_5091,N_5803);
xnor U7986 (N_7986,N_4913,N_5894);
xnor U7987 (N_7987,N_5594,N_5885);
or U7988 (N_7988,N_5468,N_4274);
and U7989 (N_7989,N_4291,N_4213);
nand U7990 (N_7990,N_4357,N_4178);
or U7991 (N_7991,N_5840,N_4428);
nor U7992 (N_7992,N_5618,N_4235);
nand U7993 (N_7993,N_5143,N_5364);
and U7994 (N_7994,N_5285,N_4670);
nor U7995 (N_7995,N_5904,N_4140);
nor U7996 (N_7996,N_5379,N_5465);
or U7997 (N_7997,N_4456,N_5113);
nand U7998 (N_7998,N_4258,N_5072);
or U7999 (N_7999,N_5323,N_5519);
and U8000 (N_8000,N_7558,N_7606);
and U8001 (N_8001,N_7226,N_7010);
and U8002 (N_8002,N_6666,N_7102);
nor U8003 (N_8003,N_7603,N_6622);
or U8004 (N_8004,N_7588,N_7928);
or U8005 (N_8005,N_7186,N_7909);
nand U8006 (N_8006,N_6383,N_6414);
or U8007 (N_8007,N_7422,N_7556);
nor U8008 (N_8008,N_7595,N_7763);
or U8009 (N_8009,N_7993,N_6095);
and U8010 (N_8010,N_6929,N_7869);
nor U8011 (N_8011,N_6957,N_7589);
and U8012 (N_8012,N_6076,N_7109);
nand U8013 (N_8013,N_7120,N_7737);
and U8014 (N_8014,N_6099,N_7584);
nor U8015 (N_8015,N_6426,N_6833);
and U8016 (N_8016,N_6198,N_6104);
nor U8017 (N_8017,N_6600,N_6521);
xor U8018 (N_8018,N_6627,N_6972);
nor U8019 (N_8019,N_6392,N_7548);
xnor U8020 (N_8020,N_6202,N_7701);
xnor U8021 (N_8021,N_6643,N_7748);
nand U8022 (N_8022,N_7175,N_6677);
nor U8023 (N_8023,N_6887,N_6967);
and U8024 (N_8024,N_6192,N_7460);
or U8025 (N_8025,N_7152,N_7797);
or U8026 (N_8026,N_7182,N_6848);
nand U8027 (N_8027,N_6518,N_6443);
nand U8028 (N_8028,N_6037,N_6434);
nor U8029 (N_8029,N_7153,N_6445);
and U8030 (N_8030,N_7276,N_6488);
or U8031 (N_8031,N_7829,N_6500);
and U8032 (N_8032,N_6422,N_6898);
nand U8033 (N_8033,N_7827,N_6781);
or U8034 (N_8034,N_6913,N_6849);
and U8035 (N_8035,N_6784,N_6910);
and U8036 (N_8036,N_6337,N_7015);
nor U8037 (N_8037,N_7106,N_6792);
and U8038 (N_8038,N_6463,N_6962);
and U8039 (N_8039,N_7773,N_7514);
or U8040 (N_8040,N_6082,N_7021);
or U8041 (N_8041,N_6002,N_6873);
nand U8042 (N_8042,N_6771,N_6812);
nor U8043 (N_8043,N_7911,N_7835);
xor U8044 (N_8044,N_6736,N_6590);
nand U8045 (N_8045,N_7967,N_7978);
or U8046 (N_8046,N_7830,N_7839);
nand U8047 (N_8047,N_7434,N_6394);
nand U8048 (N_8048,N_6330,N_6746);
xnor U8049 (N_8049,N_7012,N_6578);
or U8050 (N_8050,N_7048,N_6901);
or U8051 (N_8051,N_6757,N_6814);
or U8052 (N_8052,N_7327,N_6264);
nand U8053 (N_8053,N_6664,N_6480);
or U8054 (N_8054,N_7002,N_7008);
or U8055 (N_8055,N_7515,N_6012);
or U8056 (N_8056,N_6129,N_6190);
xnor U8057 (N_8057,N_7249,N_7426);
nor U8058 (N_8058,N_6381,N_6331);
or U8059 (N_8059,N_6689,N_7782);
or U8060 (N_8060,N_7072,N_6209);
xor U8061 (N_8061,N_7694,N_7179);
or U8062 (N_8062,N_6249,N_6834);
xnor U8063 (N_8063,N_6496,N_6562);
nand U8064 (N_8064,N_6767,N_6620);
nand U8065 (N_8065,N_6127,N_7764);
or U8066 (N_8066,N_6961,N_6183);
xor U8067 (N_8067,N_7778,N_7273);
and U8068 (N_8068,N_6280,N_6876);
or U8069 (N_8069,N_6585,N_6533);
nand U8070 (N_8070,N_7962,N_7049);
nor U8071 (N_8071,N_7977,N_6541);
or U8072 (N_8072,N_7442,N_7571);
xor U8073 (N_8073,N_6278,N_7063);
nor U8074 (N_8074,N_7724,N_6718);
xor U8075 (N_8075,N_7453,N_7683);
or U8076 (N_8076,N_7920,N_6731);
and U8077 (N_8077,N_7592,N_6173);
nor U8078 (N_8078,N_6428,N_7866);
and U8079 (N_8079,N_7148,N_7073);
or U8080 (N_8080,N_7609,N_7956);
and U8081 (N_8081,N_7343,N_7802);
or U8082 (N_8082,N_6566,N_7423);
nand U8083 (N_8083,N_6390,N_6969);
and U8084 (N_8084,N_6250,N_7893);
nor U8085 (N_8085,N_6732,N_7625);
and U8086 (N_8086,N_7346,N_6869);
xnor U8087 (N_8087,N_6884,N_7331);
xnor U8088 (N_8088,N_6213,N_7900);
and U8089 (N_8089,N_7886,N_6088);
or U8090 (N_8090,N_6226,N_7275);
xnor U8091 (N_8091,N_6885,N_7128);
xnor U8092 (N_8092,N_7812,N_6520);
and U8093 (N_8093,N_6185,N_7726);
and U8094 (N_8094,N_7583,N_6623);
and U8095 (N_8095,N_6484,N_6084);
nor U8096 (N_8096,N_7338,N_7796);
nor U8097 (N_8097,N_7542,N_6852);
nand U8098 (N_8098,N_6892,N_7104);
xor U8099 (N_8099,N_6195,N_6102);
and U8100 (N_8100,N_6719,N_6244);
or U8101 (N_8101,N_6478,N_6455);
nand U8102 (N_8102,N_7283,N_7974);
and U8103 (N_8103,N_6345,N_6860);
nand U8104 (N_8104,N_6070,N_6580);
and U8105 (N_8105,N_7727,N_6351);
and U8106 (N_8106,N_6801,N_6575);
and U8107 (N_8107,N_7711,N_6239);
or U8108 (N_8108,N_7799,N_7501);
nand U8109 (N_8109,N_7597,N_6656);
nor U8110 (N_8110,N_6167,N_6459);
xor U8111 (N_8111,N_6237,N_7766);
and U8112 (N_8112,N_6125,N_7998);
nor U8113 (N_8113,N_7167,N_6322);
or U8114 (N_8114,N_7767,N_6219);
and U8115 (N_8115,N_7375,N_6145);
and U8116 (N_8116,N_6754,N_6636);
nor U8117 (N_8117,N_7480,N_6927);
nor U8118 (N_8118,N_6633,N_7244);
and U8119 (N_8119,N_6690,N_7005);
xor U8120 (N_8120,N_7805,N_6760);
nor U8121 (N_8121,N_7599,N_7046);
and U8122 (N_8122,N_7628,N_7591);
or U8123 (N_8123,N_6602,N_7696);
xor U8124 (N_8124,N_7994,N_6995);
or U8125 (N_8125,N_6068,N_7731);
xnor U8126 (N_8126,N_7441,N_7598);
nand U8127 (N_8127,N_6487,N_6100);
or U8128 (N_8128,N_7322,N_7985);
or U8129 (N_8129,N_7769,N_6476);
nor U8130 (N_8130,N_7541,N_6758);
and U8131 (N_8131,N_6701,N_6344);
or U8132 (N_8132,N_7359,N_7947);
xor U8133 (N_8133,N_6284,N_7986);
or U8134 (N_8134,N_6672,N_7301);
and U8135 (N_8135,N_6638,N_6568);
and U8136 (N_8136,N_6624,N_6366);
nand U8137 (N_8137,N_7043,N_7242);
and U8138 (N_8138,N_6640,N_7732);
xor U8139 (N_8139,N_7365,N_6918);
xnor U8140 (N_8140,N_7674,N_6517);
nor U8141 (N_8141,N_7523,N_6515);
nand U8142 (N_8142,N_7672,N_7155);
nand U8143 (N_8143,N_6153,N_6411);
xnor U8144 (N_8144,N_7966,N_6591);
xor U8145 (N_8145,N_7897,N_7999);
and U8146 (N_8146,N_6706,N_6346);
or U8147 (N_8147,N_6039,N_7424);
xor U8148 (N_8148,N_6668,N_7573);
or U8149 (N_8149,N_7604,N_7663);
or U8150 (N_8150,N_6951,N_7945);
nor U8151 (N_8151,N_7420,N_7494);
and U8152 (N_8152,N_7381,N_6859);
nand U8153 (N_8153,N_6679,N_6214);
and U8154 (N_8154,N_6217,N_7124);
nor U8155 (N_8155,N_6400,N_7313);
xor U8156 (N_8156,N_7239,N_7702);
and U8157 (N_8157,N_7526,N_7178);
xor U8158 (N_8158,N_7544,N_6639);
nand U8159 (N_8159,N_7506,N_7093);
or U8160 (N_8160,N_7225,N_7944);
nand U8161 (N_8161,N_7478,N_7315);
nand U8162 (N_8162,N_7388,N_7872);
or U8163 (N_8163,N_7014,N_6503);
nand U8164 (N_8164,N_6742,N_6840);
nand U8165 (N_8165,N_6401,N_6641);
or U8166 (N_8166,N_6328,N_7980);
nand U8167 (N_8167,N_6112,N_7537);
xor U8168 (N_8168,N_7399,N_6948);
nor U8169 (N_8169,N_6700,N_6601);
xor U8170 (N_8170,N_6696,N_7883);
nand U8171 (N_8171,N_6115,N_7164);
or U8172 (N_8172,N_6398,N_6408);
nor U8173 (N_8173,N_6954,N_6406);
and U8174 (N_8174,N_7393,N_6276);
nor U8175 (N_8175,N_6485,N_7366);
xor U8176 (N_8176,N_6015,N_7281);
nor U8177 (N_8177,N_7658,N_6338);
xnor U8178 (N_8178,N_6493,N_6654);
and U8179 (N_8179,N_6940,N_7159);
and U8180 (N_8180,N_6291,N_6512);
or U8181 (N_8181,N_6544,N_6234);
nand U8182 (N_8182,N_7814,N_6789);
xnor U8183 (N_8183,N_6931,N_6745);
xor U8184 (N_8184,N_7925,N_6750);
and U8185 (N_8185,N_7319,N_7306);
xor U8186 (N_8186,N_6772,N_7632);
xnor U8187 (N_8187,N_6258,N_6072);
or U8188 (N_8188,N_6312,N_6551);
nor U8189 (N_8189,N_7368,N_7547);
xor U8190 (N_8190,N_7861,N_6528);
and U8191 (N_8191,N_7085,N_7117);
and U8192 (N_8192,N_6530,N_6788);
nor U8193 (N_8193,N_7130,N_7027);
nand U8194 (N_8194,N_7856,N_7286);
or U8195 (N_8195,N_7485,N_6928);
or U8196 (N_8196,N_6158,N_6371);
or U8197 (N_8197,N_6404,N_7575);
and U8198 (N_8198,N_7858,N_7788);
or U8199 (N_8199,N_7648,N_7414);
or U8200 (N_8200,N_7000,N_7750);
nand U8201 (N_8201,N_7250,N_6659);
nand U8202 (N_8202,N_7071,N_6355);
nor U8203 (N_8203,N_6085,N_7676);
nor U8204 (N_8204,N_6212,N_7919);
xor U8205 (N_8205,N_7898,N_6013);
xnor U8206 (N_8206,N_7492,N_6582);
nand U8207 (N_8207,N_7335,N_6323);
xor U8208 (N_8208,N_6681,N_6955);
or U8209 (N_8209,N_7876,N_6608);
and U8210 (N_8210,N_6595,N_7241);
nor U8211 (N_8211,N_7462,N_7620);
xnor U8212 (N_8212,N_6377,N_6157);
nand U8213 (N_8213,N_7795,N_7234);
and U8214 (N_8214,N_7188,N_6702);
nand U8215 (N_8215,N_6688,N_6610);
nor U8216 (N_8216,N_6993,N_6794);
nor U8217 (N_8217,N_7105,N_6449);
nand U8218 (N_8218,N_6866,N_6343);
or U8219 (N_8219,N_7529,N_7428);
nor U8220 (N_8220,N_6862,N_7140);
nand U8221 (N_8221,N_6150,N_6571);
or U8222 (N_8222,N_7011,N_6193);
xnor U8223 (N_8223,N_6998,N_7534);
or U8224 (N_8224,N_6041,N_6205);
or U8225 (N_8225,N_7834,N_6300);
xor U8226 (N_8226,N_6415,N_6891);
and U8227 (N_8227,N_7617,N_6534);
nor U8228 (N_8228,N_6333,N_7051);
and U8229 (N_8229,N_7636,N_6557);
nor U8230 (N_8230,N_6008,N_7964);
and U8231 (N_8231,N_6550,N_7271);
or U8232 (N_8232,N_6352,N_6589);
or U8233 (N_8233,N_6796,N_6511);
or U8234 (N_8234,N_7487,N_7577);
nand U8235 (N_8235,N_6524,N_7668);
or U8236 (N_8236,N_7357,N_7621);
or U8237 (N_8237,N_7451,N_7068);
nor U8238 (N_8238,N_7195,N_7963);
nand U8239 (N_8239,N_6175,N_7644);
and U8240 (N_8240,N_6727,N_6262);
nor U8241 (N_8241,N_7937,N_6453);
nor U8242 (N_8242,N_6603,N_6616);
nor U8243 (N_8243,N_7688,N_7895);
or U8244 (N_8244,N_6753,N_7800);
xor U8245 (N_8245,N_7154,N_6332);
or U8246 (N_8246,N_6353,N_7469);
nand U8247 (N_8247,N_6994,N_7285);
or U8248 (N_8248,N_6872,N_7934);
nor U8249 (N_8249,N_7899,N_6033);
xor U8250 (N_8250,N_7661,N_7720);
or U8251 (N_8251,N_6265,N_6695);
xnor U8252 (N_8252,N_7197,N_7561);
xor U8253 (N_8253,N_7933,N_6416);
xor U8254 (N_8254,N_7025,N_7336);
nor U8255 (N_8255,N_6966,N_7230);
nand U8256 (N_8256,N_6272,N_6935);
nand U8257 (N_8257,N_7545,N_7825);
nor U8258 (N_8258,N_6116,N_6768);
or U8259 (N_8259,N_7728,N_6900);
or U8260 (N_8260,N_7376,N_6475);
nor U8261 (N_8261,N_6106,N_7902);
or U8262 (N_8262,N_6227,N_7196);
nand U8263 (N_8263,N_6024,N_7578);
nand U8264 (N_8264,N_6501,N_6465);
xor U8265 (N_8265,N_6699,N_7077);
and U8266 (N_8266,N_7267,N_7450);
nand U8267 (N_8267,N_7781,N_7940);
xnor U8268 (N_8268,N_7259,N_7212);
nor U8269 (N_8269,N_7204,N_7983);
nor U8270 (N_8270,N_7961,N_7089);
or U8271 (N_8271,N_6724,N_7047);
or U8272 (N_8272,N_6117,N_6172);
or U8273 (N_8273,N_7679,N_6118);
or U8274 (N_8274,N_7044,N_7939);
nor U8275 (N_8275,N_7170,N_6799);
nor U8276 (N_8276,N_7303,N_6964);
or U8277 (N_8277,N_7585,N_6078);
nor U8278 (N_8278,N_7041,N_6054);
nor U8279 (N_8279,N_6271,N_6233);
and U8280 (N_8280,N_6797,N_6539);
and U8281 (N_8281,N_7502,N_7162);
and U8282 (N_8282,N_7987,N_7160);
xor U8283 (N_8283,N_7618,N_7735);
and U8284 (N_8284,N_7342,N_7166);
and U8285 (N_8285,N_7543,N_7026);
xor U8286 (N_8286,N_7832,N_6368);
nand U8287 (N_8287,N_6723,N_7486);
and U8288 (N_8288,N_7177,N_7458);
xor U8289 (N_8289,N_7060,N_6987);
xor U8290 (N_8290,N_7787,N_7408);
nor U8291 (N_8291,N_6358,N_6441);
xnor U8292 (N_8292,N_7314,N_7418);
xnor U8293 (N_8293,N_6458,N_7931);
nor U8294 (N_8294,N_7991,N_7397);
xnor U8295 (N_8295,N_7435,N_7405);
and U8296 (N_8296,N_7108,N_7670);
or U8297 (N_8297,N_7559,N_6919);
or U8298 (N_8298,N_7739,N_7427);
xor U8299 (N_8299,N_7894,N_6680);
nor U8300 (N_8300,N_7682,N_7392);
nand U8301 (N_8301,N_7740,N_6791);
xnor U8302 (N_8302,N_6785,N_6267);
and U8303 (N_8303,N_6738,N_7853);
or U8304 (N_8304,N_7891,N_7233);
xor U8305 (N_8305,N_6765,N_6747);
nand U8306 (N_8306,N_6572,N_7602);
nor U8307 (N_8307,N_6468,N_7317);
xor U8308 (N_8308,N_7804,N_6963);
or U8309 (N_8309,N_6274,N_6440);
nor U8310 (N_8310,N_7600,N_6980);
nand U8311 (N_8311,N_7174,N_7907);
xnor U8312 (N_8312,N_6467,N_6925);
nor U8313 (N_8313,N_7707,N_6035);
or U8314 (N_8314,N_7278,N_6479);
or U8315 (N_8315,N_7734,N_7332);
or U8316 (N_8316,N_6004,N_7213);
nand U8317 (N_8317,N_6141,N_6313);
nor U8318 (N_8318,N_7517,N_6399);
or U8319 (N_8319,N_6536,N_6427);
nand U8320 (N_8320,N_7190,N_6830);
and U8321 (N_8321,N_6221,N_7954);
and U8322 (N_8322,N_6230,N_6879);
nand U8323 (N_8323,N_7325,N_7084);
and U8324 (N_8324,N_7007,N_6255);
nor U8325 (N_8325,N_6336,N_7292);
nor U8326 (N_8326,N_7379,N_7386);
nand U8327 (N_8327,N_6667,N_6619);
or U8328 (N_8328,N_7490,N_6697);
and U8329 (N_8329,N_6122,N_7127);
and U8330 (N_8330,N_6321,N_7113);
nand U8331 (N_8331,N_7689,N_6548);
and U8332 (N_8332,N_6748,N_6489);
or U8333 (N_8333,N_6936,N_7813);
nand U8334 (N_8334,N_7066,N_7354);
xnor U8335 (N_8335,N_7774,N_7733);
nor U8336 (N_8336,N_7790,N_6804);
and U8337 (N_8337,N_7036,N_6093);
nor U8338 (N_8338,N_6299,N_7611);
and U8339 (N_8339,N_6637,N_7811);
or U8340 (N_8340,N_7340,N_7193);
nand U8341 (N_8341,N_7401,N_7497);
nand U8342 (N_8342,N_7345,N_7922);
and U8343 (N_8343,N_6257,N_7308);
nor U8344 (N_8344,N_6018,N_6010);
nand U8345 (N_8345,N_7771,N_6941);
nand U8346 (N_8346,N_6165,N_6692);
and U8347 (N_8347,N_7555,N_6982);
xnor U8348 (N_8348,N_7581,N_6777);
or U8349 (N_8349,N_7050,N_7474);
nand U8350 (N_8350,N_7168,N_7996);
nand U8351 (N_8351,N_6287,N_6107);
nor U8352 (N_8352,N_6334,N_6868);
xor U8353 (N_8353,N_6087,N_6974);
and U8354 (N_8354,N_6663,N_6775);
or U8355 (N_8355,N_7863,N_7151);
and U8356 (N_8356,N_6798,N_6131);
nor U8357 (N_8357,N_6315,N_6561);
or U8358 (N_8358,N_6259,N_6835);
and U8359 (N_8359,N_6581,N_6556);
and U8360 (N_8360,N_7320,N_6650);
nand U8361 (N_8361,N_6136,N_7718);
or U8362 (N_8362,N_6047,N_6770);
nor U8363 (N_8363,N_6795,N_6294);
or U8364 (N_8364,N_7318,N_7202);
nand U8365 (N_8365,N_6350,N_7350);
or U8366 (N_8366,N_7333,N_7647);
xor U8367 (N_8367,N_6335,N_6555);
nor U8368 (N_8368,N_7772,N_6450);
xnor U8369 (N_8369,N_7406,N_7307);
or U8370 (N_8370,N_6716,N_6140);
nand U8371 (N_8371,N_7293,N_7507);
or U8372 (N_8372,N_6875,N_6851);
nor U8373 (N_8373,N_7698,N_6540);
xor U8374 (N_8374,N_7496,N_7169);
and U8375 (N_8375,N_7149,N_7383);
and U8376 (N_8376,N_6722,N_6210);
and U8377 (N_8377,N_6625,N_6326);
nand U8378 (N_8378,N_7132,N_6341);
nor U8379 (N_8379,N_6020,N_7305);
or U8380 (N_8380,N_6537,N_6956);
or U8381 (N_8381,N_7471,N_6292);
and U8382 (N_8382,N_6146,N_7666);
nor U8383 (N_8383,N_6286,N_6030);
and U8384 (N_8384,N_7784,N_7892);
and U8385 (N_8385,N_7262,N_6043);
nand U8386 (N_8386,N_6992,N_7086);
and U8387 (N_8387,N_6495,N_7079);
nand U8388 (N_8388,N_7216,N_7110);
nand U8389 (N_8389,N_6403,N_7681);
and U8390 (N_8390,N_6028,N_7030);
nand U8391 (N_8391,N_7981,N_7705);
xnor U8392 (N_8392,N_7844,N_7746);
nor U8393 (N_8393,N_7957,N_6693);
nand U8394 (N_8394,N_6553,N_6514);
and U8395 (N_8395,N_7463,N_6563);
and U8396 (N_8396,N_7572,N_7614);
or U8397 (N_8397,N_7147,N_7039);
nor U8398 (N_8398,N_7712,N_7411);
nand U8399 (N_8399,N_7596,N_6171);
nor U8400 (N_8400,N_7253,N_7927);
xnor U8401 (N_8401,N_6111,N_7103);
or U8402 (N_8402,N_6604,N_7851);
nor U8403 (N_8403,N_6645,N_7633);
or U8404 (N_8404,N_7510,N_6678);
or U8405 (N_8405,N_6721,N_6743);
and U8406 (N_8406,N_6318,N_6766);
nand U8407 (N_8407,N_7006,N_6256);
or U8408 (N_8408,N_6605,N_6710);
xor U8409 (N_8409,N_6402,N_6301);
or U8410 (N_8410,N_7358,N_6184);
or U8411 (N_8411,N_6147,N_7219);
and U8412 (N_8412,N_7390,N_7982);
nand U8413 (N_8413,N_6446,N_6761);
nor U8414 (N_8414,N_7730,N_6881);
or U8415 (N_8415,N_6507,N_7513);
or U8416 (N_8416,N_6907,N_6471);
nor U8417 (N_8417,N_7252,N_6614);
or U8418 (N_8418,N_6229,N_7777);
xnor U8419 (N_8419,N_6120,N_7187);
or U8420 (N_8420,N_7107,N_6384);
xnor U8421 (N_8421,N_7031,N_7650);
xor U8422 (N_8422,N_6543,N_7037);
nand U8423 (N_8423,N_7729,N_6382);
nand U8424 (N_8424,N_7351,N_6273);
or U8425 (N_8425,N_7889,N_7521);
nor U8426 (N_8426,N_6902,N_7719);
xnor U8427 (N_8427,N_7288,N_6819);
xor U8428 (N_8428,N_7616,N_7511);
nor U8429 (N_8429,N_6389,N_6634);
and U8430 (N_8430,N_6843,N_6429);
or U8431 (N_8431,N_7367,N_6588);
nor U8432 (N_8432,N_7024,N_6660);
nor U8433 (N_8433,N_7311,N_7817);
xnor U8434 (N_8434,N_7877,N_6744);
or U8435 (N_8435,N_7316,N_6232);
or U8436 (N_8436,N_7549,N_7943);
xor U8437 (N_8437,N_7150,N_7906);
xnor U8438 (N_8438,N_6809,N_7298);
nor U8439 (N_8439,N_7783,N_7415);
nand U8440 (N_8440,N_7466,N_7531);
nand U8441 (N_8441,N_7180,N_6186);
or U8442 (N_8442,N_6413,N_6074);
or U8443 (N_8443,N_6717,N_6831);
and U8444 (N_8444,N_6546,N_6045);
and U8445 (N_8445,N_6016,N_6367);
xnor U8446 (N_8446,N_7228,N_7203);
and U8447 (N_8447,N_6741,N_6508);
and U8448 (N_8448,N_6871,N_6822);
nor U8449 (N_8449,N_7477,N_7323);
nor U8450 (N_8450,N_6565,N_7997);
and U8451 (N_8451,N_6483,N_7144);
nand U8452 (N_8452,N_6361,N_6216);
nand U8453 (N_8453,N_7083,N_7246);
nand U8454 (N_8454,N_7833,N_7004);
nor U8455 (N_8455,N_6009,N_7290);
xnor U8456 (N_8456,N_7809,N_6437);
nor U8457 (N_8457,N_6032,N_6592);
nand U8458 (N_8458,N_6535,N_6973);
xnor U8459 (N_8459,N_6740,N_7838);
and U8460 (N_8460,N_7439,N_6023);
xnor U8461 (N_8461,N_7539,N_7815);
nand U8462 (N_8462,N_6461,N_7576);
xnor U8463 (N_8463,N_7791,N_7504);
xnor U8464 (N_8464,N_7565,N_7238);
or U8465 (N_8465,N_7053,N_7129);
and U8466 (N_8466,N_7171,N_6939);
xnor U8467 (N_8467,N_6053,N_6921);
nor U8468 (N_8468,N_6498,N_6316);
xnor U8469 (N_8469,N_7657,N_6372);
xor U8470 (N_8470,N_6375,N_7377);
and U8471 (N_8471,N_6593,N_7693);
and U8472 (N_8472,N_6684,N_7461);
or U8473 (N_8473,N_7503,N_6182);
and U8474 (N_8474,N_7437,N_6225);
nor U8475 (N_8475,N_7028,N_7431);
xor U8476 (N_8476,N_6825,N_7765);
nand U8477 (N_8477,N_7257,N_6762);
nand U8478 (N_8478,N_7413,N_7873);
nor U8479 (N_8479,N_6909,N_6224);
xnor U8480 (N_8480,N_7137,N_6793);
or U8481 (N_8481,N_7236,N_6289);
or U8482 (N_8482,N_7530,N_7133);
and U8483 (N_8483,N_6162,N_7550);
and U8484 (N_8484,N_6751,N_7846);
xnor U8485 (N_8485,N_7965,N_6086);
nor U8486 (N_8486,N_7139,N_7370);
xnor U8487 (N_8487,N_6065,N_7481);
nor U8488 (N_8488,N_6223,N_7780);
and U8489 (N_8489,N_7801,N_6560);
and U8490 (N_8490,N_6132,N_7924);
and U8491 (N_8491,N_7901,N_6059);
xor U8492 (N_8492,N_6842,N_7852);
and U8493 (N_8493,N_6728,N_7634);
or U8494 (N_8494,N_6867,N_6930);
xor U8495 (N_8495,N_7867,N_7090);
and U8496 (N_8496,N_6194,N_7713);
and U8497 (N_8497,N_6857,N_7918);
xor U8498 (N_8498,N_7566,N_7652);
nand U8499 (N_8499,N_7903,N_6915);
and U8500 (N_8500,N_6924,N_6756);
and U8501 (N_8501,N_6632,N_6340);
nand U8502 (N_8502,N_7706,N_6121);
or U8503 (N_8503,N_7134,N_6252);
xor U8504 (N_8504,N_7887,N_7279);
nand U8505 (N_8505,N_7067,N_6545);
and U8506 (N_8506,N_6944,N_6466);
nor U8507 (N_8507,N_7563,N_6708);
or U8508 (N_8508,N_7018,N_7580);
xor U8509 (N_8509,N_7874,N_6405);
nor U8510 (N_8510,N_6342,N_6269);
and U8511 (N_8511,N_7254,N_7753);
xnor U8512 (N_8512,N_6947,N_6456);
nor U8513 (N_8513,N_6108,N_6469);
nor U8514 (N_8514,N_7360,N_6138);
and U8515 (N_8515,N_6370,N_6387);
and U8516 (N_8516,N_7960,N_6042);
xor U8517 (N_8517,N_7888,N_7380);
or U8518 (N_8518,N_7467,N_7988);
nor U8519 (N_8519,N_7500,N_6621);
and U8520 (N_8520,N_6726,N_7865);
nor U8521 (N_8521,N_6438,N_6737);
xnor U8522 (N_8522,N_7118,N_7936);
xor U8523 (N_8523,N_6191,N_7605);
and U8524 (N_8524,N_6110,N_6270);
nor U8525 (N_8525,N_6181,N_6522);
xnor U8526 (N_8526,N_7522,N_6044);
or U8527 (N_8527,N_7329,N_6598);
and U8528 (N_8528,N_7751,N_7324);
and U8529 (N_8529,N_6066,N_6506);
and U8530 (N_8530,N_6103,N_6526);
nor U8531 (N_8531,N_6990,N_6836);
or U8532 (N_8532,N_6497,N_6424);
and U8533 (N_8533,N_7417,N_7263);
or U8534 (N_8534,N_7384,N_7266);
nand U8535 (N_8535,N_6134,N_7594);
or U8536 (N_8536,N_7615,N_6290);
nand U8537 (N_8537,N_7157,N_7508);
or U8538 (N_8538,N_7361,N_7211);
xnor U8539 (N_8539,N_7328,N_7971);
xor U8540 (N_8540,N_6739,N_6109);
nor U8541 (N_8541,N_6457,N_6128);
xnor U8542 (N_8542,N_6714,N_6161);
nor U8543 (N_8543,N_7076,N_7921);
or U8544 (N_8544,N_7095,N_6613);
and U8545 (N_8545,N_6027,N_6492);
xor U8546 (N_8546,N_7942,N_6014);
nor U8547 (N_8547,N_6419,N_6354);
and U8548 (N_8548,N_7564,N_6686);
nor U8549 (N_8549,N_7651,N_7227);
and U8550 (N_8550,N_6832,N_7391);
nand U8551 (N_8551,N_7070,N_7116);
nand U8552 (N_8552,N_7232,N_6022);
nor U8553 (N_8553,N_6698,N_7761);
xor U8554 (N_8554,N_6609,N_7755);
nand U8555 (N_8555,N_7792,N_6655);
xor U8556 (N_8556,N_6985,N_7023);
xor U8557 (N_8557,N_7347,N_6094);
nor U8558 (N_8558,N_6943,N_6482);
or U8559 (N_8559,N_6310,N_6283);
nand U8560 (N_8560,N_7820,N_7505);
xor U8561 (N_8561,N_7612,N_7810);
nor U8562 (N_8562,N_6159,N_7348);
nor U8563 (N_8563,N_6845,N_7673);
xnor U8564 (N_8564,N_7473,N_7995);
nor U8565 (N_8565,N_6435,N_6658);
xnor U8566 (N_8566,N_7640,N_6519);
xnor U8567 (N_8567,N_6135,N_6425);
nand U8568 (N_8568,N_7287,N_6409);
nand U8569 (N_8569,N_7173,N_7289);
xor U8570 (N_8570,N_6579,N_6999);
nand U8571 (N_8571,N_7762,N_7199);
and U8572 (N_8572,N_6420,N_6914);
nand U8573 (N_8573,N_6923,N_6001);
nand U8574 (N_8574,N_6373,N_6325);
nand U8575 (N_8575,N_6268,N_6707);
and U8576 (N_8576,N_7302,N_7456);
xor U8577 (N_8577,N_6691,N_7475);
xor U8578 (N_8578,N_7926,N_7794);
or U8579 (N_8579,N_6069,N_6937);
and U8580 (N_8580,N_7912,N_6152);
and U8581 (N_8581,N_7639,N_6049);
nor U8582 (N_8582,N_7678,N_7389);
nor U8583 (N_8583,N_6155,N_7430);
xnor U8584 (N_8584,N_6975,N_7786);
and U8585 (N_8585,N_6713,N_6922);
nor U8586 (N_8586,N_6896,N_7001);
nor U8587 (N_8587,N_7258,N_6559);
nand U8588 (N_8588,N_6060,N_6811);
or U8589 (N_8589,N_6242,N_6040);
xor U8590 (N_8590,N_7627,N_6285);
and U8591 (N_8591,N_7691,N_6991);
xor U8592 (N_8592,N_7968,N_6670);
and U8593 (N_8593,N_6055,N_6648);
nand U8594 (N_8594,N_6201,N_6635);
xnor U8595 (N_8595,N_6945,N_6412);
or U8596 (N_8596,N_7823,N_6675);
xnor U8597 (N_8597,N_7775,N_6137);
or U8598 (N_8598,N_7394,N_7870);
xor U8599 (N_8599,N_7655,N_6164);
xnor U8600 (N_8600,N_6026,N_7630);
or U8601 (N_8601,N_6652,N_6596);
nor U8602 (N_8602,N_7567,N_7831);
xor U8603 (N_8603,N_7880,N_7205);
nand U8604 (N_8604,N_7123,N_7793);
nor U8605 (N_8605,N_7192,N_6308);
nor U8606 (N_8606,N_7759,N_7304);
and U8607 (N_8607,N_6393,N_7040);
or U8608 (N_8608,N_7875,N_7294);
nor U8609 (N_8609,N_6241,N_6673);
nand U8610 (N_8610,N_7953,N_7516);
nand U8611 (N_8611,N_7904,N_6959);
xnor U8612 (N_8612,N_6105,N_7760);
and U8613 (N_8613,N_7754,N_7843);
nand U8614 (N_8614,N_6711,N_7112);
or U8615 (N_8615,N_6824,N_6806);
and U8616 (N_8616,N_7194,N_7321);
nor U8617 (N_8617,N_7098,N_7088);
or U8618 (N_8618,N_7269,N_7915);
xnor U8619 (N_8619,N_7533,N_7280);
xnor U8620 (N_8620,N_7686,N_6733);
and U8621 (N_8621,N_6755,N_7992);
xnor U8622 (N_8622,N_7222,N_6611);
and U8623 (N_8623,N_6442,N_6888);
xnor U8624 (N_8624,N_6038,N_7261);
nor U8625 (N_8625,N_7525,N_7789);
and U8626 (N_8626,N_6017,N_7020);
and U8627 (N_8627,N_7349,N_7057);
xor U8628 (N_8628,N_7448,N_6631);
nand U8629 (N_8629,N_7295,N_6694);
or U8630 (N_8630,N_6302,N_6444);
or U8631 (N_8631,N_7935,N_7409);
xor U8632 (N_8632,N_7862,N_7312);
nor U8633 (N_8633,N_7009,N_7034);
nor U8634 (N_8634,N_7444,N_7013);
xnor U8635 (N_8635,N_7416,N_6653);
or U8636 (N_8636,N_7436,N_6130);
or U8637 (N_8637,N_7626,N_6567);
nor U8638 (N_8638,N_6584,N_7029);
nand U8639 (N_8639,N_6597,N_7003);
xor U8640 (N_8640,N_6749,N_7586);
nand U8641 (N_8641,N_7885,N_6397);
nand U8642 (N_8642,N_7099,N_6206);
or U8643 (N_8643,N_6187,N_7499);
xor U8644 (N_8644,N_6774,N_7622);
xor U8645 (N_8645,N_7779,N_6452);
and U8646 (N_8646,N_7770,N_7822);
nand U8647 (N_8647,N_7848,N_7532);
xor U8648 (N_8648,N_6669,N_7512);
nor U8649 (N_8649,N_6926,N_7291);
nor U8650 (N_8650,N_6570,N_6050);
or U8651 (N_8651,N_6805,N_6920);
nand U8652 (N_8652,N_6628,N_6657);
xnor U8653 (N_8653,N_6071,N_7240);
nor U8654 (N_8654,N_6558,N_6529);
xor U8655 (N_8655,N_6953,N_6858);
and U8656 (N_8656,N_6880,N_6248);
xnor U8657 (N_8657,N_6547,N_7557);
xor U8658 (N_8658,N_7806,N_7265);
xor U8659 (N_8659,N_6307,N_6436);
nor U8660 (N_8660,N_6304,N_6474);
xor U8661 (N_8661,N_7540,N_7649);
or U8662 (N_8662,N_6817,N_7270);
or U8663 (N_8663,N_6934,N_7059);
xor U8664 (N_8664,N_7950,N_7685);
and U8665 (N_8665,N_7824,N_6199);
nor U8666 (N_8666,N_7654,N_6447);
or U8667 (N_8667,N_7687,N_6246);
nor U8668 (N_8668,N_7421,N_6574);
or U8669 (N_8669,N_6079,N_6810);
xor U8670 (N_8670,N_6396,N_6779);
or U8671 (N_8671,N_7656,N_7807);
xor U8672 (N_8672,N_6776,N_6968);
and U8673 (N_8673,N_7854,N_6279);
nor U8674 (N_8674,N_6996,N_7062);
and U8675 (N_8675,N_7700,N_6339);
nor U8676 (N_8676,N_6142,N_7745);
nand U8677 (N_8677,N_6081,N_6245);
nor U8678 (N_8678,N_7100,N_7973);
xor U8679 (N_8679,N_7214,N_6599);
and U8680 (N_8680,N_6025,N_6046);
or U8681 (N_8681,N_6430,N_7955);
nand U8682 (N_8682,N_6096,N_6569);
nor U8683 (N_8683,N_6815,N_7172);
nand U8684 (N_8684,N_6861,N_6647);
and U8685 (N_8685,N_7372,N_7352);
xnor U8686 (N_8686,N_6423,N_6883);
nand U8687 (N_8687,N_6882,N_7798);
nand U8688 (N_8688,N_7837,N_6091);
nor U8689 (N_8689,N_6319,N_6895);
or U8690 (N_8690,N_6704,N_6629);
xnor U8691 (N_8691,N_7447,N_7300);
nor U8692 (N_8692,N_7785,N_7019);
xnor U8693 (N_8693,N_7749,N_6448);
or U8694 (N_8694,N_6513,N_6630);
and U8695 (N_8695,N_6494,N_6395);
nand U8696 (N_8696,N_7828,N_6838);
nand U8697 (N_8697,N_6089,N_6532);
or U8698 (N_8698,N_6006,N_6083);
and U8699 (N_8699,N_7949,N_7141);
nor U8700 (N_8700,N_7744,N_7017);
and U8701 (N_8701,N_6235,N_7989);
or U8702 (N_8702,N_6586,N_7488);
nand U8703 (N_8703,N_7245,N_7905);
xnor U8704 (N_8704,N_6769,N_6816);
nor U8705 (N_8705,N_7299,N_6908);
and U8706 (N_8706,N_6188,N_6856);
and U8707 (N_8707,N_6391,N_6365);
nor U8708 (N_8708,N_7975,N_7552);
xor U8709 (N_8709,N_7297,N_7247);
nor U8710 (N_8710,N_6965,N_7509);
nor U8711 (N_8711,N_6143,N_7121);
nand U8712 (N_8712,N_7593,N_7243);
or U8713 (N_8713,N_7446,N_7917);
or U8714 (N_8714,N_7896,N_7206);
nor U8715 (N_8715,N_7757,N_6295);
or U8716 (N_8716,N_6502,N_6826);
nor U8717 (N_8717,N_6036,N_6890);
nand U8718 (N_8718,N_7181,N_6615);
xor U8719 (N_8719,N_7163,N_6505);
nor U8720 (N_8720,N_6564,N_6178);
and U8721 (N_8721,N_6360,N_6917);
and U8722 (N_8722,N_6282,N_7476);
nor U8723 (N_8723,N_6878,N_6827);
and U8724 (N_8724,N_7703,N_6064);
nand U8725 (N_8725,N_7722,N_6486);
nor U8726 (N_8726,N_6853,N_6254);
or U8727 (N_8727,N_6029,N_6828);
and U8728 (N_8728,N_6504,N_7890);
or U8729 (N_8729,N_7970,N_6594);
and U8730 (N_8730,N_7224,N_6156);
xor U8731 (N_8731,N_7958,N_6200);
nand U8732 (N_8732,N_6075,N_6363);
or U8733 (N_8733,N_6376,N_6126);
nor U8734 (N_8734,N_6870,N_7229);
xor U8735 (N_8735,N_7484,N_6052);
and U8736 (N_8736,N_6644,N_6204);
nand U8737 (N_8737,N_7445,N_6877);
nor U8738 (N_8738,N_7396,N_6275);
and U8739 (N_8739,N_7671,N_6386);
or U8740 (N_8740,N_7468,N_6786);
nand U8741 (N_8741,N_7260,N_7184);
or U8742 (N_8742,N_6247,N_7087);
xor U8743 (N_8743,N_6821,N_6538);
and U8744 (N_8744,N_7715,N_7065);
xor U8745 (N_8745,N_7131,N_7438);
and U8746 (N_8746,N_7078,N_6144);
or U8747 (N_8747,N_7284,N_6889);
or U8748 (N_8748,N_6092,N_7951);
nand U8749 (N_8749,N_6123,N_7607);
nor U8750 (N_8750,N_6978,N_7126);
xnor U8751 (N_8751,N_6886,N_6119);
nand U8752 (N_8752,N_6952,N_6179);
nor U8753 (N_8753,N_7914,N_7158);
and U8754 (N_8754,N_6243,N_7881);
xnor U8755 (N_8755,N_7659,N_7842);
or U8756 (N_8756,N_7579,N_7952);
nor U8757 (N_8757,N_6874,N_6021);
and U8758 (N_8758,N_6349,N_7637);
or U8759 (N_8759,N_6454,N_7546);
or U8760 (N_8760,N_6823,N_6464);
nand U8761 (N_8761,N_6288,N_6617);
nand U8762 (N_8762,N_7553,N_7826);
nor U8763 (N_8763,N_6997,N_7183);
nor U8764 (N_8764,N_6780,N_6011);
nand U8765 (N_8765,N_7074,N_7353);
nor U8766 (N_8766,N_7741,N_6057);
and U8767 (N_8767,N_6470,N_7161);
or U8768 (N_8768,N_7207,N_7716);
nand U8769 (N_8769,N_7840,N_6839);
or U8770 (N_8770,N_6261,N_7404);
xnor U8771 (N_8771,N_7695,N_6950);
xnor U8772 (N_8772,N_6356,N_6139);
nor U8773 (N_8773,N_7520,N_7378);
nand U8774 (N_8774,N_6549,N_7528);
and U8775 (N_8775,N_6531,N_7551);
and U8776 (N_8776,N_7554,N_7146);
or U8777 (N_8777,N_7231,N_6583);
and U8778 (N_8778,N_7326,N_7282);
xor U8779 (N_8779,N_7337,N_6380);
nor U8780 (N_8780,N_7064,N_7610);
xor U8781 (N_8781,N_7629,N_7082);
nand U8782 (N_8782,N_7042,N_6730);
or U8783 (N_8783,N_7432,N_7491);
and U8784 (N_8784,N_7096,N_6783);
or U8785 (N_8785,N_6460,N_6687);
nor U8786 (N_8786,N_7176,N_7479);
nand U8787 (N_8787,N_7776,N_7482);
and U8788 (N_8788,N_6298,N_7054);
and U8789 (N_8789,N_7930,N_6906);
or U8790 (N_8790,N_7022,N_7198);
or U8791 (N_8791,N_6215,N_6362);
and U8792 (N_8792,N_7330,N_6916);
or U8793 (N_8793,N_6863,N_7660);
or U8794 (N_8794,N_6499,N_6646);
and U8795 (N_8795,N_6451,N_7631);
and U8796 (N_8796,N_6491,N_7092);
nand U8797 (N_8797,N_7464,N_7457);
and U8798 (N_8798,N_6782,N_6685);
and U8799 (N_8799,N_7248,N_7235);
nor U8800 (N_8800,N_6481,N_6790);
nand U8801 (N_8801,N_6808,N_6222);
xor U8802 (N_8802,N_6897,N_6329);
or U8803 (N_8803,N_7845,N_6552);
and U8804 (N_8804,N_6003,N_7680);
and U8805 (N_8805,N_6912,N_6970);
nand U8806 (N_8806,N_7111,N_7742);
nand U8807 (N_8807,N_6904,N_7268);
nand U8808 (N_8808,N_7016,N_7402);
xor U8809 (N_8809,N_6813,N_6683);
or U8810 (N_8810,N_7309,N_7662);
or U8811 (N_8811,N_6077,N_7385);
or U8812 (N_8812,N_6439,N_6170);
or U8813 (N_8813,N_7433,N_7237);
and U8814 (N_8814,N_7075,N_6062);
or U8815 (N_8815,N_7536,N_6218);
nand U8816 (N_8816,N_7362,N_7272);
xnor U8817 (N_8817,N_6364,N_7709);
nand U8818 (N_8818,N_6977,N_7221);
or U8819 (N_8819,N_6554,N_6098);
nand U8820 (N_8820,N_7941,N_6168);
nand U8821 (N_8821,N_7714,N_6705);
nor U8822 (N_8822,N_7752,N_6958);
nand U8823 (N_8823,N_7560,N_6378);
nand U8824 (N_8824,N_6421,N_6433);
nand U8825 (N_8825,N_7470,N_6573);
and U8826 (N_8826,N_6932,N_6725);
and U8827 (N_8827,N_6211,N_7419);
nand U8828 (N_8828,N_6807,N_7608);
xor U8829 (N_8829,N_6114,N_7455);
nand U8830 (N_8830,N_6418,N_7138);
and U8831 (N_8831,N_6101,N_7398);
xnor U8832 (N_8832,N_7527,N_6160);
nand U8833 (N_8833,N_6709,N_6763);
nor U8834 (N_8834,N_6734,N_7758);
and U8835 (N_8835,N_6576,N_7069);
nor U8836 (N_8836,N_6208,N_7808);
xor U8837 (N_8837,N_7818,N_7871);
nand U8838 (N_8838,N_7836,N_6063);
nor U8839 (N_8839,N_7498,N_7373);
or U8840 (N_8840,N_6979,N_6266);
and U8841 (N_8841,N_7519,N_7878);
and U8842 (N_8842,N_7518,N_7472);
nand U8843 (N_8843,N_6752,N_6846);
nand U8844 (N_8844,N_7721,N_6347);
or U8845 (N_8845,N_7699,N_7459);
nor U8846 (N_8846,N_6000,N_7723);
or U8847 (N_8847,N_7816,N_6005);
and U8848 (N_8848,N_6787,N_6618);
and U8849 (N_8849,N_7916,N_6228);
or U8850 (N_8850,N_7667,N_6516);
or U8851 (N_8851,N_6019,N_7339);
or U8852 (N_8852,N_6314,N_6240);
and U8853 (N_8853,N_7570,N_6607);
nand U8854 (N_8854,N_7908,N_7879);
and U8855 (N_8855,N_6893,N_6007);
nand U8856 (N_8856,N_7929,N_7747);
nor U8857 (N_8857,N_7125,N_6984);
and U8858 (N_8858,N_6169,N_6803);
nor U8859 (N_8859,N_7255,N_6238);
nor U8860 (N_8860,N_6197,N_6986);
nand U8861 (N_8861,N_6327,N_6818);
nand U8862 (N_8862,N_7032,N_6847);
and U8863 (N_8863,N_7624,N_7882);
nor U8864 (N_8864,N_7101,N_7923);
nor U8865 (N_8865,N_7849,N_7264);
nor U8866 (N_8866,N_6369,N_7946);
nand U8867 (N_8867,N_6676,N_6180);
nand U8868 (N_8868,N_7220,N_6703);
xor U8869 (N_8869,N_6067,N_7185);
and U8870 (N_8870,N_7708,N_6864);
or U8871 (N_8871,N_7643,N_6778);
nand U8872 (N_8872,N_6509,N_6720);
nand U8873 (N_8873,N_6988,N_6058);
nand U8874 (N_8874,N_6855,N_6933);
xnor U8875 (N_8875,N_7948,N_6665);
nand U8876 (N_8876,N_6651,N_6712);
nor U8877 (N_8877,N_6090,N_7277);
nand U8878 (N_8878,N_6263,N_6149);
and U8879 (N_8879,N_7208,N_6729);
nand U8880 (N_8880,N_7412,N_6431);
xor U8881 (N_8881,N_7189,N_7035);
and U8882 (N_8882,N_7538,N_7201);
nand U8883 (N_8883,N_7223,N_7959);
nand U8884 (N_8884,N_6073,N_7119);
and U8885 (N_8885,N_6802,N_6662);
nand U8886 (N_8886,N_7400,N_7736);
nand U8887 (N_8887,N_6960,N_6305);
xor U8888 (N_8888,N_6407,N_7884);
nor U8889 (N_8889,N_6236,N_6642);
xnor U8890 (N_8890,N_7341,N_6176);
nand U8891 (N_8891,N_7932,N_7038);
nand U8892 (N_8892,N_7156,N_6297);
nor U8893 (N_8893,N_6911,N_6983);
or U8894 (N_8894,N_7364,N_6124);
nor U8895 (N_8895,N_6177,N_7756);
and U8896 (N_8896,N_6510,N_7310);
or U8897 (N_8897,N_7058,N_7052);
or U8898 (N_8898,N_6661,N_7613);
or U8899 (N_8899,N_6682,N_7535);
and U8900 (N_8900,N_7489,N_7483);
or U8901 (N_8901,N_7642,N_6905);
nor U8902 (N_8902,N_6311,N_6759);
and U8903 (N_8903,N_7645,N_7033);
and U8904 (N_8904,N_7407,N_6357);
nand U8905 (N_8905,N_7743,N_7803);
nor U8906 (N_8906,N_6061,N_7274);
or U8907 (N_8907,N_6303,N_7410);
and U8908 (N_8908,N_7857,N_6542);
nand U8909 (N_8909,N_7425,N_7819);
or U8910 (N_8910,N_6388,N_6773);
or U8911 (N_8911,N_6899,N_6432);
and U8912 (N_8912,N_7452,N_6207);
and U8913 (N_8913,N_6281,N_7395);
nand U8914 (N_8914,N_7256,N_7403);
xnor U8915 (N_8915,N_6841,N_7142);
xor U8916 (N_8916,N_7569,N_7623);
nor U8917 (N_8917,N_6048,N_7690);
nor U8918 (N_8918,N_6097,N_7495);
and U8919 (N_8919,N_7601,N_6220);
nor U8920 (N_8920,N_7251,N_6306);
and U8921 (N_8921,N_7145,N_7717);
and U8922 (N_8922,N_7738,N_6525);
and U8923 (N_8923,N_7136,N_6293);
nand U8924 (N_8924,N_7568,N_6148);
or U8925 (N_8925,N_6971,N_7653);
xnor U8926 (N_8926,N_7115,N_7344);
or U8927 (N_8927,N_7061,N_7768);
and U8928 (N_8928,N_7091,N_7969);
or U8929 (N_8929,N_6051,N_6894);
nand U8930 (N_8930,N_7619,N_6612);
xor U8931 (N_8931,N_7692,N_7355);
nand U8932 (N_8932,N_7984,N_7465);
nand U8933 (N_8933,N_7665,N_7590);
or U8934 (N_8934,N_6348,N_7864);
nand U8935 (N_8935,N_6938,N_7382);
xnor U8936 (N_8936,N_7850,N_7369);
nor U8937 (N_8937,N_6031,N_6309);
nor U8938 (N_8938,N_6379,N_7210);
nand U8939 (N_8939,N_7821,N_7972);
xnor U8940 (N_8940,N_7217,N_6989);
or U8941 (N_8941,N_7045,N_6523);
or U8942 (N_8942,N_7524,N_7725);
nor U8943 (N_8943,N_7218,N_7859);
nor U8944 (N_8944,N_6034,N_7296);
or U8945 (N_8945,N_6473,N_6324);
or U8946 (N_8946,N_7215,N_7056);
nand U8947 (N_8947,N_6976,N_6133);
nor U8948 (N_8948,N_6477,N_6154);
xnor U8949 (N_8949,N_6166,N_6674);
xor U8950 (N_8950,N_7387,N_7374);
xnor U8951 (N_8951,N_7938,N_6174);
nor U8952 (N_8952,N_6800,N_7191);
and U8953 (N_8953,N_6080,N_6253);
or U8954 (N_8954,N_7429,N_6251);
or U8955 (N_8955,N_7641,N_7574);
xnor U8956 (N_8956,N_7664,N_7646);
nand U8957 (N_8957,N_7209,N_7080);
and U8958 (N_8958,N_6359,N_6764);
xor U8959 (N_8959,N_6949,N_7493);
or U8960 (N_8960,N_7443,N_6844);
and U8961 (N_8961,N_7913,N_7454);
and U8962 (N_8962,N_7363,N_7114);
xor U8963 (N_8963,N_6410,N_7910);
xor U8964 (N_8964,N_7855,N_7356);
xnor U8965 (N_8965,N_6837,N_7868);
or U8966 (N_8966,N_6490,N_6577);
nor U8967 (N_8967,N_6260,N_7841);
xor U8968 (N_8968,N_6829,N_7135);
and U8969 (N_8969,N_6417,N_6163);
xnor U8970 (N_8970,N_7635,N_7684);
nor U8971 (N_8971,N_7334,N_7200);
and U8972 (N_8972,N_7847,N_6903);
nand U8973 (N_8973,N_6462,N_6626);
nor U8974 (N_8974,N_6374,N_6320);
nor U8975 (N_8975,N_7669,N_6151);
xnor U8976 (N_8976,N_6587,N_7976);
xor U8977 (N_8977,N_6317,N_6189);
xnor U8978 (N_8978,N_6385,N_7860);
and U8979 (N_8979,N_7704,N_7697);
and U8980 (N_8980,N_7582,N_6850);
or U8981 (N_8981,N_6942,N_6981);
nand U8982 (N_8982,N_6649,N_6671);
nand U8983 (N_8983,N_6203,N_7165);
xnor U8984 (N_8984,N_6472,N_6865);
xor U8985 (N_8985,N_7675,N_7055);
xnor U8986 (N_8986,N_6113,N_6820);
nand U8987 (N_8987,N_6715,N_6735);
or U8988 (N_8988,N_7979,N_7677);
and U8989 (N_8989,N_7587,N_6296);
nor U8990 (N_8990,N_6854,N_7449);
nand U8991 (N_8991,N_7638,N_6196);
nor U8992 (N_8992,N_6606,N_6527);
or U8993 (N_8993,N_7710,N_7440);
or U8994 (N_8994,N_6056,N_7143);
and U8995 (N_8995,N_7122,N_7094);
and U8996 (N_8996,N_7081,N_6231);
nand U8997 (N_8997,N_6277,N_7097);
nor U8998 (N_8998,N_6946,N_7990);
nand U8999 (N_8999,N_7562,N_7371);
and U9000 (N_9000,N_6602,N_7247);
nand U9001 (N_9001,N_7794,N_7740);
nor U9002 (N_9002,N_7816,N_6865);
xnor U9003 (N_9003,N_6163,N_7269);
nor U9004 (N_9004,N_6974,N_6872);
and U9005 (N_9005,N_7304,N_6418);
nor U9006 (N_9006,N_6422,N_6266);
nor U9007 (N_9007,N_7542,N_7879);
nor U9008 (N_9008,N_6615,N_6446);
xnor U9009 (N_9009,N_6551,N_6082);
xor U9010 (N_9010,N_6838,N_6847);
nor U9011 (N_9011,N_7660,N_7579);
or U9012 (N_9012,N_6913,N_7730);
and U9013 (N_9013,N_6874,N_7862);
xnor U9014 (N_9014,N_6716,N_6725);
xnor U9015 (N_9015,N_7799,N_6984);
nand U9016 (N_9016,N_6104,N_7955);
and U9017 (N_9017,N_6085,N_7245);
nand U9018 (N_9018,N_6864,N_6447);
nor U9019 (N_9019,N_7942,N_7347);
or U9020 (N_9020,N_6718,N_7574);
and U9021 (N_9021,N_6791,N_7542);
nand U9022 (N_9022,N_7288,N_7624);
and U9023 (N_9023,N_6442,N_6886);
or U9024 (N_9024,N_7098,N_7012);
and U9025 (N_9025,N_7965,N_6907);
and U9026 (N_9026,N_7546,N_6532);
and U9027 (N_9027,N_6398,N_6992);
nand U9028 (N_9028,N_7060,N_6018);
nand U9029 (N_9029,N_7952,N_7552);
or U9030 (N_9030,N_7304,N_6965);
nand U9031 (N_9031,N_6543,N_7628);
nor U9032 (N_9032,N_7123,N_6252);
nor U9033 (N_9033,N_6752,N_7266);
or U9034 (N_9034,N_7215,N_6084);
nand U9035 (N_9035,N_7197,N_6370);
nand U9036 (N_9036,N_6845,N_7246);
nor U9037 (N_9037,N_7513,N_7361);
and U9038 (N_9038,N_6237,N_6565);
xor U9039 (N_9039,N_6296,N_6554);
or U9040 (N_9040,N_7206,N_6597);
nand U9041 (N_9041,N_7648,N_7683);
or U9042 (N_9042,N_6087,N_7498);
or U9043 (N_9043,N_6204,N_6250);
and U9044 (N_9044,N_6655,N_7715);
nor U9045 (N_9045,N_7437,N_6241);
xor U9046 (N_9046,N_6025,N_7560);
and U9047 (N_9047,N_7520,N_7790);
or U9048 (N_9048,N_7860,N_6223);
nor U9049 (N_9049,N_7043,N_6925);
and U9050 (N_9050,N_7314,N_7021);
nand U9051 (N_9051,N_6613,N_7779);
nor U9052 (N_9052,N_6690,N_6589);
nand U9053 (N_9053,N_6199,N_7346);
or U9054 (N_9054,N_6011,N_7381);
and U9055 (N_9055,N_7117,N_7579);
or U9056 (N_9056,N_6847,N_7938);
nor U9057 (N_9057,N_6718,N_6703);
and U9058 (N_9058,N_7616,N_6339);
and U9059 (N_9059,N_6968,N_7717);
and U9060 (N_9060,N_7732,N_7477);
or U9061 (N_9061,N_6390,N_7425);
nor U9062 (N_9062,N_6116,N_7673);
or U9063 (N_9063,N_7373,N_6664);
or U9064 (N_9064,N_6366,N_7333);
nand U9065 (N_9065,N_6784,N_7487);
and U9066 (N_9066,N_7288,N_7824);
and U9067 (N_9067,N_7956,N_6395);
or U9068 (N_9068,N_7036,N_7546);
or U9069 (N_9069,N_7619,N_6124);
xnor U9070 (N_9070,N_7187,N_6603);
or U9071 (N_9071,N_6381,N_6456);
and U9072 (N_9072,N_7054,N_6818);
and U9073 (N_9073,N_7711,N_6088);
nand U9074 (N_9074,N_6793,N_7046);
or U9075 (N_9075,N_7068,N_7311);
and U9076 (N_9076,N_6824,N_6620);
xor U9077 (N_9077,N_7848,N_7384);
xor U9078 (N_9078,N_7679,N_6458);
xor U9079 (N_9079,N_7574,N_7355);
and U9080 (N_9080,N_6531,N_6506);
xnor U9081 (N_9081,N_6111,N_7719);
or U9082 (N_9082,N_7173,N_7080);
or U9083 (N_9083,N_6914,N_7552);
and U9084 (N_9084,N_6121,N_6508);
nand U9085 (N_9085,N_6869,N_6694);
or U9086 (N_9086,N_7094,N_7545);
nor U9087 (N_9087,N_6209,N_7215);
or U9088 (N_9088,N_6931,N_7328);
nand U9089 (N_9089,N_6665,N_7107);
xor U9090 (N_9090,N_7350,N_6979);
nor U9091 (N_9091,N_7682,N_6267);
nand U9092 (N_9092,N_6030,N_6757);
and U9093 (N_9093,N_6736,N_7412);
and U9094 (N_9094,N_6560,N_6247);
nor U9095 (N_9095,N_6013,N_6642);
and U9096 (N_9096,N_6517,N_7868);
xor U9097 (N_9097,N_6840,N_7385);
or U9098 (N_9098,N_7123,N_6871);
nand U9099 (N_9099,N_7883,N_7440);
and U9100 (N_9100,N_6400,N_6592);
nand U9101 (N_9101,N_7674,N_7690);
nand U9102 (N_9102,N_7572,N_7075);
nor U9103 (N_9103,N_7652,N_7612);
nand U9104 (N_9104,N_7445,N_7979);
or U9105 (N_9105,N_7345,N_6153);
nand U9106 (N_9106,N_7592,N_7505);
nand U9107 (N_9107,N_6550,N_7551);
nand U9108 (N_9108,N_6219,N_7849);
xor U9109 (N_9109,N_6206,N_7457);
nand U9110 (N_9110,N_7848,N_6425);
and U9111 (N_9111,N_6523,N_6470);
xor U9112 (N_9112,N_7771,N_6451);
xor U9113 (N_9113,N_7003,N_6432);
nand U9114 (N_9114,N_7651,N_6744);
nand U9115 (N_9115,N_6237,N_7993);
or U9116 (N_9116,N_6040,N_6433);
or U9117 (N_9117,N_6464,N_6219);
nand U9118 (N_9118,N_6274,N_7107);
and U9119 (N_9119,N_7756,N_7357);
nand U9120 (N_9120,N_6706,N_7563);
and U9121 (N_9121,N_7841,N_7663);
and U9122 (N_9122,N_6571,N_7439);
and U9123 (N_9123,N_7246,N_7380);
xor U9124 (N_9124,N_7091,N_6836);
nor U9125 (N_9125,N_7070,N_6197);
and U9126 (N_9126,N_7251,N_7069);
nor U9127 (N_9127,N_6406,N_6775);
nand U9128 (N_9128,N_7182,N_6908);
xor U9129 (N_9129,N_7671,N_6625);
xnor U9130 (N_9130,N_7454,N_6018);
and U9131 (N_9131,N_7587,N_7980);
or U9132 (N_9132,N_6540,N_7781);
or U9133 (N_9133,N_6474,N_6925);
nand U9134 (N_9134,N_6348,N_6785);
nand U9135 (N_9135,N_7962,N_7293);
or U9136 (N_9136,N_7666,N_6546);
and U9137 (N_9137,N_7999,N_7719);
and U9138 (N_9138,N_6058,N_7250);
xnor U9139 (N_9139,N_7896,N_7485);
nor U9140 (N_9140,N_7978,N_7843);
nor U9141 (N_9141,N_6700,N_6119);
and U9142 (N_9142,N_7046,N_7087);
nand U9143 (N_9143,N_6072,N_6995);
nor U9144 (N_9144,N_7340,N_6760);
or U9145 (N_9145,N_6967,N_7121);
and U9146 (N_9146,N_7837,N_7964);
nand U9147 (N_9147,N_7281,N_7830);
and U9148 (N_9148,N_7542,N_7981);
xnor U9149 (N_9149,N_6598,N_6432);
xnor U9150 (N_9150,N_6915,N_6927);
xor U9151 (N_9151,N_6217,N_7217);
or U9152 (N_9152,N_6242,N_6782);
xnor U9153 (N_9153,N_7463,N_6681);
and U9154 (N_9154,N_6494,N_7712);
nand U9155 (N_9155,N_6004,N_6856);
nor U9156 (N_9156,N_7109,N_7797);
or U9157 (N_9157,N_6068,N_6497);
or U9158 (N_9158,N_6336,N_6899);
nand U9159 (N_9159,N_7188,N_6541);
or U9160 (N_9160,N_6504,N_6120);
nor U9161 (N_9161,N_6499,N_6495);
nor U9162 (N_9162,N_6720,N_6078);
xnor U9163 (N_9163,N_7211,N_7792);
nand U9164 (N_9164,N_7267,N_7747);
or U9165 (N_9165,N_7546,N_7122);
nand U9166 (N_9166,N_6319,N_6679);
nand U9167 (N_9167,N_6560,N_7927);
nor U9168 (N_9168,N_7990,N_6667);
nand U9169 (N_9169,N_6434,N_6698);
nor U9170 (N_9170,N_7342,N_6135);
xor U9171 (N_9171,N_7608,N_7308);
or U9172 (N_9172,N_6901,N_7155);
nand U9173 (N_9173,N_7847,N_6612);
nor U9174 (N_9174,N_6276,N_6827);
nor U9175 (N_9175,N_6065,N_7930);
nor U9176 (N_9176,N_6653,N_6116);
and U9177 (N_9177,N_7401,N_7279);
nor U9178 (N_9178,N_6597,N_7114);
nand U9179 (N_9179,N_7285,N_7827);
nand U9180 (N_9180,N_6215,N_7310);
nand U9181 (N_9181,N_7732,N_7747);
and U9182 (N_9182,N_7466,N_6630);
nor U9183 (N_9183,N_6162,N_6295);
and U9184 (N_9184,N_6151,N_6738);
or U9185 (N_9185,N_7148,N_7204);
nand U9186 (N_9186,N_6146,N_6777);
or U9187 (N_9187,N_7080,N_7709);
or U9188 (N_9188,N_6099,N_7700);
nor U9189 (N_9189,N_6221,N_6097);
nor U9190 (N_9190,N_6606,N_6918);
or U9191 (N_9191,N_7030,N_7198);
nor U9192 (N_9192,N_6383,N_6792);
xnor U9193 (N_9193,N_6679,N_7939);
or U9194 (N_9194,N_6800,N_7300);
or U9195 (N_9195,N_6212,N_7200);
or U9196 (N_9196,N_7149,N_6430);
xnor U9197 (N_9197,N_6147,N_7839);
xor U9198 (N_9198,N_7413,N_6718);
nand U9199 (N_9199,N_7333,N_6066);
or U9200 (N_9200,N_7483,N_7865);
and U9201 (N_9201,N_6345,N_7531);
nand U9202 (N_9202,N_7019,N_7919);
xor U9203 (N_9203,N_7968,N_7977);
or U9204 (N_9204,N_7915,N_7795);
and U9205 (N_9205,N_7808,N_7183);
or U9206 (N_9206,N_6986,N_7865);
xor U9207 (N_9207,N_7896,N_7098);
nor U9208 (N_9208,N_6959,N_7762);
and U9209 (N_9209,N_6291,N_6605);
and U9210 (N_9210,N_6326,N_6243);
xor U9211 (N_9211,N_7739,N_6661);
nor U9212 (N_9212,N_7895,N_6360);
and U9213 (N_9213,N_6434,N_6633);
or U9214 (N_9214,N_6547,N_6792);
xor U9215 (N_9215,N_7674,N_6122);
nand U9216 (N_9216,N_7763,N_6846);
and U9217 (N_9217,N_7254,N_7730);
nand U9218 (N_9218,N_7933,N_6374);
nand U9219 (N_9219,N_6632,N_6195);
nor U9220 (N_9220,N_7491,N_7095);
xnor U9221 (N_9221,N_6851,N_7099);
nor U9222 (N_9222,N_7914,N_7434);
or U9223 (N_9223,N_7089,N_6128);
and U9224 (N_9224,N_7075,N_6848);
nand U9225 (N_9225,N_6746,N_6697);
nand U9226 (N_9226,N_6089,N_7373);
nand U9227 (N_9227,N_7319,N_6443);
and U9228 (N_9228,N_6869,N_7645);
and U9229 (N_9229,N_7922,N_6469);
or U9230 (N_9230,N_7828,N_7433);
and U9231 (N_9231,N_7029,N_7154);
or U9232 (N_9232,N_7045,N_7685);
or U9233 (N_9233,N_7994,N_6046);
nand U9234 (N_9234,N_6327,N_7037);
nor U9235 (N_9235,N_6052,N_7800);
nand U9236 (N_9236,N_6129,N_7620);
nor U9237 (N_9237,N_7273,N_6655);
nor U9238 (N_9238,N_7804,N_6817);
and U9239 (N_9239,N_7375,N_6098);
xnor U9240 (N_9240,N_6444,N_7969);
xnor U9241 (N_9241,N_6308,N_7162);
xor U9242 (N_9242,N_7343,N_6610);
xnor U9243 (N_9243,N_7822,N_6413);
xnor U9244 (N_9244,N_7473,N_6765);
nand U9245 (N_9245,N_7745,N_7725);
and U9246 (N_9246,N_6826,N_7255);
nor U9247 (N_9247,N_7601,N_6627);
xor U9248 (N_9248,N_7120,N_6218);
nand U9249 (N_9249,N_6764,N_7154);
nand U9250 (N_9250,N_7891,N_7457);
nand U9251 (N_9251,N_7863,N_7137);
or U9252 (N_9252,N_7869,N_6467);
and U9253 (N_9253,N_6917,N_6727);
nor U9254 (N_9254,N_6905,N_6813);
nor U9255 (N_9255,N_6588,N_6265);
or U9256 (N_9256,N_7049,N_6908);
and U9257 (N_9257,N_7412,N_7078);
and U9258 (N_9258,N_6766,N_6427);
nor U9259 (N_9259,N_7788,N_7811);
nand U9260 (N_9260,N_7107,N_7842);
or U9261 (N_9261,N_6020,N_6968);
nor U9262 (N_9262,N_7809,N_6462);
nand U9263 (N_9263,N_6456,N_6869);
xnor U9264 (N_9264,N_7558,N_7421);
xnor U9265 (N_9265,N_6506,N_6946);
xnor U9266 (N_9266,N_7041,N_7502);
nor U9267 (N_9267,N_6456,N_6422);
nand U9268 (N_9268,N_6601,N_7054);
and U9269 (N_9269,N_7189,N_7904);
nor U9270 (N_9270,N_7395,N_7344);
nor U9271 (N_9271,N_6546,N_6676);
or U9272 (N_9272,N_7829,N_6782);
and U9273 (N_9273,N_6271,N_6956);
or U9274 (N_9274,N_6297,N_7845);
and U9275 (N_9275,N_6182,N_7710);
nand U9276 (N_9276,N_7489,N_6858);
or U9277 (N_9277,N_6235,N_7547);
nor U9278 (N_9278,N_6403,N_7453);
nor U9279 (N_9279,N_6406,N_7765);
nand U9280 (N_9280,N_7247,N_6114);
nand U9281 (N_9281,N_7393,N_6423);
or U9282 (N_9282,N_6328,N_7341);
or U9283 (N_9283,N_7761,N_6115);
and U9284 (N_9284,N_6741,N_7972);
nand U9285 (N_9285,N_6639,N_6762);
nand U9286 (N_9286,N_7442,N_7378);
and U9287 (N_9287,N_7545,N_7244);
nand U9288 (N_9288,N_7281,N_6953);
xor U9289 (N_9289,N_6167,N_7428);
nor U9290 (N_9290,N_7203,N_6065);
or U9291 (N_9291,N_7415,N_7261);
nor U9292 (N_9292,N_6376,N_6379);
xor U9293 (N_9293,N_6484,N_6017);
or U9294 (N_9294,N_7208,N_6796);
xor U9295 (N_9295,N_7981,N_7125);
nor U9296 (N_9296,N_6242,N_6151);
and U9297 (N_9297,N_7009,N_6883);
nor U9298 (N_9298,N_6580,N_6285);
xor U9299 (N_9299,N_7252,N_7389);
or U9300 (N_9300,N_6794,N_7854);
and U9301 (N_9301,N_7192,N_6671);
or U9302 (N_9302,N_7191,N_7163);
xnor U9303 (N_9303,N_6651,N_7241);
and U9304 (N_9304,N_7868,N_6188);
and U9305 (N_9305,N_6195,N_6019);
xor U9306 (N_9306,N_7390,N_6028);
and U9307 (N_9307,N_6151,N_6256);
nor U9308 (N_9308,N_7647,N_7257);
nor U9309 (N_9309,N_6936,N_6961);
nor U9310 (N_9310,N_7253,N_7470);
nor U9311 (N_9311,N_6367,N_7897);
xnor U9312 (N_9312,N_7076,N_6541);
nand U9313 (N_9313,N_6033,N_6176);
xnor U9314 (N_9314,N_7081,N_6220);
and U9315 (N_9315,N_6917,N_7306);
nand U9316 (N_9316,N_7278,N_6606);
xnor U9317 (N_9317,N_7800,N_6730);
xnor U9318 (N_9318,N_6612,N_6505);
and U9319 (N_9319,N_6254,N_6061);
and U9320 (N_9320,N_6238,N_6520);
and U9321 (N_9321,N_6513,N_7934);
nand U9322 (N_9322,N_6842,N_7137);
xor U9323 (N_9323,N_7159,N_7618);
xor U9324 (N_9324,N_7139,N_7423);
and U9325 (N_9325,N_7874,N_6377);
nor U9326 (N_9326,N_7560,N_7946);
and U9327 (N_9327,N_7693,N_7375);
nand U9328 (N_9328,N_7714,N_6424);
xnor U9329 (N_9329,N_6035,N_7562);
nand U9330 (N_9330,N_6168,N_6071);
and U9331 (N_9331,N_6841,N_6819);
and U9332 (N_9332,N_7584,N_7592);
nand U9333 (N_9333,N_7691,N_7493);
nand U9334 (N_9334,N_7744,N_7335);
and U9335 (N_9335,N_7834,N_6558);
xor U9336 (N_9336,N_7307,N_6980);
nand U9337 (N_9337,N_7511,N_7958);
or U9338 (N_9338,N_7624,N_7551);
nand U9339 (N_9339,N_7010,N_6048);
nor U9340 (N_9340,N_7308,N_7318);
xnor U9341 (N_9341,N_6206,N_6405);
xor U9342 (N_9342,N_7395,N_6292);
nand U9343 (N_9343,N_6349,N_7211);
xnor U9344 (N_9344,N_7676,N_6549);
and U9345 (N_9345,N_6128,N_6771);
xor U9346 (N_9346,N_6190,N_6495);
or U9347 (N_9347,N_7387,N_6159);
xnor U9348 (N_9348,N_6340,N_7908);
nor U9349 (N_9349,N_7790,N_7721);
or U9350 (N_9350,N_6485,N_6091);
xnor U9351 (N_9351,N_7892,N_7195);
nor U9352 (N_9352,N_6971,N_6323);
xnor U9353 (N_9353,N_7866,N_7508);
nor U9354 (N_9354,N_7699,N_6851);
xor U9355 (N_9355,N_7788,N_6569);
and U9356 (N_9356,N_6858,N_7112);
or U9357 (N_9357,N_7752,N_6181);
nor U9358 (N_9358,N_6550,N_7630);
and U9359 (N_9359,N_7797,N_6868);
and U9360 (N_9360,N_7257,N_6239);
and U9361 (N_9361,N_7205,N_7816);
and U9362 (N_9362,N_6737,N_6505);
nor U9363 (N_9363,N_6014,N_6070);
nand U9364 (N_9364,N_7131,N_6288);
or U9365 (N_9365,N_6800,N_7731);
nand U9366 (N_9366,N_6415,N_7012);
xor U9367 (N_9367,N_6365,N_6529);
nor U9368 (N_9368,N_6377,N_6479);
nor U9369 (N_9369,N_7591,N_7819);
nand U9370 (N_9370,N_7731,N_7994);
nor U9371 (N_9371,N_7821,N_7320);
xnor U9372 (N_9372,N_7237,N_6086);
or U9373 (N_9373,N_6972,N_7985);
or U9374 (N_9374,N_7379,N_6368);
and U9375 (N_9375,N_7154,N_6536);
nor U9376 (N_9376,N_6755,N_6300);
nor U9377 (N_9377,N_7999,N_6382);
and U9378 (N_9378,N_6904,N_6325);
nor U9379 (N_9379,N_6793,N_6922);
xor U9380 (N_9380,N_6708,N_6634);
xor U9381 (N_9381,N_7774,N_7528);
nor U9382 (N_9382,N_6377,N_6995);
and U9383 (N_9383,N_7207,N_6706);
xnor U9384 (N_9384,N_6470,N_7544);
xnor U9385 (N_9385,N_6800,N_7749);
nand U9386 (N_9386,N_6173,N_7972);
nand U9387 (N_9387,N_7356,N_6393);
and U9388 (N_9388,N_7186,N_6879);
and U9389 (N_9389,N_7234,N_6174);
nor U9390 (N_9390,N_6522,N_6173);
nand U9391 (N_9391,N_6665,N_6457);
xor U9392 (N_9392,N_7505,N_7152);
nor U9393 (N_9393,N_6917,N_7753);
or U9394 (N_9394,N_6170,N_6653);
or U9395 (N_9395,N_6427,N_7874);
xor U9396 (N_9396,N_7643,N_6339);
xor U9397 (N_9397,N_7391,N_6938);
and U9398 (N_9398,N_6548,N_7471);
nor U9399 (N_9399,N_6940,N_6311);
and U9400 (N_9400,N_6118,N_7083);
xor U9401 (N_9401,N_7963,N_6442);
xnor U9402 (N_9402,N_6644,N_6584);
nor U9403 (N_9403,N_6531,N_6553);
xnor U9404 (N_9404,N_7063,N_6749);
nand U9405 (N_9405,N_6981,N_6208);
or U9406 (N_9406,N_6588,N_6685);
xnor U9407 (N_9407,N_7658,N_7259);
or U9408 (N_9408,N_6534,N_6991);
nand U9409 (N_9409,N_7438,N_7748);
xor U9410 (N_9410,N_6208,N_6071);
and U9411 (N_9411,N_6944,N_7653);
nor U9412 (N_9412,N_6143,N_6823);
and U9413 (N_9413,N_6003,N_6304);
or U9414 (N_9414,N_6654,N_6842);
and U9415 (N_9415,N_7579,N_6124);
xor U9416 (N_9416,N_7130,N_7485);
or U9417 (N_9417,N_6081,N_7893);
xor U9418 (N_9418,N_7617,N_6140);
xor U9419 (N_9419,N_6197,N_6907);
nor U9420 (N_9420,N_7698,N_6803);
or U9421 (N_9421,N_7993,N_7991);
xnor U9422 (N_9422,N_6284,N_7167);
nor U9423 (N_9423,N_7500,N_7920);
nor U9424 (N_9424,N_7737,N_7445);
or U9425 (N_9425,N_6720,N_6986);
nor U9426 (N_9426,N_6994,N_7802);
and U9427 (N_9427,N_7797,N_6800);
and U9428 (N_9428,N_7758,N_7501);
xnor U9429 (N_9429,N_7339,N_6871);
nor U9430 (N_9430,N_7199,N_7246);
or U9431 (N_9431,N_7631,N_7616);
and U9432 (N_9432,N_7331,N_6645);
nor U9433 (N_9433,N_6993,N_7508);
or U9434 (N_9434,N_7075,N_6189);
nand U9435 (N_9435,N_7812,N_6962);
nand U9436 (N_9436,N_7984,N_7471);
and U9437 (N_9437,N_6762,N_6433);
and U9438 (N_9438,N_6318,N_7012);
and U9439 (N_9439,N_6600,N_6240);
xor U9440 (N_9440,N_6835,N_7015);
or U9441 (N_9441,N_6126,N_6218);
or U9442 (N_9442,N_6959,N_6313);
nor U9443 (N_9443,N_7915,N_6378);
or U9444 (N_9444,N_6198,N_7511);
nor U9445 (N_9445,N_6551,N_6498);
or U9446 (N_9446,N_7765,N_6379);
nand U9447 (N_9447,N_7208,N_6683);
nor U9448 (N_9448,N_7551,N_7533);
and U9449 (N_9449,N_6392,N_7174);
xor U9450 (N_9450,N_6812,N_7381);
xnor U9451 (N_9451,N_6317,N_6813);
nand U9452 (N_9452,N_6985,N_7663);
nor U9453 (N_9453,N_7092,N_7508);
nand U9454 (N_9454,N_6590,N_6185);
and U9455 (N_9455,N_6860,N_6932);
nor U9456 (N_9456,N_6017,N_7417);
or U9457 (N_9457,N_7885,N_6892);
nand U9458 (N_9458,N_6227,N_6618);
nor U9459 (N_9459,N_6398,N_6801);
or U9460 (N_9460,N_6665,N_7941);
and U9461 (N_9461,N_7466,N_6550);
xor U9462 (N_9462,N_7019,N_6816);
or U9463 (N_9463,N_7764,N_7207);
nor U9464 (N_9464,N_6006,N_6897);
nand U9465 (N_9465,N_6972,N_6159);
nor U9466 (N_9466,N_7936,N_7029);
or U9467 (N_9467,N_6969,N_7855);
and U9468 (N_9468,N_7310,N_6644);
nor U9469 (N_9469,N_7033,N_7390);
or U9470 (N_9470,N_7578,N_6320);
xor U9471 (N_9471,N_6627,N_6491);
xor U9472 (N_9472,N_6692,N_6614);
or U9473 (N_9473,N_7947,N_7724);
xnor U9474 (N_9474,N_7708,N_7508);
xnor U9475 (N_9475,N_6470,N_6574);
nand U9476 (N_9476,N_7128,N_6911);
or U9477 (N_9477,N_6046,N_7230);
nor U9478 (N_9478,N_6557,N_7197);
or U9479 (N_9479,N_7336,N_6461);
nor U9480 (N_9480,N_6996,N_7779);
and U9481 (N_9481,N_7179,N_7828);
nor U9482 (N_9482,N_7124,N_6834);
or U9483 (N_9483,N_7330,N_7003);
or U9484 (N_9484,N_6980,N_6474);
and U9485 (N_9485,N_6096,N_7723);
xnor U9486 (N_9486,N_6294,N_7776);
or U9487 (N_9487,N_6231,N_6821);
xor U9488 (N_9488,N_7846,N_6135);
and U9489 (N_9489,N_7261,N_6292);
and U9490 (N_9490,N_7056,N_6717);
nor U9491 (N_9491,N_6110,N_7851);
nor U9492 (N_9492,N_6657,N_6051);
nor U9493 (N_9493,N_6568,N_7586);
nand U9494 (N_9494,N_7943,N_7730);
xnor U9495 (N_9495,N_6762,N_7481);
nor U9496 (N_9496,N_7489,N_6173);
xor U9497 (N_9497,N_6437,N_6229);
nor U9498 (N_9498,N_6943,N_6944);
or U9499 (N_9499,N_7316,N_6645);
xnor U9500 (N_9500,N_6967,N_6058);
and U9501 (N_9501,N_7538,N_7468);
or U9502 (N_9502,N_6573,N_7598);
xor U9503 (N_9503,N_6679,N_6127);
nor U9504 (N_9504,N_7191,N_6069);
and U9505 (N_9505,N_7454,N_7922);
nor U9506 (N_9506,N_7968,N_7411);
and U9507 (N_9507,N_6239,N_6110);
nand U9508 (N_9508,N_7591,N_6420);
or U9509 (N_9509,N_6284,N_7832);
nor U9510 (N_9510,N_6528,N_7877);
xor U9511 (N_9511,N_7286,N_6642);
nand U9512 (N_9512,N_7986,N_6749);
nor U9513 (N_9513,N_7894,N_7613);
nand U9514 (N_9514,N_7122,N_6274);
or U9515 (N_9515,N_6263,N_7560);
or U9516 (N_9516,N_6269,N_7690);
or U9517 (N_9517,N_6260,N_7806);
xor U9518 (N_9518,N_7578,N_6594);
xor U9519 (N_9519,N_6162,N_7451);
or U9520 (N_9520,N_7127,N_6622);
nand U9521 (N_9521,N_6702,N_7051);
nand U9522 (N_9522,N_7586,N_6548);
nand U9523 (N_9523,N_7261,N_6802);
nand U9524 (N_9524,N_6539,N_7821);
nor U9525 (N_9525,N_6995,N_6475);
and U9526 (N_9526,N_6362,N_6936);
xor U9527 (N_9527,N_6667,N_7868);
and U9528 (N_9528,N_6957,N_7080);
xnor U9529 (N_9529,N_7733,N_6623);
nor U9530 (N_9530,N_7817,N_6107);
and U9531 (N_9531,N_7769,N_7231);
nor U9532 (N_9532,N_6699,N_6978);
xnor U9533 (N_9533,N_7248,N_6748);
nand U9534 (N_9534,N_6275,N_6691);
and U9535 (N_9535,N_7951,N_7131);
nor U9536 (N_9536,N_7721,N_6650);
and U9537 (N_9537,N_6356,N_6988);
nor U9538 (N_9538,N_6784,N_7103);
nor U9539 (N_9539,N_6635,N_6706);
and U9540 (N_9540,N_6990,N_7898);
and U9541 (N_9541,N_6020,N_6031);
or U9542 (N_9542,N_6399,N_6564);
or U9543 (N_9543,N_6869,N_6363);
nor U9544 (N_9544,N_7268,N_6177);
nor U9545 (N_9545,N_7234,N_7644);
or U9546 (N_9546,N_6698,N_7642);
nand U9547 (N_9547,N_7652,N_6153);
xor U9548 (N_9548,N_7281,N_7234);
nor U9549 (N_9549,N_7325,N_7725);
or U9550 (N_9550,N_6288,N_7796);
xor U9551 (N_9551,N_7218,N_6377);
and U9552 (N_9552,N_7065,N_6165);
nor U9553 (N_9553,N_6558,N_6425);
xnor U9554 (N_9554,N_7415,N_7114);
nand U9555 (N_9555,N_7080,N_6212);
nand U9556 (N_9556,N_6687,N_7299);
and U9557 (N_9557,N_6479,N_7599);
and U9558 (N_9558,N_7722,N_7114);
xnor U9559 (N_9559,N_6425,N_7904);
xor U9560 (N_9560,N_6068,N_6774);
or U9561 (N_9561,N_6265,N_7338);
xnor U9562 (N_9562,N_6874,N_6357);
nand U9563 (N_9563,N_6624,N_6662);
and U9564 (N_9564,N_6979,N_7904);
xnor U9565 (N_9565,N_6931,N_7230);
and U9566 (N_9566,N_7457,N_7771);
and U9567 (N_9567,N_6356,N_7283);
nand U9568 (N_9568,N_7152,N_6271);
xor U9569 (N_9569,N_6025,N_6146);
nand U9570 (N_9570,N_6455,N_6708);
xor U9571 (N_9571,N_6585,N_6204);
and U9572 (N_9572,N_6856,N_6993);
xor U9573 (N_9573,N_6725,N_6249);
xor U9574 (N_9574,N_7220,N_6370);
xnor U9575 (N_9575,N_6701,N_6062);
nor U9576 (N_9576,N_7369,N_7634);
nor U9577 (N_9577,N_6362,N_6182);
xor U9578 (N_9578,N_7984,N_6178);
or U9579 (N_9579,N_7689,N_6019);
xor U9580 (N_9580,N_7741,N_7572);
or U9581 (N_9581,N_6158,N_7729);
nor U9582 (N_9582,N_6189,N_7343);
xor U9583 (N_9583,N_7171,N_7023);
nand U9584 (N_9584,N_7936,N_6738);
nor U9585 (N_9585,N_6583,N_7611);
or U9586 (N_9586,N_6401,N_6643);
xor U9587 (N_9587,N_6138,N_6534);
xor U9588 (N_9588,N_7283,N_7673);
nor U9589 (N_9589,N_7795,N_6934);
or U9590 (N_9590,N_6560,N_7524);
and U9591 (N_9591,N_6510,N_7085);
or U9592 (N_9592,N_6672,N_7080);
xnor U9593 (N_9593,N_7488,N_7845);
xor U9594 (N_9594,N_7696,N_6409);
or U9595 (N_9595,N_6744,N_7294);
nor U9596 (N_9596,N_7583,N_6630);
and U9597 (N_9597,N_6709,N_6331);
and U9598 (N_9598,N_6081,N_7608);
nand U9599 (N_9599,N_7853,N_7451);
and U9600 (N_9600,N_7047,N_7159);
nand U9601 (N_9601,N_7422,N_6308);
or U9602 (N_9602,N_6535,N_6026);
xor U9603 (N_9603,N_7514,N_7965);
or U9604 (N_9604,N_7670,N_7385);
and U9605 (N_9605,N_6145,N_6272);
nand U9606 (N_9606,N_6750,N_6490);
and U9607 (N_9607,N_7974,N_6934);
or U9608 (N_9608,N_6434,N_7826);
nor U9609 (N_9609,N_7696,N_7351);
nor U9610 (N_9610,N_6813,N_7277);
and U9611 (N_9611,N_7957,N_6542);
xor U9612 (N_9612,N_7491,N_7862);
xnor U9613 (N_9613,N_6797,N_6120);
nand U9614 (N_9614,N_6872,N_6009);
xnor U9615 (N_9615,N_6388,N_6297);
nand U9616 (N_9616,N_6648,N_6603);
nor U9617 (N_9617,N_7535,N_6182);
or U9618 (N_9618,N_6533,N_7714);
xnor U9619 (N_9619,N_6888,N_6741);
and U9620 (N_9620,N_7307,N_6466);
and U9621 (N_9621,N_7149,N_7895);
nand U9622 (N_9622,N_6002,N_7231);
and U9623 (N_9623,N_6062,N_7383);
nor U9624 (N_9624,N_7952,N_7586);
xor U9625 (N_9625,N_6245,N_6285);
xnor U9626 (N_9626,N_6294,N_7934);
nor U9627 (N_9627,N_6419,N_7407);
and U9628 (N_9628,N_6127,N_6428);
xnor U9629 (N_9629,N_6022,N_6433);
xor U9630 (N_9630,N_7205,N_7113);
or U9631 (N_9631,N_6741,N_6611);
nand U9632 (N_9632,N_6621,N_6715);
xor U9633 (N_9633,N_6972,N_6694);
and U9634 (N_9634,N_6064,N_7529);
xor U9635 (N_9635,N_6380,N_6113);
nand U9636 (N_9636,N_6005,N_6286);
and U9637 (N_9637,N_6262,N_6468);
or U9638 (N_9638,N_7867,N_6907);
and U9639 (N_9639,N_6836,N_6462);
nand U9640 (N_9640,N_6765,N_6443);
xor U9641 (N_9641,N_7906,N_7885);
xnor U9642 (N_9642,N_7597,N_7584);
xor U9643 (N_9643,N_7618,N_6221);
and U9644 (N_9644,N_7188,N_7198);
nand U9645 (N_9645,N_7229,N_7930);
nor U9646 (N_9646,N_7036,N_6127);
and U9647 (N_9647,N_7005,N_6675);
and U9648 (N_9648,N_6849,N_7457);
or U9649 (N_9649,N_6510,N_7962);
nand U9650 (N_9650,N_6718,N_6475);
and U9651 (N_9651,N_7547,N_7927);
or U9652 (N_9652,N_7657,N_6196);
nand U9653 (N_9653,N_6369,N_7437);
nand U9654 (N_9654,N_6678,N_7056);
xor U9655 (N_9655,N_7528,N_6763);
nor U9656 (N_9656,N_7362,N_7319);
nor U9657 (N_9657,N_7457,N_6678);
nor U9658 (N_9658,N_7098,N_7717);
nand U9659 (N_9659,N_6872,N_7628);
nor U9660 (N_9660,N_7963,N_6413);
or U9661 (N_9661,N_7195,N_6957);
or U9662 (N_9662,N_6268,N_7960);
nor U9663 (N_9663,N_6672,N_7305);
or U9664 (N_9664,N_7237,N_6174);
and U9665 (N_9665,N_7892,N_6677);
xnor U9666 (N_9666,N_6262,N_6829);
nand U9667 (N_9667,N_7663,N_6873);
or U9668 (N_9668,N_6906,N_7042);
nand U9669 (N_9669,N_6586,N_7827);
or U9670 (N_9670,N_6696,N_6305);
nor U9671 (N_9671,N_7885,N_6255);
xnor U9672 (N_9672,N_7862,N_6797);
xor U9673 (N_9673,N_7309,N_6329);
nand U9674 (N_9674,N_7809,N_6470);
nor U9675 (N_9675,N_6304,N_7171);
xor U9676 (N_9676,N_6474,N_6705);
nand U9677 (N_9677,N_7141,N_6136);
or U9678 (N_9678,N_7207,N_7297);
or U9679 (N_9679,N_6807,N_6637);
xnor U9680 (N_9680,N_7346,N_6451);
nand U9681 (N_9681,N_6012,N_7176);
nand U9682 (N_9682,N_7289,N_7149);
or U9683 (N_9683,N_6719,N_6292);
or U9684 (N_9684,N_7679,N_6216);
xor U9685 (N_9685,N_6531,N_6218);
or U9686 (N_9686,N_6364,N_6516);
and U9687 (N_9687,N_6407,N_7366);
and U9688 (N_9688,N_6947,N_6024);
nor U9689 (N_9689,N_7654,N_7690);
and U9690 (N_9690,N_6335,N_7274);
xor U9691 (N_9691,N_7478,N_6377);
nand U9692 (N_9692,N_7375,N_6912);
or U9693 (N_9693,N_7704,N_6770);
xor U9694 (N_9694,N_6209,N_6979);
nand U9695 (N_9695,N_7478,N_6308);
nor U9696 (N_9696,N_6608,N_7162);
xor U9697 (N_9697,N_7364,N_7854);
or U9698 (N_9698,N_6907,N_7851);
or U9699 (N_9699,N_7461,N_7601);
nand U9700 (N_9700,N_7009,N_7587);
nor U9701 (N_9701,N_6876,N_6239);
nor U9702 (N_9702,N_7600,N_6233);
nand U9703 (N_9703,N_7135,N_6753);
nand U9704 (N_9704,N_6113,N_7824);
and U9705 (N_9705,N_6359,N_6896);
nand U9706 (N_9706,N_6374,N_7930);
nand U9707 (N_9707,N_6647,N_6163);
or U9708 (N_9708,N_7484,N_7766);
xnor U9709 (N_9709,N_6646,N_7395);
and U9710 (N_9710,N_6809,N_7593);
nand U9711 (N_9711,N_7696,N_7524);
or U9712 (N_9712,N_6653,N_7496);
or U9713 (N_9713,N_6148,N_6294);
xnor U9714 (N_9714,N_7717,N_6034);
and U9715 (N_9715,N_6249,N_7645);
nand U9716 (N_9716,N_6506,N_7211);
nand U9717 (N_9717,N_7228,N_7027);
nor U9718 (N_9718,N_7394,N_7112);
and U9719 (N_9719,N_7584,N_7088);
nor U9720 (N_9720,N_7606,N_7873);
and U9721 (N_9721,N_6087,N_7374);
xnor U9722 (N_9722,N_6607,N_6151);
and U9723 (N_9723,N_7483,N_6613);
nor U9724 (N_9724,N_6107,N_7712);
and U9725 (N_9725,N_6828,N_7088);
nor U9726 (N_9726,N_6729,N_6564);
nand U9727 (N_9727,N_6853,N_7294);
nor U9728 (N_9728,N_7522,N_7086);
or U9729 (N_9729,N_7068,N_7802);
or U9730 (N_9730,N_6015,N_7827);
xor U9731 (N_9731,N_7559,N_7251);
or U9732 (N_9732,N_7654,N_6595);
or U9733 (N_9733,N_7550,N_6531);
nand U9734 (N_9734,N_6514,N_6214);
xor U9735 (N_9735,N_7316,N_6975);
or U9736 (N_9736,N_7279,N_7230);
nand U9737 (N_9737,N_6713,N_7724);
xnor U9738 (N_9738,N_6078,N_6517);
or U9739 (N_9739,N_7327,N_6477);
nand U9740 (N_9740,N_7125,N_7240);
xnor U9741 (N_9741,N_6136,N_6901);
xnor U9742 (N_9742,N_7287,N_7274);
nand U9743 (N_9743,N_7499,N_7176);
nor U9744 (N_9744,N_7846,N_6061);
or U9745 (N_9745,N_7751,N_6215);
nand U9746 (N_9746,N_7611,N_7633);
nor U9747 (N_9747,N_6259,N_7937);
or U9748 (N_9748,N_6833,N_7457);
or U9749 (N_9749,N_6985,N_6601);
or U9750 (N_9750,N_6047,N_7985);
xor U9751 (N_9751,N_7717,N_6447);
or U9752 (N_9752,N_7374,N_7795);
xor U9753 (N_9753,N_6327,N_7257);
xnor U9754 (N_9754,N_7647,N_7011);
nor U9755 (N_9755,N_6477,N_7403);
or U9756 (N_9756,N_6187,N_6396);
or U9757 (N_9757,N_6467,N_7370);
xor U9758 (N_9758,N_7243,N_6162);
or U9759 (N_9759,N_7398,N_7360);
nand U9760 (N_9760,N_7487,N_6266);
or U9761 (N_9761,N_7012,N_7988);
or U9762 (N_9762,N_6269,N_7962);
nand U9763 (N_9763,N_7687,N_7363);
and U9764 (N_9764,N_7886,N_6060);
nand U9765 (N_9765,N_6902,N_6224);
or U9766 (N_9766,N_6095,N_6918);
nor U9767 (N_9767,N_6958,N_6880);
xor U9768 (N_9768,N_7401,N_7909);
nand U9769 (N_9769,N_6189,N_6613);
nor U9770 (N_9770,N_6710,N_7948);
nor U9771 (N_9771,N_6828,N_6596);
or U9772 (N_9772,N_6110,N_6343);
nand U9773 (N_9773,N_6737,N_7482);
or U9774 (N_9774,N_7155,N_7808);
and U9775 (N_9775,N_7008,N_6452);
nor U9776 (N_9776,N_7394,N_6127);
nand U9777 (N_9777,N_7379,N_6157);
xor U9778 (N_9778,N_6239,N_6722);
xor U9779 (N_9779,N_6541,N_6402);
or U9780 (N_9780,N_7040,N_7955);
nor U9781 (N_9781,N_6191,N_7765);
nor U9782 (N_9782,N_7256,N_7446);
and U9783 (N_9783,N_6607,N_6435);
nor U9784 (N_9784,N_7762,N_7235);
nor U9785 (N_9785,N_7742,N_7807);
or U9786 (N_9786,N_7084,N_7461);
and U9787 (N_9787,N_6465,N_7530);
or U9788 (N_9788,N_6758,N_7787);
xnor U9789 (N_9789,N_6400,N_6367);
nor U9790 (N_9790,N_6668,N_6895);
and U9791 (N_9791,N_6390,N_6031);
nor U9792 (N_9792,N_6093,N_7917);
xnor U9793 (N_9793,N_6336,N_6700);
nor U9794 (N_9794,N_6112,N_7268);
xor U9795 (N_9795,N_6703,N_6048);
nor U9796 (N_9796,N_7292,N_6254);
and U9797 (N_9797,N_6682,N_6501);
and U9798 (N_9798,N_6271,N_6426);
nand U9799 (N_9799,N_7089,N_7343);
and U9800 (N_9800,N_6448,N_6294);
or U9801 (N_9801,N_6305,N_7146);
and U9802 (N_9802,N_7454,N_7500);
nand U9803 (N_9803,N_6191,N_6881);
xnor U9804 (N_9804,N_7370,N_7257);
nor U9805 (N_9805,N_6418,N_6796);
xor U9806 (N_9806,N_6878,N_7096);
nand U9807 (N_9807,N_7451,N_7747);
or U9808 (N_9808,N_6320,N_6482);
xnor U9809 (N_9809,N_7241,N_7783);
nor U9810 (N_9810,N_6380,N_6331);
or U9811 (N_9811,N_6596,N_6016);
xor U9812 (N_9812,N_7063,N_6744);
nand U9813 (N_9813,N_7492,N_6044);
or U9814 (N_9814,N_6376,N_7271);
nor U9815 (N_9815,N_6081,N_6102);
and U9816 (N_9816,N_6429,N_6645);
and U9817 (N_9817,N_6245,N_6403);
or U9818 (N_9818,N_7344,N_7670);
or U9819 (N_9819,N_7964,N_6218);
nor U9820 (N_9820,N_7489,N_6021);
nand U9821 (N_9821,N_7762,N_6787);
or U9822 (N_9822,N_6775,N_7231);
nand U9823 (N_9823,N_7467,N_6525);
or U9824 (N_9824,N_7409,N_7843);
and U9825 (N_9825,N_6549,N_6099);
and U9826 (N_9826,N_6398,N_6289);
or U9827 (N_9827,N_7231,N_6691);
or U9828 (N_9828,N_7893,N_6653);
and U9829 (N_9829,N_7638,N_7545);
or U9830 (N_9830,N_6147,N_6471);
nor U9831 (N_9831,N_7691,N_6850);
and U9832 (N_9832,N_7977,N_6273);
nor U9833 (N_9833,N_7215,N_6497);
xor U9834 (N_9834,N_7084,N_6064);
xor U9835 (N_9835,N_7355,N_6817);
or U9836 (N_9836,N_6838,N_6559);
xor U9837 (N_9837,N_7709,N_7579);
xnor U9838 (N_9838,N_7435,N_6950);
or U9839 (N_9839,N_7562,N_6311);
xnor U9840 (N_9840,N_7563,N_7409);
and U9841 (N_9841,N_7576,N_6783);
or U9842 (N_9842,N_7354,N_6807);
nand U9843 (N_9843,N_6543,N_7412);
or U9844 (N_9844,N_7175,N_7956);
xor U9845 (N_9845,N_7313,N_7188);
or U9846 (N_9846,N_6424,N_6912);
nor U9847 (N_9847,N_7400,N_6371);
xnor U9848 (N_9848,N_7802,N_7280);
nor U9849 (N_9849,N_7064,N_6320);
nor U9850 (N_9850,N_7681,N_7582);
nor U9851 (N_9851,N_6566,N_6483);
or U9852 (N_9852,N_7335,N_6755);
nand U9853 (N_9853,N_7692,N_6169);
or U9854 (N_9854,N_7588,N_7572);
nand U9855 (N_9855,N_7917,N_7146);
nand U9856 (N_9856,N_7623,N_6147);
and U9857 (N_9857,N_7075,N_7408);
nor U9858 (N_9858,N_7088,N_6645);
xor U9859 (N_9859,N_7807,N_7372);
and U9860 (N_9860,N_7554,N_7850);
nand U9861 (N_9861,N_7867,N_7699);
nand U9862 (N_9862,N_6911,N_6154);
xnor U9863 (N_9863,N_6786,N_6706);
or U9864 (N_9864,N_6687,N_6898);
or U9865 (N_9865,N_6974,N_7034);
nand U9866 (N_9866,N_6543,N_7707);
or U9867 (N_9867,N_6706,N_7523);
nand U9868 (N_9868,N_6419,N_6778);
nand U9869 (N_9869,N_6978,N_7693);
and U9870 (N_9870,N_6494,N_6678);
or U9871 (N_9871,N_6130,N_7044);
nand U9872 (N_9872,N_7087,N_7474);
xor U9873 (N_9873,N_6588,N_7937);
xor U9874 (N_9874,N_7830,N_7476);
nand U9875 (N_9875,N_7989,N_7037);
or U9876 (N_9876,N_6369,N_6002);
xnor U9877 (N_9877,N_7908,N_7793);
xor U9878 (N_9878,N_6597,N_7997);
and U9879 (N_9879,N_6362,N_6064);
nor U9880 (N_9880,N_7964,N_7890);
or U9881 (N_9881,N_7614,N_7821);
xor U9882 (N_9882,N_6406,N_7379);
and U9883 (N_9883,N_7091,N_7932);
or U9884 (N_9884,N_7274,N_7260);
xor U9885 (N_9885,N_7267,N_6333);
nor U9886 (N_9886,N_7679,N_6876);
or U9887 (N_9887,N_7349,N_6896);
and U9888 (N_9888,N_7805,N_7460);
nand U9889 (N_9889,N_6280,N_6981);
and U9890 (N_9890,N_6561,N_7622);
xnor U9891 (N_9891,N_6474,N_7489);
nand U9892 (N_9892,N_7025,N_6560);
and U9893 (N_9893,N_6259,N_6661);
xnor U9894 (N_9894,N_6251,N_7320);
and U9895 (N_9895,N_6206,N_7872);
and U9896 (N_9896,N_7089,N_6793);
xnor U9897 (N_9897,N_7803,N_7899);
xor U9898 (N_9898,N_6974,N_6135);
and U9899 (N_9899,N_7243,N_7687);
xnor U9900 (N_9900,N_7831,N_6536);
nand U9901 (N_9901,N_6814,N_7963);
and U9902 (N_9902,N_6425,N_6645);
xnor U9903 (N_9903,N_7395,N_7568);
nor U9904 (N_9904,N_7745,N_7586);
or U9905 (N_9905,N_6972,N_6502);
xnor U9906 (N_9906,N_7489,N_7764);
nor U9907 (N_9907,N_6826,N_6787);
and U9908 (N_9908,N_6161,N_6796);
or U9909 (N_9909,N_7806,N_7084);
and U9910 (N_9910,N_7178,N_7544);
nor U9911 (N_9911,N_7152,N_7885);
and U9912 (N_9912,N_7015,N_6634);
and U9913 (N_9913,N_7689,N_6508);
nand U9914 (N_9914,N_7421,N_6373);
or U9915 (N_9915,N_7913,N_6703);
nand U9916 (N_9916,N_6404,N_6907);
nor U9917 (N_9917,N_7168,N_6537);
xor U9918 (N_9918,N_6791,N_7979);
nand U9919 (N_9919,N_7521,N_6090);
nor U9920 (N_9920,N_7258,N_6065);
nor U9921 (N_9921,N_7454,N_7662);
nand U9922 (N_9922,N_7679,N_6792);
xnor U9923 (N_9923,N_7948,N_6697);
nand U9924 (N_9924,N_6882,N_7860);
or U9925 (N_9925,N_6738,N_7441);
and U9926 (N_9926,N_6493,N_6628);
xor U9927 (N_9927,N_6434,N_7008);
xnor U9928 (N_9928,N_6587,N_6819);
or U9929 (N_9929,N_7386,N_6076);
or U9930 (N_9930,N_7058,N_7783);
or U9931 (N_9931,N_7442,N_7553);
or U9932 (N_9932,N_6481,N_7130);
or U9933 (N_9933,N_6733,N_7763);
nor U9934 (N_9934,N_7772,N_6013);
xor U9935 (N_9935,N_7430,N_6027);
xnor U9936 (N_9936,N_7336,N_7344);
nor U9937 (N_9937,N_6827,N_6266);
and U9938 (N_9938,N_6917,N_6146);
and U9939 (N_9939,N_6100,N_6830);
xor U9940 (N_9940,N_6762,N_7856);
and U9941 (N_9941,N_7780,N_6226);
or U9942 (N_9942,N_7667,N_6532);
nor U9943 (N_9943,N_7260,N_7884);
and U9944 (N_9944,N_6931,N_6433);
nor U9945 (N_9945,N_6498,N_7791);
xnor U9946 (N_9946,N_6894,N_7801);
and U9947 (N_9947,N_7146,N_7942);
or U9948 (N_9948,N_6113,N_6871);
and U9949 (N_9949,N_7474,N_7417);
nor U9950 (N_9950,N_6419,N_7811);
and U9951 (N_9951,N_7272,N_6038);
nand U9952 (N_9952,N_7548,N_7567);
xor U9953 (N_9953,N_6317,N_6300);
and U9954 (N_9954,N_7456,N_6427);
or U9955 (N_9955,N_7352,N_6306);
or U9956 (N_9956,N_6297,N_7428);
nand U9957 (N_9957,N_6490,N_6407);
xnor U9958 (N_9958,N_6434,N_7933);
or U9959 (N_9959,N_6404,N_6139);
xor U9960 (N_9960,N_6087,N_7014);
nor U9961 (N_9961,N_6732,N_7799);
nor U9962 (N_9962,N_6310,N_7015);
or U9963 (N_9963,N_7210,N_6307);
nor U9964 (N_9964,N_6484,N_7015);
nor U9965 (N_9965,N_6051,N_7732);
or U9966 (N_9966,N_6301,N_7800);
or U9967 (N_9967,N_6910,N_7248);
nand U9968 (N_9968,N_7922,N_7527);
nor U9969 (N_9969,N_7653,N_6356);
nand U9970 (N_9970,N_6318,N_7026);
or U9971 (N_9971,N_7149,N_7682);
nor U9972 (N_9972,N_6544,N_7434);
nor U9973 (N_9973,N_6136,N_6006);
nand U9974 (N_9974,N_6266,N_7055);
or U9975 (N_9975,N_6450,N_7162);
or U9976 (N_9976,N_7683,N_6469);
nor U9977 (N_9977,N_7335,N_7652);
xnor U9978 (N_9978,N_7456,N_7263);
nor U9979 (N_9979,N_6604,N_6970);
and U9980 (N_9980,N_6768,N_6607);
or U9981 (N_9981,N_7322,N_7627);
nand U9982 (N_9982,N_6626,N_6146);
nor U9983 (N_9983,N_6243,N_6855);
nand U9984 (N_9984,N_7769,N_6340);
xnor U9985 (N_9985,N_7918,N_7441);
and U9986 (N_9986,N_7829,N_7833);
xnor U9987 (N_9987,N_6622,N_7145);
nor U9988 (N_9988,N_6122,N_7791);
nand U9989 (N_9989,N_7983,N_6222);
or U9990 (N_9990,N_7211,N_6683);
and U9991 (N_9991,N_6866,N_6005);
or U9992 (N_9992,N_7639,N_7272);
nand U9993 (N_9993,N_6362,N_6022);
nand U9994 (N_9994,N_7412,N_6582);
and U9995 (N_9995,N_7446,N_6944);
nand U9996 (N_9996,N_7463,N_7248);
nand U9997 (N_9997,N_6234,N_7600);
and U9998 (N_9998,N_7934,N_6843);
xor U9999 (N_9999,N_6951,N_7015);
nand U10000 (N_10000,N_8194,N_9041);
or U10001 (N_10001,N_8625,N_8677);
xor U10002 (N_10002,N_9449,N_9895);
nor U10003 (N_10003,N_9297,N_8416);
nor U10004 (N_10004,N_8477,N_8041);
and U10005 (N_10005,N_8404,N_8142);
nand U10006 (N_10006,N_8736,N_8353);
nor U10007 (N_10007,N_9771,N_8853);
or U10008 (N_10008,N_8707,N_8400);
xnor U10009 (N_10009,N_9482,N_9524);
and U10010 (N_10010,N_9175,N_9243);
or U10011 (N_10011,N_9138,N_9985);
xnor U10012 (N_10012,N_8760,N_9417);
or U10013 (N_10013,N_8420,N_8044);
and U10014 (N_10014,N_9376,N_9316);
and U10015 (N_10015,N_9997,N_8585);
nand U10016 (N_10016,N_8882,N_8702);
nand U10017 (N_10017,N_8614,N_8491);
nor U10018 (N_10018,N_8822,N_9083);
xor U10019 (N_10019,N_8174,N_9195);
and U10020 (N_10020,N_9352,N_9079);
xor U10021 (N_10021,N_8465,N_9669);
nor U10022 (N_10022,N_8922,N_8438);
nand U10023 (N_10023,N_8936,N_8385);
nand U10024 (N_10024,N_9527,N_9720);
or U10025 (N_10025,N_9535,N_9672);
nor U10026 (N_10026,N_9575,N_8396);
and U10027 (N_10027,N_9455,N_8540);
nand U10028 (N_10028,N_8361,N_9748);
nor U10029 (N_10029,N_9753,N_8535);
and U10030 (N_10030,N_9387,N_8154);
xnor U10031 (N_10031,N_9300,N_8847);
nor U10032 (N_10032,N_8640,N_9879);
xnor U10033 (N_10033,N_8810,N_8428);
and U10034 (N_10034,N_9066,N_8274);
xor U10035 (N_10035,N_9270,N_8074);
nor U10036 (N_10036,N_9391,N_9882);
or U10037 (N_10037,N_8529,N_8413);
or U10038 (N_10038,N_9596,N_8160);
xor U10039 (N_10039,N_9188,N_9705);
xnor U10040 (N_10040,N_9339,N_8580);
and U10041 (N_10041,N_9980,N_8196);
nor U10042 (N_10042,N_9056,N_9650);
nor U10043 (N_10043,N_9583,N_8746);
and U10044 (N_10044,N_8077,N_8402);
and U10045 (N_10045,N_8971,N_9230);
nand U10046 (N_10046,N_8016,N_8935);
xor U10047 (N_10047,N_9335,N_8412);
nor U10048 (N_10048,N_9366,N_9479);
and U10049 (N_10049,N_8342,N_8090);
xor U10050 (N_10050,N_8229,N_8842);
nor U10051 (N_10051,N_8650,N_9186);
nand U10052 (N_10052,N_8287,N_9855);
and U10053 (N_10053,N_8674,N_9279);
nor U10054 (N_10054,N_8830,N_9866);
xor U10055 (N_10055,N_8210,N_8193);
xor U10056 (N_10056,N_9143,N_9172);
xor U10057 (N_10057,N_9151,N_8728);
xor U10058 (N_10058,N_8252,N_8458);
nand U10059 (N_10059,N_9035,N_9309);
nor U10060 (N_10060,N_8864,N_8499);
nand U10061 (N_10061,N_8500,N_8979);
nand U10062 (N_10062,N_8942,N_9989);
nor U10063 (N_10063,N_8398,N_8722);
nand U10064 (N_10064,N_9184,N_8206);
or U10065 (N_10065,N_9197,N_9369);
nand U10066 (N_10066,N_9580,N_8545);
xor U10067 (N_10067,N_9487,N_9465);
nand U10068 (N_10068,N_8275,N_8724);
or U10069 (N_10069,N_8800,N_9847);
nor U10070 (N_10070,N_8656,N_8292);
xor U10071 (N_10071,N_8629,N_8259);
and U10072 (N_10072,N_9337,N_8388);
or U10073 (N_10073,N_9735,N_8363);
nor U10074 (N_10074,N_9658,N_9639);
and U10075 (N_10075,N_9068,N_8757);
nand U10076 (N_10076,N_8321,N_9024);
nand U10077 (N_10077,N_9805,N_8845);
and U10078 (N_10078,N_9183,N_8064);
nand U10079 (N_10079,N_8272,N_8240);
nor U10080 (N_10080,N_9229,N_8813);
nand U10081 (N_10081,N_8909,N_8443);
or U10082 (N_10082,N_8870,N_9646);
nor U10083 (N_10083,N_8941,N_9137);
nor U10084 (N_10084,N_9573,N_8249);
or U10085 (N_10085,N_9690,N_8377);
nor U10086 (N_10086,N_8595,N_8097);
or U10087 (N_10087,N_9264,N_9336);
and U10088 (N_10088,N_9784,N_9221);
nand U10089 (N_10089,N_9797,N_8664);
and U10090 (N_10090,N_8589,N_9707);
and U10091 (N_10091,N_9028,N_8356);
and U10092 (N_10092,N_9237,N_8852);
or U10093 (N_10093,N_8148,N_8890);
nor U10094 (N_10094,N_9131,N_9281);
and U10095 (N_10095,N_9531,N_8308);
xnor U10096 (N_10096,N_8537,N_8043);
xor U10097 (N_10097,N_8780,N_9933);
xnor U10098 (N_10098,N_8565,N_8096);
nor U10099 (N_10099,N_9677,N_9001);
nand U10100 (N_10100,N_8668,N_9925);
xnor U10101 (N_10101,N_8246,N_9547);
xor U10102 (N_10102,N_9263,N_8091);
xnor U10103 (N_10103,N_8965,N_9841);
and U10104 (N_10104,N_9875,N_9042);
or U10105 (N_10105,N_8324,N_8029);
xor U10106 (N_10106,N_9497,N_9863);
nor U10107 (N_10107,N_8508,N_9957);
xnor U10108 (N_10108,N_8302,N_9605);
nand U10109 (N_10109,N_9610,N_8171);
xor U10110 (N_10110,N_8783,N_9528);
nand U10111 (N_10111,N_9766,N_8492);
or U10112 (N_10112,N_9200,N_8348);
nand U10113 (N_10113,N_8968,N_9890);
nor U10114 (N_10114,N_9459,N_9955);
or U10115 (N_10115,N_8118,N_8689);
nand U10116 (N_10116,N_8505,N_9511);
and U10117 (N_10117,N_9351,N_8991);
nor U10118 (N_10118,N_9679,N_9045);
xnor U10119 (N_10119,N_9832,N_8102);
nor U10120 (N_10120,N_8604,N_8989);
or U10121 (N_10121,N_8327,N_9254);
and U10122 (N_10122,N_8109,N_9262);
or U10123 (N_10123,N_8758,N_9236);
and U10124 (N_10124,N_8410,N_9947);
or U10125 (N_10125,N_9606,N_8775);
xnor U10126 (N_10126,N_8226,N_9700);
or U10127 (N_10127,N_9812,N_8141);
and U10128 (N_10128,N_9666,N_9886);
and U10129 (N_10129,N_9092,N_8312);
nand U10130 (N_10130,N_8701,N_8539);
or U10131 (N_10131,N_8378,N_8619);
and U10132 (N_10132,N_9038,N_9681);
xnor U10133 (N_10133,N_9225,N_8268);
and U10134 (N_10134,N_9116,N_9404);
nand U10135 (N_10135,N_8498,N_8352);
nor U10136 (N_10136,N_9238,N_9246);
nor U10137 (N_10137,N_9257,N_8187);
nor U10138 (N_10138,N_8506,N_8571);
nor U10139 (N_10139,N_9443,N_9872);
nand U10140 (N_10140,N_8888,N_8988);
and U10141 (N_10141,N_9394,N_9331);
xnor U10142 (N_10142,N_8713,N_9106);
nor U10143 (N_10143,N_9312,N_8161);
xnor U10144 (N_10144,N_9098,N_8738);
nor U10145 (N_10145,N_9298,N_9108);
nand U10146 (N_10146,N_9828,N_9166);
or U10147 (N_10147,N_8932,N_9570);
nor U10148 (N_10148,N_8820,N_9058);
xnor U10149 (N_10149,N_9086,N_8901);
xor U10150 (N_10150,N_9081,N_8265);
nor U10151 (N_10151,N_9785,N_9842);
or U10152 (N_10152,N_8247,N_8397);
nor U10153 (N_10153,N_9463,N_9897);
nand U10154 (N_10154,N_9428,N_8393);
and U10155 (N_10155,N_9954,N_8264);
nand U10156 (N_10156,N_8328,N_8671);
nand U10157 (N_10157,N_9839,N_8243);
nor U10158 (N_10158,N_9460,N_9619);
and U10159 (N_10159,N_9633,N_8447);
nor U10160 (N_10160,N_9966,N_9661);
xor U10161 (N_10161,N_8787,N_9598);
and U10162 (N_10162,N_8937,N_8111);
xnor U10163 (N_10163,N_8859,N_9837);
xnor U10164 (N_10164,N_8923,N_9220);
xnor U10165 (N_10165,N_9029,N_8216);
nand U10166 (N_10166,N_8086,N_8013);
nand U10167 (N_10167,N_8134,N_9719);
nor U10168 (N_10168,N_9825,N_8336);
and U10169 (N_10169,N_9458,N_9161);
nand U10170 (N_10170,N_9242,N_9003);
and U10171 (N_10171,N_9622,N_9763);
and U10172 (N_10172,N_9426,N_8591);
and U10173 (N_10173,N_9589,N_9304);
xor U10174 (N_10174,N_9268,N_8144);
nor U10175 (N_10175,N_8081,N_8290);
nor U10176 (N_10176,N_8683,N_8358);
nand U10177 (N_10177,N_9370,N_8884);
and U10178 (N_10178,N_8889,N_9569);
nand U10179 (N_10179,N_9908,N_8801);
and U10180 (N_10180,N_9587,N_8954);
xor U10181 (N_10181,N_8285,N_9836);
nand U10182 (N_10182,N_9928,N_8153);
nand U10183 (N_10183,N_9412,N_8547);
nand U10184 (N_10184,N_9416,N_8485);
nand U10185 (N_10185,N_8294,N_9330);
and U10186 (N_10186,N_9942,N_8548);
xor U10187 (N_10187,N_8222,N_9613);
and U10188 (N_10188,N_8912,N_9385);
nor U10189 (N_10189,N_8372,N_9071);
or U10190 (N_10190,N_8568,N_9711);
and U10191 (N_10191,N_9647,N_9436);
and U10192 (N_10192,N_8370,N_9961);
xor U10193 (N_10193,N_8167,N_8108);
nand U10194 (N_10194,N_9920,N_8334);
or U10195 (N_10195,N_8149,N_9571);
xnor U10196 (N_10196,N_9590,N_8362);
xor U10197 (N_10197,N_9219,N_8573);
xnor U10198 (N_10198,N_8974,N_8865);
nand U10199 (N_10199,N_8310,N_9550);
or U10200 (N_10200,N_9861,N_9602);
or U10201 (N_10201,N_8280,N_9764);
or U10202 (N_10202,N_9804,N_9102);
nand U10203 (N_10203,N_8143,N_8957);
nand U10204 (N_10204,N_9938,N_9585);
xor U10205 (N_10205,N_8073,N_9375);
nor U10206 (N_10206,N_9063,N_8110);
xnor U10207 (N_10207,N_9578,N_9181);
nor U10208 (N_10208,N_9680,N_8481);
xor U10209 (N_10209,N_8618,N_8531);
or U10210 (N_10210,N_9149,N_9537);
xnor U10211 (N_10211,N_8592,N_9781);
nand U10212 (N_10212,N_8137,N_9280);
xor U10213 (N_10213,N_9848,N_9626);
or U10214 (N_10214,N_8977,N_8791);
and U10215 (N_10215,N_9256,N_8833);
xor U10216 (N_10216,N_9457,N_8515);
or U10217 (N_10217,N_8387,N_9769);
xor U10218 (N_10218,N_9935,N_8846);
and U10219 (N_10219,N_8424,N_8964);
or U10220 (N_10220,N_8414,N_9329);
xor U10221 (N_10221,N_9860,N_9770);
and U10222 (N_10222,N_9345,N_8533);
or U10223 (N_10223,N_9683,N_9208);
or U10224 (N_10224,N_8227,N_9393);
and U10225 (N_10225,N_9233,N_8101);
nand U10226 (N_10226,N_9902,N_8215);
nor U10227 (N_10227,N_8705,N_8245);
nand U10228 (N_10228,N_9498,N_9165);
xor U10229 (N_10229,N_9651,N_8770);
nand U10230 (N_10230,N_8814,N_9155);
or U10231 (N_10231,N_9572,N_9892);
or U10232 (N_10232,N_9541,N_8475);
and U10233 (N_10233,N_8019,N_8335);
or U10234 (N_10234,N_9721,N_9378);
nor U10235 (N_10235,N_9507,N_9338);
and U10236 (N_10236,N_9654,N_9964);
and U10237 (N_10237,N_8711,N_8848);
and U10238 (N_10238,N_8927,N_8175);
xor U10239 (N_10239,N_8376,N_8703);
xor U10240 (N_10240,N_9873,N_8311);
nor U10241 (N_10241,N_9128,N_9552);
or U10242 (N_10242,N_9125,N_8751);
nor U10243 (N_10243,N_8764,N_9745);
or U10244 (N_10244,N_9868,N_9940);
or U10245 (N_10245,N_9075,N_8559);
and U10246 (N_10246,N_8960,N_9776);
and U10247 (N_10247,N_8896,N_9461);
and U10248 (N_10248,N_8777,N_8809);
or U10249 (N_10249,N_8962,N_9348);
and U10250 (N_10250,N_8762,N_9517);
or U10251 (N_10251,N_9044,N_8135);
nand U10252 (N_10252,N_8295,N_9931);
xnor U10253 (N_10253,N_9365,N_9379);
nor U10254 (N_10254,N_9704,N_9815);
or U10255 (N_10255,N_8718,N_8902);
nand U10256 (N_10256,N_9388,N_9314);
and U10257 (N_10257,N_8769,N_9693);
nor U10258 (N_10258,N_9290,N_9820);
and U10259 (N_10259,N_9010,N_8065);
nor U10260 (N_10260,N_9642,N_8596);
or U10261 (N_10261,N_8451,N_8201);
or U10262 (N_10262,N_9976,N_8433);
nand U10263 (N_10263,N_9429,N_8799);
nor U10264 (N_10264,N_9641,N_8474);
xor U10265 (N_10265,N_8798,N_9409);
or U10266 (N_10266,N_8049,N_9193);
or U10267 (N_10267,N_8928,N_8934);
nand U10268 (N_10268,N_9757,N_8919);
nor U10269 (N_10269,N_9918,N_8641);
nor U10270 (N_10270,N_8445,N_8435);
and U10271 (N_10271,N_9601,N_8234);
nand U10272 (N_10272,N_9067,N_8841);
or U10273 (N_10273,N_8033,N_8710);
nor U10274 (N_10274,N_8569,N_9134);
and U10275 (N_10275,N_8861,N_9983);
or U10276 (N_10276,N_9526,N_9085);
nand U10277 (N_10277,N_8808,N_8862);
and U10278 (N_10278,N_9147,N_9286);
xnor U10279 (N_10279,N_9939,N_9756);
xnor U10280 (N_10280,N_8634,N_9509);
and U10281 (N_10281,N_8384,N_8779);
nor U10282 (N_10282,N_8098,N_9169);
or U10283 (N_10283,N_9213,N_9525);
nand U10284 (N_10284,N_8028,N_8299);
nand U10285 (N_10285,N_9712,N_8084);
nor U10286 (N_10286,N_8686,N_9419);
nor U10287 (N_10287,N_9470,N_8784);
xnor U10288 (N_10288,N_8440,N_8891);
xnor U10289 (N_10289,N_8966,N_9854);
xor U10290 (N_10290,N_9907,N_8453);
and U10291 (N_10291,N_9791,N_8908);
nor U10292 (N_10292,N_8817,N_8341);
or U10293 (N_10293,N_8254,N_8422);
nor U10294 (N_10294,N_8078,N_9135);
xor U10295 (N_10295,N_8622,N_9826);
and U10296 (N_10296,N_9730,N_9343);
and U10297 (N_10297,N_9311,N_9456);
xor U10298 (N_10298,N_8766,N_9747);
and U10299 (N_10299,N_9414,N_8646);
or U10300 (N_10300,N_9153,N_9802);
xnor U10301 (N_10301,N_8603,N_9779);
or U10302 (N_10302,N_9054,N_8637);
nand U10303 (N_10303,N_9755,N_9951);
or U10304 (N_10304,N_8827,N_9157);
nor U10305 (N_10305,N_8442,N_8000);
or U10306 (N_10306,N_9708,N_8129);
xnor U10307 (N_10307,N_8522,N_8463);
nor U10308 (N_10308,N_9732,N_8288);
nor U10309 (N_10309,N_9126,N_9501);
and U10310 (N_10310,N_8776,N_8651);
xnor U10311 (N_10311,N_8164,N_8998);
nand U10312 (N_10312,N_8031,N_9005);
xor U10313 (N_10313,N_8690,N_8587);
and U10314 (N_10314,N_9052,N_9260);
nor U10315 (N_10315,N_9678,N_9689);
xor U10316 (N_10316,N_8552,N_8836);
nor U10317 (N_10317,N_8790,N_8553);
or U10318 (N_10318,N_8205,N_9726);
and U10319 (N_10319,N_8733,N_8649);
nand U10320 (N_10320,N_9586,N_8911);
or U10321 (N_10321,N_8200,N_8369);
xor U10322 (N_10322,N_8570,N_9555);
and U10323 (N_10323,N_8807,N_9725);
and U10324 (N_10324,N_9880,N_8642);
nand U10325 (N_10325,N_8879,N_9293);
nand U10326 (N_10326,N_9970,N_8439);
nor U10327 (N_10327,N_8743,N_8658);
xnor U10328 (N_10328,N_9364,N_8296);
and U10329 (N_10329,N_8399,N_9353);
or U10330 (N_10330,N_9673,N_9563);
and U10331 (N_10331,N_9949,N_8339);
nand U10332 (N_10332,N_8507,N_9518);
or U10333 (N_10333,N_9729,N_8150);
xnor U10334 (N_10334,N_9561,N_9333);
xnor U10335 (N_10335,N_9495,N_8693);
xor U10336 (N_10336,N_8875,N_8963);
or U10337 (N_10337,N_9798,N_8316);
xor U10338 (N_10338,N_9018,N_9473);
nand U10339 (N_10339,N_8297,N_9201);
xnor U10340 (N_10340,N_9808,N_8730);
or U10341 (N_10341,N_9354,N_9621);
and U10342 (N_10342,N_9142,N_8237);
xnor U10343 (N_10343,N_8903,N_9810);
nand U10344 (N_10344,N_8696,N_9405);
xor U10345 (N_10345,N_9255,N_8347);
xnor U10346 (N_10346,N_9205,N_9087);
and U10347 (N_10347,N_8325,N_8156);
nor U10348 (N_10348,N_9715,N_8995);
xnor U10349 (N_10349,N_8961,N_8095);
or U10350 (N_10350,N_9196,N_9272);
or U10351 (N_10351,N_9653,N_9037);
or U10352 (N_10352,N_9009,N_9752);
xnor U10353 (N_10353,N_9817,N_9656);
xnor U10354 (N_10354,N_8929,N_8030);
xor U10355 (N_10355,N_8228,N_9995);
and U10356 (N_10356,N_8250,N_9629);
nand U10357 (N_10357,N_8943,N_8262);
xor U10358 (N_10358,N_8138,N_9987);
or U10359 (N_10359,N_8546,N_8871);
nand U10360 (N_10360,N_8434,N_9556);
or U10361 (N_10361,N_8409,N_8906);
or U10362 (N_10362,N_8562,N_9581);
nor U10363 (N_10363,N_9437,N_8967);
or U10364 (N_10364,N_9988,N_8124);
or U10365 (N_10365,N_9212,N_8615);
nor U10366 (N_10366,N_9332,N_8389);
nand U10367 (N_10367,N_9099,N_9508);
xnor U10368 (N_10368,N_8613,N_9540);
xnor U10369 (N_10369,N_9624,N_9905);
nor U10370 (N_10370,N_9140,N_8804);
nor U10371 (N_10371,N_8269,N_9034);
nor U10372 (N_10372,N_9751,N_8765);
and U10373 (N_10373,N_9051,N_9662);
nor U10374 (N_10374,N_8687,N_8232);
or U10375 (N_10375,N_8876,N_9317);
or U10376 (N_10376,N_9671,N_9060);
nand U10377 (N_10377,N_8047,N_9380);
nand U10378 (N_10378,N_9840,N_9634);
nand U10379 (N_10379,N_8430,N_9289);
and U10380 (N_10380,N_8127,N_8886);
or U10381 (N_10381,N_9844,N_9883);
nand U10382 (N_10382,N_8005,N_8106);
xnor U10383 (N_10383,N_8856,N_9189);
nand U10384 (N_10384,N_8825,N_9865);
nand U10385 (N_10385,N_8218,N_9475);
or U10386 (N_10386,N_9046,N_8018);
nand U10387 (N_10387,N_9676,N_8293);
or U10388 (N_10388,N_8759,N_8555);
xor U10389 (N_10389,N_8997,N_9059);
and U10390 (N_10390,N_9522,N_8694);
or U10391 (N_10391,N_9228,N_8350);
and U10392 (N_10392,N_9386,N_9446);
nor U10393 (N_10393,N_8209,N_9418);
nand U10394 (N_10394,N_9400,N_9699);
xnor U10395 (N_10395,N_8238,N_8828);
or U10396 (N_10396,N_9340,N_8550);
nor U10397 (N_10397,N_8819,N_8415);
xnor U10398 (N_10398,N_8607,N_8744);
or U10399 (N_10399,N_8107,N_8584);
nand U10400 (N_10400,N_9623,N_8955);
or U10401 (N_10401,N_8038,N_9782);
nand U10402 (N_10402,N_8920,N_8857);
nor U10403 (N_10403,N_8147,N_9471);
xor U10404 (N_10404,N_8797,N_8305);
xnor U10405 (N_10405,N_9282,N_9628);
and U10406 (N_10406,N_9795,N_9334);
nor U10407 (N_10407,N_9870,N_8831);
or U10408 (N_10408,N_9121,N_9274);
xor U10409 (N_10409,N_8322,N_9894);
nor U10410 (N_10410,N_9834,N_8289);
nor U10411 (N_10411,N_8680,N_9991);
nand U10412 (N_10412,N_8873,N_8145);
nor U10413 (N_10413,N_8993,N_9218);
and U10414 (N_10414,N_9724,N_8382);
nor U10415 (N_10415,N_9788,N_9105);
xnor U10416 (N_10416,N_8394,N_8586);
or U10417 (N_10417,N_8843,N_8741);
and U10418 (N_10418,N_8576,N_9271);
xor U10419 (N_10419,N_9807,N_8560);
and U10420 (N_10420,N_8538,N_8661);
nand U10421 (N_10421,N_9900,N_8554);
and U10422 (N_10422,N_8682,N_9123);
nor U10423 (N_10423,N_8956,N_8978);
and U10424 (N_10424,N_9247,N_8017);
or U10425 (N_10425,N_8583,N_8307);
or U10426 (N_10426,N_9319,N_8916);
nor U10427 (N_10427,N_8300,N_9668);
nor U10428 (N_10428,N_8610,N_9911);
and U10429 (N_10429,N_9420,N_9288);
or U10430 (N_10430,N_9864,N_8103);
nand U10431 (N_10431,N_9395,N_8419);
xnor U10432 (N_10432,N_8714,N_9206);
or U10433 (N_10433,N_8893,N_8892);
nor U10434 (N_10434,N_9222,N_8020);
or U10435 (N_10435,N_8915,N_9898);
or U10436 (N_10436,N_9521,N_9554);
or U10437 (N_10437,N_9937,N_8898);
and U10438 (N_10438,N_9069,N_8128);
nand U10439 (N_10439,N_8716,N_8260);
and U10440 (N_10440,N_9148,N_8599);
nand U10441 (N_10441,N_9697,N_8931);
and U10442 (N_10442,N_8072,N_9950);
nand U10443 (N_10443,N_8944,N_8803);
and U10444 (N_10444,N_8100,N_8125);
nor U10445 (N_10445,N_8959,N_9593);
and U10446 (N_10446,N_9396,N_9091);
nand U10447 (N_10447,N_9974,N_8905);
or U10448 (N_10448,N_9434,N_8794);
nand U10449 (N_10449,N_9885,N_8623);
or U10450 (N_10450,N_8720,N_8076);
or U10451 (N_10451,N_8318,N_9506);
or U10452 (N_10452,N_9778,N_8704);
nor U10453 (N_10453,N_8345,N_9047);
nand U10454 (N_10454,N_9454,N_8126);
or U10455 (N_10455,N_9122,N_9287);
and U10456 (N_10456,N_8326,N_8725);
and U10457 (N_10457,N_9248,N_9292);
nor U10458 (N_10458,N_9793,N_9551);
xor U10459 (N_10459,N_9179,N_9941);
nor U10460 (N_10460,N_8910,N_9849);
and U10461 (N_10461,N_9965,N_8364);
or U10462 (N_10462,N_9407,N_9829);
or U10463 (N_10463,N_9856,N_9533);
or U10464 (N_10464,N_9273,N_9294);
nor U10465 (N_10465,N_8981,N_8717);
nor U10466 (N_10466,N_8904,N_8181);
nand U10467 (N_10467,N_9207,N_9644);
nor U10468 (N_10468,N_8510,N_9096);
nand U10469 (N_10469,N_8631,N_9484);
nor U10470 (N_10470,N_8391,N_9100);
nand U10471 (N_10471,N_8368,N_8926);
nor U10472 (N_10472,N_9927,N_9660);
xor U10473 (N_10473,N_8130,N_9000);
and U10474 (N_10474,N_8781,N_9251);
and U10475 (N_10475,N_8566,N_9768);
and U10476 (N_10476,N_8869,N_9504);
nor U10477 (N_10477,N_8365,N_8407);
nand U10478 (N_10478,N_9692,N_8745);
or U10479 (N_10479,N_9845,N_8627);
nand U10480 (N_10480,N_9478,N_9210);
xor U10481 (N_10481,N_8444,N_9015);
and U10482 (N_10482,N_8528,N_9969);
nor U10483 (N_10483,N_8858,N_9869);
and U10484 (N_10484,N_8574,N_9984);
and U10485 (N_10485,N_8040,N_9211);
and U10486 (N_10486,N_9916,N_9967);
nand U10487 (N_10487,N_9891,N_8740);
and U10488 (N_10488,N_8773,N_8582);
nor U10489 (N_10489,N_8524,N_8520);
and U10490 (N_10490,N_9761,N_9406);
nor U10491 (N_10491,N_9496,N_8454);
nand U10492 (N_10492,N_9801,N_9141);
nand U10493 (N_10493,N_8752,N_9536);
or U10494 (N_10494,N_9235,N_9819);
and U10495 (N_10495,N_9538,N_9408);
xnor U10496 (N_10496,N_8511,N_9686);
nor U10497 (N_10497,N_9452,N_9190);
nand U10498 (N_10498,N_8806,N_9026);
xnor U10499 (N_10499,N_9162,N_8421);
nor U10500 (N_10500,N_8700,N_8980);
or U10501 (N_10501,N_8006,N_9846);
nand U10502 (N_10502,N_9088,N_9367);
nor U10503 (N_10503,N_9636,N_8277);
or U10504 (N_10504,N_9505,N_9652);
or U10505 (N_10505,N_9901,N_9737);
and U10506 (N_10506,N_8344,N_8159);
and U10507 (N_10507,N_8390,N_9982);
and U10508 (N_10508,N_8180,N_8832);
nand U10509 (N_10509,N_9553,N_9565);
nand U10510 (N_10510,N_8986,N_9226);
and U10511 (N_10511,N_8225,N_8854);
nor U10512 (N_10512,N_8530,N_8542);
nor U10513 (N_10513,N_9953,N_8633);
xnor U10514 (N_10514,N_8496,N_9800);
nor U10515 (N_10515,N_8881,N_9684);
and U10516 (N_10516,N_8897,N_8406);
nor U10517 (N_10517,N_8329,N_9117);
and U10518 (N_10518,N_9382,N_8835);
nor U10519 (N_10519,N_9932,N_8900);
nor U10520 (N_10520,N_9291,N_8793);
or U10521 (N_10521,N_8802,N_9604);
xor U10522 (N_10522,N_8557,N_9811);
nand U10523 (N_10523,N_9564,N_9410);
and U10524 (N_10524,N_9780,N_9082);
nand U10525 (N_10525,N_8785,N_9363);
nor U10526 (N_10526,N_9609,N_9612);
nand U10527 (N_10527,N_8315,N_8467);
and U10528 (N_10528,N_9577,N_9914);
or U10529 (N_10529,N_8611,N_9874);
and U10530 (N_10530,N_9835,N_8155);
nor U10531 (N_10531,N_8208,N_8374);
nand U10532 (N_10532,N_9285,N_8089);
or U10533 (N_10533,N_8670,N_9198);
nand U10534 (N_10534,N_9906,N_8712);
and U10535 (N_10535,N_8617,N_9002);
nor U10536 (N_10536,N_9948,N_9742);
or U10537 (N_10537,N_8612,N_8070);
or U10538 (N_10538,N_9635,N_8829);
and U10539 (N_10539,N_8340,N_9614);
nand U10540 (N_10540,N_8534,N_9853);
nor U10541 (N_10541,N_9607,N_8184);
xnor U10542 (N_10542,N_8476,N_8645);
xnor U10543 (N_10543,N_8355,N_8025);
xor U10544 (N_10544,N_8446,N_8958);
nor U10545 (N_10545,N_9040,N_8450);
nor U10546 (N_10546,N_8590,N_9266);
and U10547 (N_10547,N_9451,N_8068);
nor U10548 (N_10548,N_9350,N_9532);
nor U10549 (N_10549,N_9231,N_8742);
or U10550 (N_10550,N_8037,N_8952);
nand U10551 (N_10551,N_8004,N_8114);
or U10552 (N_10552,N_8009,N_8244);
or U10553 (N_10553,N_8053,N_9008);
or U10554 (N_10554,N_9960,N_8449);
nor U10555 (N_10555,N_9594,N_8452);
nor U10556 (N_10556,N_9232,N_8314);
xor U10557 (N_10557,N_9489,N_9741);
or U10558 (N_10558,N_8213,N_8202);
nand U10559 (N_10559,N_8046,N_9944);
and U10560 (N_10560,N_9031,N_8189);
or U10561 (N_10561,N_8563,N_9084);
nor U10562 (N_10562,N_8039,N_8940);
or U10563 (N_10563,N_8578,N_8121);
or U10564 (N_10564,N_8052,N_9758);
and U10565 (N_10565,N_9978,N_9315);
xnor U10566 (N_10566,N_9664,N_9341);
nand U10567 (N_10567,N_9772,N_9549);
and U10568 (N_10568,N_8605,N_9512);
nor U10569 (N_10569,N_8544,N_8480);
xor U10570 (N_10570,N_8644,N_9267);
nor U10571 (N_10571,N_9011,N_9740);
nand U10572 (N_10572,N_9548,N_9346);
nand U10573 (N_10573,N_9464,N_9881);
and U10574 (N_10574,N_9284,N_8178);
nand U10575 (N_10575,N_9145,N_8839);
or U10576 (N_10576,N_8036,N_9381);
or U10577 (N_10577,N_9278,N_8251);
nor U10578 (N_10578,N_9033,N_8373);
nor U10579 (N_10579,N_8723,N_9558);
xor U10580 (N_10580,N_9321,N_8976);
nor U10581 (N_10581,N_9822,N_8165);
nand U10582 (N_10582,N_9307,N_8085);
nor U10583 (N_10583,N_9023,N_8063);
and U10584 (N_10584,N_9713,N_9889);
and U10585 (N_10585,N_9515,N_9792);
and U10586 (N_10586,N_9696,N_9775);
or U10587 (N_10587,N_9996,N_9803);
or U10588 (N_10588,N_8431,N_8183);
or U10589 (N_10589,N_9185,N_9600);
and U10590 (N_10590,N_8306,N_9727);
or U10591 (N_10591,N_9127,N_8045);
nand U10592 (N_10592,N_9733,N_8197);
and U10593 (N_10593,N_8732,N_9477);
nand U10594 (N_10594,N_9994,N_9783);
or U10595 (N_10595,N_9717,N_8392);
or U10596 (N_10596,N_9576,N_9513);
and U10597 (N_10597,N_8338,N_9592);
nand U10598 (N_10598,N_8756,N_9422);
nor U10599 (N_10599,N_9357,N_8495);
nand U10600 (N_10600,N_8666,N_9017);
nor U10601 (N_10601,N_8456,N_9912);
nand U10602 (N_10602,N_9224,N_9530);
nor U10603 (N_10603,N_9180,N_8172);
or U10604 (N_10604,N_8517,N_8973);
or U10605 (N_10605,N_8750,N_9899);
and U10606 (N_10606,N_8709,N_9397);
nor U10607 (N_10607,N_8080,N_8291);
nand U10608 (N_10608,N_8034,N_9915);
nand U10609 (N_10609,N_8556,N_8731);
xnor U10610 (N_10610,N_9129,N_8581);
or U10611 (N_10611,N_8518,N_9234);
nor U10612 (N_10612,N_8448,N_9977);
nand U10613 (N_10613,N_9492,N_9615);
and U10614 (N_10614,N_9425,N_9992);
or U10615 (N_10615,N_9631,N_9637);
nor U10616 (N_10616,N_8092,N_8163);
nor U10617 (N_10617,N_8608,N_8620);
or U10618 (N_10618,N_8015,N_8488);
or U10619 (N_10619,N_8279,N_9261);
xnor U10620 (N_10620,N_9486,N_8616);
or U10621 (N_10621,N_9043,N_8951);
or U10622 (N_10622,N_9318,N_9209);
nand U10623 (N_10623,N_9119,N_9356);
nor U10624 (N_10624,N_9358,N_8918);
nor U10625 (N_10625,N_8117,N_8636);
nand U10626 (N_10626,N_9245,N_9675);
nor U10627 (N_10627,N_9476,N_9302);
nor U10628 (N_10628,N_9144,N_8665);
nand U10629 (N_10629,N_8504,N_9736);
nor U10630 (N_10630,N_9919,N_9738);
and U10631 (N_10631,N_9199,N_8685);
or U10632 (N_10632,N_9373,N_9794);
nor U10633 (N_10633,N_8459,N_9691);
nand U10634 (N_10634,N_9990,N_9164);
nand U10635 (N_10635,N_9130,N_9702);
and U10636 (N_10636,N_8598,N_9986);
xnor U10637 (N_10637,N_8628,N_9467);
nor U10638 (N_10638,N_9076,N_9862);
and U10639 (N_10639,N_9444,N_9584);
nand U10640 (N_10640,N_9057,N_8014);
or U10641 (N_10641,N_8708,N_8002);
nor U10642 (N_10642,N_8643,N_8333);
nor U10643 (N_10643,N_8432,N_9021);
nand U10644 (N_10644,N_9665,N_9731);
nand U10645 (N_10645,N_9006,N_9152);
xnor U10646 (N_10646,N_9275,N_9399);
nand U10647 (N_10647,N_8478,N_8008);
nand U10648 (N_10648,N_9830,N_9722);
nor U10649 (N_10649,N_9176,N_8286);
and U10650 (N_10650,N_9806,N_8648);
and U10651 (N_10651,N_9620,N_9217);
nor U10652 (N_10652,N_9714,N_9299);
nor U10653 (N_10653,N_9616,N_9560);
or U10654 (N_10654,N_9946,N_8626);
or U10655 (N_10655,N_8177,N_8913);
and U10656 (N_10656,N_8460,N_9439);
nor U10657 (N_10657,N_8021,N_8660);
nand U10658 (N_10658,N_8071,N_8173);
xnor U10659 (N_10659,N_8236,N_9061);
or U10660 (N_10660,N_8099,N_9502);
or U10661 (N_10661,N_9158,N_8734);
xor U10662 (N_10662,N_8868,N_9080);
nor U10663 (N_10663,N_9643,N_9111);
or U10664 (N_10664,N_9566,N_8022);
nor U10665 (N_10665,N_8461,N_8921);
and U10666 (N_10666,N_8470,N_9789);
nand U10667 (N_10667,N_8663,N_8561);
nor U10668 (N_10668,N_8055,N_8152);
nand U10669 (N_10669,N_9625,N_9999);
nand U10670 (N_10670,N_9754,N_9136);
nand U10671 (N_10671,N_9240,N_9706);
or U10672 (N_10672,N_8657,N_9962);
and U10673 (N_10673,N_9481,N_8468);
nand U10674 (N_10674,N_8270,N_9402);
xor U10675 (N_10675,N_9790,N_9632);
xor U10676 (N_10676,N_9368,N_9638);
nand U10677 (N_10677,N_8168,N_9545);
xnor U10678 (N_10678,N_9124,N_8749);
nor U10679 (N_10679,N_9876,N_8681);
nand U10680 (N_10680,N_8985,N_8987);
and U10681 (N_10681,N_9816,N_8190);
or U10682 (N_10682,N_8471,N_8123);
or U10683 (N_10683,N_9952,N_8692);
nor U10684 (N_10684,N_8990,N_9973);
or U10685 (N_10685,N_8675,N_9253);
or U10686 (N_10686,N_8472,N_9739);
and U10687 (N_10687,N_9909,N_9214);
xnor U10688 (N_10688,N_9173,N_9688);
xor U10689 (N_10689,N_8360,N_8982);
nor U10690 (N_10690,N_8624,N_8838);
nand U10691 (N_10691,N_9546,N_9039);
or U10692 (N_10692,N_9469,N_8812);
nor U10693 (N_10693,N_8261,N_9617);
or U10694 (N_10694,N_9759,N_9359);
or U10695 (N_10695,N_9320,N_9384);
nand U10696 (N_10696,N_9904,N_8217);
nor U10697 (N_10697,N_9857,N_8371);
nand U10698 (N_10698,N_9159,N_9579);
or U10699 (N_10699,N_9283,N_9433);
nor U10700 (N_10700,N_8188,N_8815);
and U10701 (N_10701,N_8179,N_8062);
nand U10702 (N_10702,N_9361,N_8659);
or U10703 (N_10703,N_8753,N_9659);
nand U10704 (N_10704,N_8069,N_9910);
nand U10705 (N_10705,N_8309,N_8662);
or U10706 (N_10706,N_8087,N_8354);
nor U10707 (N_10707,N_9120,N_9597);
and U10708 (N_10708,N_9215,N_8054);
nor U10709 (N_10709,N_9389,N_8536);
xnor U10710 (N_10710,N_9055,N_9171);
nor U10711 (N_10711,N_8494,N_8051);
nor U10712 (N_10712,N_8204,N_8593);
xor U10713 (N_10713,N_9796,N_8357);
nand U10714 (N_10714,N_9743,N_8737);
nor U10715 (N_10715,N_9520,N_9833);
nor U10716 (N_10716,N_8575,N_8317);
xor U10717 (N_10717,N_9250,N_8747);
or U10718 (N_10718,N_8023,N_9663);
nand U10719 (N_10719,N_9377,N_8771);
and U10720 (N_10720,N_9956,N_8320);
xor U10721 (N_10721,N_9030,N_8116);
or U10722 (N_10722,N_8375,N_8304);
xnor U10723 (N_10723,N_8949,N_8198);
nand U10724 (N_10724,N_9649,N_8950);
nand U10725 (N_10725,N_8332,N_8169);
and U10726 (N_10726,N_9252,N_8816);
and U10727 (N_10727,N_9390,N_8899);
and U10728 (N_10728,N_8525,N_9095);
and U10729 (N_10729,N_9971,N_8667);
and U10730 (N_10730,N_8104,N_8170);
or U10731 (N_10731,N_9296,N_9827);
xor U10732 (N_10732,N_8464,N_9202);
or U10733 (N_10733,N_8429,N_9070);
and U10734 (N_10734,N_8767,N_9981);
nand U10735 (N_10735,N_8241,N_9327);
or U10736 (N_10736,N_8684,N_8239);
nor U10737 (N_10737,N_9878,N_9744);
nand U10738 (N_10738,N_9322,N_8067);
nor U10739 (N_10739,N_9588,N_8735);
and U10740 (N_10740,N_9611,N_9896);
nor U10741 (N_10741,N_9884,N_8782);
and U10742 (N_10742,N_8012,N_9328);
and U10743 (N_10743,N_8359,N_8248);
nand U10744 (N_10744,N_9618,N_8418);
xor U10745 (N_10745,N_8214,N_9993);
and U10746 (N_10746,N_8509,N_9277);
nor U10747 (N_10747,N_8706,N_8632);
nand U10748 (N_10748,N_8223,N_9746);
or U10749 (N_10749,N_8242,N_9773);
nand U10750 (N_10750,N_9851,N_9723);
nor U10751 (N_10751,N_9227,N_9074);
or U10752 (N_10752,N_9648,N_9716);
and U10753 (N_10753,N_9645,N_9667);
nand U10754 (N_10754,N_8946,N_8878);
nor U10755 (N_10755,N_8818,N_8441);
or U10756 (N_10756,N_9118,N_8212);
nand U10757 (N_10757,N_8423,N_9582);
nor U10758 (N_10758,N_9929,N_9774);
or U10759 (N_10759,N_9191,N_8652);
xor U10760 (N_10760,N_9424,N_9466);
and U10761 (N_10761,N_9401,N_8337);
or U10762 (N_10762,N_8513,N_8796);
or U10763 (N_10763,N_9787,N_9073);
and U10764 (N_10764,N_9187,N_8602);
or U10765 (N_10765,N_9813,N_8778);
nor U10766 (N_10766,N_8609,N_9170);
nand U10767 (N_10767,N_9194,N_8883);
or U10768 (N_10768,N_8379,N_8930);
and U10769 (N_10769,N_8276,N_8403);
or U10770 (N_10770,N_9877,N_8748);
or U10771 (N_10771,N_8343,N_9265);
xnor U10772 (N_10772,N_9519,N_8366);
nand U10773 (N_10773,N_8754,N_9305);
and U10774 (N_10774,N_9510,N_9818);
or U10775 (N_10775,N_9921,N_8837);
nor U10776 (N_10776,N_9146,N_8486);
or U10777 (N_10777,N_8131,N_8866);
and U10778 (N_10778,N_8219,N_8011);
or U10779 (N_10779,N_9657,N_8466);
and U10780 (N_10780,N_8235,N_9523);
and U10781 (N_10781,N_8427,N_8877);
and U10782 (N_10782,N_8256,N_8933);
xor U10783 (N_10783,N_8093,N_8655);
nor U10784 (N_10784,N_8514,N_8729);
xor U10785 (N_10785,N_8113,N_8082);
nor U10786 (N_10786,N_8411,N_8319);
or U10787 (N_10787,N_9403,N_8597);
nor U10788 (N_10788,N_8146,N_9216);
and U10789 (N_10789,N_9514,N_9362);
xnor U10790 (N_10790,N_8855,N_9934);
and U10791 (N_10791,N_9103,N_9843);
and U10792 (N_10792,N_8698,N_8255);
nor U10793 (N_10793,N_8405,N_9809);
nand U10794 (N_10794,N_8887,N_8695);
nand U10795 (N_10795,N_9703,N_8699);
nor U10796 (N_10796,N_8715,N_8437);
nor U10797 (N_10797,N_9415,N_9421);
xnor U10798 (N_10798,N_8726,N_9821);
and U10799 (N_10799,N_8283,N_8349);
and U10800 (N_10800,N_9344,N_9603);
nor U10801 (N_10801,N_9930,N_9310);
xnor U10802 (N_10802,N_8795,N_8323);
nor U10803 (N_10803,N_9326,N_8298);
xnor U10804 (N_10804,N_8947,N_8455);
nand U10805 (N_10805,N_9640,N_9490);
nor U10806 (N_10806,N_9968,N_9871);
and U10807 (N_10807,N_8768,N_8805);
or U10808 (N_10808,N_8301,N_8057);
xor U10809 (N_10809,N_8840,N_9922);
nor U10810 (N_10810,N_8523,N_9445);
xnor U10811 (N_10811,N_9539,N_9064);
xor U10812 (N_10812,N_8482,N_8351);
xnor U10813 (N_10813,N_9019,N_8639);
xor U10814 (N_10814,N_8874,N_8024);
or U10815 (N_10815,N_9695,N_9867);
and U10816 (N_10816,N_9674,N_9072);
and U10817 (N_10817,N_9823,N_9516);
xor U10818 (N_10818,N_9053,N_9500);
xor U10819 (N_10819,N_9132,N_9347);
and U10820 (N_10820,N_8691,N_9503);
xnor U10821 (N_10821,N_8233,N_8151);
or U10822 (N_10822,N_8638,N_9483);
or U10823 (N_10823,N_9112,N_8948);
or U10824 (N_10824,N_9150,N_9110);
nor U10825 (N_10825,N_8823,N_8983);
or U10826 (N_10826,N_8772,N_8939);
nand U10827 (N_10827,N_8469,N_8195);
nor U10828 (N_10828,N_8792,N_8221);
or U10829 (N_10829,N_9423,N_8001);
nor U10830 (N_10830,N_9480,N_8789);
nand U10831 (N_10831,N_9655,N_9694);
or U10832 (N_10832,N_8426,N_8266);
or U10833 (N_10833,N_8493,N_9027);
nor U10834 (N_10834,N_9852,N_8122);
or U10835 (N_10835,N_9160,N_8501);
xor U10836 (N_10836,N_9687,N_8678);
nand U10837 (N_10837,N_8157,N_9682);
xnor U10838 (N_10838,N_8516,N_8140);
nand U10839 (N_10839,N_8061,N_8761);
or U10840 (N_10840,N_8577,N_9430);
xnor U10841 (N_10841,N_9192,N_8996);
xnor U10842 (N_10842,N_9427,N_9168);
and U10843 (N_10843,N_9371,N_9308);
xor U10844 (N_10844,N_9411,N_9133);
and U10845 (N_10845,N_8083,N_9392);
and U10846 (N_10846,N_8386,N_9050);
nand U10847 (N_10847,N_8924,N_9831);
nand U10848 (N_10848,N_9670,N_8673);
xnor U10849 (N_10849,N_8588,N_9355);
or U10850 (N_10850,N_8331,N_8786);
nor U10851 (N_10851,N_8105,N_9453);
xor U10852 (N_10852,N_8938,N_8497);
xor U10853 (N_10853,N_9917,N_9438);
and U10854 (N_10854,N_8278,N_9777);
xnor U10855 (N_10855,N_9107,N_9499);
and U10856 (N_10856,N_8558,N_9824);
nand U10857 (N_10857,N_9204,N_8088);
xnor U10858 (N_10858,N_8925,N_9007);
nand U10859 (N_10859,N_9959,N_9269);
nor U10860 (N_10860,N_8479,N_9032);
xnor U10861 (N_10861,N_9077,N_9474);
nand U10862 (N_10862,N_8543,N_8526);
nand U10863 (N_10863,N_8788,N_9016);
or U10864 (N_10864,N_8056,N_8600);
xor U10865 (N_10865,N_8273,N_8885);
xor U10866 (N_10866,N_8824,N_9698);
nor U10867 (N_10867,N_8192,N_8721);
and U10868 (N_10868,N_8872,N_8303);
or U10869 (N_10869,N_9462,N_9276);
xnor U10870 (N_10870,N_8257,N_9924);
xor U10871 (N_10871,N_9013,N_9435);
nor U10872 (N_10872,N_8503,N_8211);
xor U10873 (N_10873,N_8263,N_8763);
nor U10874 (N_10874,N_8203,N_9440);
nand U10875 (N_10875,N_8462,N_9599);
and U10876 (N_10876,N_8672,N_9945);
nor U10877 (N_10877,N_9114,N_9529);
nor U10878 (N_10878,N_8042,N_9244);
nor U10879 (N_10879,N_9090,N_9078);
and U10880 (N_10880,N_9383,N_9223);
or U10881 (N_10881,N_9557,N_8688);
xnor U10882 (N_10882,N_8953,N_8473);
or U10883 (N_10883,N_8572,N_9295);
or U10884 (N_10884,N_9089,N_8880);
xnor U10885 (N_10885,N_9494,N_8253);
nand U10886 (N_10886,N_9259,N_9441);
nor U10887 (N_10887,N_9432,N_9448);
and U10888 (N_10888,N_9562,N_9313);
xnor U10889 (N_10889,N_8647,N_8635);
and U10890 (N_10890,N_9249,N_8630);
nor U10891 (N_10891,N_9154,N_9442);
and U10892 (N_10892,N_8035,N_9710);
or U10893 (N_10893,N_9893,N_8182);
and U10894 (N_10894,N_8207,N_9025);
xor U10895 (N_10895,N_9963,N_9786);
and U10896 (N_10896,N_9709,N_8026);
and U10897 (N_10897,N_9923,N_9022);
or U10898 (N_10898,N_9542,N_9591);
and U10899 (N_10899,N_8519,N_9850);
xor U10900 (N_10900,N_8119,N_8914);
or U10901 (N_10901,N_8601,N_8727);
nor U10902 (N_10902,N_8676,N_9858);
or U10903 (N_10903,N_8564,N_9488);
xor U10904 (N_10904,N_9012,N_8975);
nor U10905 (N_10905,N_8821,N_8436);
nor U10906 (N_10906,N_8972,N_8621);
xor U10907 (N_10907,N_8999,N_9113);
nor U10908 (N_10908,N_9979,N_9728);
nor U10909 (N_10909,N_8579,N_8267);
and U10910 (N_10910,N_8527,N_8079);
and U10911 (N_10911,N_9325,N_9372);
nand U10912 (N_10912,N_9750,N_8220);
or U10913 (N_10913,N_9701,N_9749);
nand U10914 (N_10914,N_9324,N_8380);
and U10915 (N_10915,N_9139,N_8512);
or U10916 (N_10916,N_9718,N_8060);
or U10917 (N_10917,N_8115,N_8281);
or U10918 (N_10918,N_9972,N_9468);
nor U10919 (N_10919,N_8231,N_8484);
and U10920 (N_10920,N_8185,N_8487);
xor U10921 (N_10921,N_8606,N_8120);
and U10922 (N_10922,N_8401,N_8850);
nor U10923 (N_10923,N_8970,N_9049);
xor U10924 (N_10924,N_8408,N_8313);
and U10925 (N_10925,N_8521,N_8050);
xor U10926 (N_10926,N_8059,N_8112);
and U10927 (N_10927,N_8191,N_9342);
or U10928 (N_10928,N_8653,N_9608);
and U10929 (N_10929,N_8383,N_9349);
xnor U10930 (N_10930,N_8271,N_9913);
nand U10931 (N_10931,N_9258,N_9115);
or U10932 (N_10932,N_9374,N_9799);
and U10933 (N_10933,N_8058,N_8532);
nor U10934 (N_10934,N_8007,N_8346);
or U10935 (N_10935,N_9943,N_8844);
nand U10936 (N_10936,N_9859,N_9020);
and U10937 (N_10937,N_9036,N_9360);
and U10938 (N_10938,N_8186,N_8425);
nand U10939 (N_10939,N_9760,N_8003);
or U10940 (N_10940,N_9838,N_9413);
xnor U10941 (N_10941,N_9101,N_9447);
xor U10942 (N_10942,N_9567,N_8162);
or U10943 (N_10943,N_9685,N_8139);
or U10944 (N_10944,N_9493,N_8199);
xor U10945 (N_10945,N_9323,N_8860);
nand U10946 (N_10946,N_9177,N_8994);
or U10947 (N_10947,N_9174,N_8417);
or U10948 (N_10948,N_8330,N_8282);
nand U10949 (N_10949,N_8739,N_9574);
nand U10950 (N_10950,N_8755,N_9450);
and U10951 (N_10951,N_8654,N_9203);
or U10952 (N_10952,N_8851,N_9301);
or U10953 (N_10953,N_8284,N_8945);
or U10954 (N_10954,N_8811,N_8230);
nor U10955 (N_10955,N_8395,N_8367);
xnor U10956 (N_10956,N_8176,N_9104);
and U10957 (N_10957,N_8027,N_8094);
nor U10958 (N_10958,N_8381,N_9975);
nand U10959 (N_10959,N_9630,N_9814);
and U10960 (N_10960,N_8457,N_9065);
nor U10961 (N_10961,N_8136,N_8826);
nor U10962 (N_10962,N_9048,N_8541);
xnor U10963 (N_10963,N_8224,N_8867);
xnor U10964 (N_10964,N_9094,N_9998);
xnor U10965 (N_10965,N_9241,N_8166);
nand U10966 (N_10966,N_9167,N_8984);
or U10967 (N_10967,N_8066,N_9926);
nor U10968 (N_10968,N_8917,N_9182);
nor U10969 (N_10969,N_8679,N_9178);
nor U10970 (N_10970,N_8774,N_8719);
and U10971 (N_10971,N_9491,N_8834);
and U10972 (N_10972,N_9431,N_8158);
nand U10973 (N_10973,N_8907,N_8258);
xor U10974 (N_10974,N_9303,N_9627);
xnor U10975 (N_10975,N_8849,N_9062);
nand U10976 (N_10976,N_9097,N_9239);
xor U10977 (N_10977,N_9156,N_8132);
or U10978 (N_10978,N_8551,N_9595);
and U10979 (N_10979,N_8075,N_9936);
nand U10980 (N_10980,N_9568,N_9014);
nand U10981 (N_10981,N_8133,N_8048);
nor U10982 (N_10982,N_9306,N_9903);
nor U10983 (N_10983,N_8567,N_9093);
and U10984 (N_10984,N_9472,N_9887);
xnor U10985 (N_10985,N_9398,N_8010);
nor U10986 (N_10986,N_9109,N_8863);
xnor U10987 (N_10987,N_9734,N_8894);
nor U10988 (N_10988,N_9765,N_8490);
nor U10989 (N_10989,N_9559,N_9958);
xor U10990 (N_10990,N_8697,N_9163);
or U10991 (N_10991,N_8549,N_9485);
nor U10992 (N_10992,N_8489,N_8969);
nor U10993 (N_10993,N_9543,N_8483);
nor U10994 (N_10994,N_9544,N_9004);
xor U10995 (N_10995,N_8895,N_9888);
xor U10996 (N_10996,N_8032,N_9767);
or U10997 (N_10997,N_8669,N_8594);
nand U10998 (N_10998,N_9762,N_8502);
and U10999 (N_10999,N_8992,N_9534);
nand U11000 (N_11000,N_8822,N_8347);
nand U11001 (N_11001,N_9483,N_8256);
xor U11002 (N_11002,N_9343,N_8903);
nand U11003 (N_11003,N_9519,N_8071);
and U11004 (N_11004,N_9530,N_9192);
and U11005 (N_11005,N_9359,N_9028);
nor U11006 (N_11006,N_9721,N_8343);
nor U11007 (N_11007,N_9901,N_9211);
nand U11008 (N_11008,N_9700,N_9831);
nor U11009 (N_11009,N_8583,N_8834);
nor U11010 (N_11010,N_9071,N_8302);
nand U11011 (N_11011,N_8370,N_8144);
nand U11012 (N_11012,N_8158,N_8101);
xnor U11013 (N_11013,N_8879,N_9506);
xor U11014 (N_11014,N_9399,N_9710);
xor U11015 (N_11015,N_9504,N_9034);
nor U11016 (N_11016,N_8952,N_9633);
nand U11017 (N_11017,N_8580,N_9791);
or U11018 (N_11018,N_9303,N_8289);
or U11019 (N_11019,N_9707,N_8023);
and U11020 (N_11020,N_9500,N_9290);
xor U11021 (N_11021,N_9008,N_8406);
nand U11022 (N_11022,N_9210,N_9397);
and U11023 (N_11023,N_9386,N_8808);
nor U11024 (N_11024,N_9562,N_9118);
xnor U11025 (N_11025,N_9237,N_8481);
and U11026 (N_11026,N_9966,N_9990);
xor U11027 (N_11027,N_9323,N_9144);
or U11028 (N_11028,N_8189,N_9082);
nand U11029 (N_11029,N_8741,N_8152);
nor U11030 (N_11030,N_8511,N_8864);
nand U11031 (N_11031,N_9080,N_9289);
and U11032 (N_11032,N_9634,N_8986);
xnor U11033 (N_11033,N_9730,N_8574);
nor U11034 (N_11034,N_9889,N_8412);
nor U11035 (N_11035,N_9472,N_9309);
or U11036 (N_11036,N_8257,N_9620);
and U11037 (N_11037,N_9035,N_8139);
and U11038 (N_11038,N_8694,N_9120);
nand U11039 (N_11039,N_8398,N_8528);
xor U11040 (N_11040,N_9166,N_9757);
nor U11041 (N_11041,N_9595,N_8191);
nor U11042 (N_11042,N_8333,N_9081);
nor U11043 (N_11043,N_8803,N_8505);
xnor U11044 (N_11044,N_8720,N_8734);
xnor U11045 (N_11045,N_8752,N_8842);
nand U11046 (N_11046,N_8495,N_9845);
xnor U11047 (N_11047,N_9859,N_9634);
nand U11048 (N_11048,N_9714,N_9189);
or U11049 (N_11049,N_9491,N_9675);
or U11050 (N_11050,N_8122,N_9817);
and U11051 (N_11051,N_9159,N_8442);
or U11052 (N_11052,N_8448,N_8615);
xor U11053 (N_11053,N_9891,N_9947);
or U11054 (N_11054,N_9098,N_9255);
and U11055 (N_11055,N_9370,N_8875);
or U11056 (N_11056,N_8484,N_8110);
nor U11057 (N_11057,N_8859,N_8916);
or U11058 (N_11058,N_8812,N_9180);
xnor U11059 (N_11059,N_8219,N_8205);
nand U11060 (N_11060,N_9337,N_9853);
nand U11061 (N_11061,N_8695,N_9448);
and U11062 (N_11062,N_9867,N_9841);
or U11063 (N_11063,N_8408,N_9237);
xnor U11064 (N_11064,N_9531,N_9997);
and U11065 (N_11065,N_8871,N_9669);
nand U11066 (N_11066,N_9427,N_9061);
or U11067 (N_11067,N_9232,N_9412);
or U11068 (N_11068,N_9112,N_8031);
nand U11069 (N_11069,N_8431,N_8826);
or U11070 (N_11070,N_9001,N_8290);
and U11071 (N_11071,N_9927,N_9509);
and U11072 (N_11072,N_9617,N_9594);
xnor U11073 (N_11073,N_9185,N_8333);
nor U11074 (N_11074,N_8643,N_9689);
and U11075 (N_11075,N_8048,N_9441);
nand U11076 (N_11076,N_8344,N_8405);
xor U11077 (N_11077,N_9200,N_8985);
nand U11078 (N_11078,N_8436,N_9111);
and U11079 (N_11079,N_9122,N_9572);
nand U11080 (N_11080,N_9434,N_8415);
or U11081 (N_11081,N_8923,N_9714);
nor U11082 (N_11082,N_8116,N_9648);
nand U11083 (N_11083,N_9375,N_9129);
xor U11084 (N_11084,N_8332,N_8929);
nor U11085 (N_11085,N_9174,N_9566);
xor U11086 (N_11086,N_8772,N_9570);
nor U11087 (N_11087,N_9928,N_9416);
or U11088 (N_11088,N_9954,N_8936);
or U11089 (N_11089,N_9740,N_9711);
and U11090 (N_11090,N_9702,N_9822);
nor U11091 (N_11091,N_9722,N_9185);
nand U11092 (N_11092,N_8332,N_9056);
xor U11093 (N_11093,N_9635,N_9600);
and U11094 (N_11094,N_9395,N_9604);
xnor U11095 (N_11095,N_8752,N_9211);
nor U11096 (N_11096,N_8806,N_8596);
xnor U11097 (N_11097,N_8170,N_8532);
xor U11098 (N_11098,N_9439,N_8533);
nor U11099 (N_11099,N_9414,N_8884);
nor U11100 (N_11100,N_8831,N_8551);
nand U11101 (N_11101,N_9143,N_9762);
nor U11102 (N_11102,N_8934,N_9062);
xor U11103 (N_11103,N_9599,N_9846);
nor U11104 (N_11104,N_9167,N_9950);
and U11105 (N_11105,N_8282,N_9084);
and U11106 (N_11106,N_8153,N_9887);
or U11107 (N_11107,N_9181,N_9679);
and U11108 (N_11108,N_8371,N_9936);
xnor U11109 (N_11109,N_8260,N_9079);
or U11110 (N_11110,N_8085,N_9346);
nand U11111 (N_11111,N_9527,N_8257);
nor U11112 (N_11112,N_8181,N_8585);
or U11113 (N_11113,N_8918,N_8270);
nor U11114 (N_11114,N_9405,N_9718);
xor U11115 (N_11115,N_9708,N_8080);
and U11116 (N_11116,N_8323,N_8828);
or U11117 (N_11117,N_9034,N_9653);
nor U11118 (N_11118,N_8375,N_9143);
or U11119 (N_11119,N_8405,N_9781);
nand U11120 (N_11120,N_8253,N_9275);
nor U11121 (N_11121,N_8668,N_8187);
or U11122 (N_11122,N_9390,N_9208);
xnor U11123 (N_11123,N_8686,N_9500);
or U11124 (N_11124,N_8096,N_8035);
nor U11125 (N_11125,N_9272,N_9173);
nor U11126 (N_11126,N_9883,N_8442);
nand U11127 (N_11127,N_8242,N_9402);
and U11128 (N_11128,N_9378,N_8328);
nor U11129 (N_11129,N_8548,N_9514);
nor U11130 (N_11130,N_9809,N_8387);
nor U11131 (N_11131,N_9253,N_9497);
nand U11132 (N_11132,N_9338,N_8529);
or U11133 (N_11133,N_9283,N_9865);
xor U11134 (N_11134,N_8213,N_9311);
or U11135 (N_11135,N_8633,N_9814);
or U11136 (N_11136,N_9278,N_9350);
and U11137 (N_11137,N_9822,N_9470);
or U11138 (N_11138,N_8267,N_9009);
and U11139 (N_11139,N_9560,N_8301);
nor U11140 (N_11140,N_8611,N_8143);
nor U11141 (N_11141,N_8682,N_9660);
xor U11142 (N_11142,N_9411,N_8342);
nor U11143 (N_11143,N_8474,N_9886);
nand U11144 (N_11144,N_8106,N_9010);
and U11145 (N_11145,N_8816,N_9036);
and U11146 (N_11146,N_8802,N_8769);
and U11147 (N_11147,N_8201,N_9138);
and U11148 (N_11148,N_9010,N_9349);
or U11149 (N_11149,N_8243,N_8887);
or U11150 (N_11150,N_9043,N_8799);
nand U11151 (N_11151,N_8665,N_9669);
nor U11152 (N_11152,N_8705,N_8569);
or U11153 (N_11153,N_8408,N_9803);
xnor U11154 (N_11154,N_9479,N_8360);
and U11155 (N_11155,N_8568,N_9299);
or U11156 (N_11156,N_9795,N_9090);
nand U11157 (N_11157,N_8360,N_8203);
or U11158 (N_11158,N_8021,N_9726);
or U11159 (N_11159,N_8687,N_8472);
or U11160 (N_11160,N_8127,N_8024);
nor U11161 (N_11161,N_8430,N_9789);
xor U11162 (N_11162,N_9141,N_8383);
and U11163 (N_11163,N_8663,N_9281);
or U11164 (N_11164,N_9831,N_8910);
and U11165 (N_11165,N_9972,N_8335);
nand U11166 (N_11166,N_8605,N_9456);
and U11167 (N_11167,N_8953,N_8199);
or U11168 (N_11168,N_8451,N_9261);
and U11169 (N_11169,N_9695,N_8116);
or U11170 (N_11170,N_8695,N_9749);
or U11171 (N_11171,N_8803,N_8535);
nor U11172 (N_11172,N_9493,N_9663);
xnor U11173 (N_11173,N_9542,N_8361);
nor U11174 (N_11174,N_9384,N_9956);
nor U11175 (N_11175,N_8367,N_9464);
xnor U11176 (N_11176,N_9595,N_8549);
or U11177 (N_11177,N_9629,N_8239);
or U11178 (N_11178,N_9152,N_9102);
nor U11179 (N_11179,N_9222,N_8054);
nor U11180 (N_11180,N_9892,N_9642);
nand U11181 (N_11181,N_8309,N_9169);
or U11182 (N_11182,N_9057,N_9788);
nand U11183 (N_11183,N_9405,N_9276);
nand U11184 (N_11184,N_8776,N_8698);
nor U11185 (N_11185,N_9520,N_8265);
xor U11186 (N_11186,N_9921,N_9574);
and U11187 (N_11187,N_9759,N_9150);
nor U11188 (N_11188,N_8336,N_8544);
or U11189 (N_11189,N_9700,N_8391);
nand U11190 (N_11190,N_8912,N_9942);
nand U11191 (N_11191,N_9302,N_8252);
or U11192 (N_11192,N_8806,N_9165);
or U11193 (N_11193,N_9821,N_9485);
xnor U11194 (N_11194,N_8956,N_8461);
or U11195 (N_11195,N_9661,N_9483);
nor U11196 (N_11196,N_8448,N_8469);
nor U11197 (N_11197,N_9102,N_9343);
nand U11198 (N_11198,N_8689,N_8900);
or U11199 (N_11199,N_9793,N_8156);
or U11200 (N_11200,N_8654,N_8703);
nor U11201 (N_11201,N_8662,N_9172);
or U11202 (N_11202,N_9772,N_8053);
or U11203 (N_11203,N_9823,N_8729);
xnor U11204 (N_11204,N_9751,N_9511);
and U11205 (N_11205,N_8978,N_9017);
nor U11206 (N_11206,N_9807,N_8418);
and U11207 (N_11207,N_8116,N_9366);
nand U11208 (N_11208,N_8102,N_8190);
nand U11209 (N_11209,N_9108,N_8452);
xor U11210 (N_11210,N_8064,N_9161);
nor U11211 (N_11211,N_9212,N_9977);
nand U11212 (N_11212,N_9949,N_8292);
or U11213 (N_11213,N_8058,N_8959);
xor U11214 (N_11214,N_9991,N_9512);
and U11215 (N_11215,N_8839,N_8994);
nand U11216 (N_11216,N_9900,N_8055);
or U11217 (N_11217,N_9811,N_8253);
xnor U11218 (N_11218,N_9624,N_8672);
xor U11219 (N_11219,N_8820,N_9740);
xor U11220 (N_11220,N_9142,N_9529);
nor U11221 (N_11221,N_8462,N_8778);
nand U11222 (N_11222,N_9571,N_9189);
nor U11223 (N_11223,N_9452,N_9819);
or U11224 (N_11224,N_8701,N_9719);
and U11225 (N_11225,N_9020,N_8156);
nand U11226 (N_11226,N_8075,N_9262);
nor U11227 (N_11227,N_9938,N_8276);
and U11228 (N_11228,N_9732,N_9006);
nand U11229 (N_11229,N_9543,N_9638);
and U11230 (N_11230,N_9794,N_8442);
nor U11231 (N_11231,N_9554,N_8707);
or U11232 (N_11232,N_9682,N_8141);
and U11233 (N_11233,N_9733,N_9845);
and U11234 (N_11234,N_8514,N_8900);
xor U11235 (N_11235,N_9433,N_9667);
xnor U11236 (N_11236,N_8911,N_8164);
xor U11237 (N_11237,N_8703,N_8145);
or U11238 (N_11238,N_9310,N_8795);
or U11239 (N_11239,N_9807,N_9976);
or U11240 (N_11240,N_8565,N_9243);
nor U11241 (N_11241,N_8905,N_9404);
nor U11242 (N_11242,N_9978,N_9201);
and U11243 (N_11243,N_8523,N_8976);
nor U11244 (N_11244,N_8863,N_8612);
nand U11245 (N_11245,N_8915,N_8938);
or U11246 (N_11246,N_8845,N_8536);
xor U11247 (N_11247,N_8767,N_8923);
xor U11248 (N_11248,N_8588,N_9808);
or U11249 (N_11249,N_9515,N_9090);
and U11250 (N_11250,N_9057,N_8066);
xnor U11251 (N_11251,N_8712,N_9124);
xnor U11252 (N_11252,N_9885,N_8939);
nand U11253 (N_11253,N_8405,N_9525);
and U11254 (N_11254,N_8389,N_8243);
and U11255 (N_11255,N_9427,N_8561);
nor U11256 (N_11256,N_9931,N_8686);
nor U11257 (N_11257,N_9322,N_9382);
and U11258 (N_11258,N_8109,N_8945);
xor U11259 (N_11259,N_9167,N_8341);
xnor U11260 (N_11260,N_8003,N_9726);
nor U11261 (N_11261,N_9129,N_9502);
and U11262 (N_11262,N_8986,N_9722);
nand U11263 (N_11263,N_9205,N_8626);
or U11264 (N_11264,N_9281,N_8994);
nor U11265 (N_11265,N_9883,N_8017);
nor U11266 (N_11266,N_8093,N_8645);
xnor U11267 (N_11267,N_8756,N_8574);
nand U11268 (N_11268,N_9139,N_8177);
and U11269 (N_11269,N_8023,N_8129);
and U11270 (N_11270,N_8768,N_8823);
nand U11271 (N_11271,N_9949,N_8333);
or U11272 (N_11272,N_8598,N_9240);
nand U11273 (N_11273,N_8906,N_9211);
nand U11274 (N_11274,N_8976,N_8096);
or U11275 (N_11275,N_8503,N_9999);
and U11276 (N_11276,N_8908,N_8395);
nor U11277 (N_11277,N_8505,N_9666);
nand U11278 (N_11278,N_8457,N_9020);
and U11279 (N_11279,N_9022,N_8212);
nand U11280 (N_11280,N_8101,N_9114);
or U11281 (N_11281,N_9763,N_9892);
and U11282 (N_11282,N_9870,N_8257);
nand U11283 (N_11283,N_8490,N_9167);
and U11284 (N_11284,N_9500,N_8460);
nand U11285 (N_11285,N_9704,N_9597);
and U11286 (N_11286,N_9246,N_8520);
and U11287 (N_11287,N_9724,N_9619);
nor U11288 (N_11288,N_8394,N_8370);
or U11289 (N_11289,N_8029,N_9895);
and U11290 (N_11290,N_9199,N_8050);
nor U11291 (N_11291,N_8746,N_8162);
and U11292 (N_11292,N_8771,N_8466);
nor U11293 (N_11293,N_8501,N_9515);
nand U11294 (N_11294,N_8958,N_9178);
or U11295 (N_11295,N_8334,N_8920);
nor U11296 (N_11296,N_9559,N_8530);
xnor U11297 (N_11297,N_8249,N_8924);
and U11298 (N_11298,N_9336,N_9910);
xnor U11299 (N_11299,N_8368,N_9972);
and U11300 (N_11300,N_8443,N_9981);
nor U11301 (N_11301,N_8044,N_8622);
nor U11302 (N_11302,N_8021,N_8370);
xor U11303 (N_11303,N_9308,N_9699);
or U11304 (N_11304,N_9926,N_9785);
and U11305 (N_11305,N_8118,N_8449);
nor U11306 (N_11306,N_8925,N_9703);
or U11307 (N_11307,N_9362,N_8186);
nor U11308 (N_11308,N_9140,N_9595);
xor U11309 (N_11309,N_8691,N_8195);
and U11310 (N_11310,N_8836,N_9818);
nor U11311 (N_11311,N_9069,N_8327);
nor U11312 (N_11312,N_8878,N_8971);
nor U11313 (N_11313,N_9361,N_8248);
or U11314 (N_11314,N_9853,N_9334);
and U11315 (N_11315,N_8082,N_9865);
nand U11316 (N_11316,N_9173,N_9235);
nor U11317 (N_11317,N_8719,N_9952);
nor U11318 (N_11318,N_8114,N_9349);
or U11319 (N_11319,N_9681,N_9853);
and U11320 (N_11320,N_8681,N_9973);
and U11321 (N_11321,N_9188,N_9280);
nand U11322 (N_11322,N_9916,N_9855);
nor U11323 (N_11323,N_8412,N_9569);
nor U11324 (N_11324,N_8547,N_8706);
nor U11325 (N_11325,N_9515,N_9958);
and U11326 (N_11326,N_8599,N_9262);
and U11327 (N_11327,N_9145,N_8882);
xnor U11328 (N_11328,N_9977,N_9996);
nand U11329 (N_11329,N_8021,N_9399);
xnor U11330 (N_11330,N_9741,N_8342);
xnor U11331 (N_11331,N_8032,N_8192);
nand U11332 (N_11332,N_8899,N_9461);
xor U11333 (N_11333,N_8275,N_9817);
and U11334 (N_11334,N_8560,N_8612);
and U11335 (N_11335,N_8410,N_9095);
or U11336 (N_11336,N_9044,N_9472);
or U11337 (N_11337,N_8705,N_9874);
nand U11338 (N_11338,N_8959,N_8531);
xor U11339 (N_11339,N_9446,N_9783);
or U11340 (N_11340,N_9765,N_9114);
nor U11341 (N_11341,N_8878,N_8588);
or U11342 (N_11342,N_8589,N_9098);
and U11343 (N_11343,N_9992,N_9379);
xnor U11344 (N_11344,N_9247,N_8049);
nand U11345 (N_11345,N_9728,N_9601);
xnor U11346 (N_11346,N_9702,N_9755);
or U11347 (N_11347,N_8664,N_9735);
nor U11348 (N_11348,N_8479,N_8517);
nand U11349 (N_11349,N_9301,N_9160);
xor U11350 (N_11350,N_9516,N_8043);
nor U11351 (N_11351,N_8302,N_8063);
nand U11352 (N_11352,N_9537,N_8107);
or U11353 (N_11353,N_9111,N_8506);
or U11354 (N_11354,N_8644,N_8574);
xor U11355 (N_11355,N_9549,N_9354);
xor U11356 (N_11356,N_9538,N_8744);
and U11357 (N_11357,N_8338,N_9920);
and U11358 (N_11358,N_9787,N_9478);
and U11359 (N_11359,N_8334,N_9421);
or U11360 (N_11360,N_8356,N_9351);
or U11361 (N_11361,N_9712,N_8712);
nor U11362 (N_11362,N_9728,N_9627);
and U11363 (N_11363,N_9033,N_8823);
or U11364 (N_11364,N_8260,N_9198);
or U11365 (N_11365,N_8080,N_8950);
nor U11366 (N_11366,N_8845,N_9763);
and U11367 (N_11367,N_8720,N_9711);
xor U11368 (N_11368,N_9382,N_8363);
xor U11369 (N_11369,N_8710,N_9909);
nor U11370 (N_11370,N_9061,N_9109);
xor U11371 (N_11371,N_8814,N_8464);
xnor U11372 (N_11372,N_9491,N_9329);
xor U11373 (N_11373,N_9602,N_9024);
xor U11374 (N_11374,N_9447,N_9288);
or U11375 (N_11375,N_9170,N_8251);
xnor U11376 (N_11376,N_9528,N_8380);
nor U11377 (N_11377,N_8336,N_8364);
xnor U11378 (N_11378,N_8091,N_9201);
nand U11379 (N_11379,N_9268,N_8880);
xnor U11380 (N_11380,N_9024,N_9560);
nand U11381 (N_11381,N_8208,N_8041);
xnor U11382 (N_11382,N_8197,N_9242);
nor U11383 (N_11383,N_9634,N_8276);
and U11384 (N_11384,N_9578,N_9226);
and U11385 (N_11385,N_8304,N_9860);
nand U11386 (N_11386,N_9673,N_9163);
nand U11387 (N_11387,N_8622,N_8230);
and U11388 (N_11388,N_8270,N_9641);
nand U11389 (N_11389,N_9121,N_8077);
xnor U11390 (N_11390,N_8255,N_8504);
nor U11391 (N_11391,N_9099,N_9991);
nand U11392 (N_11392,N_9656,N_9788);
and U11393 (N_11393,N_8817,N_9820);
nand U11394 (N_11394,N_9515,N_9204);
and U11395 (N_11395,N_9435,N_8467);
nor U11396 (N_11396,N_8417,N_9416);
xnor U11397 (N_11397,N_8210,N_8686);
xnor U11398 (N_11398,N_8691,N_8187);
nand U11399 (N_11399,N_8551,N_9554);
nand U11400 (N_11400,N_8807,N_8470);
or U11401 (N_11401,N_9871,N_8112);
or U11402 (N_11402,N_8427,N_9845);
or U11403 (N_11403,N_9583,N_8983);
nand U11404 (N_11404,N_9716,N_8308);
nor U11405 (N_11405,N_9273,N_9330);
or U11406 (N_11406,N_9891,N_8694);
xnor U11407 (N_11407,N_8148,N_9806);
xnor U11408 (N_11408,N_8216,N_8235);
or U11409 (N_11409,N_8479,N_9418);
and U11410 (N_11410,N_8853,N_8608);
and U11411 (N_11411,N_9295,N_8845);
or U11412 (N_11412,N_9997,N_8566);
nor U11413 (N_11413,N_8641,N_9950);
or U11414 (N_11414,N_8534,N_8167);
xnor U11415 (N_11415,N_9946,N_8224);
nor U11416 (N_11416,N_8255,N_9556);
nor U11417 (N_11417,N_8184,N_9947);
nand U11418 (N_11418,N_8698,N_9243);
xnor U11419 (N_11419,N_9610,N_8350);
nor U11420 (N_11420,N_9247,N_8504);
or U11421 (N_11421,N_9967,N_9719);
and U11422 (N_11422,N_9471,N_9534);
nand U11423 (N_11423,N_9922,N_8998);
or U11424 (N_11424,N_8373,N_8816);
xnor U11425 (N_11425,N_8071,N_8640);
nand U11426 (N_11426,N_9280,N_8676);
or U11427 (N_11427,N_9229,N_9859);
and U11428 (N_11428,N_8839,N_8908);
and U11429 (N_11429,N_8421,N_9524);
xor U11430 (N_11430,N_9691,N_9520);
nand U11431 (N_11431,N_8716,N_9428);
nand U11432 (N_11432,N_8971,N_9809);
or U11433 (N_11433,N_9507,N_9296);
nor U11434 (N_11434,N_9311,N_9202);
nand U11435 (N_11435,N_9565,N_8960);
nor U11436 (N_11436,N_8746,N_9077);
xor U11437 (N_11437,N_8890,N_9628);
xnor U11438 (N_11438,N_8570,N_9547);
and U11439 (N_11439,N_9605,N_9593);
and U11440 (N_11440,N_9824,N_8105);
nor U11441 (N_11441,N_9171,N_8301);
and U11442 (N_11442,N_9370,N_9986);
and U11443 (N_11443,N_8226,N_8962);
and U11444 (N_11444,N_9403,N_9831);
or U11445 (N_11445,N_9113,N_9943);
or U11446 (N_11446,N_8755,N_9287);
nor U11447 (N_11447,N_9217,N_8954);
and U11448 (N_11448,N_8184,N_9596);
or U11449 (N_11449,N_9694,N_9589);
and U11450 (N_11450,N_8311,N_9769);
or U11451 (N_11451,N_9314,N_8323);
nor U11452 (N_11452,N_9778,N_8437);
nand U11453 (N_11453,N_9674,N_9021);
xnor U11454 (N_11454,N_8866,N_9139);
nor U11455 (N_11455,N_9567,N_9666);
nor U11456 (N_11456,N_8958,N_8587);
nor U11457 (N_11457,N_8816,N_8471);
xnor U11458 (N_11458,N_9948,N_8886);
xnor U11459 (N_11459,N_9316,N_9665);
or U11460 (N_11460,N_9522,N_8740);
xor U11461 (N_11461,N_9411,N_9700);
nor U11462 (N_11462,N_9234,N_9454);
and U11463 (N_11463,N_8966,N_8719);
nand U11464 (N_11464,N_9416,N_8389);
nor U11465 (N_11465,N_8701,N_9231);
and U11466 (N_11466,N_9745,N_8552);
xnor U11467 (N_11467,N_8612,N_9056);
xnor U11468 (N_11468,N_9200,N_9126);
nor U11469 (N_11469,N_8773,N_9879);
and U11470 (N_11470,N_9115,N_8317);
nor U11471 (N_11471,N_8150,N_8858);
xor U11472 (N_11472,N_8187,N_9773);
nand U11473 (N_11473,N_9585,N_8736);
nand U11474 (N_11474,N_8644,N_9331);
and U11475 (N_11475,N_8912,N_9956);
or U11476 (N_11476,N_8887,N_8060);
nor U11477 (N_11477,N_8169,N_9205);
nand U11478 (N_11478,N_9420,N_8182);
and U11479 (N_11479,N_8035,N_9459);
or U11480 (N_11480,N_9261,N_8276);
and U11481 (N_11481,N_8993,N_8446);
or U11482 (N_11482,N_8460,N_8329);
nor U11483 (N_11483,N_8359,N_9988);
nand U11484 (N_11484,N_9939,N_8782);
nand U11485 (N_11485,N_9404,N_8329);
or U11486 (N_11486,N_8539,N_9378);
nand U11487 (N_11487,N_8411,N_9255);
nand U11488 (N_11488,N_9323,N_8341);
or U11489 (N_11489,N_8906,N_9044);
nor U11490 (N_11490,N_8886,N_9116);
nand U11491 (N_11491,N_9155,N_9315);
or U11492 (N_11492,N_8615,N_9400);
and U11493 (N_11493,N_9848,N_9251);
xor U11494 (N_11494,N_8818,N_8990);
nand U11495 (N_11495,N_9562,N_9997);
xnor U11496 (N_11496,N_8708,N_8017);
or U11497 (N_11497,N_9693,N_8449);
and U11498 (N_11498,N_9437,N_9608);
nor U11499 (N_11499,N_9173,N_8743);
xnor U11500 (N_11500,N_8893,N_9544);
nor U11501 (N_11501,N_8124,N_8216);
nand U11502 (N_11502,N_8079,N_8460);
or U11503 (N_11503,N_9633,N_9856);
nand U11504 (N_11504,N_8040,N_8051);
xnor U11505 (N_11505,N_9452,N_8565);
nor U11506 (N_11506,N_8402,N_9395);
or U11507 (N_11507,N_9287,N_8629);
nor U11508 (N_11508,N_9077,N_9312);
nand U11509 (N_11509,N_9107,N_8837);
and U11510 (N_11510,N_8435,N_8515);
nor U11511 (N_11511,N_8582,N_9258);
or U11512 (N_11512,N_9702,N_9423);
nor U11513 (N_11513,N_8179,N_9421);
and U11514 (N_11514,N_9579,N_9491);
or U11515 (N_11515,N_9452,N_8139);
xor U11516 (N_11516,N_9146,N_8384);
xor U11517 (N_11517,N_8830,N_8008);
nor U11518 (N_11518,N_9820,N_9533);
nand U11519 (N_11519,N_9942,N_8083);
nand U11520 (N_11520,N_8741,N_9368);
or U11521 (N_11521,N_9711,N_8680);
xor U11522 (N_11522,N_8988,N_8701);
nand U11523 (N_11523,N_8375,N_8283);
nor U11524 (N_11524,N_9727,N_8024);
xor U11525 (N_11525,N_9421,N_8728);
and U11526 (N_11526,N_9542,N_9097);
or U11527 (N_11527,N_8660,N_9864);
nand U11528 (N_11528,N_9996,N_8013);
xor U11529 (N_11529,N_9418,N_8444);
xor U11530 (N_11530,N_9290,N_9066);
or U11531 (N_11531,N_9533,N_9398);
nor U11532 (N_11532,N_9414,N_9848);
xnor U11533 (N_11533,N_8620,N_9319);
or U11534 (N_11534,N_9780,N_8512);
xnor U11535 (N_11535,N_8737,N_8018);
xnor U11536 (N_11536,N_9783,N_8605);
or U11537 (N_11537,N_8155,N_9047);
xnor U11538 (N_11538,N_9093,N_9403);
or U11539 (N_11539,N_8543,N_9461);
nor U11540 (N_11540,N_9540,N_9794);
xor U11541 (N_11541,N_9009,N_8095);
or U11542 (N_11542,N_8063,N_9951);
and U11543 (N_11543,N_9306,N_9305);
and U11544 (N_11544,N_9885,N_9933);
and U11545 (N_11545,N_9320,N_9722);
nand U11546 (N_11546,N_9845,N_8902);
and U11547 (N_11547,N_9266,N_8327);
xnor U11548 (N_11548,N_9610,N_8413);
and U11549 (N_11549,N_8746,N_8803);
or U11550 (N_11550,N_8652,N_8775);
nand U11551 (N_11551,N_8508,N_9072);
nand U11552 (N_11552,N_8017,N_8619);
and U11553 (N_11553,N_8966,N_9104);
or U11554 (N_11554,N_8653,N_9711);
nand U11555 (N_11555,N_8045,N_8519);
nand U11556 (N_11556,N_9871,N_8435);
nand U11557 (N_11557,N_9314,N_8168);
and U11558 (N_11558,N_8245,N_8276);
nand U11559 (N_11559,N_8419,N_9201);
xnor U11560 (N_11560,N_8916,N_9270);
and U11561 (N_11561,N_8301,N_8466);
xnor U11562 (N_11562,N_9002,N_9335);
xor U11563 (N_11563,N_8054,N_9294);
nand U11564 (N_11564,N_9451,N_8583);
and U11565 (N_11565,N_9178,N_8699);
xnor U11566 (N_11566,N_9687,N_8357);
nand U11567 (N_11567,N_9224,N_8585);
xnor U11568 (N_11568,N_8947,N_8526);
nand U11569 (N_11569,N_8646,N_8421);
nand U11570 (N_11570,N_9283,N_9026);
xor U11571 (N_11571,N_9151,N_8952);
nor U11572 (N_11572,N_8385,N_8331);
or U11573 (N_11573,N_9141,N_8281);
or U11574 (N_11574,N_9343,N_9174);
nand U11575 (N_11575,N_9029,N_8640);
nor U11576 (N_11576,N_9470,N_8723);
and U11577 (N_11577,N_8369,N_9383);
xor U11578 (N_11578,N_9652,N_8347);
nor U11579 (N_11579,N_8637,N_8220);
and U11580 (N_11580,N_9964,N_8616);
nor U11581 (N_11581,N_8082,N_8308);
and U11582 (N_11582,N_8615,N_9958);
xor U11583 (N_11583,N_8182,N_8441);
and U11584 (N_11584,N_8306,N_8808);
nor U11585 (N_11585,N_9134,N_8128);
and U11586 (N_11586,N_9566,N_9437);
nand U11587 (N_11587,N_8013,N_9042);
and U11588 (N_11588,N_9386,N_9823);
or U11589 (N_11589,N_8946,N_9993);
or U11590 (N_11590,N_9268,N_8233);
nor U11591 (N_11591,N_9574,N_9925);
nor U11592 (N_11592,N_8063,N_8182);
xnor U11593 (N_11593,N_9309,N_8009);
xor U11594 (N_11594,N_8293,N_9718);
nor U11595 (N_11595,N_9912,N_9745);
nor U11596 (N_11596,N_9756,N_8878);
xnor U11597 (N_11597,N_9044,N_8948);
xnor U11598 (N_11598,N_8730,N_8316);
xnor U11599 (N_11599,N_8559,N_8008);
or U11600 (N_11600,N_9048,N_8105);
xor U11601 (N_11601,N_9848,N_8405);
and U11602 (N_11602,N_8504,N_9069);
nand U11603 (N_11603,N_8255,N_8938);
nand U11604 (N_11604,N_9191,N_9451);
or U11605 (N_11605,N_8957,N_9111);
or U11606 (N_11606,N_8882,N_9194);
nand U11607 (N_11607,N_9886,N_8458);
and U11608 (N_11608,N_9120,N_8853);
xnor U11609 (N_11609,N_9589,N_8901);
or U11610 (N_11610,N_8991,N_8856);
or U11611 (N_11611,N_9436,N_9172);
xor U11612 (N_11612,N_8949,N_9025);
xnor U11613 (N_11613,N_9600,N_9975);
nor U11614 (N_11614,N_9856,N_9774);
xor U11615 (N_11615,N_8373,N_8913);
or U11616 (N_11616,N_8453,N_9837);
or U11617 (N_11617,N_8019,N_9295);
or U11618 (N_11618,N_9670,N_8413);
and U11619 (N_11619,N_9769,N_8287);
xnor U11620 (N_11620,N_8035,N_9849);
or U11621 (N_11621,N_8623,N_8052);
or U11622 (N_11622,N_8831,N_9087);
and U11623 (N_11623,N_8312,N_9013);
nand U11624 (N_11624,N_8757,N_8556);
and U11625 (N_11625,N_8823,N_8729);
nor U11626 (N_11626,N_9674,N_9275);
or U11627 (N_11627,N_8832,N_9616);
and U11628 (N_11628,N_8191,N_8177);
nor U11629 (N_11629,N_9246,N_9516);
and U11630 (N_11630,N_8700,N_9773);
xor U11631 (N_11631,N_9549,N_9156);
nor U11632 (N_11632,N_8815,N_8607);
or U11633 (N_11633,N_8846,N_8470);
and U11634 (N_11634,N_9491,N_9144);
nand U11635 (N_11635,N_8095,N_8787);
or U11636 (N_11636,N_9161,N_8297);
xor U11637 (N_11637,N_8584,N_8792);
nor U11638 (N_11638,N_9204,N_8355);
and U11639 (N_11639,N_8927,N_9215);
xor U11640 (N_11640,N_8227,N_9551);
nand U11641 (N_11641,N_8596,N_9627);
nand U11642 (N_11642,N_8907,N_8601);
or U11643 (N_11643,N_8949,N_8328);
xnor U11644 (N_11644,N_8359,N_8558);
xnor U11645 (N_11645,N_8590,N_9032);
nor U11646 (N_11646,N_8516,N_9737);
nand U11647 (N_11647,N_9646,N_8183);
nor U11648 (N_11648,N_9468,N_9177);
and U11649 (N_11649,N_8178,N_8643);
and U11650 (N_11650,N_8379,N_8356);
nand U11651 (N_11651,N_9781,N_9480);
and U11652 (N_11652,N_9369,N_8026);
nor U11653 (N_11653,N_8671,N_9196);
xor U11654 (N_11654,N_8657,N_9313);
nor U11655 (N_11655,N_9115,N_9563);
and U11656 (N_11656,N_8322,N_9871);
or U11657 (N_11657,N_9096,N_8377);
nand U11658 (N_11658,N_9192,N_9251);
nor U11659 (N_11659,N_9523,N_8290);
xor U11660 (N_11660,N_9743,N_8101);
or U11661 (N_11661,N_8330,N_9165);
xnor U11662 (N_11662,N_8922,N_8192);
xor U11663 (N_11663,N_8174,N_9899);
or U11664 (N_11664,N_9949,N_8653);
nor U11665 (N_11665,N_8778,N_8144);
xnor U11666 (N_11666,N_9071,N_8735);
and U11667 (N_11667,N_9572,N_9765);
or U11668 (N_11668,N_9635,N_9226);
and U11669 (N_11669,N_9027,N_8613);
and U11670 (N_11670,N_9889,N_8749);
and U11671 (N_11671,N_9219,N_9253);
or U11672 (N_11672,N_9154,N_8984);
nor U11673 (N_11673,N_8642,N_8594);
nand U11674 (N_11674,N_9439,N_8380);
and U11675 (N_11675,N_8138,N_9205);
and U11676 (N_11676,N_8006,N_8970);
xnor U11677 (N_11677,N_9511,N_9131);
nand U11678 (N_11678,N_9803,N_8389);
nand U11679 (N_11679,N_9744,N_9714);
xnor U11680 (N_11680,N_8726,N_8230);
and U11681 (N_11681,N_8864,N_8928);
nand U11682 (N_11682,N_9376,N_8611);
and U11683 (N_11683,N_9432,N_8454);
xor U11684 (N_11684,N_9196,N_9965);
nor U11685 (N_11685,N_9428,N_8143);
nor U11686 (N_11686,N_9267,N_9068);
and U11687 (N_11687,N_9977,N_9475);
nor U11688 (N_11688,N_9374,N_8726);
nor U11689 (N_11689,N_8224,N_8755);
nand U11690 (N_11690,N_8454,N_9004);
xor U11691 (N_11691,N_9270,N_8412);
nand U11692 (N_11692,N_9810,N_8425);
xnor U11693 (N_11693,N_8411,N_8315);
and U11694 (N_11694,N_8041,N_9875);
or U11695 (N_11695,N_9348,N_8085);
and U11696 (N_11696,N_9627,N_8276);
or U11697 (N_11697,N_8271,N_8959);
and U11698 (N_11698,N_9495,N_9406);
nand U11699 (N_11699,N_8193,N_8012);
nor U11700 (N_11700,N_8734,N_9151);
or U11701 (N_11701,N_8377,N_8370);
or U11702 (N_11702,N_9526,N_9070);
and U11703 (N_11703,N_9311,N_8563);
nor U11704 (N_11704,N_9410,N_8774);
nand U11705 (N_11705,N_9255,N_9154);
or U11706 (N_11706,N_9531,N_9836);
and U11707 (N_11707,N_8395,N_8375);
and U11708 (N_11708,N_9696,N_9883);
nor U11709 (N_11709,N_8958,N_9408);
and U11710 (N_11710,N_8937,N_9575);
and U11711 (N_11711,N_9399,N_9158);
nand U11712 (N_11712,N_9522,N_9363);
nand U11713 (N_11713,N_9557,N_8330);
nand U11714 (N_11714,N_8200,N_8616);
nand U11715 (N_11715,N_8577,N_9671);
nor U11716 (N_11716,N_8367,N_9154);
nor U11717 (N_11717,N_8164,N_9109);
nor U11718 (N_11718,N_9071,N_9651);
nor U11719 (N_11719,N_8960,N_8949);
or U11720 (N_11720,N_8923,N_8602);
and U11721 (N_11721,N_9623,N_9842);
and U11722 (N_11722,N_9619,N_8221);
or U11723 (N_11723,N_9924,N_8779);
nor U11724 (N_11724,N_9727,N_8717);
or U11725 (N_11725,N_8812,N_9594);
nor U11726 (N_11726,N_8848,N_8648);
nor U11727 (N_11727,N_9057,N_8289);
nand U11728 (N_11728,N_8168,N_8252);
or U11729 (N_11729,N_9234,N_9840);
nand U11730 (N_11730,N_9402,N_8510);
nand U11731 (N_11731,N_9615,N_8563);
nor U11732 (N_11732,N_9447,N_9738);
or U11733 (N_11733,N_8412,N_9395);
and U11734 (N_11734,N_8551,N_9183);
xnor U11735 (N_11735,N_9130,N_9446);
or U11736 (N_11736,N_8167,N_8164);
or U11737 (N_11737,N_9850,N_9044);
nor U11738 (N_11738,N_9974,N_9633);
nand U11739 (N_11739,N_9038,N_9843);
or U11740 (N_11740,N_8829,N_9649);
and U11741 (N_11741,N_9122,N_8686);
xor U11742 (N_11742,N_9779,N_8333);
nor U11743 (N_11743,N_9546,N_9046);
xor U11744 (N_11744,N_9328,N_8323);
xnor U11745 (N_11745,N_8071,N_8577);
xnor U11746 (N_11746,N_9388,N_9431);
or U11747 (N_11747,N_8043,N_9441);
nor U11748 (N_11748,N_8841,N_8964);
nand U11749 (N_11749,N_8387,N_8882);
nor U11750 (N_11750,N_9496,N_9165);
nand U11751 (N_11751,N_8309,N_8840);
and U11752 (N_11752,N_8581,N_9185);
or U11753 (N_11753,N_8899,N_8231);
xor U11754 (N_11754,N_9178,N_9961);
xor U11755 (N_11755,N_8457,N_8989);
and U11756 (N_11756,N_8064,N_9540);
and U11757 (N_11757,N_9635,N_8732);
and U11758 (N_11758,N_9953,N_9428);
nor U11759 (N_11759,N_8522,N_9105);
and U11760 (N_11760,N_8406,N_9704);
and U11761 (N_11761,N_9831,N_8085);
or U11762 (N_11762,N_8662,N_8303);
nand U11763 (N_11763,N_9410,N_9882);
nor U11764 (N_11764,N_9754,N_9503);
nand U11765 (N_11765,N_8880,N_8459);
or U11766 (N_11766,N_8718,N_8903);
or U11767 (N_11767,N_8772,N_9685);
nor U11768 (N_11768,N_8022,N_9922);
and U11769 (N_11769,N_9583,N_8896);
and U11770 (N_11770,N_9816,N_9872);
and U11771 (N_11771,N_9156,N_9662);
nor U11772 (N_11772,N_9213,N_9276);
nand U11773 (N_11773,N_9698,N_8559);
nor U11774 (N_11774,N_8427,N_8223);
or U11775 (N_11775,N_9719,N_8738);
or U11776 (N_11776,N_8618,N_8504);
xnor U11777 (N_11777,N_9476,N_9268);
nor U11778 (N_11778,N_8191,N_9861);
nand U11779 (N_11779,N_9805,N_9941);
and U11780 (N_11780,N_8834,N_9889);
nand U11781 (N_11781,N_9668,N_9769);
xnor U11782 (N_11782,N_9315,N_8846);
or U11783 (N_11783,N_9224,N_8990);
xor U11784 (N_11784,N_9673,N_9391);
nand U11785 (N_11785,N_9883,N_8830);
xnor U11786 (N_11786,N_9260,N_8663);
nor U11787 (N_11787,N_9189,N_9124);
and U11788 (N_11788,N_9856,N_9585);
nand U11789 (N_11789,N_8316,N_9002);
or U11790 (N_11790,N_9792,N_9208);
or U11791 (N_11791,N_8209,N_8378);
or U11792 (N_11792,N_9066,N_8878);
xnor U11793 (N_11793,N_9869,N_8183);
xnor U11794 (N_11794,N_8081,N_8439);
xnor U11795 (N_11795,N_8372,N_8594);
nor U11796 (N_11796,N_8680,N_9920);
nor U11797 (N_11797,N_9184,N_8879);
or U11798 (N_11798,N_9992,N_9609);
and U11799 (N_11799,N_8826,N_9192);
and U11800 (N_11800,N_8008,N_9643);
nand U11801 (N_11801,N_8901,N_8917);
nand U11802 (N_11802,N_8939,N_9998);
and U11803 (N_11803,N_8907,N_9053);
and U11804 (N_11804,N_8381,N_8045);
nor U11805 (N_11805,N_8104,N_8006);
xnor U11806 (N_11806,N_8051,N_8305);
nand U11807 (N_11807,N_9353,N_8538);
nor U11808 (N_11808,N_9845,N_9986);
and U11809 (N_11809,N_9753,N_8764);
or U11810 (N_11810,N_8294,N_9198);
nor U11811 (N_11811,N_8158,N_8593);
nand U11812 (N_11812,N_9141,N_8700);
xor U11813 (N_11813,N_8796,N_9107);
nand U11814 (N_11814,N_9891,N_9791);
or U11815 (N_11815,N_8446,N_9671);
or U11816 (N_11816,N_9244,N_9075);
xnor U11817 (N_11817,N_8147,N_9431);
or U11818 (N_11818,N_8261,N_8825);
and U11819 (N_11819,N_8036,N_9986);
nor U11820 (N_11820,N_9768,N_8971);
nand U11821 (N_11821,N_9306,N_8173);
xor U11822 (N_11822,N_8287,N_9705);
nand U11823 (N_11823,N_9668,N_9200);
or U11824 (N_11824,N_9503,N_8283);
nand U11825 (N_11825,N_8711,N_8137);
or U11826 (N_11826,N_8048,N_9243);
and U11827 (N_11827,N_9136,N_9780);
and U11828 (N_11828,N_8177,N_9170);
nor U11829 (N_11829,N_9690,N_8635);
xnor U11830 (N_11830,N_8983,N_9834);
nor U11831 (N_11831,N_9775,N_9046);
or U11832 (N_11832,N_9653,N_9078);
nand U11833 (N_11833,N_9019,N_9463);
nor U11834 (N_11834,N_9542,N_9327);
and U11835 (N_11835,N_9703,N_8572);
and U11836 (N_11836,N_8549,N_9533);
and U11837 (N_11837,N_8409,N_8572);
xnor U11838 (N_11838,N_8698,N_8321);
or U11839 (N_11839,N_9123,N_9321);
or U11840 (N_11840,N_9341,N_8478);
and U11841 (N_11841,N_8788,N_8406);
nand U11842 (N_11842,N_8384,N_8667);
and U11843 (N_11843,N_8975,N_8987);
or U11844 (N_11844,N_9491,N_8930);
xnor U11845 (N_11845,N_9145,N_8664);
nor U11846 (N_11846,N_8893,N_9365);
and U11847 (N_11847,N_8472,N_8632);
nor U11848 (N_11848,N_8029,N_8083);
nand U11849 (N_11849,N_8603,N_9105);
nand U11850 (N_11850,N_8648,N_8049);
or U11851 (N_11851,N_8992,N_9484);
nand U11852 (N_11852,N_9978,N_8469);
or U11853 (N_11853,N_9290,N_8696);
nand U11854 (N_11854,N_8706,N_9247);
xor U11855 (N_11855,N_8935,N_8482);
and U11856 (N_11856,N_9774,N_8218);
nand U11857 (N_11857,N_9353,N_8426);
nor U11858 (N_11858,N_9644,N_9243);
and U11859 (N_11859,N_8233,N_8884);
nand U11860 (N_11860,N_8464,N_9307);
nor U11861 (N_11861,N_8059,N_9256);
xnor U11862 (N_11862,N_9744,N_8633);
nor U11863 (N_11863,N_9528,N_8420);
xor U11864 (N_11864,N_9829,N_9445);
nand U11865 (N_11865,N_8219,N_8534);
or U11866 (N_11866,N_9924,N_8639);
nand U11867 (N_11867,N_9116,N_9552);
and U11868 (N_11868,N_9042,N_8450);
or U11869 (N_11869,N_9773,N_8088);
and U11870 (N_11870,N_9616,N_9449);
or U11871 (N_11871,N_8610,N_8719);
nor U11872 (N_11872,N_8541,N_8241);
xor U11873 (N_11873,N_8981,N_9240);
nand U11874 (N_11874,N_9529,N_8455);
xor U11875 (N_11875,N_9081,N_8283);
or U11876 (N_11876,N_9030,N_9174);
or U11877 (N_11877,N_8229,N_9786);
and U11878 (N_11878,N_8883,N_8112);
nor U11879 (N_11879,N_9830,N_8775);
nor U11880 (N_11880,N_8650,N_8013);
nor U11881 (N_11881,N_9298,N_9671);
and U11882 (N_11882,N_9803,N_8804);
nor U11883 (N_11883,N_8658,N_9974);
xnor U11884 (N_11884,N_9691,N_8633);
xor U11885 (N_11885,N_9712,N_8406);
or U11886 (N_11886,N_9217,N_9638);
xor U11887 (N_11887,N_8527,N_9649);
xnor U11888 (N_11888,N_9341,N_9373);
or U11889 (N_11889,N_9882,N_8169);
or U11890 (N_11890,N_8668,N_8304);
nand U11891 (N_11891,N_8465,N_8668);
nand U11892 (N_11892,N_8310,N_9023);
or U11893 (N_11893,N_9365,N_9129);
xor U11894 (N_11894,N_9765,N_9863);
and U11895 (N_11895,N_8859,N_8004);
xor U11896 (N_11896,N_8525,N_8495);
xnor U11897 (N_11897,N_8748,N_8777);
nor U11898 (N_11898,N_8641,N_9910);
or U11899 (N_11899,N_9470,N_9724);
or U11900 (N_11900,N_9242,N_9446);
nand U11901 (N_11901,N_8680,N_9041);
nor U11902 (N_11902,N_8943,N_8790);
and U11903 (N_11903,N_8662,N_8888);
nand U11904 (N_11904,N_8670,N_8789);
or U11905 (N_11905,N_9746,N_9673);
xnor U11906 (N_11906,N_9014,N_8589);
and U11907 (N_11907,N_8151,N_8217);
or U11908 (N_11908,N_8211,N_9819);
or U11909 (N_11909,N_9872,N_9959);
and U11910 (N_11910,N_8346,N_8436);
xor U11911 (N_11911,N_9411,N_9875);
nand U11912 (N_11912,N_8633,N_8166);
or U11913 (N_11913,N_8712,N_9078);
xnor U11914 (N_11914,N_9683,N_8922);
nor U11915 (N_11915,N_9762,N_8824);
nand U11916 (N_11916,N_9838,N_8067);
and U11917 (N_11917,N_9875,N_8268);
xor U11918 (N_11918,N_8163,N_8624);
nand U11919 (N_11919,N_9663,N_8016);
nand U11920 (N_11920,N_8897,N_9567);
xnor U11921 (N_11921,N_9885,N_9268);
and U11922 (N_11922,N_9294,N_9849);
or U11923 (N_11923,N_8656,N_8667);
nand U11924 (N_11924,N_8070,N_8775);
xnor U11925 (N_11925,N_8379,N_8201);
and U11926 (N_11926,N_8710,N_9428);
and U11927 (N_11927,N_8775,N_8194);
and U11928 (N_11928,N_8058,N_8900);
xor U11929 (N_11929,N_8983,N_8328);
nand U11930 (N_11930,N_8698,N_9006);
nand U11931 (N_11931,N_8238,N_8577);
and U11932 (N_11932,N_9946,N_8816);
nor U11933 (N_11933,N_9571,N_9495);
nor U11934 (N_11934,N_9824,N_8433);
nand U11935 (N_11935,N_9394,N_8799);
nor U11936 (N_11936,N_9036,N_9603);
or U11937 (N_11937,N_9261,N_9466);
nor U11938 (N_11938,N_9122,N_9806);
nand U11939 (N_11939,N_8948,N_8900);
nor U11940 (N_11940,N_9955,N_8884);
nand U11941 (N_11941,N_8127,N_9671);
or U11942 (N_11942,N_8821,N_9327);
xnor U11943 (N_11943,N_8301,N_8082);
nand U11944 (N_11944,N_9472,N_9578);
nand U11945 (N_11945,N_8886,N_8340);
and U11946 (N_11946,N_8183,N_9364);
nor U11947 (N_11947,N_8701,N_8959);
nor U11948 (N_11948,N_9984,N_8306);
xor U11949 (N_11949,N_9959,N_8254);
nor U11950 (N_11950,N_8456,N_9233);
nand U11951 (N_11951,N_8326,N_8976);
nand U11952 (N_11952,N_8450,N_9666);
or U11953 (N_11953,N_8800,N_8137);
nor U11954 (N_11954,N_9684,N_9359);
nand U11955 (N_11955,N_9502,N_8186);
xor U11956 (N_11956,N_9186,N_8873);
or U11957 (N_11957,N_8458,N_8446);
xor U11958 (N_11958,N_9006,N_9223);
nor U11959 (N_11959,N_9541,N_8343);
xor U11960 (N_11960,N_8342,N_8515);
nand U11961 (N_11961,N_9617,N_8294);
or U11962 (N_11962,N_9354,N_8525);
nor U11963 (N_11963,N_8407,N_8096);
or U11964 (N_11964,N_9883,N_8169);
xor U11965 (N_11965,N_9880,N_9724);
and U11966 (N_11966,N_8456,N_8892);
or U11967 (N_11967,N_8724,N_9843);
or U11968 (N_11968,N_8753,N_8006);
or U11969 (N_11969,N_8607,N_9921);
xnor U11970 (N_11970,N_8098,N_9827);
xnor U11971 (N_11971,N_8474,N_9190);
nand U11972 (N_11972,N_8505,N_8299);
and U11973 (N_11973,N_8397,N_8563);
nand U11974 (N_11974,N_9343,N_9264);
nor U11975 (N_11975,N_8304,N_9251);
xnor U11976 (N_11976,N_9420,N_8745);
nand U11977 (N_11977,N_9343,N_8366);
nand U11978 (N_11978,N_9778,N_9708);
nand U11979 (N_11979,N_9924,N_8702);
xnor U11980 (N_11980,N_8646,N_8432);
or U11981 (N_11981,N_9835,N_9900);
nor U11982 (N_11982,N_9387,N_8678);
and U11983 (N_11983,N_8030,N_8374);
or U11984 (N_11984,N_8357,N_8987);
nor U11985 (N_11985,N_8049,N_8551);
xnor U11986 (N_11986,N_8331,N_9637);
and U11987 (N_11987,N_9256,N_9904);
or U11988 (N_11988,N_8283,N_8708);
xor U11989 (N_11989,N_9928,N_8756);
or U11990 (N_11990,N_8360,N_9835);
xor U11991 (N_11991,N_9337,N_9532);
nor U11992 (N_11992,N_8879,N_9343);
xor U11993 (N_11993,N_9894,N_8526);
or U11994 (N_11994,N_9590,N_9483);
xor U11995 (N_11995,N_8862,N_8301);
and U11996 (N_11996,N_9952,N_8273);
or U11997 (N_11997,N_9518,N_9849);
xnor U11998 (N_11998,N_9421,N_9734);
or U11999 (N_11999,N_9355,N_9337);
nor U12000 (N_12000,N_10763,N_11914);
nor U12001 (N_12001,N_11484,N_10781);
or U12002 (N_12002,N_11593,N_10179);
or U12003 (N_12003,N_11241,N_11079);
nand U12004 (N_12004,N_11600,N_10320);
nand U12005 (N_12005,N_11985,N_11024);
xnor U12006 (N_12006,N_10548,N_11367);
nand U12007 (N_12007,N_11181,N_10856);
and U12008 (N_12008,N_11917,N_10576);
and U12009 (N_12009,N_11143,N_10828);
or U12010 (N_12010,N_10500,N_10916);
or U12011 (N_12011,N_11696,N_11651);
or U12012 (N_12012,N_10988,N_10526);
nand U12013 (N_12013,N_11277,N_11062);
nor U12014 (N_12014,N_10051,N_11787);
and U12015 (N_12015,N_10744,N_11773);
and U12016 (N_12016,N_11476,N_10274);
or U12017 (N_12017,N_10951,N_11782);
xor U12018 (N_12018,N_11247,N_11388);
or U12019 (N_12019,N_11092,N_11950);
and U12020 (N_12020,N_10260,N_10296);
and U12021 (N_12021,N_10643,N_11621);
and U12022 (N_12022,N_10058,N_11262);
or U12023 (N_12023,N_10886,N_10559);
and U12024 (N_12024,N_10146,N_10417);
xor U12025 (N_12025,N_11995,N_11620);
or U12026 (N_12026,N_10242,N_11123);
or U12027 (N_12027,N_11330,N_11242);
or U12028 (N_12028,N_10771,N_10852);
and U12029 (N_12029,N_11137,N_10780);
or U12030 (N_12030,N_10101,N_10129);
nor U12031 (N_12031,N_10564,N_11148);
and U12032 (N_12032,N_10449,N_11477);
nor U12033 (N_12033,N_10419,N_10445);
xor U12034 (N_12034,N_11341,N_10271);
nor U12035 (N_12035,N_11231,N_11552);
or U12036 (N_12036,N_11912,N_10261);
or U12037 (N_12037,N_10008,N_10117);
xor U12038 (N_12038,N_10055,N_10778);
or U12039 (N_12039,N_11580,N_10741);
xnor U12040 (N_12040,N_10562,N_11776);
xnor U12041 (N_12041,N_11847,N_10821);
nand U12042 (N_12042,N_10357,N_11276);
or U12043 (N_12043,N_10048,N_10790);
nand U12044 (N_12044,N_10710,N_11035);
xnor U12045 (N_12045,N_11564,N_10577);
nor U12046 (N_12046,N_11952,N_11350);
and U12047 (N_12047,N_10388,N_11984);
or U12048 (N_12048,N_10553,N_10441);
nor U12049 (N_12049,N_11465,N_10703);
nand U12050 (N_12050,N_11257,N_11043);
nand U12051 (N_12051,N_11415,N_10334);
nor U12052 (N_12052,N_11097,N_10869);
nor U12053 (N_12053,N_11106,N_11141);
xor U12054 (N_12054,N_11509,N_11044);
xnor U12055 (N_12055,N_11048,N_10862);
xnor U12056 (N_12056,N_11941,N_11969);
nor U12057 (N_12057,N_10481,N_11215);
and U12058 (N_12058,N_10620,N_10226);
and U12059 (N_12059,N_10606,N_11925);
xor U12060 (N_12060,N_11358,N_10377);
xnor U12061 (N_12061,N_11523,N_10695);
or U12062 (N_12062,N_10994,N_11928);
nor U12063 (N_12063,N_10541,N_11757);
nor U12064 (N_12064,N_10599,N_10372);
nor U12065 (N_12065,N_11189,N_11193);
nand U12066 (N_12066,N_11260,N_10955);
nor U12067 (N_12067,N_11034,N_10996);
nand U12068 (N_12068,N_10777,N_10196);
nor U12069 (N_12069,N_11646,N_10454);
nand U12070 (N_12070,N_10718,N_11308);
nand U12071 (N_12071,N_11582,N_11938);
nor U12072 (N_12072,N_10857,N_11485);
nand U12073 (N_12073,N_10642,N_11986);
nand U12074 (N_12074,N_11012,N_11404);
and U12075 (N_12075,N_10505,N_11587);
and U12076 (N_12076,N_10430,N_10939);
or U12077 (N_12077,N_11864,N_11547);
nor U12078 (N_12078,N_11921,N_11820);
or U12079 (N_12079,N_10268,N_11434);
or U12080 (N_12080,N_10975,N_10211);
or U12081 (N_12081,N_10387,N_10344);
or U12082 (N_12082,N_10640,N_11529);
xor U12083 (N_12083,N_10265,N_11220);
or U12084 (N_12084,N_10518,N_11296);
nand U12085 (N_12085,N_10414,N_10169);
and U12086 (N_12086,N_10085,N_11674);
nor U12087 (N_12087,N_11566,N_10880);
nand U12088 (N_12088,N_10711,N_11441);
xor U12089 (N_12089,N_11899,N_10890);
nor U12090 (N_12090,N_10533,N_10561);
nand U12091 (N_12091,N_10183,N_11882);
and U12092 (N_12092,N_11433,N_11107);
nor U12093 (N_12093,N_11115,N_10749);
xor U12094 (N_12094,N_11307,N_10650);
nand U12095 (N_12095,N_11890,N_11119);
nor U12096 (N_12096,N_10484,N_11187);
xor U12097 (N_12097,N_10495,N_10425);
nand U12098 (N_12098,N_10941,N_10927);
or U12099 (N_12099,N_10760,N_10090);
and U12100 (N_12100,N_10841,N_10231);
or U12101 (N_12101,N_11069,N_10701);
and U12102 (N_12102,N_11480,N_11692);
xor U12103 (N_12103,N_10350,N_11759);
nand U12104 (N_12104,N_11709,N_11101);
or U12105 (N_12105,N_10486,N_10240);
xnor U12106 (N_12106,N_10670,N_10096);
xor U12107 (N_12107,N_11020,N_11103);
and U12108 (N_12108,N_11936,N_10970);
or U12109 (N_12109,N_11660,N_10367);
and U12110 (N_12110,N_11518,N_11526);
nand U12111 (N_12111,N_10833,N_10250);
and U12112 (N_12112,N_11364,N_11629);
nand U12113 (N_12113,N_11288,N_10931);
and U12114 (N_12114,N_10433,N_10194);
nor U12115 (N_12115,N_11573,N_10865);
or U12116 (N_12116,N_10012,N_11511);
or U12117 (N_12117,N_11769,N_10832);
or U12118 (N_12118,N_11129,N_11727);
nand U12119 (N_12119,N_11852,N_10903);
nor U12120 (N_12120,N_10630,N_11319);
and U12121 (N_12121,N_10379,N_10013);
nor U12122 (N_12122,N_10794,N_11033);
nor U12123 (N_12123,N_10732,N_11205);
nand U12124 (N_12124,N_11647,N_10512);
nor U12125 (N_12125,N_11948,N_11046);
nor U12126 (N_12126,N_11027,N_10788);
nor U12127 (N_12127,N_10629,N_11344);
xor U12128 (N_12128,N_11543,N_11520);
nor U12129 (N_12129,N_11963,N_11091);
nand U12130 (N_12130,N_10646,N_11830);
nor U12131 (N_12131,N_10950,N_11156);
xor U12132 (N_12132,N_10390,N_10340);
nand U12133 (N_12133,N_11184,N_10587);
nor U12134 (N_12134,N_10581,N_10727);
and U12135 (N_12135,N_11720,N_10607);
xor U12136 (N_12136,N_11779,N_11318);
nand U12137 (N_12137,N_11239,N_10256);
nor U12138 (N_12138,N_10913,N_11606);
nand U12139 (N_12139,N_11849,N_10847);
and U12140 (N_12140,N_11562,N_10397);
xnor U12141 (N_12141,N_11083,N_10990);
nor U12142 (N_12142,N_10259,N_11706);
nand U12143 (N_12143,N_10917,N_11152);
nor U12144 (N_12144,N_10353,N_10187);
and U12145 (N_12145,N_11267,N_10122);
xnor U12146 (N_12146,N_11322,N_10653);
or U12147 (N_12147,N_11366,N_11530);
and U12148 (N_12148,N_11884,N_11352);
and U12149 (N_12149,N_11274,N_11466);
xnor U12150 (N_12150,N_10336,N_10962);
and U12151 (N_12151,N_11351,N_11596);
xnor U12152 (N_12152,N_11841,N_10195);
xnor U12153 (N_12153,N_10509,N_11142);
nor U12154 (N_12154,N_10470,N_10567);
xnor U12155 (N_12155,N_10027,N_11817);
or U12156 (N_12156,N_10635,N_10068);
or U12157 (N_12157,N_10172,N_11204);
or U12158 (N_12158,N_11462,N_10074);
nand U12159 (N_12159,N_10306,N_10693);
xnor U12160 (N_12160,N_10210,N_10091);
nand U12161 (N_12161,N_11336,N_11812);
xor U12162 (N_12162,N_11805,N_10991);
nor U12163 (N_12163,N_11694,N_10522);
nor U12164 (N_12164,N_11829,N_10477);
and U12165 (N_12165,N_11569,N_10901);
and U12166 (N_12166,N_11872,N_11022);
and U12167 (N_12167,N_11042,N_11321);
and U12168 (N_12168,N_10099,N_11784);
xnor U12169 (N_12169,N_10382,N_11377);
and U12170 (N_12170,N_10675,N_10077);
nand U12171 (N_12171,N_11512,N_11655);
or U12172 (N_12172,N_10300,N_10983);
and U12173 (N_12173,N_11454,N_10097);
and U12174 (N_12174,N_11954,N_11290);
or U12175 (N_12175,N_11907,N_11471);
and U12176 (N_12176,N_11677,N_11447);
or U12177 (N_12177,N_11634,N_10656);
nand U12178 (N_12178,N_10582,N_11534);
or U12179 (N_12179,N_10960,N_10060);
or U12180 (N_12180,N_10621,N_10592);
and U12181 (N_12181,N_11117,N_11036);
xnor U12182 (N_12182,N_10685,N_11831);
or U12183 (N_12183,N_11394,N_11765);
nand U12184 (N_12184,N_10396,N_10283);
and U12185 (N_12185,N_10861,N_11836);
nor U12186 (N_12186,N_10839,N_11889);
nand U12187 (N_12187,N_10918,N_11126);
and U12188 (N_12188,N_11935,N_11924);
xnor U12189 (N_12189,N_11312,N_11113);
nor U12190 (N_12190,N_10779,N_11934);
or U12191 (N_12191,N_11329,N_11082);
or U12192 (N_12192,N_10059,N_11370);
xnor U12193 (N_12193,N_10128,N_11248);
or U12194 (N_12194,N_11088,N_11704);
nor U12195 (N_12195,N_11521,N_10978);
nand U12196 (N_12196,N_11541,N_11444);
or U12197 (N_12197,N_11347,N_11681);
or U12198 (N_12198,N_11056,N_11893);
xor U12199 (N_12199,N_11631,N_10932);
nor U12200 (N_12200,N_10520,N_11000);
nor U12201 (N_12201,N_11977,N_11237);
nor U12202 (N_12202,N_10020,N_10885);
xor U12203 (N_12203,N_10747,N_10733);
or U12204 (N_12204,N_11616,N_10722);
or U12205 (N_12205,N_10514,N_10007);
nand U12206 (N_12206,N_11284,N_10258);
and U12207 (N_12207,N_10282,N_10787);
nor U12208 (N_12208,N_10106,N_11653);
nand U12209 (N_12209,N_11008,N_11559);
nor U12210 (N_12210,N_11942,N_10442);
or U12211 (N_12211,N_11363,N_11640);
nand U12212 (N_12212,N_11980,N_11240);
nor U12213 (N_12213,N_11075,N_11609);
nand U12214 (N_12214,N_11275,N_10603);
or U12215 (N_12215,N_11424,N_10228);
xor U12216 (N_12216,N_10114,N_11806);
nor U12217 (N_12217,N_10536,N_10174);
and U12218 (N_12218,N_10017,N_10806);
or U12219 (N_12219,N_11158,N_10203);
and U12220 (N_12220,N_11125,N_11268);
nand U12221 (N_12221,N_10432,N_10384);
or U12222 (N_12222,N_10023,N_10318);
xnor U12223 (N_12223,N_11081,N_10827);
nand U12224 (N_12224,N_10698,N_10699);
or U12225 (N_12225,N_11865,N_10768);
nor U12226 (N_12226,N_11226,N_11737);
or U12227 (N_12227,N_10288,N_11555);
and U12228 (N_12228,N_11315,N_10123);
and U12229 (N_12229,N_11598,N_10598);
and U12230 (N_12230,N_10467,N_11228);
nand U12231 (N_12231,N_11061,N_10403);
nor U12232 (N_12232,N_11910,N_10823);
xor U12233 (N_12233,N_11168,N_11519);
or U12234 (N_12234,N_11915,N_11497);
xnor U12235 (N_12235,N_11554,N_10108);
nand U12236 (N_12236,N_10801,N_10895);
nor U12237 (N_12237,N_10785,N_11293);
xnor U12238 (N_12238,N_10907,N_10158);
nand U12239 (N_12239,N_11828,N_11725);
nand U12240 (N_12240,N_10112,N_11084);
nor U12241 (N_12241,N_11111,N_10444);
and U12242 (N_12242,N_11968,N_11197);
and U12243 (N_12243,N_10623,N_10399);
or U12244 (N_12244,N_11902,N_10906);
xnor U12245 (N_12245,N_10767,N_10748);
nand U12246 (N_12246,N_11099,N_10715);
or U12247 (N_12247,N_11846,N_11507);
xor U12248 (N_12248,N_11861,N_11951);
or U12249 (N_12249,N_11064,N_11823);
xnor U12250 (N_12250,N_10596,N_11933);
xnor U12251 (N_12251,N_11104,N_11513);
or U12252 (N_12252,N_11208,N_11906);
xor U12253 (N_12253,N_11987,N_10042);
nor U12254 (N_12254,N_11516,N_11316);
nand U12255 (N_12255,N_11926,N_10424);
or U12256 (N_12256,N_10914,N_11567);
nand U12257 (N_12257,N_10070,N_10871);
nor U12258 (N_12258,N_11793,N_10947);
xor U12259 (N_12259,N_11649,N_11203);
and U12260 (N_12260,N_10443,N_11261);
xnor U12261 (N_12261,N_10651,N_10859);
xnor U12262 (N_12262,N_10659,N_11401);
nor U12263 (N_12263,N_11147,N_10759);
nand U12264 (N_12264,N_10578,N_10864);
or U12265 (N_12265,N_11071,N_11362);
or U12266 (N_12266,N_10073,N_11353);
nand U12267 (N_12267,N_10648,N_10243);
xnor U12268 (N_12268,N_10052,N_10595);
or U12269 (N_12269,N_11688,N_11916);
xor U12270 (N_12270,N_10873,N_11630);
and U12271 (N_12271,N_11739,N_10753);
xnor U12272 (N_12272,N_11488,N_10440);
nand U12273 (N_12273,N_11932,N_10661);
nor U12274 (N_12274,N_10611,N_11810);
xnor U12275 (N_12275,N_10363,N_11764);
nand U12276 (N_12276,N_11221,N_11473);
nor U12277 (N_12277,N_11689,N_10180);
xor U12278 (N_12278,N_11334,N_10339);
nand U12279 (N_12279,N_11929,N_10963);
or U12280 (N_12280,N_10789,N_10819);
or U12281 (N_12281,N_10290,N_10930);
xnor U12282 (N_12282,N_10157,N_10152);
nand U12283 (N_12283,N_11326,N_11604);
xnor U12284 (N_12284,N_11964,N_11051);
nor U12285 (N_12285,N_11379,N_11775);
and U12286 (N_12286,N_11766,N_11427);
and U12287 (N_12287,N_11338,N_11668);
or U12288 (N_12288,N_10757,N_10908);
and U12289 (N_12289,N_11430,N_11486);
nand U12290 (N_12290,N_10116,N_11032);
nor U12291 (N_12291,N_11273,N_10884);
xnor U12292 (N_12292,N_10280,N_10657);
and U12293 (N_12293,N_11230,N_10186);
nor U12294 (N_12294,N_10079,N_10984);
xnor U12295 (N_12295,N_10507,N_11762);
xor U12296 (N_12296,N_10791,N_11632);
or U12297 (N_12297,N_10054,N_11007);
or U12298 (N_12298,N_10673,N_10126);
xor U12299 (N_12299,N_11687,N_11816);
or U12300 (N_12300,N_11613,N_10050);
nor U12301 (N_12301,N_11368,N_10198);
nor U12302 (N_12302,N_11713,N_10822);
xnor U12303 (N_12303,N_11992,N_10310);
and U12304 (N_12304,N_11186,N_10022);
xnor U12305 (N_12305,N_10949,N_11154);
or U12306 (N_12306,N_10549,N_11654);
nor U12307 (N_12307,N_10893,N_10145);
and U12308 (N_12308,N_10010,N_11055);
and U12309 (N_12309,N_10076,N_10540);
nor U12310 (N_12310,N_10330,N_11741);
or U12311 (N_12311,N_11063,N_10229);
nand U12312 (N_12312,N_11461,N_10478);
or U12313 (N_12313,N_10537,N_10874);
xor U12314 (N_12314,N_11973,N_10800);
nor U12315 (N_12315,N_10840,N_11381);
nor U12316 (N_12316,N_11839,N_10406);
xor U12317 (N_12317,N_10824,N_11525);
and U12318 (N_12318,N_10876,N_11417);
nand U12319 (N_12319,N_11858,N_10503);
or U12320 (N_12320,N_10115,N_10466);
or U12321 (N_12321,N_11535,N_10804);
and U12322 (N_12322,N_10735,N_10795);
or U12323 (N_12323,N_11392,N_11191);
nor U12324 (N_12324,N_11149,N_10737);
nor U12325 (N_12325,N_10053,N_10622);
nor U12326 (N_12326,N_10143,N_10047);
nor U12327 (N_12327,N_11328,N_11978);
or U12328 (N_12328,N_11445,N_10121);
xor U12329 (N_12329,N_11223,N_10181);
or U12330 (N_12330,N_10161,N_11999);
nor U12331 (N_12331,N_10566,N_10929);
nand U12332 (N_12332,N_10545,N_11734);
nor U12333 (N_12333,N_11845,N_11502);
xnor U12334 (N_12334,N_10867,N_10408);
or U12335 (N_12335,N_11908,N_10401);
xor U12336 (N_12336,N_11834,N_10057);
and U12337 (N_12337,N_11481,N_10738);
nand U12338 (N_12338,N_10304,N_10437);
and U12339 (N_12339,N_11021,N_11431);
nand U12340 (N_12340,N_10998,N_10750);
nand U12341 (N_12341,N_10168,N_10618);
and U12342 (N_12342,N_10029,N_10345);
and U12343 (N_12343,N_11570,N_10402);
nand U12344 (N_12344,N_10523,N_10257);
or U12345 (N_12345,N_10585,N_10579);
xnor U12346 (N_12346,N_10035,N_11626);
xor U12347 (N_12347,N_11453,N_11232);
or U12348 (N_12348,N_11015,N_11278);
and U12349 (N_12349,N_11151,N_11642);
or U12350 (N_12350,N_11238,N_11174);
and U12351 (N_12351,N_10617,N_10217);
nand U12352 (N_12352,N_10634,N_11699);
xnor U12353 (N_12353,N_10391,N_10316);
nand U12354 (N_12354,N_10993,N_11023);
nor U12355 (N_12355,N_10758,N_10667);
or U12356 (N_12356,N_10594,N_11648);
xnor U12357 (N_12357,N_10851,N_11542);
nand U12358 (N_12358,N_11611,N_10359);
xor U12359 (N_12359,N_10665,N_11073);
nor U12360 (N_12360,N_11196,N_10574);
xnor U12361 (N_12361,N_11505,N_10644);
nor U12362 (N_12362,N_10527,N_10797);
xnor U12363 (N_12363,N_10385,N_11300);
nor U12364 (N_12364,N_10669,N_11735);
nand U12365 (N_12365,N_11059,N_11705);
nand U12366 (N_12366,N_11931,N_10080);
and U12367 (N_12367,N_10016,N_11877);
xor U12368 (N_12368,N_11470,N_10696);
xnor U12369 (N_12369,N_11072,N_10153);
and U12370 (N_12370,N_10775,N_11639);
nand U12371 (N_12371,N_11801,N_11691);
nor U12372 (N_12372,N_11803,N_11819);
and U12373 (N_12373,N_10515,N_11774);
and U12374 (N_12374,N_11335,N_11900);
and U12375 (N_12375,N_10506,N_11393);
and U12376 (N_12376,N_11905,N_10365);
and U12377 (N_12377,N_11491,N_11815);
or U12378 (N_12378,N_11291,N_11718);
nor U12379 (N_12379,N_10393,N_11348);
xnor U12380 (N_12380,N_10147,N_10191);
nor U12381 (N_12381,N_10275,N_11991);
nand U12382 (N_12382,N_10909,N_11665);
xnor U12383 (N_12383,N_10784,N_10429);
and U12384 (N_12384,N_11961,N_10590);
or U12385 (N_12385,N_10378,N_10376);
nor U12386 (N_12386,N_11545,N_10298);
or U12387 (N_12387,N_10660,N_11589);
nor U12388 (N_12388,N_11749,N_10739);
xor U12389 (N_12389,N_11965,N_10683);
or U12390 (N_12390,N_10754,N_11904);
nand U12391 (N_12391,N_11792,N_11711);
or U12392 (N_12392,N_10586,N_10619);
nor U12393 (N_12393,N_11093,N_10473);
nand U12394 (N_12394,N_10149,N_10654);
or U12395 (N_12395,N_11493,N_11678);
and U12396 (N_12396,N_11057,N_10138);
nand U12397 (N_12397,N_11324,N_11575);
nand U12398 (N_12398,N_10065,N_11994);
and U12399 (N_12399,N_11478,N_11854);
and U12400 (N_12400,N_11612,N_11435);
and U12401 (N_12401,N_11795,N_11294);
nand U12402 (N_12402,N_10912,N_10166);
nand U12403 (N_12403,N_10421,N_10597);
and U12404 (N_12404,N_11423,N_11586);
nand U12405 (N_12405,N_11579,N_11039);
and U12406 (N_12406,N_11581,N_10647);
nand U12407 (N_12407,N_11550,N_11971);
nor U12408 (N_12408,N_11661,N_10286);
or U12409 (N_12409,N_10066,N_10766);
nor U12410 (N_12410,N_11199,N_11474);
nor U12411 (N_12411,N_10850,N_10986);
nor U12412 (N_12412,N_10360,N_11332);
nand U12413 (N_12413,N_11558,N_10462);
and U12414 (N_12414,N_10538,N_10207);
nor U12415 (N_12415,N_11594,N_11871);
xor U12416 (N_12416,N_10616,N_11498);
xor U12417 (N_12417,N_11078,N_10628);
nand U12418 (N_12418,N_11159,N_11745);
nor U12419 (N_12419,N_11826,N_10571);
and U12420 (N_12420,N_11420,N_11878);
nor U12421 (N_12421,N_10273,N_11173);
and U12422 (N_12422,N_10381,N_11644);
nor U12423 (N_12423,N_10105,N_11369);
and U12424 (N_12424,N_10302,N_10689);
or U12425 (N_12425,N_10413,N_11599);
xnor U12426 (N_12426,N_10252,N_10206);
and U12427 (N_12427,N_11967,N_10019);
xor U12428 (N_12428,N_10362,N_11627);
xnor U12429 (N_12429,N_10925,N_10093);
nor U12430 (N_12430,N_10992,N_10855);
nor U12431 (N_12431,N_11058,N_10463);
nand U12432 (N_12432,N_11708,N_10854);
nor U12433 (N_12433,N_10171,N_10033);
and U12434 (N_12434,N_10151,N_11443);
xor U12435 (N_12435,N_10528,N_10919);
nor U12436 (N_12436,N_10036,N_11391);
and U12437 (N_12437,N_10610,N_11998);
and U12438 (N_12438,N_10411,N_10317);
and U12439 (N_12439,N_10863,N_11120);
and U12440 (N_12440,N_10144,N_11747);
nor U12441 (N_12441,N_10793,N_10087);
xnor U12442 (N_12442,N_11376,N_11279);
and U12443 (N_12443,N_11402,N_11337);
nor U12444 (N_12444,N_10072,N_11508);
nand U12445 (N_12445,N_10104,N_11074);
xor U12446 (N_12446,N_11659,N_11603);
xnor U12447 (N_12447,N_11755,N_10835);
and U12448 (N_12448,N_11625,N_11956);
or U12449 (N_12449,N_10573,N_11047);
xor U12450 (N_12450,N_11177,N_10707);
nand U12451 (N_12451,N_11780,N_11359);
xnor U12452 (N_12452,N_11601,N_10636);
nand U12453 (N_12453,N_10083,N_11354);
xnor U12454 (N_12454,N_10358,N_11517);
nor U12455 (N_12455,N_10215,N_10038);
nor U12456 (N_12456,N_10327,N_10428);
nand U12457 (N_12457,N_11456,N_11698);
or U12458 (N_12458,N_10740,N_11732);
xnor U12459 (N_12459,N_11450,N_11229);
and U12460 (N_12460,N_10879,N_11763);
nor U12461 (N_12461,N_11894,N_11982);
xor U12462 (N_12462,N_11467,N_11683);
nor U12463 (N_12463,N_11669,N_10844);
nor U12464 (N_12464,N_11179,N_10551);
nor U12465 (N_12465,N_10124,N_10255);
or U12466 (N_12466,N_11038,N_10380);
nand U12467 (N_12467,N_11306,N_11459);
nor U12468 (N_12468,N_10434,N_11707);
nor U12469 (N_12469,N_11853,N_11213);
or U12470 (N_12470,N_10221,N_11145);
or U12471 (N_12471,N_10631,N_10245);
or U12472 (N_12472,N_10026,N_10920);
nor U12473 (N_12473,N_10639,N_10713);
nand U12474 (N_12474,N_11198,N_10882);
and U12475 (N_12475,N_10468,N_10067);
nand U12476 (N_12476,N_10614,N_11469);
and U12477 (N_12477,N_10349,N_10281);
nor U12478 (N_12478,N_11472,N_11052);
nand U12479 (N_12479,N_10728,N_11325);
nand U12480 (N_12480,N_10626,N_10770);
xor U12481 (N_12481,N_10973,N_10830);
nor U12482 (N_12482,N_10453,N_10299);
nor U12483 (N_12483,N_10731,N_10405);
nand U12484 (N_12484,N_10891,N_10209);
nand U12485 (N_12485,N_11524,N_11676);
nand U12486 (N_12486,N_10006,N_10570);
and U12487 (N_12487,N_11373,N_11730);
and U12488 (N_12488,N_11037,N_10447);
xnor U12489 (N_12489,N_11605,N_10716);
xor U12490 (N_12490,N_10637,N_10246);
xnor U12491 (N_12491,N_10489,N_10589);
xnor U12492 (N_12492,N_11153,N_10999);
nor U12493 (N_12493,N_10849,N_11452);
nand U12494 (N_12494,N_11522,N_11096);
or U12495 (N_12495,N_11797,N_11723);
nand U12496 (N_12496,N_11251,N_11721);
nor U12497 (N_12497,N_10009,N_11527);
and U12498 (N_12498,N_10510,N_11372);
nor U12499 (N_12499,N_10164,N_11114);
and U12500 (N_12500,N_10061,N_11049);
or U12501 (N_12501,N_11822,N_11761);
nor U12502 (N_12502,N_10534,N_10782);
or U12503 (N_12503,N_10276,N_10346);
nand U12504 (N_12504,N_11976,N_10269);
nand U12505 (N_12505,N_10089,N_10294);
nand U12506 (N_12506,N_11411,N_11943);
xnor U12507 (N_12507,N_11171,N_11118);
xnor U12508 (N_12508,N_11395,N_11832);
nor U12509 (N_12509,N_10508,N_10469);
or U12510 (N_12510,N_11662,N_11259);
nor U12511 (N_12511,N_10724,N_11009);
nor U12512 (N_12512,N_10312,N_11164);
nand U12513 (N_12513,N_11975,N_11421);
and U12514 (N_12514,N_10039,N_11657);
and U12515 (N_12515,N_11843,N_11619);
xnor U12516 (N_12516,N_10702,N_11501);
and U12517 (N_12517,N_10981,N_11583);
nand U12518 (N_12518,N_10860,N_10452);
or U12519 (N_12519,N_11771,N_11162);
nor U12520 (N_12520,N_10723,N_10799);
nor U12521 (N_12521,N_11170,N_10450);
and U12522 (N_12522,N_10001,N_11419);
xor U12523 (N_12523,N_11413,N_11576);
or U12524 (N_12524,N_11743,N_11384);
or U12525 (N_12525,N_10292,N_11297);
nor U12526 (N_12526,N_11442,N_11235);
nand U12527 (N_12527,N_11610,N_11207);
nand U12528 (N_12528,N_10132,N_10974);
and U12529 (N_12529,N_10501,N_11989);
xnor U12530 (N_12530,N_10783,N_11236);
or U12531 (N_12531,N_11192,N_11637);
nand U12532 (N_12532,N_11243,N_11272);
or U12533 (N_12533,N_11310,N_11615);
xor U12534 (N_12534,N_11496,N_10488);
xor U12535 (N_12535,N_10805,N_10765);
or U12536 (N_12536,N_11225,N_11155);
or U12537 (N_12537,N_11770,N_10193);
and U12538 (N_12538,N_11201,N_11887);
or U12539 (N_12539,N_11695,N_10892);
nor U12540 (N_12540,N_10746,N_10369);
nand U12541 (N_12541,N_10264,N_10730);
nand U12542 (N_12542,N_11731,N_11342);
xnor U12543 (N_12543,N_10943,N_10655);
xor U12544 (N_12544,N_10810,N_11463);
or U12545 (N_12545,N_11790,N_11136);
or U12546 (N_12546,N_11077,N_11190);
nor U12547 (N_12547,N_11188,N_10905);
nor U12548 (N_12548,N_11537,N_11622);
and U12549 (N_12549,N_11227,N_11139);
and U12550 (N_12550,N_11783,N_10633);
nand U12551 (N_12551,N_11693,N_11458);
xnor U12552 (N_12552,N_10342,N_10812);
and U12553 (N_12553,N_10940,N_11269);
nand U12554 (N_12554,N_10201,N_10709);
xnor U12555 (N_12555,N_10690,N_11133);
xnor U12556 (N_12556,N_10137,N_10600);
and U12557 (N_12557,N_10959,N_10645);
or U12558 (N_12558,N_10965,N_11768);
xor U12559 (N_12559,N_11014,N_11753);
nor U12560 (N_12560,N_10110,N_11671);
and U12561 (N_12561,N_10546,N_11636);
nor U12562 (N_12562,N_10237,N_11796);
nand U12563 (N_12563,N_11135,N_10448);
nand U12564 (N_12564,N_10130,N_11446);
nand U12565 (N_12565,N_11495,N_11355);
nand U12566 (N_12566,N_10177,N_11249);
xor U12567 (N_12567,N_10813,N_11289);
xnor U12568 (N_12568,N_11311,N_10688);
and U12569 (N_12569,N_10714,N_10375);
nand U12570 (N_12570,N_10531,N_10224);
or U12571 (N_12571,N_11360,N_11788);
nor U12572 (N_12572,N_10910,N_10543);
and U12573 (N_12573,N_11426,N_10223);
nand U12574 (N_12574,N_11838,N_11608);
or U12575 (N_12575,N_11175,N_10625);
nand U12576 (N_12576,N_11019,N_10989);
nor U12577 (N_12577,N_11436,N_11959);
and U12578 (N_12578,N_10609,N_10846);
or U12579 (N_12579,N_11758,N_10355);
nand U12580 (N_12580,N_11429,N_10311);
nand U12581 (N_12581,N_10926,N_11881);
nand U12582 (N_12582,N_11303,N_10658);
nand U12583 (N_12583,N_10624,N_11209);
nand U12584 (N_12584,N_11210,N_11219);
xnor U12585 (N_12585,N_11736,N_11744);
nand U12586 (N_12586,N_11002,N_10687);
and U12587 (N_12587,N_11200,N_11005);
or U12588 (N_12588,N_10303,N_10704);
or U12589 (N_12589,N_11087,N_11286);
nor U12590 (N_12590,N_11112,N_11891);
and U12591 (N_12591,N_11403,N_10935);
nand U12592 (N_12592,N_11214,N_10967);
xnor U12593 (N_12593,N_10389,N_10208);
or U12594 (N_12594,N_11781,N_10141);
nor U12595 (N_12595,N_10325,N_10455);
xnor U12596 (N_12596,N_10572,N_10423);
xor U12597 (N_12597,N_11180,N_11528);
xor U12598 (N_12598,N_11918,N_10025);
nand U12599 (N_12599,N_11281,N_11375);
xnor U12600 (N_12600,N_11875,N_11920);
xnor U12601 (N_12601,N_11031,N_11252);
xor U12602 (N_12602,N_11652,N_11911);
nand U12603 (N_12603,N_11343,N_10118);
and U12604 (N_12604,N_10762,N_10708);
nor U12605 (N_12605,N_11825,N_11957);
nand U12606 (N_12606,N_10752,N_11479);
xor U12607 (N_12607,N_11638,N_11835);
or U12608 (N_12608,N_11538,N_11108);
nand U12609 (N_12609,N_10476,N_10555);
xnor U12610 (N_12610,N_11949,N_11799);
and U12611 (N_12611,N_11011,N_11080);
nand U12612 (N_12612,N_11658,N_11785);
xor U12613 (N_12613,N_11146,N_11110);
or U12614 (N_12614,N_10964,N_10547);
xnor U12615 (N_12615,N_10502,N_10968);
nor U12616 (N_12616,N_10911,N_11680);
nor U12617 (N_12617,N_11414,N_10313);
nand U12618 (N_12618,N_10524,N_11988);
nand U12619 (N_12619,N_11714,N_11958);
nand U12620 (N_12620,N_10004,N_10238);
and U12621 (N_12621,N_11390,N_10605);
or U12622 (N_12622,N_11396,N_10580);
or U12623 (N_12623,N_10786,N_11357);
nor U12624 (N_12624,N_10332,N_11500);
nor U12625 (N_12625,N_10485,N_10024);
or U12626 (N_12626,N_10338,N_10270);
and U12627 (N_12627,N_11244,N_10542);
or U12628 (N_12628,N_10921,N_10899);
or U12629 (N_12629,N_11161,N_11282);
nor U12630 (N_12630,N_10000,N_10808);
or U12631 (N_12631,N_11656,N_11752);
and U12632 (N_12632,N_10820,N_11844);
nand U12633 (N_12633,N_11686,N_10952);
or U12634 (N_12634,N_10836,N_10475);
nand U12635 (N_12635,N_11320,N_11955);
nor U12636 (N_12636,N_11167,N_10218);
or U12637 (N_12637,N_11025,N_10100);
and U12638 (N_12638,N_10831,N_11412);
nor U12639 (N_12639,N_11667,N_11777);
and U12640 (N_12640,N_10497,N_11449);
nor U12641 (N_12641,N_10848,N_11266);
nand U12642 (N_12642,N_10021,N_10185);
nand U12643 (N_12643,N_10769,N_10870);
xor U12644 (N_12644,N_10439,N_10818);
or U12645 (N_12645,N_10953,N_10465);
and U12646 (N_12646,N_11086,N_10889);
nand U12647 (N_12647,N_10743,N_11645);
xnor U12648 (N_12648,N_11557,N_10591);
xor U12649 (N_12649,N_11510,N_10329);
nor U12650 (N_12650,N_11880,N_11285);
xnor U12651 (N_12651,N_10162,N_10734);
and U12652 (N_12652,N_11253,N_10825);
and U12653 (N_12653,N_11217,N_11896);
and U12654 (N_12654,N_10482,N_10078);
xor U12655 (N_12655,N_10002,N_11536);
xnor U12656 (N_12656,N_10948,N_10386);
nor U12657 (N_12657,N_11848,N_11333);
and U12658 (N_12658,N_10163,N_11563);
xor U12659 (N_12659,N_11532,N_10056);
or U12660 (N_12660,N_11597,N_10904);
nand U12661 (N_12661,N_11772,N_11150);
nand U12662 (N_12662,N_10343,N_11295);
and U12663 (N_12663,N_10946,N_11487);
nor U12664 (N_12664,N_10139,N_11623);
xnor U12665 (N_12665,N_10961,N_10184);
nand U12666 (N_12666,N_10111,N_11568);
nor U12667 (N_12667,N_10471,N_11050);
and U12668 (N_12668,N_10938,N_11211);
nor U12669 (N_12669,N_10900,N_10588);
nor U12670 (N_12670,N_10392,N_10666);
or U12671 (N_12671,N_10107,N_10084);
xor U12672 (N_12672,N_11874,N_10575);
and U12673 (N_12673,N_11178,N_10664);
or U12674 (N_12674,N_11382,N_11163);
nand U12675 (N_12675,N_11719,N_11791);
or U12676 (N_12676,N_11483,N_10321);
or U12677 (N_12677,N_11584,N_10774);
or U12678 (N_12678,N_11913,N_11876);
or U12679 (N_12679,N_10409,N_11144);
nand U12680 (N_12680,N_10811,N_10755);
and U12681 (N_12681,N_10881,N_11789);
xnor U12682 (N_12682,N_10772,N_10326);
nor U12683 (N_12683,N_10705,N_11842);
nand U12684 (N_12684,N_10511,N_11944);
nand U12685 (N_12685,N_11729,N_10898);
or U12686 (N_12686,N_10082,N_11383);
xnor U12687 (N_12687,N_11624,N_11361);
xor U12688 (N_12688,N_11561,N_11482);
xnor U12689 (N_12689,N_11405,N_10018);
nor U12690 (N_12690,N_10680,N_10802);
nand U12691 (N_12691,N_10525,N_10426);
nor U12692 (N_12692,N_10092,N_11824);
nand U12693 (N_12693,N_11748,N_10337);
and U12694 (N_12694,N_11054,N_10190);
nor U12695 (N_12695,N_10368,N_11553);
nand U12696 (N_12696,N_10315,N_11122);
and U12697 (N_12697,N_11577,N_10842);
nand U12698 (N_12698,N_10233,N_10915);
or U12699 (N_12699,N_10356,N_11265);
or U12700 (N_12700,N_11246,N_10075);
nand U12701 (N_12701,N_11804,N_11400);
or U12702 (N_12702,N_10295,N_10043);
and U12703 (N_12703,N_10251,N_11076);
and U12704 (N_12704,N_10165,N_10985);
or U12705 (N_12705,N_11746,N_10464);
nor U12706 (N_12706,N_11218,N_10291);
nand U12707 (N_12707,N_11492,N_10954);
and U12708 (N_12708,N_11990,N_10127);
or U12709 (N_12709,N_10373,N_11428);
and U12710 (N_12710,N_10249,N_11250);
and U12711 (N_12711,N_10235,N_11945);
xor U12712 (N_12712,N_11365,N_10241);
xnor U12713 (N_12713,N_10796,N_10216);
or U12714 (N_12714,N_11722,N_11224);
nor U12715 (N_12715,N_10924,N_10608);
nor U12716 (N_12716,N_10219,N_11818);
nor U12717 (N_12717,N_10370,N_10535);
or U12718 (N_12718,N_10040,N_11733);
or U12719 (N_12719,N_10494,N_11641);
xnor U12720 (N_12720,N_10700,N_11947);
or U12721 (N_12721,N_10697,N_10558);
nand U12722 (N_12722,N_10225,N_11166);
nor U12723 (N_12723,N_10176,N_10532);
or U12724 (N_12724,N_10230,N_10322);
nor U12725 (N_12725,N_10601,N_10150);
xor U12726 (N_12726,N_11919,N_10936);
nor U12727 (N_12727,N_10456,N_11182);
xor U12728 (N_12728,N_11176,N_11590);
xnor U12729 (N_12729,N_11425,N_11258);
nand U12730 (N_12730,N_10736,N_10875);
and U12731 (N_12731,N_10014,N_10671);
and U12732 (N_12732,N_11160,N_11397);
or U12733 (N_12733,N_10415,N_10593);
nand U12734 (N_12734,N_10119,N_10479);
nand U12735 (N_12735,N_11873,N_11664);
and U12736 (N_12736,N_10568,N_11132);
xor U12737 (N_12737,N_11760,N_10005);
nand U12738 (N_12738,N_10498,N_11128);
and U12739 (N_12739,N_10289,N_11888);
xnor U12740 (N_12740,N_11700,N_11283);
xnor U12741 (N_12741,N_11305,N_10140);
and U12742 (N_12742,N_11602,N_11703);
or U12743 (N_12743,N_10742,N_11592);
xnor U12744 (N_12744,N_11506,N_10113);
nor U12745 (N_12745,N_11591,N_11001);
and U12746 (N_12746,N_11030,N_10254);
and U12747 (N_12747,N_10175,N_11617);
nor U12748 (N_12748,N_11909,N_10063);
nor U12749 (N_12749,N_11821,N_10987);
or U12750 (N_12750,N_10803,N_11172);
or U12751 (N_12751,N_10247,N_10807);
or U12752 (N_12752,N_11216,N_10279);
xnor U12753 (N_12753,N_11939,N_10490);
and U12754 (N_12754,N_11029,N_10335);
xor U12755 (N_12755,N_11808,N_11751);
and U12756 (N_12756,N_10301,N_11879);
nand U12757 (N_12757,N_11670,N_10154);
nor U12758 (N_12758,N_11131,N_10160);
nor U12759 (N_12759,N_11851,N_11716);
nor U12760 (N_12760,N_10897,N_11475);
nand U12761 (N_12761,N_10529,N_11406);
xnor U12762 (N_12762,N_10922,N_10333);
nor U12763 (N_12763,N_11560,N_11974);
nor U12764 (N_12764,N_11551,N_10277);
nor U12765 (N_12765,N_10398,N_10632);
nor U12766 (N_12766,N_10662,N_10461);
nor U12767 (N_12767,N_10451,N_11868);
nor U12768 (N_12768,N_10519,N_10761);
nand U12769 (N_12769,N_11464,N_11409);
nor U12770 (N_12770,N_10098,N_11407);
nor U12771 (N_12771,N_11065,N_10971);
nand U12772 (N_12772,N_10366,N_11859);
and U12773 (N_12773,N_10721,N_10095);
or U12774 (N_12774,N_11979,N_10267);
nor U12775 (N_12775,N_10676,N_10982);
and U12776 (N_12776,N_10866,N_11116);
nand U12777 (N_12777,N_11298,N_11940);
or U12778 (N_12778,N_11130,N_10557);
nor U12779 (N_12779,N_11717,N_10817);
and U12780 (N_12780,N_11572,N_11548);
nand U12781 (N_12781,N_10244,N_11457);
or U12782 (N_12782,N_11514,N_11018);
xnor U12783 (N_12783,N_11833,N_10957);
nand U12784 (N_12784,N_11697,N_10416);
or U12785 (N_12785,N_11371,N_10937);
nor U12786 (N_12786,N_10809,N_11618);
nand U12787 (N_12787,N_11448,N_10155);
or U12788 (N_12788,N_10232,N_11202);
or U12789 (N_12789,N_10888,N_11885);
and U12790 (N_12790,N_11302,N_11993);
nor U12791 (N_12791,N_10263,N_10563);
xor U12792 (N_12792,N_11264,N_10997);
or U12793 (N_12793,N_10285,N_11800);
xor U12794 (N_12794,N_11862,N_10319);
nor U12795 (N_12795,N_10638,N_11313);
nand U12796 (N_12796,N_11006,N_10120);
xnor U12797 (N_12797,N_11234,N_10142);
xor U12798 (N_12798,N_11673,N_10678);
and U12799 (N_12799,N_10297,N_11724);
xor U12800 (N_12800,N_11323,N_10612);
and U12801 (N_12801,N_10565,N_10395);
and U12802 (N_12802,N_10976,N_10725);
and U12803 (N_12803,N_10371,N_10487);
nor U12804 (N_12804,N_10248,N_11565);
or U12805 (N_12805,N_11595,N_11378);
or U12806 (N_12806,N_10435,N_11533);
nand U12807 (N_12807,N_11539,N_11663);
nand U12808 (N_12808,N_11685,N_10726);
nor U12809 (N_12809,N_11937,N_11898);
nand U12810 (N_12810,N_10686,N_10492);
nor U12811 (N_12811,N_10513,N_11194);
nor U12812 (N_12812,N_10192,N_11850);
and U12813 (N_12813,N_10798,N_11578);
xnor U12814 (N_12814,N_11095,N_11157);
nor U12815 (N_12815,N_10041,N_11287);
and U12816 (N_12816,N_10979,N_10189);
or U12817 (N_12817,N_10135,N_10499);
nand U12818 (N_12818,N_10125,N_10200);
nor U12819 (N_12819,N_10584,N_11422);
or U12820 (N_12820,N_11327,N_11966);
xnor U12821 (N_12821,N_11185,N_10552);
nor U12822 (N_12822,N_11017,N_10845);
xnor U12823 (N_12823,N_11045,N_11715);
or U12824 (N_12824,N_11255,N_10604);
nand U12825 (N_12825,N_11455,N_10028);
nor U12826 (N_12826,N_10202,N_11756);
or U12827 (N_12827,N_11222,N_10692);
nor U12828 (N_12828,N_10928,N_10776);
nor U12829 (N_12829,N_11607,N_11280);
xnor U12830 (N_12830,N_11867,N_11750);
nand U12831 (N_12831,N_11041,N_11270);
and U12832 (N_12832,N_10878,N_11040);
or U12833 (N_12833,N_11922,N_11675);
nand U12834 (N_12834,N_11794,N_10472);
and U12835 (N_12835,N_11679,N_10167);
or U12836 (N_12836,N_10308,N_10015);
and U12837 (N_12837,N_10679,N_10834);
nand U12838 (N_12838,N_10284,N_11883);
nand U12839 (N_12839,N_10556,N_11494);
and U12840 (N_12840,N_10958,N_11490);
xor U12841 (N_12841,N_10459,N_10034);
or U12842 (N_12842,N_10483,N_11245);
and U12843 (N_12843,N_10011,N_11386);
nand U12844 (N_12844,N_10815,N_10560);
and U12845 (N_12845,N_10868,N_10227);
nor U12846 (N_12846,N_11340,N_11398);
nor U12847 (N_12847,N_10496,N_10214);
nor U12848 (N_12848,N_11996,N_11070);
xor U12849 (N_12849,N_10672,N_10969);
or U12850 (N_12850,N_10037,N_10412);
and U12851 (N_12851,N_11684,N_10213);
xor U12852 (N_12852,N_11098,N_11385);
or U12853 (N_12853,N_11233,N_11953);
nor U12854 (N_12854,N_10438,N_10418);
nor U12855 (N_12855,N_10980,N_10945);
nor U12856 (N_12856,N_10843,N_11016);
and U12857 (N_12857,N_10374,N_10530);
or U12858 (N_12858,N_10204,N_11183);
nand U12859 (N_12859,N_10995,N_10934);
xnor U12860 (N_12860,N_11946,N_10427);
or U12861 (N_12861,N_11840,N_11299);
or U12862 (N_12862,N_11515,N_10493);
xor U12863 (N_12863,N_10923,N_10049);
nand U12864 (N_12864,N_11356,N_11432);
and U12865 (N_12865,N_10148,N_10977);
nor U12866 (N_12866,N_11927,N_11053);
nand U12867 (N_12867,N_10691,N_10480);
and U12868 (N_12868,N_10539,N_10613);
or U12869 (N_12869,N_11399,N_10956);
or U12870 (N_12870,N_11813,N_10170);
or U12871 (N_12871,N_11380,N_11489);
xnor U12872 (N_12872,N_11416,N_10641);
nand U12873 (N_12873,N_10197,N_11140);
nand U12874 (N_12874,N_11304,N_10677);
and U12875 (N_12875,N_10182,N_11588);
xnor U12876 (N_12876,N_10420,N_10069);
nand U12877 (N_12877,N_10156,N_10729);
nor U12878 (N_12878,N_10081,N_10460);
or U12879 (N_12879,N_11089,N_10838);
nand U12880 (N_12880,N_11802,N_11798);
xnor U12881 (N_12881,N_11742,N_11930);
or U12882 (N_12882,N_10933,N_10972);
and U12883 (N_12883,N_10814,N_10136);
and U12884 (N_12884,N_10309,N_11060);
and U12885 (N_12885,N_11374,N_10615);
nor U12886 (N_12886,N_11856,N_11628);
nand U12887 (N_12887,N_11827,N_10681);
xnor U12888 (N_12888,N_10044,N_10877);
and U12889 (N_12889,N_11013,N_11468);
and U12890 (N_12890,N_11387,N_11544);
nor U12891 (N_12891,N_11212,N_10902);
nor U12892 (N_12892,N_10086,N_11556);
xor U12893 (N_12893,N_11635,N_11460);
and U12894 (N_12894,N_10436,N_11701);
and U12895 (N_12895,N_10348,N_11085);
nand U12896 (N_12896,N_11811,N_11923);
xnor U12897 (N_12897,N_10694,N_11728);
xnor U12898 (N_12898,N_10253,N_10046);
nand U12899 (N_12899,N_10569,N_11169);
xnor U12900 (N_12900,N_10674,N_11121);
nand U12901 (N_12901,N_11254,N_11504);
nor U12902 (N_12902,N_11292,N_10272);
nand U12903 (N_12903,N_11026,N_11860);
and U12904 (N_12904,N_11786,N_10829);
xor U12905 (N_12905,N_10720,N_10030);
nand U12906 (N_12906,N_11165,N_11837);
and U12907 (N_12907,N_11726,N_10652);
nand U12908 (N_12908,N_10474,N_10328);
or U12909 (N_12909,N_10410,N_11712);
and U12910 (N_12910,N_10663,N_10351);
nand U12911 (N_12911,N_11418,N_10756);
nand U12912 (N_12912,N_10331,N_10751);
nor U12913 (N_12913,N_10188,N_11702);
nor U12914 (N_12914,N_10887,N_11124);
nand U12915 (N_12915,N_10719,N_11127);
xor U12916 (N_12916,N_10088,N_10212);
xor U12917 (N_12917,N_11134,N_11809);
and U12918 (N_12918,N_10278,N_10896);
and U12919 (N_12919,N_11068,N_11738);
nand U12920 (N_12920,N_10341,N_11499);
and U12921 (N_12921,N_10773,N_11540);
xor U12922 (N_12922,N_10407,N_11901);
nand U12923 (N_12923,N_10816,N_10134);
or U12924 (N_12924,N_11410,N_11643);
nand U12925 (N_12925,N_10031,N_10668);
xor U12926 (N_12926,N_10550,N_10062);
and U12927 (N_12927,N_11206,N_11094);
and U12928 (N_12928,N_10102,N_11740);
and U12929 (N_12929,N_10173,N_10944);
xor U12930 (N_12930,N_10103,N_11331);
and U12931 (N_12931,N_11574,N_11897);
nor U12932 (N_12932,N_10094,N_10649);
xnor U12933 (N_12933,N_10682,N_11997);
and U12934 (N_12934,N_10516,N_10457);
or U12935 (N_12935,N_11650,N_10287);
xnor U12936 (N_12936,N_11105,N_10858);
nand U12937 (N_12937,N_10422,N_10003);
xor U12938 (N_12938,N_11256,N_10446);
and U12939 (N_12939,N_10872,N_10045);
nor U12940 (N_12940,N_11263,N_10032);
nand U12941 (N_12941,N_10894,N_10205);
xor U12942 (N_12942,N_11138,N_11869);
xnor U12943 (N_12943,N_10314,N_10307);
xor U12944 (N_12944,N_11895,N_11807);
nor U12945 (N_12945,N_11317,N_11585);
or U12946 (N_12946,N_10347,N_11503);
nor U12947 (N_12947,N_10159,N_11438);
or U12948 (N_12948,N_10364,N_11301);
nor U12949 (N_12949,N_10554,N_11531);
and U12950 (N_12950,N_10745,N_11389);
xor U12951 (N_12951,N_11345,N_10837);
and U12952 (N_12952,N_10133,N_11633);
xnor U12953 (N_12953,N_10352,N_10361);
xor U12954 (N_12954,N_11754,N_10266);
or U12955 (N_12955,N_10305,N_10234);
nand U12956 (N_12956,N_11109,N_10431);
or U12957 (N_12957,N_10764,N_11857);
or U12958 (N_12958,N_10394,N_10400);
nand U12959 (N_12959,N_10262,N_11710);
and U12960 (N_12960,N_10064,N_10883);
or U12961 (N_12961,N_11682,N_10293);
or U12962 (N_12962,N_11778,N_10491);
or U12963 (N_12963,N_11100,N_10706);
and U12964 (N_12964,N_10239,N_11346);
nand U12965 (N_12965,N_10109,N_10717);
nor U12966 (N_12966,N_10826,N_10458);
nand U12967 (N_12967,N_11960,N_11666);
nand U12968 (N_12968,N_10517,N_11549);
and U12969 (N_12969,N_11690,N_10602);
and U12970 (N_12970,N_10942,N_10178);
nor U12971 (N_12971,N_10131,N_11309);
or U12972 (N_12972,N_11102,N_10504);
nor U12973 (N_12973,N_11672,N_11903);
xnor U12974 (N_12974,N_11863,N_11090);
nor U12975 (N_12975,N_11440,N_11451);
xnor U12976 (N_12976,N_11970,N_11349);
nand U12977 (N_12977,N_11962,N_11010);
nand U12978 (N_12978,N_11339,N_11981);
xnor U12979 (N_12979,N_11067,N_11767);
or U12980 (N_12980,N_10684,N_10236);
and U12981 (N_12981,N_10404,N_11271);
and U12982 (N_12982,N_10354,N_11814);
xor U12983 (N_12983,N_10220,N_11408);
or U12984 (N_12984,N_10071,N_10199);
xor U12985 (N_12985,N_11004,N_11314);
nor U12986 (N_12986,N_10966,N_10853);
nor U12987 (N_12987,N_11886,N_11066);
nor U12988 (N_12988,N_10583,N_11028);
xor U12989 (N_12989,N_11195,N_10383);
or U12990 (N_12990,N_11439,N_11437);
xor U12991 (N_12991,N_11892,N_11870);
and U12992 (N_12992,N_10324,N_10792);
xor U12993 (N_12993,N_11546,N_11855);
or U12994 (N_12994,N_10544,N_11972);
and U12995 (N_12995,N_11614,N_10323);
nor U12996 (N_12996,N_10627,N_10521);
nand U12997 (N_12997,N_11571,N_10712);
xor U12998 (N_12998,N_10222,N_11003);
xor U12999 (N_12999,N_11866,N_11983);
and U13000 (N_13000,N_10826,N_11903);
xnor U13001 (N_13001,N_10822,N_10760);
and U13002 (N_13002,N_10652,N_11995);
nand U13003 (N_13003,N_11336,N_11654);
xnor U13004 (N_13004,N_11211,N_11038);
or U13005 (N_13005,N_11047,N_10353);
and U13006 (N_13006,N_11043,N_11880);
xnor U13007 (N_13007,N_11212,N_10848);
nor U13008 (N_13008,N_10648,N_10848);
xor U13009 (N_13009,N_10400,N_11095);
xor U13010 (N_13010,N_11181,N_10800);
or U13011 (N_13011,N_10552,N_11484);
or U13012 (N_13012,N_10724,N_10728);
and U13013 (N_13013,N_11423,N_11279);
or U13014 (N_13014,N_11980,N_10301);
nor U13015 (N_13015,N_11500,N_10314);
nand U13016 (N_13016,N_11670,N_11068);
xor U13017 (N_13017,N_10836,N_11618);
and U13018 (N_13018,N_10112,N_10808);
or U13019 (N_13019,N_10404,N_10556);
xor U13020 (N_13020,N_11874,N_11622);
and U13021 (N_13021,N_10367,N_10171);
nor U13022 (N_13022,N_11239,N_10207);
nor U13023 (N_13023,N_10515,N_10932);
nor U13024 (N_13024,N_11570,N_11910);
and U13025 (N_13025,N_10106,N_11514);
or U13026 (N_13026,N_10338,N_10815);
nor U13027 (N_13027,N_11035,N_11205);
and U13028 (N_13028,N_10614,N_11981);
or U13029 (N_13029,N_10169,N_10046);
or U13030 (N_13030,N_10102,N_10929);
or U13031 (N_13031,N_11415,N_11273);
and U13032 (N_13032,N_11529,N_10844);
or U13033 (N_13033,N_10770,N_10699);
nor U13034 (N_13034,N_11982,N_10936);
or U13035 (N_13035,N_11783,N_11987);
xnor U13036 (N_13036,N_10309,N_11517);
xnor U13037 (N_13037,N_11495,N_10724);
and U13038 (N_13038,N_10063,N_10263);
nand U13039 (N_13039,N_11765,N_11270);
nor U13040 (N_13040,N_10243,N_11868);
nand U13041 (N_13041,N_10992,N_10506);
nor U13042 (N_13042,N_11967,N_11022);
nor U13043 (N_13043,N_11884,N_11355);
xor U13044 (N_13044,N_10617,N_11538);
xor U13045 (N_13045,N_10459,N_11890);
xor U13046 (N_13046,N_10835,N_11746);
xnor U13047 (N_13047,N_11540,N_11249);
nor U13048 (N_13048,N_10742,N_11734);
xor U13049 (N_13049,N_11519,N_11491);
and U13050 (N_13050,N_10069,N_11989);
or U13051 (N_13051,N_11623,N_11021);
and U13052 (N_13052,N_10538,N_10492);
or U13053 (N_13053,N_10966,N_10528);
nor U13054 (N_13054,N_10803,N_10659);
and U13055 (N_13055,N_11980,N_11633);
nor U13056 (N_13056,N_11618,N_11319);
nand U13057 (N_13057,N_10646,N_10556);
xnor U13058 (N_13058,N_11254,N_11259);
nor U13059 (N_13059,N_11642,N_10392);
nor U13060 (N_13060,N_10639,N_10551);
or U13061 (N_13061,N_11307,N_10175);
nor U13062 (N_13062,N_11956,N_10714);
nand U13063 (N_13063,N_11027,N_11669);
nand U13064 (N_13064,N_11824,N_11171);
nand U13065 (N_13065,N_10169,N_11183);
nand U13066 (N_13066,N_10277,N_10542);
nor U13067 (N_13067,N_10496,N_10959);
nand U13068 (N_13068,N_10432,N_10313);
and U13069 (N_13069,N_11505,N_10800);
or U13070 (N_13070,N_11073,N_10202);
nand U13071 (N_13071,N_11031,N_10654);
nor U13072 (N_13072,N_11339,N_11737);
xor U13073 (N_13073,N_11455,N_11257);
and U13074 (N_13074,N_10407,N_11383);
xor U13075 (N_13075,N_10167,N_11345);
or U13076 (N_13076,N_11754,N_10861);
xor U13077 (N_13077,N_11984,N_11956);
and U13078 (N_13078,N_10742,N_11156);
and U13079 (N_13079,N_10147,N_11170);
or U13080 (N_13080,N_10663,N_11405);
and U13081 (N_13081,N_10222,N_11939);
nand U13082 (N_13082,N_11240,N_11619);
xor U13083 (N_13083,N_11273,N_11777);
nand U13084 (N_13084,N_11021,N_10780);
xor U13085 (N_13085,N_10149,N_11363);
nor U13086 (N_13086,N_10784,N_10151);
and U13087 (N_13087,N_11147,N_10624);
or U13088 (N_13088,N_10569,N_11226);
xor U13089 (N_13089,N_10856,N_11100);
xor U13090 (N_13090,N_10015,N_10593);
xor U13091 (N_13091,N_11804,N_10379);
nand U13092 (N_13092,N_11393,N_10401);
xnor U13093 (N_13093,N_11312,N_10782);
nand U13094 (N_13094,N_10609,N_10319);
nand U13095 (N_13095,N_10834,N_11333);
nand U13096 (N_13096,N_10654,N_10666);
and U13097 (N_13097,N_11501,N_11499);
nand U13098 (N_13098,N_10819,N_10437);
and U13099 (N_13099,N_11107,N_11117);
nand U13100 (N_13100,N_10499,N_11895);
nor U13101 (N_13101,N_11161,N_11009);
nand U13102 (N_13102,N_11021,N_10989);
nor U13103 (N_13103,N_11571,N_10811);
nand U13104 (N_13104,N_10022,N_10568);
or U13105 (N_13105,N_11250,N_10146);
xor U13106 (N_13106,N_11955,N_10123);
and U13107 (N_13107,N_10660,N_11288);
nand U13108 (N_13108,N_10487,N_10812);
nand U13109 (N_13109,N_11511,N_11524);
xnor U13110 (N_13110,N_10635,N_11060);
xor U13111 (N_13111,N_10059,N_10631);
nor U13112 (N_13112,N_11590,N_10115);
and U13113 (N_13113,N_10087,N_10257);
xor U13114 (N_13114,N_11235,N_11225);
xnor U13115 (N_13115,N_11069,N_10411);
and U13116 (N_13116,N_11067,N_10562);
or U13117 (N_13117,N_10906,N_10004);
or U13118 (N_13118,N_10770,N_10165);
and U13119 (N_13119,N_10935,N_10083);
and U13120 (N_13120,N_11519,N_11200);
or U13121 (N_13121,N_11662,N_10018);
xor U13122 (N_13122,N_10612,N_10053);
and U13123 (N_13123,N_11564,N_10970);
xnor U13124 (N_13124,N_11485,N_10081);
nor U13125 (N_13125,N_10428,N_10255);
or U13126 (N_13126,N_11842,N_10217);
and U13127 (N_13127,N_11101,N_10593);
or U13128 (N_13128,N_11185,N_11593);
xnor U13129 (N_13129,N_10407,N_10869);
nor U13130 (N_13130,N_11473,N_10267);
nor U13131 (N_13131,N_10431,N_10759);
nor U13132 (N_13132,N_10551,N_10972);
or U13133 (N_13133,N_10115,N_11505);
nor U13134 (N_13134,N_10848,N_11062);
nor U13135 (N_13135,N_10246,N_10464);
or U13136 (N_13136,N_10930,N_11037);
nand U13137 (N_13137,N_11485,N_11943);
nand U13138 (N_13138,N_10296,N_10819);
and U13139 (N_13139,N_10580,N_10836);
and U13140 (N_13140,N_10313,N_11820);
nand U13141 (N_13141,N_11865,N_11035);
nor U13142 (N_13142,N_11032,N_11553);
xnor U13143 (N_13143,N_10420,N_11563);
nand U13144 (N_13144,N_11699,N_11619);
and U13145 (N_13145,N_10663,N_11593);
nand U13146 (N_13146,N_10143,N_10489);
or U13147 (N_13147,N_11993,N_10844);
nand U13148 (N_13148,N_10379,N_10000);
nor U13149 (N_13149,N_10564,N_10121);
or U13150 (N_13150,N_10299,N_11323);
and U13151 (N_13151,N_11633,N_11816);
xnor U13152 (N_13152,N_11407,N_11679);
nand U13153 (N_13153,N_10659,N_11828);
xnor U13154 (N_13154,N_11113,N_10647);
nor U13155 (N_13155,N_11101,N_11503);
xnor U13156 (N_13156,N_10580,N_10005);
xnor U13157 (N_13157,N_10523,N_11229);
or U13158 (N_13158,N_10426,N_10129);
xnor U13159 (N_13159,N_10714,N_10932);
or U13160 (N_13160,N_10644,N_10586);
and U13161 (N_13161,N_11794,N_10350);
or U13162 (N_13162,N_10019,N_10791);
xor U13163 (N_13163,N_10054,N_10770);
nor U13164 (N_13164,N_10127,N_11225);
and U13165 (N_13165,N_10961,N_11191);
nor U13166 (N_13166,N_11538,N_11649);
and U13167 (N_13167,N_11978,N_10062);
nand U13168 (N_13168,N_11871,N_10132);
nand U13169 (N_13169,N_11662,N_10215);
or U13170 (N_13170,N_11872,N_10883);
nor U13171 (N_13171,N_10340,N_10860);
nor U13172 (N_13172,N_10127,N_11824);
or U13173 (N_13173,N_11406,N_11412);
nor U13174 (N_13174,N_11721,N_10877);
xor U13175 (N_13175,N_10517,N_11662);
xor U13176 (N_13176,N_10416,N_11182);
nor U13177 (N_13177,N_11360,N_11076);
or U13178 (N_13178,N_10171,N_11530);
xnor U13179 (N_13179,N_10955,N_11043);
xnor U13180 (N_13180,N_10468,N_11504);
nand U13181 (N_13181,N_10610,N_10637);
nor U13182 (N_13182,N_11494,N_11748);
xor U13183 (N_13183,N_10386,N_11168);
nand U13184 (N_13184,N_11246,N_10461);
and U13185 (N_13185,N_11431,N_11026);
or U13186 (N_13186,N_10479,N_11988);
and U13187 (N_13187,N_11958,N_10942);
and U13188 (N_13188,N_10041,N_10036);
nand U13189 (N_13189,N_10588,N_10337);
nand U13190 (N_13190,N_11748,N_10639);
and U13191 (N_13191,N_10250,N_11890);
xnor U13192 (N_13192,N_10785,N_11847);
or U13193 (N_13193,N_11841,N_11298);
or U13194 (N_13194,N_11887,N_11744);
nor U13195 (N_13195,N_11743,N_11132);
and U13196 (N_13196,N_10517,N_10977);
nand U13197 (N_13197,N_10394,N_10815);
xnor U13198 (N_13198,N_11846,N_11056);
nor U13199 (N_13199,N_11801,N_11312);
or U13200 (N_13200,N_11525,N_11456);
or U13201 (N_13201,N_10955,N_10136);
or U13202 (N_13202,N_10668,N_11484);
or U13203 (N_13203,N_11294,N_11099);
nand U13204 (N_13204,N_10512,N_10019);
nor U13205 (N_13205,N_10988,N_11446);
xor U13206 (N_13206,N_10446,N_10462);
nor U13207 (N_13207,N_10793,N_11653);
or U13208 (N_13208,N_10120,N_10346);
nand U13209 (N_13209,N_11035,N_11860);
xor U13210 (N_13210,N_11755,N_11884);
xor U13211 (N_13211,N_10063,N_10183);
nor U13212 (N_13212,N_10493,N_11522);
and U13213 (N_13213,N_11615,N_11543);
or U13214 (N_13214,N_10356,N_11211);
or U13215 (N_13215,N_10455,N_10715);
xnor U13216 (N_13216,N_11394,N_10422);
nand U13217 (N_13217,N_11692,N_11888);
and U13218 (N_13218,N_10645,N_10002);
and U13219 (N_13219,N_10574,N_10655);
nor U13220 (N_13220,N_10213,N_10411);
xor U13221 (N_13221,N_10147,N_11463);
nand U13222 (N_13222,N_11916,N_10309);
or U13223 (N_13223,N_10383,N_10784);
nor U13224 (N_13224,N_10727,N_10038);
xor U13225 (N_13225,N_10048,N_11596);
nand U13226 (N_13226,N_11409,N_11093);
xnor U13227 (N_13227,N_11345,N_11677);
nand U13228 (N_13228,N_11072,N_11530);
nand U13229 (N_13229,N_11190,N_10656);
nor U13230 (N_13230,N_11134,N_10386);
and U13231 (N_13231,N_11626,N_10061);
xnor U13232 (N_13232,N_10472,N_11156);
nor U13233 (N_13233,N_11295,N_10737);
nand U13234 (N_13234,N_11585,N_10292);
nand U13235 (N_13235,N_11535,N_10991);
or U13236 (N_13236,N_11291,N_10569);
xor U13237 (N_13237,N_10362,N_10007);
xor U13238 (N_13238,N_10339,N_10561);
nor U13239 (N_13239,N_10749,N_11298);
xnor U13240 (N_13240,N_10223,N_10778);
xor U13241 (N_13241,N_10065,N_10646);
and U13242 (N_13242,N_11112,N_11990);
and U13243 (N_13243,N_11859,N_11187);
nor U13244 (N_13244,N_11470,N_10232);
xor U13245 (N_13245,N_11234,N_11726);
nand U13246 (N_13246,N_10430,N_11889);
nand U13247 (N_13247,N_11384,N_10119);
and U13248 (N_13248,N_10301,N_11041);
nor U13249 (N_13249,N_10875,N_11886);
and U13250 (N_13250,N_11942,N_11541);
xor U13251 (N_13251,N_10670,N_10049);
and U13252 (N_13252,N_10540,N_11672);
xor U13253 (N_13253,N_10358,N_11094);
xor U13254 (N_13254,N_10894,N_11410);
or U13255 (N_13255,N_11121,N_10159);
or U13256 (N_13256,N_11961,N_10774);
xor U13257 (N_13257,N_11708,N_10416);
xnor U13258 (N_13258,N_11073,N_11207);
nand U13259 (N_13259,N_10990,N_10579);
nand U13260 (N_13260,N_10710,N_10911);
xnor U13261 (N_13261,N_10403,N_11457);
xnor U13262 (N_13262,N_11852,N_11277);
xnor U13263 (N_13263,N_11847,N_10692);
and U13264 (N_13264,N_10340,N_11936);
and U13265 (N_13265,N_10073,N_10254);
or U13266 (N_13266,N_11480,N_10274);
nand U13267 (N_13267,N_11914,N_11968);
and U13268 (N_13268,N_10604,N_10160);
or U13269 (N_13269,N_11390,N_10162);
or U13270 (N_13270,N_11597,N_11068);
nand U13271 (N_13271,N_10608,N_11564);
and U13272 (N_13272,N_11412,N_11183);
nand U13273 (N_13273,N_11940,N_11117);
nand U13274 (N_13274,N_11988,N_10928);
and U13275 (N_13275,N_10912,N_11215);
nor U13276 (N_13276,N_11120,N_11134);
nand U13277 (N_13277,N_10407,N_11501);
nand U13278 (N_13278,N_11715,N_10789);
xnor U13279 (N_13279,N_10096,N_10572);
xor U13280 (N_13280,N_10731,N_11480);
xnor U13281 (N_13281,N_10893,N_11857);
and U13282 (N_13282,N_11378,N_11353);
nor U13283 (N_13283,N_10402,N_10939);
or U13284 (N_13284,N_10164,N_11556);
xnor U13285 (N_13285,N_11000,N_10508);
and U13286 (N_13286,N_10283,N_11366);
or U13287 (N_13287,N_10157,N_11949);
or U13288 (N_13288,N_11293,N_11125);
nand U13289 (N_13289,N_10230,N_11732);
or U13290 (N_13290,N_10724,N_10312);
or U13291 (N_13291,N_11504,N_11270);
or U13292 (N_13292,N_11005,N_11817);
nor U13293 (N_13293,N_10173,N_11570);
nor U13294 (N_13294,N_11615,N_10896);
xor U13295 (N_13295,N_11911,N_10602);
nand U13296 (N_13296,N_11003,N_10488);
or U13297 (N_13297,N_11255,N_11048);
or U13298 (N_13298,N_11664,N_11584);
and U13299 (N_13299,N_10261,N_11366);
nor U13300 (N_13300,N_11813,N_11147);
or U13301 (N_13301,N_11705,N_11979);
or U13302 (N_13302,N_10365,N_10307);
or U13303 (N_13303,N_11942,N_11831);
or U13304 (N_13304,N_11642,N_10102);
nand U13305 (N_13305,N_11242,N_11266);
and U13306 (N_13306,N_11094,N_11181);
xnor U13307 (N_13307,N_10233,N_10903);
xor U13308 (N_13308,N_11205,N_11862);
or U13309 (N_13309,N_10750,N_11938);
xor U13310 (N_13310,N_10808,N_10827);
or U13311 (N_13311,N_11812,N_10041);
or U13312 (N_13312,N_11843,N_10635);
nand U13313 (N_13313,N_11285,N_11226);
or U13314 (N_13314,N_10726,N_10750);
nor U13315 (N_13315,N_11472,N_11835);
xnor U13316 (N_13316,N_10069,N_11246);
or U13317 (N_13317,N_10207,N_11973);
nor U13318 (N_13318,N_11036,N_11378);
and U13319 (N_13319,N_11459,N_11852);
xnor U13320 (N_13320,N_11636,N_11310);
or U13321 (N_13321,N_10882,N_10016);
and U13322 (N_13322,N_11599,N_10943);
nor U13323 (N_13323,N_10573,N_11758);
nand U13324 (N_13324,N_10319,N_10713);
nand U13325 (N_13325,N_11110,N_10885);
nor U13326 (N_13326,N_10408,N_10290);
nand U13327 (N_13327,N_11767,N_10294);
xnor U13328 (N_13328,N_10628,N_10763);
or U13329 (N_13329,N_10735,N_11504);
nor U13330 (N_13330,N_11279,N_10678);
and U13331 (N_13331,N_10920,N_11452);
nor U13332 (N_13332,N_10813,N_10514);
or U13333 (N_13333,N_10417,N_10278);
xnor U13334 (N_13334,N_11127,N_10794);
xnor U13335 (N_13335,N_11023,N_10630);
xor U13336 (N_13336,N_10642,N_10787);
xor U13337 (N_13337,N_11712,N_10627);
nand U13338 (N_13338,N_11526,N_11473);
xor U13339 (N_13339,N_10100,N_11523);
or U13340 (N_13340,N_11967,N_10007);
nand U13341 (N_13341,N_10597,N_11230);
or U13342 (N_13342,N_10307,N_10851);
or U13343 (N_13343,N_10153,N_10878);
or U13344 (N_13344,N_11076,N_11839);
and U13345 (N_13345,N_11920,N_11967);
and U13346 (N_13346,N_11395,N_10503);
xor U13347 (N_13347,N_10097,N_10661);
nor U13348 (N_13348,N_10201,N_11074);
and U13349 (N_13349,N_11206,N_10778);
and U13350 (N_13350,N_11279,N_11164);
or U13351 (N_13351,N_10557,N_10371);
or U13352 (N_13352,N_11680,N_10283);
nand U13353 (N_13353,N_11986,N_11905);
nand U13354 (N_13354,N_10880,N_11935);
xnor U13355 (N_13355,N_10659,N_10459);
and U13356 (N_13356,N_11819,N_11143);
and U13357 (N_13357,N_10895,N_10162);
nor U13358 (N_13358,N_11024,N_11832);
and U13359 (N_13359,N_11339,N_10357);
nand U13360 (N_13360,N_10994,N_11422);
nor U13361 (N_13361,N_10440,N_11111);
or U13362 (N_13362,N_10891,N_10872);
nand U13363 (N_13363,N_11235,N_11142);
nor U13364 (N_13364,N_11788,N_11036);
or U13365 (N_13365,N_10201,N_10280);
nor U13366 (N_13366,N_10808,N_10332);
xnor U13367 (N_13367,N_10631,N_11523);
nand U13368 (N_13368,N_10229,N_11948);
or U13369 (N_13369,N_11940,N_11414);
xnor U13370 (N_13370,N_10867,N_10822);
or U13371 (N_13371,N_10550,N_11589);
xor U13372 (N_13372,N_11744,N_11875);
or U13373 (N_13373,N_11548,N_10664);
nand U13374 (N_13374,N_11817,N_10586);
and U13375 (N_13375,N_10215,N_11044);
nand U13376 (N_13376,N_10054,N_11543);
and U13377 (N_13377,N_11762,N_11402);
or U13378 (N_13378,N_11878,N_11149);
or U13379 (N_13379,N_10372,N_10873);
or U13380 (N_13380,N_11279,N_11306);
nor U13381 (N_13381,N_11235,N_11285);
and U13382 (N_13382,N_10913,N_10170);
xor U13383 (N_13383,N_11327,N_10884);
xnor U13384 (N_13384,N_11286,N_11437);
xnor U13385 (N_13385,N_10193,N_10414);
nand U13386 (N_13386,N_11283,N_10095);
and U13387 (N_13387,N_11971,N_10154);
nor U13388 (N_13388,N_10584,N_11461);
nand U13389 (N_13389,N_10139,N_11200);
nor U13390 (N_13390,N_11254,N_11220);
or U13391 (N_13391,N_11096,N_11314);
or U13392 (N_13392,N_11600,N_11140);
nand U13393 (N_13393,N_11852,N_11047);
xor U13394 (N_13394,N_11477,N_11074);
and U13395 (N_13395,N_11985,N_11957);
and U13396 (N_13396,N_11932,N_10915);
nand U13397 (N_13397,N_11288,N_10605);
nand U13398 (N_13398,N_11382,N_11584);
nand U13399 (N_13399,N_10473,N_10963);
or U13400 (N_13400,N_10453,N_10188);
or U13401 (N_13401,N_10926,N_10462);
xor U13402 (N_13402,N_11286,N_10326);
xnor U13403 (N_13403,N_11034,N_11254);
nand U13404 (N_13404,N_10619,N_11460);
nor U13405 (N_13405,N_11889,N_11009);
or U13406 (N_13406,N_10426,N_11806);
nand U13407 (N_13407,N_11830,N_11135);
nor U13408 (N_13408,N_11389,N_11073);
nor U13409 (N_13409,N_10270,N_10784);
nand U13410 (N_13410,N_11456,N_10027);
xnor U13411 (N_13411,N_10258,N_10715);
nand U13412 (N_13412,N_11126,N_11426);
and U13413 (N_13413,N_10142,N_10319);
xnor U13414 (N_13414,N_10401,N_10149);
xor U13415 (N_13415,N_10628,N_11844);
or U13416 (N_13416,N_11398,N_11169);
and U13417 (N_13417,N_10139,N_10001);
nand U13418 (N_13418,N_10444,N_11548);
or U13419 (N_13419,N_11188,N_10908);
or U13420 (N_13420,N_11763,N_11037);
nand U13421 (N_13421,N_10382,N_11902);
and U13422 (N_13422,N_10564,N_10956);
or U13423 (N_13423,N_10399,N_11177);
and U13424 (N_13424,N_11499,N_10889);
xnor U13425 (N_13425,N_11068,N_10508);
or U13426 (N_13426,N_10608,N_11332);
or U13427 (N_13427,N_11511,N_10858);
nand U13428 (N_13428,N_11340,N_10294);
or U13429 (N_13429,N_10401,N_10845);
nand U13430 (N_13430,N_11010,N_11591);
and U13431 (N_13431,N_11586,N_10125);
and U13432 (N_13432,N_11005,N_10641);
xnor U13433 (N_13433,N_10530,N_11798);
and U13434 (N_13434,N_10100,N_11676);
nand U13435 (N_13435,N_11401,N_11247);
nor U13436 (N_13436,N_10341,N_11862);
and U13437 (N_13437,N_11440,N_10608);
nand U13438 (N_13438,N_10220,N_11903);
xnor U13439 (N_13439,N_10478,N_11895);
nor U13440 (N_13440,N_10336,N_10691);
and U13441 (N_13441,N_11834,N_10881);
nor U13442 (N_13442,N_11633,N_11004);
and U13443 (N_13443,N_10139,N_11721);
xnor U13444 (N_13444,N_11104,N_10993);
nor U13445 (N_13445,N_11071,N_10748);
nand U13446 (N_13446,N_11729,N_11275);
or U13447 (N_13447,N_10438,N_10160);
nand U13448 (N_13448,N_11949,N_11550);
xnor U13449 (N_13449,N_11100,N_11610);
or U13450 (N_13450,N_11909,N_10396);
nor U13451 (N_13451,N_10636,N_11182);
nor U13452 (N_13452,N_11935,N_10689);
or U13453 (N_13453,N_11800,N_10493);
nor U13454 (N_13454,N_10403,N_10316);
nor U13455 (N_13455,N_11324,N_10788);
or U13456 (N_13456,N_10450,N_10989);
or U13457 (N_13457,N_11368,N_10399);
xnor U13458 (N_13458,N_11756,N_10465);
or U13459 (N_13459,N_11898,N_10968);
nand U13460 (N_13460,N_10468,N_10562);
xnor U13461 (N_13461,N_10862,N_10734);
nand U13462 (N_13462,N_10518,N_11966);
xnor U13463 (N_13463,N_10720,N_10593);
xnor U13464 (N_13464,N_11576,N_11881);
or U13465 (N_13465,N_10360,N_10228);
nand U13466 (N_13466,N_11475,N_10289);
nand U13467 (N_13467,N_11218,N_10979);
nand U13468 (N_13468,N_11657,N_10591);
xor U13469 (N_13469,N_11161,N_10172);
or U13470 (N_13470,N_10402,N_10520);
xnor U13471 (N_13471,N_11688,N_10667);
and U13472 (N_13472,N_11491,N_11673);
xor U13473 (N_13473,N_11705,N_10835);
nor U13474 (N_13474,N_11106,N_11624);
nand U13475 (N_13475,N_10643,N_11708);
or U13476 (N_13476,N_11242,N_10352);
nand U13477 (N_13477,N_11338,N_10147);
xor U13478 (N_13478,N_11615,N_11050);
or U13479 (N_13479,N_11707,N_10521);
xor U13480 (N_13480,N_11221,N_10491);
xor U13481 (N_13481,N_10166,N_11225);
nand U13482 (N_13482,N_11021,N_10263);
nand U13483 (N_13483,N_11436,N_10994);
nand U13484 (N_13484,N_11053,N_11083);
or U13485 (N_13485,N_11701,N_11493);
nand U13486 (N_13486,N_11117,N_11876);
xnor U13487 (N_13487,N_11772,N_10213);
xor U13488 (N_13488,N_10115,N_10617);
and U13489 (N_13489,N_11384,N_11993);
nand U13490 (N_13490,N_11597,N_10946);
xor U13491 (N_13491,N_11058,N_11369);
and U13492 (N_13492,N_11686,N_11543);
and U13493 (N_13493,N_11985,N_10236);
nand U13494 (N_13494,N_10583,N_11564);
nand U13495 (N_13495,N_10822,N_11962);
nand U13496 (N_13496,N_11013,N_10558);
nor U13497 (N_13497,N_11152,N_11038);
nor U13498 (N_13498,N_11939,N_10593);
nor U13499 (N_13499,N_10013,N_10081);
xnor U13500 (N_13500,N_11974,N_10692);
or U13501 (N_13501,N_10999,N_10296);
nor U13502 (N_13502,N_10022,N_10249);
and U13503 (N_13503,N_10385,N_11589);
nand U13504 (N_13504,N_10965,N_10246);
nor U13505 (N_13505,N_11695,N_11206);
xnor U13506 (N_13506,N_11712,N_11017);
nand U13507 (N_13507,N_10664,N_11593);
or U13508 (N_13508,N_10548,N_10846);
nand U13509 (N_13509,N_11342,N_10990);
and U13510 (N_13510,N_11227,N_10770);
or U13511 (N_13511,N_10853,N_11078);
nor U13512 (N_13512,N_10678,N_10770);
xnor U13513 (N_13513,N_10655,N_10507);
xor U13514 (N_13514,N_10991,N_11633);
xnor U13515 (N_13515,N_10126,N_10781);
or U13516 (N_13516,N_10977,N_11331);
and U13517 (N_13517,N_11823,N_11487);
and U13518 (N_13518,N_11366,N_10556);
nor U13519 (N_13519,N_10114,N_10952);
nand U13520 (N_13520,N_10840,N_10682);
and U13521 (N_13521,N_10281,N_10261);
xnor U13522 (N_13522,N_10110,N_11677);
nor U13523 (N_13523,N_11326,N_11185);
and U13524 (N_13524,N_10202,N_10162);
or U13525 (N_13525,N_10592,N_11955);
xnor U13526 (N_13526,N_10330,N_11213);
or U13527 (N_13527,N_11583,N_11311);
nand U13528 (N_13528,N_10205,N_11476);
or U13529 (N_13529,N_11760,N_11120);
or U13530 (N_13530,N_11235,N_11743);
and U13531 (N_13531,N_10089,N_11495);
or U13532 (N_13532,N_10349,N_10245);
xor U13533 (N_13533,N_11594,N_10753);
or U13534 (N_13534,N_11014,N_11683);
and U13535 (N_13535,N_10751,N_10616);
nor U13536 (N_13536,N_10787,N_11386);
and U13537 (N_13537,N_10007,N_11857);
nor U13538 (N_13538,N_10919,N_11693);
nor U13539 (N_13539,N_11188,N_10563);
or U13540 (N_13540,N_10410,N_10186);
nand U13541 (N_13541,N_10894,N_11500);
xor U13542 (N_13542,N_10231,N_10915);
nor U13543 (N_13543,N_11443,N_11695);
and U13544 (N_13544,N_10863,N_11521);
or U13545 (N_13545,N_11316,N_10173);
xor U13546 (N_13546,N_11419,N_11556);
nand U13547 (N_13547,N_11259,N_11471);
or U13548 (N_13548,N_10067,N_10767);
xor U13549 (N_13549,N_11823,N_10015);
and U13550 (N_13550,N_10260,N_11172);
and U13551 (N_13551,N_11498,N_10859);
nor U13552 (N_13552,N_11406,N_10841);
and U13553 (N_13553,N_11726,N_11574);
nand U13554 (N_13554,N_11271,N_11442);
nand U13555 (N_13555,N_11834,N_11548);
and U13556 (N_13556,N_10825,N_10392);
nor U13557 (N_13557,N_10748,N_11669);
and U13558 (N_13558,N_10682,N_11085);
xor U13559 (N_13559,N_11666,N_10659);
and U13560 (N_13560,N_11852,N_11120);
nor U13561 (N_13561,N_11641,N_10427);
or U13562 (N_13562,N_11092,N_11301);
nand U13563 (N_13563,N_10662,N_11311);
and U13564 (N_13564,N_11869,N_10883);
nand U13565 (N_13565,N_10684,N_11401);
or U13566 (N_13566,N_10674,N_10580);
and U13567 (N_13567,N_10172,N_11315);
and U13568 (N_13568,N_10344,N_11336);
nand U13569 (N_13569,N_10950,N_10168);
nor U13570 (N_13570,N_10956,N_10146);
and U13571 (N_13571,N_11895,N_10775);
and U13572 (N_13572,N_10172,N_11411);
xnor U13573 (N_13573,N_10225,N_11046);
nand U13574 (N_13574,N_11140,N_11567);
or U13575 (N_13575,N_11916,N_10956);
or U13576 (N_13576,N_10710,N_10221);
or U13577 (N_13577,N_10451,N_11041);
and U13578 (N_13578,N_11402,N_11875);
nor U13579 (N_13579,N_10572,N_10275);
xnor U13580 (N_13580,N_10686,N_11829);
or U13581 (N_13581,N_11469,N_11188);
xor U13582 (N_13582,N_10697,N_10463);
nand U13583 (N_13583,N_10676,N_10799);
and U13584 (N_13584,N_11685,N_10312);
and U13585 (N_13585,N_10415,N_11277);
or U13586 (N_13586,N_10875,N_11349);
nand U13587 (N_13587,N_11789,N_11355);
nor U13588 (N_13588,N_10357,N_10482);
xnor U13589 (N_13589,N_11764,N_11232);
or U13590 (N_13590,N_11778,N_11046);
nor U13591 (N_13591,N_11119,N_10093);
nand U13592 (N_13592,N_10723,N_10004);
xnor U13593 (N_13593,N_10174,N_10933);
nor U13594 (N_13594,N_10011,N_10182);
nand U13595 (N_13595,N_10786,N_11996);
or U13596 (N_13596,N_11211,N_10622);
or U13597 (N_13597,N_10676,N_10965);
xnor U13598 (N_13598,N_11723,N_10358);
nor U13599 (N_13599,N_10985,N_10642);
nor U13600 (N_13600,N_11127,N_11542);
nand U13601 (N_13601,N_11098,N_11796);
nor U13602 (N_13602,N_10610,N_10314);
nand U13603 (N_13603,N_11545,N_11487);
nor U13604 (N_13604,N_11891,N_11147);
nand U13605 (N_13605,N_11234,N_11917);
nor U13606 (N_13606,N_11059,N_10043);
and U13607 (N_13607,N_11177,N_11443);
or U13608 (N_13608,N_10968,N_11449);
nor U13609 (N_13609,N_11315,N_10000);
or U13610 (N_13610,N_10270,N_11203);
xnor U13611 (N_13611,N_11804,N_11696);
nor U13612 (N_13612,N_11352,N_10774);
nor U13613 (N_13613,N_10856,N_10621);
nand U13614 (N_13614,N_11927,N_10694);
and U13615 (N_13615,N_10442,N_11259);
nor U13616 (N_13616,N_10244,N_11692);
or U13617 (N_13617,N_11428,N_10947);
xnor U13618 (N_13618,N_10390,N_10871);
and U13619 (N_13619,N_10648,N_11551);
nand U13620 (N_13620,N_11682,N_11070);
and U13621 (N_13621,N_10051,N_10916);
nor U13622 (N_13622,N_10757,N_11098);
or U13623 (N_13623,N_10814,N_11495);
and U13624 (N_13624,N_10971,N_11218);
xnor U13625 (N_13625,N_10515,N_11129);
or U13626 (N_13626,N_11615,N_10998);
nand U13627 (N_13627,N_10323,N_11178);
nor U13628 (N_13628,N_11505,N_10348);
nor U13629 (N_13629,N_11912,N_11229);
nor U13630 (N_13630,N_10968,N_10036);
nand U13631 (N_13631,N_10270,N_11750);
or U13632 (N_13632,N_10915,N_11571);
or U13633 (N_13633,N_11244,N_10441);
or U13634 (N_13634,N_10269,N_10004);
and U13635 (N_13635,N_10872,N_11843);
nor U13636 (N_13636,N_10500,N_10414);
xor U13637 (N_13637,N_11779,N_11794);
xnor U13638 (N_13638,N_10622,N_11147);
or U13639 (N_13639,N_11145,N_11005);
and U13640 (N_13640,N_11443,N_10360);
and U13641 (N_13641,N_10943,N_10351);
or U13642 (N_13642,N_10385,N_11607);
nor U13643 (N_13643,N_10799,N_10870);
xnor U13644 (N_13644,N_10210,N_10154);
nor U13645 (N_13645,N_10453,N_11385);
nand U13646 (N_13646,N_11047,N_11698);
xnor U13647 (N_13647,N_11141,N_11720);
and U13648 (N_13648,N_11070,N_11419);
nand U13649 (N_13649,N_11999,N_10909);
nand U13650 (N_13650,N_10435,N_11882);
and U13651 (N_13651,N_10640,N_11227);
or U13652 (N_13652,N_11997,N_11113);
xnor U13653 (N_13653,N_11009,N_10278);
or U13654 (N_13654,N_11718,N_11733);
nor U13655 (N_13655,N_10511,N_10501);
nor U13656 (N_13656,N_10372,N_11367);
and U13657 (N_13657,N_11684,N_10521);
or U13658 (N_13658,N_10993,N_10557);
or U13659 (N_13659,N_11283,N_10372);
and U13660 (N_13660,N_10184,N_10625);
and U13661 (N_13661,N_11734,N_10077);
nor U13662 (N_13662,N_10995,N_11182);
nor U13663 (N_13663,N_10827,N_11216);
and U13664 (N_13664,N_10690,N_10967);
or U13665 (N_13665,N_11593,N_11516);
and U13666 (N_13666,N_10405,N_10306);
xor U13667 (N_13667,N_11432,N_10022);
nor U13668 (N_13668,N_10043,N_10774);
xnor U13669 (N_13669,N_11770,N_11426);
nor U13670 (N_13670,N_10910,N_11397);
nand U13671 (N_13671,N_10682,N_11155);
or U13672 (N_13672,N_10140,N_10427);
nand U13673 (N_13673,N_10651,N_11806);
xnor U13674 (N_13674,N_11943,N_11000);
and U13675 (N_13675,N_11108,N_10443);
and U13676 (N_13676,N_11364,N_10278);
or U13677 (N_13677,N_10957,N_11291);
nor U13678 (N_13678,N_11373,N_11139);
nor U13679 (N_13679,N_11926,N_11343);
nand U13680 (N_13680,N_11922,N_11865);
nor U13681 (N_13681,N_10305,N_10181);
xnor U13682 (N_13682,N_10963,N_10254);
or U13683 (N_13683,N_10281,N_11753);
nand U13684 (N_13684,N_11718,N_11542);
xor U13685 (N_13685,N_10706,N_10322);
and U13686 (N_13686,N_10259,N_10888);
nor U13687 (N_13687,N_11274,N_10421);
or U13688 (N_13688,N_10288,N_10770);
and U13689 (N_13689,N_10803,N_10329);
nand U13690 (N_13690,N_11605,N_11481);
and U13691 (N_13691,N_10363,N_11441);
nor U13692 (N_13692,N_10297,N_10946);
and U13693 (N_13693,N_11797,N_11500);
xor U13694 (N_13694,N_11952,N_11663);
nand U13695 (N_13695,N_11452,N_11068);
and U13696 (N_13696,N_11630,N_11966);
and U13697 (N_13697,N_11852,N_11725);
xnor U13698 (N_13698,N_11802,N_11346);
nor U13699 (N_13699,N_10808,N_11946);
xor U13700 (N_13700,N_11175,N_11332);
nand U13701 (N_13701,N_11703,N_11464);
nand U13702 (N_13702,N_11394,N_10536);
or U13703 (N_13703,N_10590,N_11282);
or U13704 (N_13704,N_10411,N_10811);
nand U13705 (N_13705,N_10116,N_10946);
and U13706 (N_13706,N_10263,N_11919);
or U13707 (N_13707,N_10444,N_11812);
nand U13708 (N_13708,N_11659,N_10645);
nand U13709 (N_13709,N_10238,N_10895);
xor U13710 (N_13710,N_11252,N_11841);
nand U13711 (N_13711,N_11174,N_11910);
and U13712 (N_13712,N_11096,N_10799);
or U13713 (N_13713,N_11546,N_10530);
xor U13714 (N_13714,N_10560,N_10758);
or U13715 (N_13715,N_10163,N_11777);
nand U13716 (N_13716,N_11591,N_11383);
and U13717 (N_13717,N_11338,N_10376);
xor U13718 (N_13718,N_11250,N_10320);
nor U13719 (N_13719,N_11848,N_11057);
and U13720 (N_13720,N_10030,N_11388);
xor U13721 (N_13721,N_10525,N_11879);
or U13722 (N_13722,N_10771,N_11021);
xor U13723 (N_13723,N_10886,N_10829);
nor U13724 (N_13724,N_11412,N_10562);
xor U13725 (N_13725,N_11059,N_10333);
and U13726 (N_13726,N_10648,N_11092);
nand U13727 (N_13727,N_11558,N_11461);
and U13728 (N_13728,N_10793,N_10201);
or U13729 (N_13729,N_10336,N_11192);
nand U13730 (N_13730,N_10555,N_10889);
nor U13731 (N_13731,N_11018,N_11591);
nor U13732 (N_13732,N_10762,N_11177);
nand U13733 (N_13733,N_10126,N_11008);
and U13734 (N_13734,N_10425,N_11433);
or U13735 (N_13735,N_10679,N_11072);
or U13736 (N_13736,N_11809,N_11479);
and U13737 (N_13737,N_10969,N_10885);
and U13738 (N_13738,N_11442,N_11320);
xnor U13739 (N_13739,N_10769,N_11524);
and U13740 (N_13740,N_10100,N_10437);
and U13741 (N_13741,N_10931,N_11451);
nand U13742 (N_13742,N_10403,N_11912);
and U13743 (N_13743,N_10873,N_11447);
or U13744 (N_13744,N_10901,N_11539);
nand U13745 (N_13745,N_10471,N_11493);
or U13746 (N_13746,N_10888,N_11755);
and U13747 (N_13747,N_11626,N_11042);
nor U13748 (N_13748,N_11368,N_11671);
nor U13749 (N_13749,N_10052,N_11511);
nor U13750 (N_13750,N_10829,N_11718);
and U13751 (N_13751,N_11125,N_10624);
and U13752 (N_13752,N_10562,N_10273);
xnor U13753 (N_13753,N_10496,N_11614);
nor U13754 (N_13754,N_11828,N_10804);
nor U13755 (N_13755,N_10101,N_10004);
nand U13756 (N_13756,N_11184,N_10539);
or U13757 (N_13757,N_11445,N_11838);
nor U13758 (N_13758,N_11290,N_11126);
nand U13759 (N_13759,N_10411,N_10055);
nor U13760 (N_13760,N_10769,N_10580);
xor U13761 (N_13761,N_11924,N_10530);
or U13762 (N_13762,N_11784,N_11273);
nor U13763 (N_13763,N_10242,N_10114);
nor U13764 (N_13764,N_11487,N_11747);
and U13765 (N_13765,N_11883,N_10613);
nor U13766 (N_13766,N_11482,N_11039);
or U13767 (N_13767,N_10355,N_11948);
nand U13768 (N_13768,N_10990,N_10570);
nand U13769 (N_13769,N_11439,N_11853);
xnor U13770 (N_13770,N_10754,N_11372);
nand U13771 (N_13771,N_10237,N_11935);
or U13772 (N_13772,N_10527,N_11838);
or U13773 (N_13773,N_10951,N_11508);
nor U13774 (N_13774,N_11292,N_11731);
nand U13775 (N_13775,N_10117,N_10043);
nor U13776 (N_13776,N_11238,N_10890);
nor U13777 (N_13777,N_11356,N_10484);
and U13778 (N_13778,N_10456,N_10531);
or U13779 (N_13779,N_11344,N_11991);
and U13780 (N_13780,N_10488,N_10894);
nor U13781 (N_13781,N_11573,N_11238);
or U13782 (N_13782,N_11190,N_11377);
nor U13783 (N_13783,N_11676,N_10493);
and U13784 (N_13784,N_11535,N_10669);
xor U13785 (N_13785,N_11569,N_10239);
nor U13786 (N_13786,N_11589,N_11191);
nor U13787 (N_13787,N_11890,N_10139);
nand U13788 (N_13788,N_10918,N_11527);
nand U13789 (N_13789,N_10517,N_10207);
xor U13790 (N_13790,N_10018,N_10563);
nor U13791 (N_13791,N_11830,N_11176);
or U13792 (N_13792,N_11958,N_11543);
and U13793 (N_13793,N_10838,N_11754);
or U13794 (N_13794,N_10186,N_10761);
nor U13795 (N_13795,N_10743,N_11467);
nand U13796 (N_13796,N_10834,N_11726);
xor U13797 (N_13797,N_11504,N_10056);
or U13798 (N_13798,N_11394,N_11508);
xor U13799 (N_13799,N_11985,N_10424);
and U13800 (N_13800,N_10713,N_11136);
nand U13801 (N_13801,N_10434,N_10507);
xor U13802 (N_13802,N_11794,N_10874);
xor U13803 (N_13803,N_11981,N_10083);
nor U13804 (N_13804,N_10664,N_11673);
xnor U13805 (N_13805,N_10923,N_10690);
xor U13806 (N_13806,N_10402,N_11700);
and U13807 (N_13807,N_11645,N_10269);
or U13808 (N_13808,N_11636,N_11314);
nand U13809 (N_13809,N_11172,N_10561);
or U13810 (N_13810,N_11966,N_11290);
or U13811 (N_13811,N_10866,N_10186);
xor U13812 (N_13812,N_11275,N_10691);
nor U13813 (N_13813,N_11752,N_10284);
or U13814 (N_13814,N_11236,N_11406);
nor U13815 (N_13815,N_11534,N_11718);
or U13816 (N_13816,N_10181,N_11754);
or U13817 (N_13817,N_10251,N_11314);
and U13818 (N_13818,N_10462,N_10455);
nor U13819 (N_13819,N_11917,N_11762);
or U13820 (N_13820,N_10489,N_11809);
xor U13821 (N_13821,N_10184,N_10107);
or U13822 (N_13822,N_11805,N_11692);
nand U13823 (N_13823,N_11097,N_11866);
xor U13824 (N_13824,N_10146,N_10831);
xnor U13825 (N_13825,N_11559,N_10537);
xnor U13826 (N_13826,N_11382,N_10868);
or U13827 (N_13827,N_11270,N_10814);
and U13828 (N_13828,N_11238,N_10661);
or U13829 (N_13829,N_10049,N_10438);
nand U13830 (N_13830,N_11053,N_10544);
or U13831 (N_13831,N_11749,N_10488);
xor U13832 (N_13832,N_11272,N_10375);
and U13833 (N_13833,N_11375,N_11350);
nor U13834 (N_13834,N_11176,N_10179);
or U13835 (N_13835,N_11604,N_11881);
nor U13836 (N_13836,N_11168,N_10970);
and U13837 (N_13837,N_10181,N_10511);
xnor U13838 (N_13838,N_11701,N_10704);
xnor U13839 (N_13839,N_11523,N_10168);
and U13840 (N_13840,N_11669,N_11866);
nand U13841 (N_13841,N_10470,N_11747);
and U13842 (N_13842,N_10977,N_10106);
and U13843 (N_13843,N_10298,N_10073);
xnor U13844 (N_13844,N_11288,N_10051);
nand U13845 (N_13845,N_11457,N_11383);
and U13846 (N_13846,N_11326,N_11954);
and U13847 (N_13847,N_10012,N_11983);
or U13848 (N_13848,N_10981,N_10736);
nor U13849 (N_13849,N_11201,N_11973);
nand U13850 (N_13850,N_10651,N_11439);
xor U13851 (N_13851,N_10639,N_11196);
nand U13852 (N_13852,N_11660,N_11098);
nor U13853 (N_13853,N_10420,N_11688);
xnor U13854 (N_13854,N_10067,N_11625);
and U13855 (N_13855,N_11999,N_11101);
or U13856 (N_13856,N_11189,N_11078);
and U13857 (N_13857,N_10832,N_10574);
xnor U13858 (N_13858,N_10632,N_10266);
or U13859 (N_13859,N_10053,N_10772);
and U13860 (N_13860,N_10754,N_11231);
nand U13861 (N_13861,N_11826,N_11184);
and U13862 (N_13862,N_11815,N_10581);
and U13863 (N_13863,N_11639,N_10027);
and U13864 (N_13864,N_11686,N_10039);
nand U13865 (N_13865,N_10642,N_11068);
or U13866 (N_13866,N_10917,N_10862);
xor U13867 (N_13867,N_10460,N_11218);
nand U13868 (N_13868,N_11642,N_10841);
or U13869 (N_13869,N_10314,N_10587);
or U13870 (N_13870,N_10381,N_11925);
xor U13871 (N_13871,N_10190,N_11384);
and U13872 (N_13872,N_11094,N_11756);
or U13873 (N_13873,N_10413,N_11137);
nand U13874 (N_13874,N_11734,N_11944);
or U13875 (N_13875,N_10367,N_11599);
or U13876 (N_13876,N_11922,N_11382);
or U13877 (N_13877,N_11733,N_11879);
and U13878 (N_13878,N_10137,N_11196);
nor U13879 (N_13879,N_11437,N_11222);
and U13880 (N_13880,N_11469,N_10485);
nand U13881 (N_13881,N_10142,N_11645);
nand U13882 (N_13882,N_10927,N_11344);
and U13883 (N_13883,N_10943,N_10388);
nor U13884 (N_13884,N_11757,N_11150);
and U13885 (N_13885,N_11749,N_10530);
and U13886 (N_13886,N_10355,N_10915);
and U13887 (N_13887,N_11053,N_10291);
and U13888 (N_13888,N_10342,N_10166);
nor U13889 (N_13889,N_10374,N_11456);
or U13890 (N_13890,N_11482,N_11421);
or U13891 (N_13891,N_10881,N_10727);
and U13892 (N_13892,N_10305,N_10300);
nor U13893 (N_13893,N_11875,N_10210);
xor U13894 (N_13894,N_10117,N_11993);
or U13895 (N_13895,N_10411,N_11366);
nor U13896 (N_13896,N_10359,N_11867);
nand U13897 (N_13897,N_11214,N_11601);
and U13898 (N_13898,N_10047,N_11532);
nor U13899 (N_13899,N_10287,N_11821);
nor U13900 (N_13900,N_10910,N_11359);
nand U13901 (N_13901,N_10100,N_10119);
xor U13902 (N_13902,N_11458,N_10844);
xor U13903 (N_13903,N_10795,N_10404);
nor U13904 (N_13904,N_11962,N_11825);
and U13905 (N_13905,N_11257,N_10414);
and U13906 (N_13906,N_11202,N_11672);
nand U13907 (N_13907,N_11459,N_11585);
xnor U13908 (N_13908,N_10166,N_11437);
nand U13909 (N_13909,N_10049,N_10640);
or U13910 (N_13910,N_10890,N_11177);
nand U13911 (N_13911,N_10550,N_11231);
nor U13912 (N_13912,N_10503,N_10473);
and U13913 (N_13913,N_11105,N_10631);
and U13914 (N_13914,N_10651,N_10981);
or U13915 (N_13915,N_10145,N_11310);
nand U13916 (N_13916,N_11036,N_11589);
xor U13917 (N_13917,N_10700,N_11672);
nand U13918 (N_13918,N_10302,N_10556);
or U13919 (N_13919,N_11511,N_11778);
nand U13920 (N_13920,N_11878,N_10234);
nand U13921 (N_13921,N_10192,N_11754);
nor U13922 (N_13922,N_11219,N_10318);
nor U13923 (N_13923,N_11879,N_11202);
xnor U13924 (N_13924,N_10141,N_11664);
and U13925 (N_13925,N_11831,N_10077);
xnor U13926 (N_13926,N_11247,N_11111);
and U13927 (N_13927,N_10399,N_10552);
and U13928 (N_13928,N_10707,N_11096);
and U13929 (N_13929,N_11618,N_11889);
xor U13930 (N_13930,N_11116,N_10478);
xor U13931 (N_13931,N_10388,N_11668);
and U13932 (N_13932,N_11629,N_11931);
nor U13933 (N_13933,N_10613,N_10126);
xnor U13934 (N_13934,N_11249,N_11729);
nand U13935 (N_13935,N_11072,N_10619);
or U13936 (N_13936,N_10222,N_10910);
nor U13937 (N_13937,N_11968,N_11906);
or U13938 (N_13938,N_11034,N_11823);
nand U13939 (N_13939,N_10749,N_10782);
nand U13940 (N_13940,N_11091,N_10508);
xor U13941 (N_13941,N_10718,N_11517);
xnor U13942 (N_13942,N_11432,N_10149);
xor U13943 (N_13943,N_10033,N_10867);
and U13944 (N_13944,N_11386,N_11118);
or U13945 (N_13945,N_10673,N_10670);
or U13946 (N_13946,N_10118,N_11389);
nor U13947 (N_13947,N_10833,N_10504);
xor U13948 (N_13948,N_11949,N_10389);
nand U13949 (N_13949,N_11179,N_11855);
xor U13950 (N_13950,N_11965,N_11557);
and U13951 (N_13951,N_11817,N_10890);
nand U13952 (N_13952,N_10936,N_11426);
nor U13953 (N_13953,N_10108,N_11407);
nor U13954 (N_13954,N_10080,N_10445);
nand U13955 (N_13955,N_10981,N_11564);
xor U13956 (N_13956,N_11479,N_11498);
nor U13957 (N_13957,N_11464,N_11750);
nand U13958 (N_13958,N_11180,N_11646);
xor U13959 (N_13959,N_10655,N_11332);
xor U13960 (N_13960,N_11566,N_11663);
xnor U13961 (N_13961,N_10733,N_11881);
xnor U13962 (N_13962,N_11385,N_10075);
or U13963 (N_13963,N_10162,N_11292);
nand U13964 (N_13964,N_11545,N_11149);
nand U13965 (N_13965,N_10254,N_10369);
or U13966 (N_13966,N_11034,N_11730);
nor U13967 (N_13967,N_10341,N_10437);
nand U13968 (N_13968,N_10305,N_10188);
xor U13969 (N_13969,N_11377,N_11422);
or U13970 (N_13970,N_10585,N_10752);
and U13971 (N_13971,N_11969,N_11181);
and U13972 (N_13972,N_10404,N_11129);
nor U13973 (N_13973,N_10377,N_11526);
xor U13974 (N_13974,N_11264,N_11347);
and U13975 (N_13975,N_10659,N_10555);
nand U13976 (N_13976,N_10181,N_10304);
and U13977 (N_13977,N_11896,N_10696);
xnor U13978 (N_13978,N_10769,N_10355);
nand U13979 (N_13979,N_11444,N_11063);
nand U13980 (N_13980,N_10589,N_11451);
xnor U13981 (N_13981,N_11920,N_11010);
and U13982 (N_13982,N_11529,N_10449);
nor U13983 (N_13983,N_10916,N_10082);
xor U13984 (N_13984,N_10754,N_11973);
and U13985 (N_13985,N_10607,N_11886);
xnor U13986 (N_13986,N_11752,N_11569);
and U13987 (N_13987,N_10657,N_11111);
nor U13988 (N_13988,N_11677,N_10886);
or U13989 (N_13989,N_11239,N_11172);
nand U13990 (N_13990,N_11869,N_11355);
and U13991 (N_13991,N_10595,N_11423);
or U13992 (N_13992,N_10071,N_11401);
or U13993 (N_13993,N_10060,N_11806);
xor U13994 (N_13994,N_11320,N_10842);
xor U13995 (N_13995,N_10355,N_11716);
xnor U13996 (N_13996,N_10685,N_10944);
nand U13997 (N_13997,N_10387,N_11471);
nor U13998 (N_13998,N_10752,N_11709);
and U13999 (N_13999,N_11026,N_10375);
or U14000 (N_14000,N_12632,N_13747);
nand U14001 (N_14001,N_12439,N_12811);
and U14002 (N_14002,N_12651,N_12927);
xor U14003 (N_14003,N_13280,N_13829);
or U14004 (N_14004,N_13940,N_12943);
xor U14005 (N_14005,N_12199,N_12914);
xnor U14006 (N_14006,N_12595,N_12638);
xor U14007 (N_14007,N_13188,N_13096);
nand U14008 (N_14008,N_13852,N_13804);
xnor U14009 (N_14009,N_12664,N_13507);
nand U14010 (N_14010,N_13077,N_12331);
nor U14011 (N_14011,N_13473,N_12428);
and U14012 (N_14012,N_13437,N_12018);
xnor U14013 (N_14013,N_13351,N_12585);
nor U14014 (N_14014,N_12765,N_13838);
xnor U14015 (N_14015,N_12644,N_12621);
or U14016 (N_14016,N_12965,N_13156);
and U14017 (N_14017,N_13134,N_13956);
or U14018 (N_14018,N_12752,N_13180);
and U14019 (N_14019,N_12564,N_12838);
nand U14020 (N_14020,N_13249,N_12633);
or U14021 (N_14021,N_13432,N_13759);
xor U14022 (N_14022,N_13035,N_12556);
and U14023 (N_14023,N_12101,N_12722);
nor U14024 (N_14024,N_13092,N_12923);
nor U14025 (N_14025,N_12951,N_13282);
and U14026 (N_14026,N_12495,N_13807);
nor U14027 (N_14027,N_12590,N_13052);
or U14028 (N_14028,N_12151,N_12374);
nor U14029 (N_14029,N_13319,N_12306);
nor U14030 (N_14030,N_12853,N_13532);
and U14031 (N_14031,N_13542,N_13118);
or U14032 (N_14032,N_13775,N_12142);
xnor U14033 (N_14033,N_13205,N_12614);
nand U14034 (N_14034,N_13619,N_12033);
and U14035 (N_14035,N_13192,N_12265);
nor U14036 (N_14036,N_13495,N_13251);
and U14037 (N_14037,N_12011,N_13826);
or U14038 (N_14038,N_12711,N_13292);
nor U14039 (N_14039,N_13164,N_12852);
nor U14040 (N_14040,N_13915,N_12121);
and U14041 (N_14041,N_12322,N_12190);
nand U14042 (N_14042,N_13451,N_13030);
and U14043 (N_14043,N_12936,N_13571);
nand U14044 (N_14044,N_13376,N_13399);
nor U14045 (N_14045,N_13259,N_12065);
and U14046 (N_14046,N_13355,N_13086);
nand U14047 (N_14047,N_13177,N_12820);
xor U14048 (N_14048,N_13873,N_12764);
or U14049 (N_14049,N_13230,N_13402);
xnor U14050 (N_14050,N_13763,N_13293);
nor U14051 (N_14051,N_13862,N_12582);
and U14052 (N_14052,N_13950,N_12677);
nand U14053 (N_14053,N_13048,N_13544);
or U14054 (N_14054,N_13124,N_13746);
nand U14055 (N_14055,N_13037,N_12946);
nor U14056 (N_14056,N_13558,N_13132);
xnor U14057 (N_14057,N_13817,N_12004);
nor U14058 (N_14058,N_12436,N_13444);
nor U14059 (N_14059,N_13988,N_12920);
nand U14060 (N_14060,N_13548,N_12997);
nand U14061 (N_14061,N_12160,N_13635);
xor U14062 (N_14062,N_12482,N_13466);
and U14063 (N_14063,N_12840,N_13816);
nand U14064 (N_14064,N_13993,N_12432);
nor U14065 (N_14065,N_13499,N_13799);
and U14066 (N_14066,N_12640,N_13452);
and U14067 (N_14067,N_12587,N_12201);
nand U14068 (N_14068,N_12691,N_13889);
nand U14069 (N_14069,N_13369,N_13331);
or U14070 (N_14070,N_13933,N_12387);
xor U14071 (N_14071,N_12808,N_13069);
nor U14072 (N_14072,N_13498,N_13574);
nand U14073 (N_14073,N_12348,N_12545);
or U14074 (N_14074,N_13729,N_13485);
xor U14075 (N_14075,N_12252,N_12657);
nand U14076 (N_14076,N_13700,N_12817);
and U14077 (N_14077,N_12412,N_13684);
nor U14078 (N_14078,N_13263,N_12938);
nor U14079 (N_14079,N_13411,N_12406);
and U14080 (N_14080,N_12656,N_12672);
xor U14081 (N_14081,N_13347,N_13670);
nor U14082 (N_14082,N_12944,N_13461);
or U14083 (N_14083,N_12518,N_13624);
nor U14084 (N_14084,N_13527,N_13632);
or U14085 (N_14085,N_12675,N_13952);
nand U14086 (N_14086,N_13934,N_12708);
xnor U14087 (N_14087,N_12670,N_12593);
nor U14088 (N_14088,N_12122,N_13051);
or U14089 (N_14089,N_13029,N_13577);
nor U14090 (N_14090,N_12441,N_12816);
nand U14091 (N_14091,N_12897,N_12976);
xnor U14092 (N_14092,N_12703,N_13623);
nor U14093 (N_14093,N_12391,N_13935);
nand U14094 (N_14094,N_12193,N_13598);
nand U14095 (N_14095,N_12224,N_12480);
xor U14096 (N_14096,N_13459,N_12110);
nand U14097 (N_14097,N_13036,N_13478);
xnor U14098 (N_14098,N_13782,N_13133);
xnor U14099 (N_14099,N_13801,N_12512);
or U14100 (N_14100,N_13825,N_13394);
xor U14101 (N_14101,N_12502,N_13438);
and U14102 (N_14102,N_12673,N_13242);
and U14103 (N_14103,N_13496,N_12909);
nand U14104 (N_14104,N_13716,N_13137);
and U14105 (N_14105,N_13543,N_13892);
nor U14106 (N_14106,N_13206,N_13207);
nor U14107 (N_14107,N_12723,N_12431);
and U14108 (N_14108,N_13784,N_12574);
nand U14109 (N_14109,N_12351,N_13645);
or U14110 (N_14110,N_13117,N_12460);
nor U14111 (N_14111,N_12639,N_13880);
nor U14112 (N_14112,N_12197,N_12696);
and U14113 (N_14113,N_12850,N_13406);
and U14114 (N_14114,N_13240,N_12119);
nand U14115 (N_14115,N_13278,N_13553);
xor U14116 (N_14116,N_12172,N_12051);
or U14117 (N_14117,N_13665,N_12453);
xor U14118 (N_14118,N_13354,N_12269);
and U14119 (N_14119,N_12916,N_13304);
or U14120 (N_14120,N_12216,N_12841);
or U14121 (N_14121,N_12520,N_12753);
nand U14122 (N_14122,N_13016,N_13013);
or U14123 (N_14123,N_13014,N_12885);
or U14124 (N_14124,N_13267,N_13503);
xnor U14125 (N_14125,N_13870,N_13919);
nand U14126 (N_14126,N_12855,N_12097);
and U14127 (N_14127,N_13162,N_12266);
nor U14128 (N_14128,N_13615,N_13458);
nand U14129 (N_14129,N_13359,N_12392);
or U14130 (N_14130,N_12140,N_13150);
and U14131 (N_14131,N_12859,N_13981);
nand U14132 (N_14132,N_13223,N_12034);
nand U14133 (N_14133,N_12583,N_12293);
xnor U14134 (N_14134,N_12731,N_12036);
and U14135 (N_14135,N_13813,N_12655);
nor U14136 (N_14136,N_13701,N_12833);
nor U14137 (N_14137,N_13294,N_12434);
nand U14138 (N_14138,N_12327,N_12356);
and U14139 (N_14139,N_12230,N_13634);
nor U14140 (N_14140,N_12438,N_13216);
and U14141 (N_14141,N_12718,N_13165);
or U14142 (N_14142,N_12894,N_13455);
or U14143 (N_14143,N_12769,N_13812);
or U14144 (N_14144,N_12493,N_13239);
or U14145 (N_14145,N_13937,N_12321);
nor U14146 (N_14146,N_13612,N_13403);
nor U14147 (N_14147,N_12008,N_12598);
xnor U14148 (N_14148,N_12009,N_12246);
or U14149 (N_14149,N_13017,N_13297);
xor U14150 (N_14150,N_13885,N_12109);
nor U14151 (N_14151,N_13640,N_12187);
nor U14152 (N_14152,N_13751,N_13334);
nor U14153 (N_14153,N_12861,N_12262);
xnor U14154 (N_14154,N_13616,N_12364);
nor U14155 (N_14155,N_12061,N_12044);
nand U14156 (N_14156,N_13814,N_12043);
and U14157 (N_14157,N_12342,N_13894);
xnor U14158 (N_14158,N_12272,N_12697);
and U14159 (N_14159,N_13991,N_12608);
or U14160 (N_14160,N_13637,N_12782);
and U14161 (N_14161,N_12551,N_13606);
nand U14162 (N_14162,N_13877,N_13677);
nor U14163 (N_14163,N_12473,N_12295);
xnor U14164 (N_14164,N_12700,N_13038);
or U14165 (N_14165,N_13520,N_13979);
nand U14166 (N_14166,N_12251,N_13453);
and U14167 (N_14167,N_13450,N_12604);
xnor U14168 (N_14168,N_13815,N_12531);
nand U14169 (N_14169,N_12826,N_12735);
nand U14170 (N_14170,N_12645,N_12258);
nand U14171 (N_14171,N_13725,N_12329);
nand U14172 (N_14172,N_12002,N_12468);
nand U14173 (N_14173,N_12452,N_13323);
nand U14174 (N_14174,N_12071,N_13288);
nor U14175 (N_14175,N_12161,N_13345);
and U14176 (N_14176,N_12413,N_12733);
xor U14177 (N_14177,N_12537,N_13744);
xnor U14178 (N_14178,N_12973,N_13776);
and U14179 (N_14179,N_12601,N_13078);
nor U14180 (N_14180,N_12757,N_12991);
nand U14181 (N_14181,N_12501,N_13456);
or U14182 (N_14182,N_12966,N_13925);
and U14183 (N_14183,N_13788,N_12040);
nand U14184 (N_14184,N_13088,N_12899);
xnor U14185 (N_14185,N_13022,N_13113);
and U14186 (N_14186,N_13413,N_13248);
and U14187 (N_14187,N_13254,N_13941);
xnor U14188 (N_14188,N_12876,N_12661);
xnor U14189 (N_14189,N_12509,N_12416);
and U14190 (N_14190,N_13899,N_13435);
nand U14191 (N_14191,N_12194,N_12349);
or U14192 (N_14192,N_13228,N_12877);
xor U14193 (N_14193,N_13045,N_12345);
or U14194 (N_14194,N_13390,N_12114);
xnor U14195 (N_14195,N_13146,N_12381);
or U14196 (N_14196,N_12622,N_13955);
nor U14197 (N_14197,N_13704,N_13696);
nor U14198 (N_14198,N_13342,N_12420);
nand U14199 (N_14199,N_12546,N_12910);
xor U14200 (N_14200,N_12450,N_12609);
or U14201 (N_14201,N_13514,N_12292);
and U14202 (N_14202,N_13839,N_13060);
xor U14203 (N_14203,N_13631,N_12568);
xnor U14204 (N_14204,N_12344,N_12611);
xnor U14205 (N_14205,N_13739,N_13064);
and U14206 (N_14206,N_13440,N_13380);
and U14207 (N_14207,N_12027,N_12143);
nand U14208 (N_14208,N_13987,N_13869);
nor U14209 (N_14209,N_13734,N_12892);
or U14210 (N_14210,N_12298,N_13457);
nand U14211 (N_14211,N_13591,N_12830);
xor U14212 (N_14212,N_12744,N_13678);
and U14213 (N_14213,N_13913,N_13592);
xnor U14214 (N_14214,N_13115,N_13600);
nand U14215 (N_14215,N_12162,N_13810);
nand U14216 (N_14216,N_12815,N_12549);
or U14217 (N_14217,N_13718,N_13143);
nand U14218 (N_14218,N_12929,N_13252);
xnor U14219 (N_14219,N_12414,N_12357);
and U14220 (N_14220,N_12496,N_13502);
or U14221 (N_14221,N_13486,N_13126);
and U14222 (N_14222,N_12103,N_12834);
nand U14223 (N_14223,N_12831,N_12083);
nor U14224 (N_14224,N_13525,N_12784);
nor U14225 (N_14225,N_12869,N_13214);
and U14226 (N_14226,N_13443,N_12257);
nor U14227 (N_14227,N_13295,N_13673);
and U14228 (N_14228,N_13794,N_13447);
and U14229 (N_14229,N_13774,N_12543);
or U14230 (N_14230,N_13985,N_12993);
and U14231 (N_14231,N_12934,N_12014);
nand U14232 (N_14232,N_12302,N_12000);
or U14233 (N_14233,N_12147,N_13924);
or U14234 (N_14234,N_13743,N_13803);
xnor U14235 (N_14235,N_12163,N_13266);
nand U14236 (N_14236,N_12280,N_12760);
or U14237 (N_14237,N_13489,N_12205);
xnor U14238 (N_14238,N_12023,N_13479);
nand U14239 (N_14239,N_13408,N_12271);
and U14240 (N_14240,N_12681,N_13856);
nor U14241 (N_14241,N_12353,N_12182);
or U14242 (N_14242,N_13875,N_12042);
and U14243 (N_14243,N_12523,N_12129);
or U14244 (N_14244,N_13805,N_13573);
xnor U14245 (N_14245,N_12317,N_12049);
and U14246 (N_14246,N_13594,N_13256);
nor U14247 (N_14247,N_12303,N_12717);
nand U14248 (N_14248,N_12297,N_13510);
xor U14249 (N_14249,N_12365,N_12594);
xor U14250 (N_14250,N_12307,N_13127);
nor U14251 (N_14251,N_12961,N_12519);
nand U14252 (N_14252,N_12339,N_12481);
or U14253 (N_14253,N_13557,N_13806);
xnor U14254 (N_14254,N_12825,N_12940);
xnor U14255 (N_14255,N_13383,N_12120);
nor U14256 (N_14256,N_12690,N_12950);
xnor U14257 (N_14257,N_13714,N_12912);
or U14258 (N_14258,N_13145,N_13170);
nor U14259 (N_14259,N_12309,N_13008);
or U14260 (N_14260,N_12851,N_13578);
or U14261 (N_14261,N_12807,N_13238);
and U14262 (N_14262,N_13027,N_12806);
xor U14263 (N_14263,N_13693,N_12746);
xor U14264 (N_14264,N_13785,N_13861);
nand U14265 (N_14265,N_13850,N_12971);
xnor U14266 (N_14266,N_13951,N_12157);
or U14267 (N_14267,N_13823,N_13664);
xor U14268 (N_14268,N_12602,N_12076);
and U14269 (N_14269,N_12024,N_12962);
xor U14270 (N_14270,N_13015,N_13681);
xnor U14271 (N_14271,N_12171,N_12898);
and U14272 (N_14272,N_13446,N_12795);
and U14273 (N_14273,N_12107,N_12067);
nor U14274 (N_14274,N_12975,N_13909);
nor U14275 (N_14275,N_12095,N_13575);
nand U14276 (N_14276,N_12062,N_12457);
and U14277 (N_14277,N_12400,N_13268);
and U14278 (N_14278,N_12591,N_12694);
and U14279 (N_14279,N_13655,N_13626);
or U14280 (N_14280,N_12259,N_13983);
or U14281 (N_14281,N_13367,N_12900);
nor U14282 (N_14282,N_12487,N_12243);
nand U14283 (N_14283,N_13586,N_12492);
nand U14284 (N_14284,N_13686,N_12176);
nand U14285 (N_14285,N_13795,N_13057);
and U14286 (N_14286,N_12278,N_12641);
and U14287 (N_14287,N_12276,N_12111);
nand U14288 (N_14288,N_13777,N_13787);
xnor U14289 (N_14289,N_13083,N_12300);
nand U14290 (N_14290,N_13003,N_13625);
or U14291 (N_14291,N_12394,N_12433);
xor U14292 (N_14292,N_13296,N_12072);
or U14293 (N_14293,N_12872,N_13313);
nand U14294 (N_14294,N_13521,N_12207);
xor U14295 (N_14295,N_13610,N_13650);
or U14296 (N_14296,N_13647,N_12476);
nor U14297 (N_14297,N_13358,N_13427);
xor U14298 (N_14298,N_13968,N_12650);
nand U14299 (N_14299,N_13727,N_13872);
nor U14300 (N_14300,N_13175,N_13505);
xor U14301 (N_14301,N_13439,N_12783);
nand U14302 (N_14302,N_13093,N_13781);
xnor U14303 (N_14303,N_13771,N_13471);
and U14304 (N_14304,N_12557,N_12294);
nor U14305 (N_14305,N_12378,N_12754);
nand U14306 (N_14306,N_13998,N_13707);
and U14307 (N_14307,N_13318,N_12737);
xnor U14308 (N_14308,N_12165,N_12709);
or U14309 (N_14309,N_13595,N_12469);
nand U14310 (N_14310,N_13247,N_12385);
nand U14311 (N_14311,N_13199,N_13546);
nand U14312 (N_14312,N_12893,N_12925);
nor U14313 (N_14313,N_12542,N_12268);
nor U14314 (N_14314,N_13196,N_12889);
and U14315 (N_14315,N_13195,N_12146);
xor U14316 (N_14316,N_12016,N_12627);
nand U14317 (N_14317,N_12430,N_13762);
nor U14318 (N_14318,N_12710,N_12352);
and U14319 (N_14319,N_12256,N_12895);
and U14320 (N_14320,N_13912,N_13928);
nor U14321 (N_14321,N_13703,N_13808);
and U14322 (N_14322,N_12813,N_13965);
nor U14323 (N_14323,N_12497,N_12053);
and U14324 (N_14324,N_13299,N_13041);
nand U14325 (N_14325,N_12462,N_12776);
xor U14326 (N_14326,N_13627,N_13225);
xor U14327 (N_14327,N_13141,N_12333);
and U14328 (N_14328,N_13617,N_12210);
xnor U14329 (N_14329,N_12706,N_12793);
and U14330 (N_14330,N_12836,N_13533);
nor U14331 (N_14331,N_13745,N_13153);
and U14332 (N_14332,N_12461,N_13379);
or U14333 (N_14333,N_13072,N_12138);
nor U14334 (N_14334,N_13215,N_13720);
or U14335 (N_14335,N_12686,N_13377);
nor U14336 (N_14336,N_12631,N_12941);
xor U14337 (N_14337,N_12446,N_13392);
or U14338 (N_14338,N_12569,N_13613);
or U14339 (N_14339,N_12939,N_12167);
and U14340 (N_14340,N_13602,N_13648);
xor U14341 (N_14341,N_12408,N_12522);
nor U14342 (N_14342,N_13980,N_12283);
nor U14343 (N_14343,N_12637,N_12313);
xor U14344 (N_14344,N_13085,N_12144);
or U14345 (N_14345,N_13706,N_13436);
nand U14346 (N_14346,N_13000,N_12041);
or U14347 (N_14347,N_13348,N_13140);
xnor U14348 (N_14348,N_13608,N_13897);
or U14349 (N_14349,N_13680,N_12248);
nor U14350 (N_14350,N_12241,N_12483);
and U14351 (N_14351,N_12514,N_13584);
nand U14352 (N_14352,N_13308,N_13246);
nand U14353 (N_14353,N_12228,N_13154);
nor U14354 (N_14354,N_12619,N_12766);
xor U14355 (N_14355,N_12756,N_13112);
and U14356 (N_14356,N_13949,N_12541);
nor U14357 (N_14357,N_12104,N_12277);
nand U14358 (N_14358,N_13986,N_13152);
and U14359 (N_14359,N_13357,N_13531);
or U14360 (N_14360,N_12328,N_12935);
nand U14361 (N_14361,N_13537,N_13136);
nand U14362 (N_14362,N_12242,N_12864);
xnor U14363 (N_14363,N_13375,N_13820);
nor U14364 (N_14364,N_13683,N_13786);
nor U14365 (N_14365,N_13149,N_13321);
xnor U14366 (N_14366,N_13559,N_12857);
xnor U14367 (N_14367,N_13961,N_12687);
nor U14368 (N_14368,N_12001,N_13837);
or U14369 (N_14369,N_12134,N_13477);
nor U14370 (N_14370,N_13234,N_12013);
nor U14371 (N_14371,N_13960,N_13066);
and U14372 (N_14372,N_12038,N_12652);
and U14373 (N_14373,N_12994,N_13135);
nor U14374 (N_14374,N_12156,N_12918);
or U14375 (N_14375,N_13504,N_12311);
and U14376 (N_14376,N_12505,N_13530);
nor U14377 (N_14377,N_12603,N_13235);
and U14378 (N_14378,N_12674,N_12159);
nand U14379 (N_14379,N_13901,N_12287);
or U14380 (N_14380,N_13522,N_12704);
nor U14381 (N_14381,N_12084,N_12273);
xnor U14382 (N_14382,N_12695,N_13824);
and U14383 (N_14383,N_12646,N_13846);
or U14384 (N_14384,N_13047,N_12498);
nand U14385 (N_14385,N_12048,N_13350);
and U14386 (N_14386,N_13310,N_12548);
xnor U14387 (N_14387,N_13517,N_12382);
nor U14388 (N_14388,N_13419,N_12981);
xnor U14389 (N_14389,N_13738,N_12139);
and U14390 (N_14390,N_12663,N_13766);
nand U14391 (N_14391,N_13942,N_13974);
nor U14392 (N_14392,N_13001,N_12239);
xnor U14393 (N_14393,N_12456,N_12534);
nor U14394 (N_14394,N_13876,N_12029);
xnor U14395 (N_14395,N_13087,N_12800);
or U14396 (N_14396,N_13679,N_13844);
and U14397 (N_14397,N_13211,N_13976);
nand U14398 (N_14398,N_12858,N_12070);
nand U14399 (N_14399,N_12102,N_13198);
or U14400 (N_14400,N_12837,N_13589);
and U14401 (N_14401,N_12599,N_12136);
and U14402 (N_14402,N_13340,N_12113);
nor U14403 (N_14403,N_13075,N_13204);
xor U14404 (N_14404,N_12253,N_13285);
and U14405 (N_14405,N_12781,N_13868);
nor U14406 (N_14406,N_13420,N_13081);
nand U14407 (N_14407,N_13190,N_12592);
or U14408 (N_14408,N_13539,N_13653);
or U14409 (N_14409,N_13271,N_13274);
nor U14410 (N_14410,N_13506,N_13791);
xor U14411 (N_14411,N_13668,N_12238);
or U14412 (N_14412,N_13131,N_13611);
nand U14413 (N_14413,N_13138,N_12959);
xor U14414 (N_14414,N_13094,N_12131);
and U14415 (N_14415,N_13732,N_13042);
nand U14416 (N_14416,N_12445,N_12092);
nand U14417 (N_14417,N_12491,N_13765);
nor U14418 (N_14418,N_13270,N_13519);
nor U14419 (N_14419,N_12977,N_12422);
or U14420 (N_14420,N_13301,N_13984);
xnor U14421 (N_14421,N_12558,N_13058);
or U14422 (N_14422,N_12485,N_13374);
or U14423 (N_14423,N_13835,N_13621);
xor U14424 (N_14424,N_13434,N_12570);
or U14425 (N_14425,N_13480,N_12472);
nor U14426 (N_14426,N_13307,N_13494);
or U14427 (N_14427,N_13863,N_12901);
nor U14428 (N_14428,N_13167,N_12748);
nor U14429 (N_14429,N_12179,N_13418);
and U14430 (N_14430,N_12533,N_13091);
nand U14431 (N_14431,N_12643,N_13883);
and U14432 (N_14432,N_13638,N_12478);
and U14433 (N_14433,N_12540,N_13995);
and U14434 (N_14434,N_12740,N_12600);
nor U14435 (N_14435,N_13338,N_13726);
nor U14436 (N_14436,N_13373,N_12220);
nand U14437 (N_14437,N_13740,N_13298);
nand U14438 (N_14438,N_12347,N_13277);
xor U14439 (N_14439,N_13713,N_12196);
and U14440 (N_14440,N_12906,N_12589);
nand U14441 (N_14441,N_12073,N_13958);
nor U14442 (N_14442,N_13019,N_12372);
nand U14443 (N_14443,N_12863,N_12435);
or U14444 (N_14444,N_12979,N_12931);
xnor U14445 (N_14445,N_13541,N_12117);
xnor U14446 (N_14446,N_12891,N_13848);
and U14447 (N_14447,N_12026,N_12279);
nand U14448 (N_14448,N_12818,N_12218);
nor U14449 (N_14449,N_13258,N_12343);
xnor U14450 (N_14450,N_12792,N_13040);
nor U14451 (N_14451,N_13929,N_12449);
and U14452 (N_14452,N_12383,N_13107);
and U14453 (N_14453,N_12954,N_12318);
or U14454 (N_14454,N_13874,N_12281);
nand U14455 (N_14455,N_13100,N_12181);
nand U14456 (N_14456,N_13953,N_12921);
or U14457 (N_14457,N_13741,N_13202);
nand U14458 (N_14458,N_13121,N_13472);
or U14459 (N_14459,N_12596,N_12046);
nor U14460 (N_14460,N_13967,N_13853);
nor U14461 (N_14461,N_13341,N_12668);
and U14462 (N_14462,N_13903,N_13629);
xor U14463 (N_14463,N_12775,N_12928);
xnor U14464 (N_14464,N_13330,N_12970);
nor U14465 (N_14465,N_12154,N_12719);
and U14466 (N_14466,N_13628,N_13265);
nor U14467 (N_14467,N_12955,N_12559);
nor U14468 (N_14468,N_13948,N_12320);
xnor U14469 (N_14469,N_12057,N_12698);
xnor U14470 (N_14470,N_12884,N_12986);
or U14471 (N_14471,N_13320,N_12508);
nor U14472 (N_14472,N_13409,N_12126);
nor U14473 (N_14473,N_13865,N_12094);
xor U14474 (N_14474,N_13857,N_13702);
nand U14475 (N_14475,N_12079,N_13328);
and U14476 (N_14476,N_12903,N_12573);
or U14477 (N_14477,N_12960,N_13695);
and U14478 (N_14478,N_13099,N_12286);
and U14479 (N_14479,N_12085,N_12770);
xor U14480 (N_14480,N_13333,N_13315);
and U14481 (N_14481,N_13119,N_12237);
nand U14482 (N_14482,N_12226,N_12787);
xnor U14483 (N_14483,N_12610,N_13316);
nand U14484 (N_14484,N_13372,N_12566);
and U14485 (N_14485,N_13737,N_12701);
nand U14486 (N_14486,N_13335,N_12032);
nand U14487 (N_14487,N_12411,N_13034);
and U14488 (N_14488,N_13054,N_12688);
and U14489 (N_14489,N_12919,N_13104);
nand U14490 (N_14490,N_13212,N_12209);
or U14491 (N_14491,N_13387,N_13144);
nand U14492 (N_14492,N_13061,N_12847);
nor U14493 (N_14493,N_12552,N_13364);
nor U14494 (N_14494,N_13609,N_12093);
xor U14495 (N_14495,N_13605,N_12184);
xnor U14496 (N_14496,N_12249,N_13855);
or U14497 (N_14497,N_13893,N_12953);
nand U14498 (N_14498,N_12059,N_13360);
nor U14499 (N_14499,N_12440,N_12069);
or U14500 (N_14500,N_12538,N_12035);
or U14501 (N_14501,N_13245,N_13555);
or U14502 (N_14502,N_12949,N_13428);
or U14503 (N_14503,N_12405,N_13840);
or U14504 (N_14504,N_12123,N_13906);
and U14505 (N_14505,N_12204,N_13690);
nor U14506 (N_14506,N_13866,N_12799);
nor U14507 (N_14507,N_12749,N_12198);
and U14508 (N_14508,N_13314,N_13491);
nor U14509 (N_14509,N_12789,N_12264);
nand U14510 (N_14510,N_12370,N_13898);
xnor U14511 (N_14511,N_13276,N_12562);
xnor U14512 (N_14512,N_12447,N_13849);
xor U14513 (N_14513,N_12060,N_13157);
or U14514 (N_14514,N_12550,N_13148);
and U14515 (N_14515,N_12010,N_13286);
nor U14516 (N_14516,N_12212,N_13658);
nor U14517 (N_14517,N_13881,N_13705);
xnor U14518 (N_14518,N_13200,N_13032);
xor U14519 (N_14519,N_12584,N_13910);
xor U14520 (N_14520,N_12424,N_13395);
xor U14521 (N_14521,N_13864,N_13487);
nor U14522 (N_14522,N_12750,N_13604);
and U14523 (N_14523,N_12458,N_13067);
nor U14524 (N_14524,N_13526,N_13977);
and U14525 (N_14525,N_12532,N_12289);
nand U14526 (N_14526,N_12354,N_13346);
and U14527 (N_14527,N_13513,N_12705);
nand U14528 (N_14528,N_13750,N_13847);
xor U14529 (N_14529,N_12796,N_13076);
and U14530 (N_14530,N_13073,N_12425);
nand U14531 (N_14531,N_13173,N_12835);
nand U14532 (N_14532,N_13063,N_13719);
or U14533 (N_14533,N_13469,N_13709);
nor U14534 (N_14534,N_12995,N_12178);
and U14535 (N_14535,N_12200,N_13197);
nor U14536 (N_14536,N_13349,N_13708);
nor U14537 (N_14537,N_12628,N_13540);
and U14538 (N_14538,N_12845,N_12626);
and U14539 (N_14539,N_12494,N_13975);
nor U14540 (N_14540,N_12235,N_13462);
nor U14541 (N_14541,N_12856,N_12319);
nand U14542 (N_14542,N_12888,N_13226);
nand U14543 (N_14543,N_12108,N_13449);
xor U14544 (N_14544,N_13026,N_12056);
nand U14545 (N_14545,N_12100,N_12219);
xor U14546 (N_14546,N_12525,N_13493);
and U14547 (N_14547,N_12527,N_13155);
nor U14548 (N_14548,N_12539,N_13070);
nor U14549 (N_14549,N_12788,N_13065);
and U14550 (N_14550,N_12653,N_13780);
nor U14551 (N_14551,N_12854,N_13770);
and U14552 (N_14552,N_12135,N_12255);
and U14553 (N_14553,N_12772,N_12571);
xnor U14554 (N_14554,N_13569,N_13516);
nand U14555 (N_14555,N_12515,N_12455);
xnor U14556 (N_14556,N_12310,N_13689);
and U14557 (N_14557,N_13264,N_13186);
nor U14558 (N_14558,N_13191,N_13879);
nor U14559 (N_14559,N_13769,N_12667);
or U14560 (N_14560,N_13698,N_13858);
nor U14561 (N_14561,N_13822,N_13642);
xor U14562 (N_14562,N_13109,N_12250);
nand U14563 (N_14563,N_13685,N_12964);
nor U14564 (N_14564,N_13261,N_12213);
or U14565 (N_14565,N_13189,N_12526);
xor U14566 (N_14566,N_13767,N_12443);
or U14567 (N_14567,N_13970,N_12106);
and U14568 (N_14568,N_13179,N_12809);
and U14569 (N_14569,N_13962,N_13311);
and U14570 (N_14570,N_13867,N_12225);
or U14571 (N_14571,N_13760,N_12880);
or U14572 (N_14572,N_12606,N_12822);
and U14573 (N_14573,N_12082,N_12517);
or U14574 (N_14574,N_12802,N_12285);
xor U14575 (N_14575,N_12148,N_13992);
xnor U14576 (N_14576,N_13400,N_13515);
and U14577 (N_14577,N_12911,N_12177);
xnor U14578 (N_14578,N_12702,N_12867);
nor U14579 (N_14579,N_12952,N_13959);
nand U14580 (N_14580,N_12658,N_12074);
xor U14581 (N_14581,N_12730,N_13753);
or U14582 (N_14582,N_13071,N_13423);
nor U14583 (N_14583,N_12399,N_13585);
xnor U14584 (N_14584,N_13662,N_12890);
nand U14585 (N_14585,N_13474,N_13229);
and U14586 (N_14586,N_12350,N_12335);
nand U14587 (N_14587,N_12747,N_12426);
xor U14588 (N_14588,N_13227,N_13887);
xor U14589 (N_14589,N_13550,N_13587);
nor U14590 (N_14590,N_13902,N_12716);
or U14591 (N_14591,N_12671,N_13878);
nor U14592 (N_14592,N_12827,N_12742);
nand U14593 (N_14593,N_12214,N_13994);
nand U14594 (N_14594,N_13244,N_13208);
and U14595 (N_14595,N_13819,N_13217);
and U14596 (N_14596,N_12474,N_13920);
and U14597 (N_14597,N_13731,N_12798);
nor U14598 (N_14598,N_12222,N_13931);
and U14599 (N_14599,N_12774,N_12985);
nand U14600 (N_14600,N_13442,N_12448);
nor U14601 (N_14601,N_12878,N_12149);
and U14602 (N_14602,N_13943,N_13445);
nand U14603 (N_14603,N_13568,N_12510);
nor U14604 (N_14604,N_12341,N_12992);
nor U14605 (N_14605,N_12284,N_13467);
nand U14606 (N_14606,N_13581,N_13010);
and U14607 (N_14607,N_13715,N_12907);
nand U14608 (N_14608,N_12124,N_12922);
and U14609 (N_14609,N_12586,N_12945);
nor U14610 (N_14610,N_12908,N_12296);
xnor U14611 (N_14611,N_12797,N_13033);
nor U14612 (N_14612,N_12503,N_13882);
and U14613 (N_14613,N_12019,N_13969);
xnor U14614 (N_14614,N_13344,N_12254);
or U14615 (N_14615,N_12990,N_13554);
nor U14616 (N_14616,N_12947,N_12804);
nor U14617 (N_14617,N_13222,N_13329);
xor U14618 (N_14618,N_13821,N_13833);
nand U14619 (N_14619,N_12409,N_12873);
xnor U14620 (N_14620,N_13111,N_13666);
nand U14621 (N_14621,N_13352,N_12366);
xor U14622 (N_14622,N_12314,N_13936);
nand U14623 (N_14623,N_12087,N_13798);
nand U14624 (N_14624,N_13921,N_12407);
nor U14625 (N_14625,N_13062,N_12725);
or U14626 (N_14626,N_13756,N_13106);
xor U14627 (N_14627,N_12524,N_12183);
and U14628 (N_14628,N_12058,N_13957);
and U14629 (N_14629,N_13300,N_13224);
xnor U14630 (N_14630,N_13724,N_13772);
nand U14631 (N_14631,N_13989,N_12654);
and U14632 (N_14632,N_13305,N_12470);
and U14633 (N_14633,N_12616,N_12128);
or U14634 (N_14634,N_13710,N_12488);
nand U14635 (N_14635,N_12575,N_13778);
nor U14636 (N_14636,N_12007,N_13095);
and U14637 (N_14637,N_12301,N_13185);
or U14638 (N_14638,N_13371,N_13488);
and U14639 (N_14639,N_12516,N_13108);
or U14640 (N_14640,N_12227,N_13939);
xnor U14641 (N_14641,N_12739,N_13643);
and U14642 (N_14642,N_13580,N_12917);
nor U14643 (N_14643,N_13021,N_12437);
and U14644 (N_14644,N_13945,N_13535);
xor U14645 (N_14645,N_12150,N_12395);
nor U14646 (N_14646,N_13006,N_12332);
nor U14647 (N_14647,N_12490,N_13828);
nor U14648 (N_14648,N_12915,N_12232);
or U14649 (N_14649,N_13098,N_12682);
or U14650 (N_14650,N_12022,N_13272);
xor U14651 (N_14651,N_13068,N_12299);
and U14652 (N_14652,N_13291,N_13614);
nand U14653 (N_14653,N_12786,N_12377);
xnor U14654 (N_14654,N_13018,N_12588);
or U14655 (N_14655,N_13669,N_13147);
and U14656 (N_14656,N_13790,N_13549);
nor U14657 (N_14657,N_12507,N_12844);
and U14658 (N_14658,N_12153,N_13923);
xnor U14659 (N_14659,N_13796,N_13187);
nand U14660 (N_14660,N_12189,N_13233);
nor U14661 (N_14661,N_13888,N_13890);
nor U14662 (N_14662,N_13389,N_12417);
xor U14663 (N_14663,N_12086,N_13663);
xnor U14664 (N_14664,N_12389,N_12099);
xnor U14665 (N_14665,N_13009,N_12623);
or U14666 (N_14666,N_13529,N_12359);
or U14667 (N_14667,N_13545,N_12132);
or U14668 (N_14668,N_12063,N_13570);
xor U14669 (N_14669,N_13536,N_12423);
and U14670 (N_14670,N_13023,N_13944);
and U14671 (N_14671,N_12741,N_12629);
or U14672 (N_14672,N_13797,N_12089);
nand U14673 (N_14673,N_13281,N_13674);
or U14674 (N_14674,N_12031,N_13105);
nand U14675 (N_14675,N_12761,N_13220);
xor U14676 (N_14676,N_13084,N_13916);
and U14677 (N_14677,N_12988,N_12270);
xor U14678 (N_14678,N_12553,N_13260);
and U14679 (N_14679,N_13845,N_12360);
nand U14680 (N_14680,N_13914,N_12486);
nor U14681 (N_14681,N_12875,N_13414);
nand U14682 (N_14682,N_12234,N_12466);
xor U14683 (N_14683,N_13163,N_12913);
or U14684 (N_14684,N_12229,N_13891);
or U14685 (N_14685,N_12555,N_13748);
xor U14686 (N_14686,N_13930,N_13652);
and U14687 (N_14687,N_13151,N_12942);
or U14688 (N_14688,N_13908,N_13723);
nand U14689 (N_14689,N_12173,N_12020);
xnor U14690 (N_14690,N_13365,N_12767);
xnor U14691 (N_14691,N_12615,N_12170);
or U14692 (N_14692,N_12684,N_12839);
nand U14693 (N_14693,N_13044,N_12355);
nor U14694 (N_14694,N_13337,N_12267);
nand U14695 (N_14695,N_12052,N_12721);
and U14696 (N_14696,N_12208,N_12115);
or U14697 (N_14697,N_13332,N_12367);
xnor U14698 (N_14698,N_13509,N_12477);
xnor U14699 (N_14699,N_12967,N_12137);
nor U14700 (N_14700,N_12883,N_13004);
and U14701 (N_14701,N_13393,N_12972);
or U14702 (N_14702,N_13900,N_12904);
nand U14703 (N_14703,N_13166,N_12777);
nor U14704 (N_14704,N_13181,N_13031);
nor U14705 (N_14705,N_13221,N_12489);
and U14706 (N_14706,N_13871,N_12081);
xor U14707 (N_14707,N_13468,N_13596);
nand U14708 (N_14708,N_13454,N_12091);
nand U14709 (N_14709,N_13236,N_13269);
nor U14710 (N_14710,N_13896,N_12152);
nand U14711 (N_14711,N_13682,N_13213);
nand U14712 (N_14712,N_12155,N_13564);
and U14713 (N_14713,N_12386,N_12418);
nand U14714 (N_14714,N_13938,N_13429);
nand U14715 (N_14715,N_13327,N_13460);
xnor U14716 (N_14716,N_13182,N_12169);
nor U14717 (N_14717,N_13560,N_13511);
and U14718 (N_14718,N_12419,N_12785);
nor U14719 (N_14719,N_12404,N_13809);
or U14720 (N_14720,N_13620,N_12678);
xnor U14721 (N_14721,N_12771,N_13500);
nand U14722 (N_14722,N_13290,N_12451);
xor U14723 (N_14723,N_12685,N_12164);
nand U14724 (N_14724,N_12231,N_12755);
nand U14725 (N_14725,N_13733,N_12005);
or U14726 (N_14726,N_13792,N_13385);
nand U14727 (N_14727,N_12535,N_12832);
or U14728 (N_14728,N_13667,N_12479);
nor U14729 (N_14729,N_12261,N_12398);
nor U14730 (N_14730,N_13243,N_13911);
nand U14731 (N_14731,N_12726,N_12186);
xnor U14732 (N_14732,N_13241,N_12734);
and U14733 (N_14733,N_12824,N_13687);
or U14734 (N_14734,N_13309,N_12127);
xor U14735 (N_14735,N_13325,N_13465);
or U14736 (N_14736,N_12998,N_13688);
nand U14737 (N_14737,N_12828,N_12736);
or U14738 (N_14738,N_13056,N_13717);
xor U14739 (N_14739,N_12580,N_13080);
xor U14740 (N_14740,N_13721,N_12634);
and U14741 (N_14741,N_12315,N_13492);
nand U14742 (N_14742,N_12617,N_12896);
and U14743 (N_14743,N_13842,N_13178);
and U14744 (N_14744,N_13742,N_12030);
xor U14745 (N_14745,N_12363,N_12871);
and U14746 (N_14746,N_12846,N_13572);
and U14747 (N_14747,N_12624,N_13947);
and U14748 (N_14748,N_13441,N_13607);
nand U14749 (N_14749,N_13128,N_13370);
xnor U14750 (N_14750,N_13275,N_13830);
or U14751 (N_14751,N_12980,N_13169);
nor U14752 (N_14752,N_12037,N_13524);
nor U14753 (N_14753,N_13361,N_13562);
xor U14754 (N_14754,N_12511,N_12006);
nand U14755 (N_14755,N_12978,N_12215);
xnor U14756 (N_14756,N_13827,N_12689);
xor U14757 (N_14757,N_13884,N_13490);
nor U14758 (N_14758,N_12015,N_13074);
or U14759 (N_14759,N_12791,N_13210);
nor U14760 (N_14760,N_13851,N_13583);
nor U14761 (N_14761,N_12105,N_12471);
xnor U14762 (N_14762,N_12429,N_13386);
nor U14763 (N_14763,N_12373,N_13971);
or U14764 (N_14764,N_13999,N_13886);
and U14765 (N_14765,N_13255,N_12751);
and U14766 (N_14766,N_12958,N_12948);
xnor U14767 (N_14767,N_12393,N_13356);
and U14768 (N_14768,N_13028,N_12554);
nor U14769 (N_14769,N_12096,N_13425);
and U14770 (N_14770,N_13818,N_13317);
and U14771 (N_14771,N_12762,N_12865);
xnor U14772 (N_14772,N_12968,N_12727);
nor U14773 (N_14773,N_12660,N_12801);
nor U14774 (N_14774,N_13159,N_12338);
nand U14775 (N_14775,N_13161,N_12759);
and U14776 (N_14776,N_13430,N_12605);
or U14777 (N_14777,N_12375,N_13176);
xnor U14778 (N_14778,N_13907,N_13381);
nor U14779 (N_14779,N_12368,N_12565);
xnor U14780 (N_14780,N_12166,N_12371);
nor U14781 (N_14781,N_12984,N_13656);
and U14782 (N_14782,N_12388,N_13582);
or U14783 (N_14783,N_12956,N_13757);
or U14784 (N_14784,N_12064,N_13972);
nor U14785 (N_14785,N_13566,N_13590);
nand U14786 (N_14786,N_12078,N_12054);
and U14787 (N_14787,N_12221,N_12195);
nand U14788 (N_14788,N_13482,N_12499);
nand U14789 (N_14789,N_12974,N_12879);
or U14790 (N_14790,N_12475,N_12669);
or U14791 (N_14791,N_13534,N_13407);
or U14792 (N_14792,N_12848,N_12484);
and U14793 (N_14793,N_13257,N_12464);
xor U14794 (N_14794,N_12763,N_12247);
or U14795 (N_14795,N_13966,N_12459);
nand U14796 (N_14796,N_12713,N_13694);
nor U14797 (N_14797,N_13597,N_13997);
xor U14798 (N_14798,N_12088,N_12098);
and U14799 (N_14799,N_13752,N_12810);
nor U14800 (N_14800,N_13501,N_13287);
and U14801 (N_14801,N_13676,N_12340);
or U14802 (N_14802,N_13836,N_13834);
nand U14803 (N_14803,N_12513,N_13917);
xor U14804 (N_14804,N_12886,N_12665);
and U14805 (N_14805,N_12547,N_12790);
nor U14806 (N_14806,N_12116,N_12068);
nand U14807 (N_14807,N_12745,N_13779);
and U14808 (N_14808,N_13384,N_12882);
nor U14809 (N_14809,N_13363,N_12648);
xnor U14810 (N_14810,N_13843,N_13672);
xnor U14811 (N_14811,N_12028,N_12185);
and U14812 (N_14812,N_12612,N_13722);
and U14813 (N_14813,N_13284,N_13926);
or U14814 (N_14814,N_13250,N_12233);
nand U14815 (N_14815,N_12729,N_13978);
xnor U14816 (N_14816,N_12803,N_12738);
nor U14817 (N_14817,N_13476,N_13905);
nand U14818 (N_14818,N_13523,N_13927);
or U14819 (N_14819,N_13283,N_12390);
nand U14820 (N_14820,N_13654,N_12812);
and U14821 (N_14821,N_12402,N_13946);
and U14822 (N_14822,N_12397,N_13463);
nand U14823 (N_14823,N_12282,N_13758);
nor U14824 (N_14824,N_12969,N_13618);
xor U14825 (N_14825,N_13007,N_12125);
nand U14826 (N_14826,N_13755,N_13129);
or U14827 (N_14827,N_13593,N_12870);
xnor U14828 (N_14828,N_13860,N_12724);
nor U14829 (N_14829,N_13262,N_12647);
nor U14830 (N_14830,N_13353,N_13730);
nand U14831 (N_14831,N_13831,N_13046);
nand U14832 (N_14832,N_12707,N_12275);
xor U14833 (N_14833,N_13551,N_13172);
nor U14834 (N_14834,N_13661,N_13005);
and U14835 (N_14835,N_13339,N_12130);
or U14836 (N_14836,N_12223,N_12467);
nor U14837 (N_14837,N_12017,N_12659);
nor U14838 (N_14838,N_12819,N_13538);
xnor U14839 (N_14839,N_13055,N_13518);
xor U14840 (N_14840,N_12773,N_13324);
nor U14841 (N_14841,N_13711,N_12561);
nand U14842 (N_14842,N_13193,N_12989);
xnor U14843 (N_14843,N_12563,N_12500);
or U14844 (N_14844,N_13547,N_13728);
xnor U14845 (N_14845,N_12203,N_12090);
or U14846 (N_14846,N_13789,N_13416);
xnor U14847 (N_14847,N_12794,N_12823);
and U14848 (N_14848,N_13556,N_13484);
or U14849 (N_14849,N_13649,N_12642);
nand U14850 (N_14850,N_13859,N_13512);
nor U14851 (N_14851,N_12025,N_13079);
nor U14852 (N_14852,N_12504,N_13398);
and U14853 (N_14853,N_13388,N_13783);
xor U14854 (N_14854,N_12358,N_13168);
xor U14855 (N_14855,N_13561,N_12630);
or U14856 (N_14856,N_13059,N_13563);
nor U14857 (N_14857,N_13712,N_12649);
or U14858 (N_14858,N_13139,N_13644);
or U14859 (N_14859,N_12323,N_12401);
and U14860 (N_14860,N_12175,N_13336);
or U14861 (N_14861,N_12732,N_12683);
and U14862 (N_14862,N_12560,N_13125);
or U14863 (N_14863,N_12410,N_13160);
or U14864 (N_14864,N_13089,N_13675);
nor U14865 (N_14865,N_13417,N_12403);
xor U14866 (N_14866,N_13378,N_13761);
and U14867 (N_14867,N_13483,N_12236);
xnor U14868 (N_14868,N_12003,N_12263);
xor U14869 (N_14869,N_13382,N_13918);
or U14870 (N_14870,N_13343,N_13973);
xor U14871 (N_14871,N_13422,N_13012);
nand U14872 (N_14872,N_12260,N_13904);
or U14873 (N_14873,N_13481,N_13552);
or U14874 (N_14874,N_12983,N_13657);
and U14875 (N_14875,N_13424,N_13768);
or U14876 (N_14876,N_13426,N_12528);
nor U14877 (N_14877,N_12308,N_13289);
xnor U14878 (N_14878,N_13312,N_13954);
xnor U14879 (N_14879,N_13603,N_13630);
nor U14880 (N_14880,N_12168,N_12380);
nor U14881 (N_14881,N_12712,N_12932);
or U14882 (N_14882,N_13231,N_12240);
xor U14883 (N_14883,N_13218,N_12521);
or U14884 (N_14884,N_13203,N_13053);
or U14885 (N_14885,N_13405,N_12180);
or U14886 (N_14886,N_12578,N_13497);
and U14887 (N_14887,N_13641,N_12607);
and U14888 (N_14888,N_12743,N_13366);
or U14889 (N_14889,N_12330,N_13431);
or U14890 (N_14890,N_12191,N_12780);
xor U14891 (N_14891,N_12805,N_12715);
or U14892 (N_14892,N_13391,N_12666);
xnor U14893 (N_14893,N_13588,N_12572);
nor U14894 (N_14894,N_12924,N_12758);
nand U14895 (N_14895,N_12933,N_13002);
nor U14896 (N_14896,N_12312,N_12618);
and U14897 (N_14897,N_12544,N_12112);
nor U14898 (N_14898,N_13764,N_13024);
and U14899 (N_14899,N_12047,N_12821);
xor U14900 (N_14900,N_13692,N_12699);
or U14901 (N_14901,N_12720,N_12369);
nor U14902 (N_14902,N_12530,N_13097);
nand U14903 (N_14903,N_13464,N_12957);
nand U14904 (N_14904,N_13174,N_13802);
and U14905 (N_14905,N_13433,N_13011);
xnor U14906 (N_14906,N_13567,N_13749);
and U14907 (N_14907,N_12679,N_12874);
and U14908 (N_14908,N_12379,N_13050);
and U14909 (N_14909,N_12075,N_13932);
nand U14910 (N_14910,N_13636,N_12577);
nor U14911 (N_14911,N_12304,N_12174);
or U14912 (N_14912,N_13671,N_13579);
and U14913 (N_14913,N_12188,N_12996);
nand U14914 (N_14914,N_13025,N_13120);
and U14915 (N_14915,N_13996,N_12465);
and U14916 (N_14916,N_13130,N_13622);
or U14917 (N_14917,N_12325,N_13102);
nor U14918 (N_14918,N_13773,N_12118);
or U14919 (N_14919,N_13101,N_13800);
nor U14920 (N_14920,N_13183,N_12999);
and U14921 (N_14921,N_12536,N_12396);
xor U14922 (N_14922,N_13123,N_12427);
xnor U14923 (N_14923,N_12768,N_12244);
and U14924 (N_14924,N_12576,N_13090);
xor U14925 (N_14925,N_12039,N_13982);
nor U14926 (N_14926,N_12778,N_12291);
nor U14927 (N_14927,N_12905,N_12887);
nand U14928 (N_14928,N_13697,N_12714);
nand U14929 (N_14929,N_13114,N_12926);
nand U14930 (N_14930,N_12982,N_13116);
or U14931 (N_14931,N_13362,N_12862);
nand U14932 (N_14932,N_13660,N_12077);
xnor U14933 (N_14933,N_12693,N_13158);
xor U14934 (N_14934,N_12021,N_12829);
nand U14935 (N_14935,N_13326,N_12326);
nor U14936 (N_14936,N_13237,N_12866);
or U14937 (N_14937,N_12842,N_12635);
and U14938 (N_14938,N_13232,N_13322);
xnor U14939 (N_14939,N_13401,N_12055);
nor U14940 (N_14940,N_12567,N_13184);
and U14941 (N_14941,N_13049,N_12625);
nand U14942 (N_14942,N_12336,N_12636);
nand U14943 (N_14943,N_12362,N_13302);
xor U14944 (N_14944,N_12274,N_13599);
xnor U14945 (N_14945,N_13811,N_13171);
nor U14946 (N_14946,N_13421,N_13368);
nor U14947 (N_14947,N_13396,N_12692);
xor U14948 (N_14948,N_12444,N_12987);
nor U14949 (N_14949,N_12158,N_13279);
xor U14950 (N_14950,N_12930,N_13735);
xnor U14951 (N_14951,N_13122,N_12288);
or U14952 (N_14952,N_13576,N_13854);
nor U14953 (N_14953,N_13306,N_13964);
nor U14954 (N_14954,N_12620,N_12579);
xnor U14955 (N_14955,N_12581,N_13691);
and U14956 (N_14956,N_12045,N_12080);
nand U14957 (N_14957,N_13253,N_12211);
and U14958 (N_14958,N_13646,N_13832);
and U14959 (N_14959,N_12728,N_13475);
or U14960 (N_14960,N_12963,N_12814);
xor U14961 (N_14961,N_12506,N_12337);
nand U14962 (N_14962,N_12937,N_13103);
nor U14963 (N_14963,N_12529,N_12454);
and U14964 (N_14964,N_13020,N_12202);
or U14965 (N_14965,N_13565,N_12384);
xor U14966 (N_14966,N_12217,N_13201);
nor U14967 (N_14967,N_13736,N_12133);
and U14968 (N_14968,N_13793,N_13142);
nand U14969 (N_14969,N_12849,N_13841);
nor U14970 (N_14970,N_13082,N_12421);
nand U14971 (N_14971,N_13470,N_13412);
nor U14972 (N_14972,N_13963,N_13448);
nand U14973 (N_14973,N_12050,N_12361);
nor U14974 (N_14974,N_12012,N_12662);
and U14975 (N_14975,N_13754,N_13273);
nor U14976 (N_14976,N_13528,N_13209);
nand U14977 (N_14977,N_13043,N_13639);
or U14978 (N_14978,N_12290,N_13633);
xnor U14979 (N_14979,N_12779,N_13699);
or U14980 (N_14980,N_12141,N_13039);
xor U14981 (N_14981,N_13601,N_12902);
nor U14982 (N_14982,N_13415,N_12597);
and U14983 (N_14983,N_12680,N_12442);
nor U14984 (N_14984,N_12316,N_13651);
nor U14985 (N_14985,N_12868,N_13659);
or U14986 (N_14986,N_12881,N_12192);
or U14987 (N_14987,N_12305,N_13110);
nand U14988 (N_14988,N_13194,N_13508);
or U14989 (N_14989,N_13410,N_13219);
nand U14990 (N_14990,N_13303,N_13895);
or U14991 (N_14991,N_12145,N_12334);
or U14992 (N_14992,N_13922,N_12415);
and U14993 (N_14993,N_12463,N_12860);
and U14994 (N_14994,N_12676,N_12324);
nor U14995 (N_14995,N_12376,N_13404);
nor U14996 (N_14996,N_12843,N_12346);
xor U14997 (N_14997,N_12245,N_12066);
nor U14998 (N_14998,N_13990,N_12206);
xor U14999 (N_14999,N_13397,N_12613);
and U15000 (N_15000,N_13985,N_13651);
nand U15001 (N_15001,N_12406,N_12002);
or U15002 (N_15002,N_13533,N_12721);
xor U15003 (N_15003,N_12225,N_13660);
or U15004 (N_15004,N_12508,N_12009);
and U15005 (N_15005,N_12498,N_12196);
or U15006 (N_15006,N_13352,N_13942);
nor U15007 (N_15007,N_12778,N_13745);
nand U15008 (N_15008,N_12386,N_13913);
nor U15009 (N_15009,N_12641,N_13465);
and U15010 (N_15010,N_13068,N_13195);
and U15011 (N_15011,N_12200,N_13331);
nand U15012 (N_15012,N_12328,N_12989);
nor U15013 (N_15013,N_13518,N_13612);
nand U15014 (N_15014,N_13736,N_12765);
nand U15015 (N_15015,N_13759,N_12651);
or U15016 (N_15016,N_13113,N_13883);
xor U15017 (N_15017,N_12935,N_12055);
and U15018 (N_15018,N_12535,N_12201);
nand U15019 (N_15019,N_12427,N_12769);
nand U15020 (N_15020,N_13164,N_13141);
nand U15021 (N_15021,N_13213,N_13211);
and U15022 (N_15022,N_13521,N_12522);
nor U15023 (N_15023,N_13859,N_13224);
and U15024 (N_15024,N_13432,N_13683);
nor U15025 (N_15025,N_13464,N_12057);
nand U15026 (N_15026,N_13642,N_12070);
nand U15027 (N_15027,N_12572,N_12507);
nor U15028 (N_15028,N_12150,N_12506);
nand U15029 (N_15029,N_12891,N_13911);
or U15030 (N_15030,N_12899,N_13367);
xnor U15031 (N_15031,N_13640,N_12028);
xor U15032 (N_15032,N_12985,N_13632);
and U15033 (N_15033,N_12210,N_12066);
nand U15034 (N_15034,N_13365,N_13066);
or U15035 (N_15035,N_12477,N_12930);
and U15036 (N_15036,N_12055,N_13486);
nand U15037 (N_15037,N_12605,N_12904);
and U15038 (N_15038,N_12554,N_13886);
nand U15039 (N_15039,N_13803,N_12280);
or U15040 (N_15040,N_13321,N_12064);
nand U15041 (N_15041,N_13228,N_13028);
or U15042 (N_15042,N_13853,N_13696);
or U15043 (N_15043,N_12962,N_12611);
or U15044 (N_15044,N_13036,N_13961);
or U15045 (N_15045,N_13325,N_12327);
and U15046 (N_15046,N_12018,N_12483);
and U15047 (N_15047,N_12840,N_12402);
or U15048 (N_15048,N_13993,N_13486);
nand U15049 (N_15049,N_13856,N_13936);
nand U15050 (N_15050,N_12269,N_13991);
xor U15051 (N_15051,N_13277,N_12801);
and U15052 (N_15052,N_13706,N_13877);
and U15053 (N_15053,N_12772,N_13340);
xor U15054 (N_15054,N_12129,N_13734);
xnor U15055 (N_15055,N_13086,N_12464);
nand U15056 (N_15056,N_13712,N_13967);
and U15057 (N_15057,N_13679,N_12935);
or U15058 (N_15058,N_12865,N_13849);
or U15059 (N_15059,N_12208,N_13707);
nand U15060 (N_15060,N_13477,N_12129);
or U15061 (N_15061,N_12402,N_13514);
xnor U15062 (N_15062,N_13421,N_12992);
nand U15063 (N_15063,N_12000,N_12099);
nand U15064 (N_15064,N_12578,N_13557);
nand U15065 (N_15065,N_13928,N_13031);
or U15066 (N_15066,N_12336,N_13354);
nand U15067 (N_15067,N_12391,N_12988);
and U15068 (N_15068,N_12594,N_12734);
and U15069 (N_15069,N_12921,N_12413);
nor U15070 (N_15070,N_13360,N_12371);
xnor U15071 (N_15071,N_13903,N_12326);
nor U15072 (N_15072,N_12758,N_13645);
xor U15073 (N_15073,N_12915,N_13219);
and U15074 (N_15074,N_13625,N_12603);
or U15075 (N_15075,N_13041,N_12157);
xnor U15076 (N_15076,N_13273,N_12997);
nand U15077 (N_15077,N_12142,N_13192);
and U15078 (N_15078,N_12705,N_12514);
xnor U15079 (N_15079,N_12006,N_13732);
nor U15080 (N_15080,N_12705,N_13255);
nand U15081 (N_15081,N_12944,N_12625);
nor U15082 (N_15082,N_13065,N_13586);
nand U15083 (N_15083,N_13287,N_13776);
nand U15084 (N_15084,N_12070,N_12501);
and U15085 (N_15085,N_12795,N_12306);
nand U15086 (N_15086,N_13418,N_13051);
nor U15087 (N_15087,N_13764,N_13782);
nand U15088 (N_15088,N_12859,N_12257);
xor U15089 (N_15089,N_12349,N_13709);
or U15090 (N_15090,N_13339,N_12730);
and U15091 (N_15091,N_12774,N_12296);
nor U15092 (N_15092,N_13506,N_12578);
and U15093 (N_15093,N_13588,N_13734);
xnor U15094 (N_15094,N_13929,N_12057);
nand U15095 (N_15095,N_13255,N_12284);
nor U15096 (N_15096,N_13558,N_13928);
or U15097 (N_15097,N_13051,N_13273);
nand U15098 (N_15098,N_12349,N_13224);
nor U15099 (N_15099,N_13661,N_12823);
or U15100 (N_15100,N_13520,N_13371);
and U15101 (N_15101,N_12543,N_12697);
nor U15102 (N_15102,N_12245,N_13036);
nand U15103 (N_15103,N_12524,N_13769);
and U15104 (N_15104,N_13632,N_13522);
xnor U15105 (N_15105,N_13643,N_12388);
xnor U15106 (N_15106,N_12499,N_13381);
or U15107 (N_15107,N_12046,N_12337);
or U15108 (N_15108,N_12302,N_12828);
and U15109 (N_15109,N_12472,N_12637);
or U15110 (N_15110,N_13774,N_13802);
or U15111 (N_15111,N_13692,N_13563);
nand U15112 (N_15112,N_12256,N_13605);
or U15113 (N_15113,N_13181,N_12543);
or U15114 (N_15114,N_13258,N_13636);
nand U15115 (N_15115,N_13204,N_13402);
and U15116 (N_15116,N_12556,N_12855);
and U15117 (N_15117,N_13805,N_12208);
or U15118 (N_15118,N_13488,N_13916);
nor U15119 (N_15119,N_12066,N_12120);
xor U15120 (N_15120,N_12774,N_13910);
nand U15121 (N_15121,N_12782,N_13712);
and U15122 (N_15122,N_13953,N_13792);
and U15123 (N_15123,N_12023,N_12440);
and U15124 (N_15124,N_12982,N_13468);
nand U15125 (N_15125,N_12839,N_13296);
nor U15126 (N_15126,N_12096,N_13331);
nor U15127 (N_15127,N_13537,N_12944);
xor U15128 (N_15128,N_13467,N_12213);
nand U15129 (N_15129,N_12231,N_13856);
xor U15130 (N_15130,N_12615,N_13206);
or U15131 (N_15131,N_13695,N_12215);
nand U15132 (N_15132,N_12475,N_13017);
and U15133 (N_15133,N_12005,N_12948);
or U15134 (N_15134,N_13133,N_13480);
nor U15135 (N_15135,N_12025,N_12998);
nand U15136 (N_15136,N_13912,N_13612);
and U15137 (N_15137,N_13772,N_13798);
or U15138 (N_15138,N_13965,N_12472);
nor U15139 (N_15139,N_13972,N_13297);
nor U15140 (N_15140,N_13591,N_13048);
nand U15141 (N_15141,N_13487,N_12783);
nand U15142 (N_15142,N_12204,N_12259);
or U15143 (N_15143,N_13622,N_12705);
and U15144 (N_15144,N_12927,N_13566);
nand U15145 (N_15145,N_12640,N_13443);
nor U15146 (N_15146,N_13063,N_13872);
xor U15147 (N_15147,N_13033,N_13463);
and U15148 (N_15148,N_13041,N_12095);
xor U15149 (N_15149,N_13519,N_12504);
nand U15150 (N_15150,N_13727,N_12156);
nor U15151 (N_15151,N_12840,N_13079);
xnor U15152 (N_15152,N_13343,N_12843);
or U15153 (N_15153,N_12480,N_13745);
nand U15154 (N_15154,N_12684,N_13154);
and U15155 (N_15155,N_12877,N_13560);
and U15156 (N_15156,N_12690,N_13172);
nor U15157 (N_15157,N_12022,N_13982);
nand U15158 (N_15158,N_12448,N_12966);
and U15159 (N_15159,N_12218,N_13134);
nor U15160 (N_15160,N_12554,N_12662);
and U15161 (N_15161,N_12910,N_12075);
and U15162 (N_15162,N_12197,N_13413);
xor U15163 (N_15163,N_13549,N_13843);
nor U15164 (N_15164,N_12329,N_13739);
nand U15165 (N_15165,N_13218,N_13574);
or U15166 (N_15166,N_12970,N_13794);
nor U15167 (N_15167,N_12766,N_13131);
nand U15168 (N_15168,N_13727,N_13717);
nor U15169 (N_15169,N_13751,N_13934);
nor U15170 (N_15170,N_12549,N_12580);
nor U15171 (N_15171,N_13934,N_13886);
nor U15172 (N_15172,N_13156,N_13971);
nand U15173 (N_15173,N_13847,N_12598);
xnor U15174 (N_15174,N_13351,N_13196);
nor U15175 (N_15175,N_13856,N_12996);
nor U15176 (N_15176,N_12744,N_13929);
nor U15177 (N_15177,N_12968,N_13834);
nor U15178 (N_15178,N_12129,N_12310);
or U15179 (N_15179,N_12565,N_13699);
or U15180 (N_15180,N_12484,N_13991);
nor U15181 (N_15181,N_13452,N_13426);
xor U15182 (N_15182,N_12418,N_13424);
xor U15183 (N_15183,N_13426,N_12697);
and U15184 (N_15184,N_12655,N_12847);
xnor U15185 (N_15185,N_12892,N_12429);
nor U15186 (N_15186,N_12550,N_13554);
nor U15187 (N_15187,N_13296,N_13672);
nand U15188 (N_15188,N_12324,N_13835);
nor U15189 (N_15189,N_12712,N_12510);
or U15190 (N_15190,N_13576,N_13484);
nor U15191 (N_15191,N_13324,N_13797);
nor U15192 (N_15192,N_13959,N_13323);
xor U15193 (N_15193,N_13135,N_12343);
or U15194 (N_15194,N_12241,N_12962);
nand U15195 (N_15195,N_12681,N_12388);
xnor U15196 (N_15196,N_12581,N_12822);
and U15197 (N_15197,N_13397,N_12528);
xnor U15198 (N_15198,N_12527,N_13529);
nor U15199 (N_15199,N_12263,N_13561);
xnor U15200 (N_15200,N_13029,N_12703);
nand U15201 (N_15201,N_13299,N_12586);
or U15202 (N_15202,N_12528,N_13643);
and U15203 (N_15203,N_12163,N_13470);
and U15204 (N_15204,N_12207,N_13091);
or U15205 (N_15205,N_12422,N_13411);
nand U15206 (N_15206,N_12205,N_12588);
or U15207 (N_15207,N_12811,N_13068);
xor U15208 (N_15208,N_12166,N_13828);
or U15209 (N_15209,N_12397,N_12877);
nand U15210 (N_15210,N_12549,N_13355);
or U15211 (N_15211,N_12860,N_13120);
xnor U15212 (N_15212,N_12710,N_12445);
or U15213 (N_15213,N_13282,N_13270);
nand U15214 (N_15214,N_12447,N_13651);
and U15215 (N_15215,N_12013,N_12207);
or U15216 (N_15216,N_13711,N_13685);
and U15217 (N_15217,N_12377,N_13187);
nand U15218 (N_15218,N_12436,N_12655);
or U15219 (N_15219,N_13133,N_12775);
nand U15220 (N_15220,N_12084,N_13704);
xor U15221 (N_15221,N_13762,N_12798);
and U15222 (N_15222,N_12112,N_12707);
and U15223 (N_15223,N_13659,N_12371);
or U15224 (N_15224,N_12857,N_12714);
nor U15225 (N_15225,N_12427,N_13422);
or U15226 (N_15226,N_12181,N_13657);
nand U15227 (N_15227,N_12419,N_13049);
nor U15228 (N_15228,N_12995,N_13884);
nand U15229 (N_15229,N_13860,N_12601);
and U15230 (N_15230,N_12765,N_13800);
xor U15231 (N_15231,N_12819,N_12868);
and U15232 (N_15232,N_12162,N_12311);
xor U15233 (N_15233,N_12950,N_13580);
xnor U15234 (N_15234,N_12674,N_12905);
or U15235 (N_15235,N_13511,N_12774);
xor U15236 (N_15236,N_12462,N_12089);
and U15237 (N_15237,N_12433,N_13033);
xnor U15238 (N_15238,N_13230,N_13575);
xor U15239 (N_15239,N_13113,N_13519);
or U15240 (N_15240,N_12252,N_12468);
nor U15241 (N_15241,N_13623,N_12508);
or U15242 (N_15242,N_13957,N_13638);
or U15243 (N_15243,N_12597,N_13790);
nand U15244 (N_15244,N_12197,N_13061);
nor U15245 (N_15245,N_13687,N_13905);
nor U15246 (N_15246,N_12931,N_12098);
nor U15247 (N_15247,N_13284,N_12016);
and U15248 (N_15248,N_12006,N_12943);
nand U15249 (N_15249,N_13738,N_12805);
and U15250 (N_15250,N_13835,N_13063);
nor U15251 (N_15251,N_12978,N_12299);
nor U15252 (N_15252,N_12505,N_12848);
nor U15253 (N_15253,N_12110,N_12082);
nand U15254 (N_15254,N_13150,N_13351);
or U15255 (N_15255,N_12586,N_13851);
or U15256 (N_15256,N_13255,N_12952);
nand U15257 (N_15257,N_13024,N_12657);
nand U15258 (N_15258,N_12007,N_13068);
xor U15259 (N_15259,N_13143,N_13915);
nand U15260 (N_15260,N_13360,N_12715);
nor U15261 (N_15261,N_13973,N_12043);
nor U15262 (N_15262,N_12988,N_13961);
or U15263 (N_15263,N_12683,N_13851);
nor U15264 (N_15264,N_12495,N_13197);
or U15265 (N_15265,N_13109,N_13997);
or U15266 (N_15266,N_12220,N_12276);
or U15267 (N_15267,N_13474,N_13083);
xnor U15268 (N_15268,N_12967,N_13716);
or U15269 (N_15269,N_12182,N_12716);
xnor U15270 (N_15270,N_13833,N_13297);
and U15271 (N_15271,N_12558,N_13559);
and U15272 (N_15272,N_13341,N_13802);
nand U15273 (N_15273,N_13812,N_12941);
and U15274 (N_15274,N_13941,N_13862);
or U15275 (N_15275,N_12522,N_13196);
nand U15276 (N_15276,N_13590,N_12301);
xor U15277 (N_15277,N_12768,N_13526);
nand U15278 (N_15278,N_12587,N_13724);
xnor U15279 (N_15279,N_13825,N_13475);
and U15280 (N_15280,N_12555,N_13766);
and U15281 (N_15281,N_12162,N_12899);
nand U15282 (N_15282,N_12390,N_13229);
xnor U15283 (N_15283,N_13657,N_12546);
nor U15284 (N_15284,N_13970,N_13726);
xnor U15285 (N_15285,N_12903,N_12706);
nor U15286 (N_15286,N_13467,N_12989);
xor U15287 (N_15287,N_13943,N_13822);
nand U15288 (N_15288,N_12137,N_13546);
nand U15289 (N_15289,N_12581,N_12593);
nor U15290 (N_15290,N_13085,N_13395);
nor U15291 (N_15291,N_13990,N_12016);
xnor U15292 (N_15292,N_13974,N_13748);
xor U15293 (N_15293,N_13148,N_13496);
and U15294 (N_15294,N_12179,N_13376);
xor U15295 (N_15295,N_13822,N_13964);
xnor U15296 (N_15296,N_13065,N_12970);
nand U15297 (N_15297,N_12832,N_13479);
xnor U15298 (N_15298,N_13104,N_12897);
xnor U15299 (N_15299,N_12132,N_12692);
and U15300 (N_15300,N_12123,N_13010);
nand U15301 (N_15301,N_13612,N_12276);
or U15302 (N_15302,N_13366,N_13273);
nand U15303 (N_15303,N_12613,N_12096);
and U15304 (N_15304,N_13779,N_13240);
or U15305 (N_15305,N_13278,N_13856);
and U15306 (N_15306,N_12604,N_13809);
nand U15307 (N_15307,N_13824,N_12618);
xnor U15308 (N_15308,N_13841,N_13835);
and U15309 (N_15309,N_12364,N_12246);
and U15310 (N_15310,N_12184,N_12164);
nor U15311 (N_15311,N_12611,N_12903);
or U15312 (N_15312,N_13207,N_13083);
and U15313 (N_15313,N_13214,N_12892);
xnor U15314 (N_15314,N_12696,N_13134);
nor U15315 (N_15315,N_13273,N_13207);
nor U15316 (N_15316,N_12482,N_12220);
and U15317 (N_15317,N_13193,N_13038);
xor U15318 (N_15318,N_12080,N_12758);
and U15319 (N_15319,N_12236,N_12507);
and U15320 (N_15320,N_12079,N_12910);
nor U15321 (N_15321,N_13363,N_13950);
or U15322 (N_15322,N_12629,N_12680);
and U15323 (N_15323,N_13797,N_12441);
or U15324 (N_15324,N_13703,N_12081);
and U15325 (N_15325,N_13559,N_13311);
nand U15326 (N_15326,N_13604,N_12517);
xnor U15327 (N_15327,N_12225,N_13939);
nor U15328 (N_15328,N_12902,N_13786);
nor U15329 (N_15329,N_12078,N_13994);
nor U15330 (N_15330,N_13603,N_12454);
and U15331 (N_15331,N_12035,N_12950);
and U15332 (N_15332,N_12734,N_12091);
nor U15333 (N_15333,N_12609,N_12351);
nand U15334 (N_15334,N_13086,N_13448);
xnor U15335 (N_15335,N_12162,N_13470);
xor U15336 (N_15336,N_12865,N_13239);
nand U15337 (N_15337,N_12288,N_13900);
and U15338 (N_15338,N_12682,N_12269);
or U15339 (N_15339,N_12354,N_13886);
nand U15340 (N_15340,N_13285,N_13480);
and U15341 (N_15341,N_13550,N_13403);
xnor U15342 (N_15342,N_12816,N_12057);
and U15343 (N_15343,N_13846,N_13261);
nor U15344 (N_15344,N_12507,N_13031);
or U15345 (N_15345,N_13235,N_13892);
xnor U15346 (N_15346,N_12825,N_13880);
xnor U15347 (N_15347,N_12529,N_13613);
nand U15348 (N_15348,N_13539,N_13935);
xnor U15349 (N_15349,N_12384,N_13628);
and U15350 (N_15350,N_13221,N_12848);
and U15351 (N_15351,N_12915,N_13023);
xnor U15352 (N_15352,N_13310,N_13163);
nand U15353 (N_15353,N_13458,N_12267);
and U15354 (N_15354,N_12488,N_13818);
xnor U15355 (N_15355,N_12861,N_12867);
nand U15356 (N_15356,N_13017,N_12989);
nand U15357 (N_15357,N_12715,N_12901);
and U15358 (N_15358,N_13823,N_13276);
nor U15359 (N_15359,N_13032,N_12589);
xor U15360 (N_15360,N_13171,N_12226);
or U15361 (N_15361,N_12680,N_13033);
or U15362 (N_15362,N_12249,N_12606);
nand U15363 (N_15363,N_13680,N_13868);
and U15364 (N_15364,N_12797,N_12618);
and U15365 (N_15365,N_13997,N_12986);
nand U15366 (N_15366,N_13968,N_13487);
or U15367 (N_15367,N_13381,N_12417);
xnor U15368 (N_15368,N_12241,N_12079);
and U15369 (N_15369,N_13920,N_13061);
or U15370 (N_15370,N_13292,N_12626);
nand U15371 (N_15371,N_12211,N_12966);
or U15372 (N_15372,N_13724,N_12262);
nor U15373 (N_15373,N_13616,N_13404);
and U15374 (N_15374,N_12927,N_13445);
nand U15375 (N_15375,N_12589,N_13954);
nor U15376 (N_15376,N_13529,N_13588);
or U15377 (N_15377,N_12182,N_12341);
or U15378 (N_15378,N_12606,N_13989);
or U15379 (N_15379,N_12876,N_12105);
nand U15380 (N_15380,N_13577,N_12108);
or U15381 (N_15381,N_12428,N_12618);
xnor U15382 (N_15382,N_12687,N_12262);
and U15383 (N_15383,N_13913,N_12951);
nor U15384 (N_15384,N_13349,N_12843);
nor U15385 (N_15385,N_12701,N_13159);
or U15386 (N_15386,N_13631,N_12099);
xor U15387 (N_15387,N_12222,N_13096);
nor U15388 (N_15388,N_12058,N_12567);
xor U15389 (N_15389,N_13753,N_13131);
nor U15390 (N_15390,N_13141,N_13058);
nor U15391 (N_15391,N_12306,N_13887);
nand U15392 (N_15392,N_12616,N_13268);
and U15393 (N_15393,N_13835,N_13274);
nor U15394 (N_15394,N_13353,N_13393);
xnor U15395 (N_15395,N_12731,N_13855);
or U15396 (N_15396,N_12588,N_12676);
and U15397 (N_15397,N_13074,N_12123);
or U15398 (N_15398,N_13275,N_13945);
or U15399 (N_15399,N_13077,N_12813);
or U15400 (N_15400,N_13604,N_13429);
nor U15401 (N_15401,N_13131,N_13548);
and U15402 (N_15402,N_12421,N_12424);
xor U15403 (N_15403,N_12043,N_12071);
and U15404 (N_15404,N_13378,N_12913);
xnor U15405 (N_15405,N_13417,N_12264);
xor U15406 (N_15406,N_12753,N_13257);
nor U15407 (N_15407,N_12779,N_12763);
and U15408 (N_15408,N_13004,N_13055);
nand U15409 (N_15409,N_12395,N_13698);
xor U15410 (N_15410,N_12313,N_12354);
and U15411 (N_15411,N_13482,N_12795);
nor U15412 (N_15412,N_12845,N_13512);
nand U15413 (N_15413,N_12857,N_13631);
or U15414 (N_15414,N_12252,N_13328);
nand U15415 (N_15415,N_13211,N_13487);
nand U15416 (N_15416,N_12540,N_12908);
nor U15417 (N_15417,N_13564,N_13282);
or U15418 (N_15418,N_13658,N_12369);
or U15419 (N_15419,N_13393,N_12550);
nor U15420 (N_15420,N_13683,N_12466);
nor U15421 (N_15421,N_12557,N_13453);
or U15422 (N_15422,N_13848,N_12136);
or U15423 (N_15423,N_13736,N_12771);
nand U15424 (N_15424,N_13014,N_12308);
and U15425 (N_15425,N_13291,N_13173);
and U15426 (N_15426,N_13379,N_12421);
xnor U15427 (N_15427,N_12586,N_13771);
nor U15428 (N_15428,N_13701,N_13800);
nand U15429 (N_15429,N_13263,N_12259);
xnor U15430 (N_15430,N_13341,N_12928);
and U15431 (N_15431,N_12398,N_13663);
or U15432 (N_15432,N_13068,N_13875);
and U15433 (N_15433,N_13879,N_13203);
and U15434 (N_15434,N_12255,N_12736);
nor U15435 (N_15435,N_12070,N_12377);
xor U15436 (N_15436,N_13284,N_13616);
nand U15437 (N_15437,N_12286,N_13874);
and U15438 (N_15438,N_13262,N_13370);
nand U15439 (N_15439,N_13965,N_12109);
nor U15440 (N_15440,N_12349,N_12806);
and U15441 (N_15441,N_13536,N_13143);
xor U15442 (N_15442,N_13174,N_12647);
nand U15443 (N_15443,N_12106,N_12682);
and U15444 (N_15444,N_12060,N_13633);
nand U15445 (N_15445,N_12754,N_12476);
xor U15446 (N_15446,N_12093,N_12310);
or U15447 (N_15447,N_13060,N_13669);
or U15448 (N_15448,N_12681,N_13505);
xor U15449 (N_15449,N_12036,N_12819);
nand U15450 (N_15450,N_13508,N_13951);
nand U15451 (N_15451,N_12464,N_12326);
and U15452 (N_15452,N_12565,N_13444);
xnor U15453 (N_15453,N_12096,N_12563);
and U15454 (N_15454,N_12958,N_12093);
and U15455 (N_15455,N_13081,N_12242);
xor U15456 (N_15456,N_12351,N_13584);
or U15457 (N_15457,N_12494,N_12979);
and U15458 (N_15458,N_13734,N_12346);
or U15459 (N_15459,N_12562,N_13184);
nand U15460 (N_15460,N_12246,N_12131);
xor U15461 (N_15461,N_12092,N_12013);
xor U15462 (N_15462,N_12007,N_12289);
or U15463 (N_15463,N_13986,N_12759);
and U15464 (N_15464,N_12983,N_12369);
or U15465 (N_15465,N_12749,N_13228);
nand U15466 (N_15466,N_12362,N_13214);
xor U15467 (N_15467,N_12143,N_13360);
nand U15468 (N_15468,N_13066,N_13715);
xor U15469 (N_15469,N_13001,N_13391);
nand U15470 (N_15470,N_12991,N_13775);
or U15471 (N_15471,N_13331,N_12988);
nor U15472 (N_15472,N_13732,N_13104);
nand U15473 (N_15473,N_12765,N_12293);
xor U15474 (N_15474,N_13691,N_12308);
nor U15475 (N_15475,N_12601,N_12567);
xnor U15476 (N_15476,N_12316,N_12136);
and U15477 (N_15477,N_13627,N_12087);
and U15478 (N_15478,N_12809,N_12966);
nand U15479 (N_15479,N_13126,N_12293);
and U15480 (N_15480,N_13822,N_12834);
or U15481 (N_15481,N_12523,N_13342);
xnor U15482 (N_15482,N_13414,N_12934);
or U15483 (N_15483,N_12835,N_12061);
or U15484 (N_15484,N_12317,N_13576);
xnor U15485 (N_15485,N_12882,N_13754);
nor U15486 (N_15486,N_13028,N_13180);
and U15487 (N_15487,N_13692,N_13497);
and U15488 (N_15488,N_12501,N_13181);
or U15489 (N_15489,N_12459,N_13368);
nand U15490 (N_15490,N_12809,N_12838);
xnor U15491 (N_15491,N_13474,N_13785);
and U15492 (N_15492,N_13328,N_13270);
and U15493 (N_15493,N_12678,N_13296);
or U15494 (N_15494,N_12229,N_12539);
nand U15495 (N_15495,N_12187,N_12877);
nand U15496 (N_15496,N_13131,N_13281);
nand U15497 (N_15497,N_13208,N_12201);
or U15498 (N_15498,N_13972,N_12137);
nand U15499 (N_15499,N_13785,N_12934);
nand U15500 (N_15500,N_12499,N_12194);
xnor U15501 (N_15501,N_12697,N_12918);
nor U15502 (N_15502,N_12451,N_12792);
or U15503 (N_15503,N_13321,N_13998);
xor U15504 (N_15504,N_12095,N_13003);
and U15505 (N_15505,N_12897,N_12589);
and U15506 (N_15506,N_13699,N_12441);
nand U15507 (N_15507,N_13346,N_12941);
or U15508 (N_15508,N_12561,N_12724);
nor U15509 (N_15509,N_12644,N_12356);
xnor U15510 (N_15510,N_12978,N_13200);
nand U15511 (N_15511,N_13689,N_12268);
or U15512 (N_15512,N_13660,N_12624);
nor U15513 (N_15513,N_13236,N_13644);
and U15514 (N_15514,N_13683,N_12633);
nand U15515 (N_15515,N_13657,N_12950);
xnor U15516 (N_15516,N_13556,N_12634);
nor U15517 (N_15517,N_13629,N_13446);
xnor U15518 (N_15518,N_13342,N_13080);
xnor U15519 (N_15519,N_12685,N_12177);
xor U15520 (N_15520,N_12237,N_13075);
nand U15521 (N_15521,N_12660,N_13109);
nand U15522 (N_15522,N_13741,N_13454);
nor U15523 (N_15523,N_13107,N_12308);
xor U15524 (N_15524,N_12792,N_13876);
xor U15525 (N_15525,N_12539,N_12960);
nand U15526 (N_15526,N_13108,N_12851);
or U15527 (N_15527,N_12475,N_12040);
xnor U15528 (N_15528,N_12928,N_12487);
nor U15529 (N_15529,N_13530,N_13928);
xor U15530 (N_15530,N_12304,N_13653);
nor U15531 (N_15531,N_12798,N_13963);
nand U15532 (N_15532,N_13740,N_12585);
xnor U15533 (N_15533,N_12302,N_12830);
nand U15534 (N_15534,N_13554,N_13825);
nand U15535 (N_15535,N_13741,N_13354);
nand U15536 (N_15536,N_13907,N_13261);
and U15537 (N_15537,N_12652,N_12090);
nor U15538 (N_15538,N_12519,N_12882);
or U15539 (N_15539,N_12180,N_12332);
nand U15540 (N_15540,N_13067,N_12363);
and U15541 (N_15541,N_13771,N_13971);
nand U15542 (N_15542,N_13881,N_13274);
or U15543 (N_15543,N_12699,N_12212);
or U15544 (N_15544,N_12196,N_12703);
xor U15545 (N_15545,N_13821,N_13687);
nor U15546 (N_15546,N_13125,N_13498);
or U15547 (N_15547,N_12796,N_13285);
or U15548 (N_15548,N_13070,N_13558);
and U15549 (N_15549,N_12530,N_13729);
and U15550 (N_15550,N_12171,N_13553);
and U15551 (N_15551,N_12555,N_13204);
and U15552 (N_15552,N_13289,N_12817);
or U15553 (N_15553,N_13944,N_13637);
or U15554 (N_15554,N_13201,N_13886);
nor U15555 (N_15555,N_12577,N_13778);
and U15556 (N_15556,N_12127,N_13207);
nand U15557 (N_15557,N_13682,N_13149);
xor U15558 (N_15558,N_13506,N_13904);
nand U15559 (N_15559,N_12044,N_13411);
nor U15560 (N_15560,N_12085,N_13548);
or U15561 (N_15561,N_12332,N_12152);
xnor U15562 (N_15562,N_12741,N_12881);
and U15563 (N_15563,N_13570,N_13971);
nor U15564 (N_15564,N_12233,N_12017);
nor U15565 (N_15565,N_12058,N_13650);
or U15566 (N_15566,N_13862,N_13001);
and U15567 (N_15567,N_12700,N_12578);
nand U15568 (N_15568,N_13380,N_13175);
nor U15569 (N_15569,N_12769,N_13481);
nand U15570 (N_15570,N_12572,N_13187);
or U15571 (N_15571,N_12639,N_12361);
xor U15572 (N_15572,N_13929,N_12180);
or U15573 (N_15573,N_13175,N_13141);
nand U15574 (N_15574,N_12792,N_13317);
nand U15575 (N_15575,N_13740,N_12424);
nor U15576 (N_15576,N_13456,N_12051);
nand U15577 (N_15577,N_12014,N_13435);
and U15578 (N_15578,N_13817,N_12639);
nand U15579 (N_15579,N_13827,N_13465);
xnor U15580 (N_15580,N_13771,N_12706);
nand U15581 (N_15581,N_12698,N_12976);
or U15582 (N_15582,N_12937,N_13204);
and U15583 (N_15583,N_12392,N_13227);
xnor U15584 (N_15584,N_13947,N_13050);
and U15585 (N_15585,N_12426,N_13318);
nand U15586 (N_15586,N_13471,N_13016);
nor U15587 (N_15587,N_13411,N_13378);
and U15588 (N_15588,N_13067,N_13314);
xnor U15589 (N_15589,N_12496,N_13599);
or U15590 (N_15590,N_12496,N_13797);
nand U15591 (N_15591,N_12374,N_13083);
or U15592 (N_15592,N_13779,N_12377);
xor U15593 (N_15593,N_12440,N_12115);
and U15594 (N_15594,N_13267,N_13663);
nand U15595 (N_15595,N_12711,N_12363);
or U15596 (N_15596,N_13520,N_13617);
nand U15597 (N_15597,N_13427,N_12027);
nor U15598 (N_15598,N_13214,N_12785);
and U15599 (N_15599,N_13628,N_12658);
or U15600 (N_15600,N_13177,N_13086);
and U15601 (N_15601,N_12223,N_13500);
and U15602 (N_15602,N_12339,N_12616);
or U15603 (N_15603,N_12488,N_12614);
xnor U15604 (N_15604,N_12768,N_12596);
and U15605 (N_15605,N_12416,N_12848);
xor U15606 (N_15606,N_13299,N_12896);
nor U15607 (N_15607,N_12446,N_12900);
xor U15608 (N_15608,N_12245,N_12911);
or U15609 (N_15609,N_12422,N_13823);
nand U15610 (N_15610,N_12817,N_12763);
or U15611 (N_15611,N_13567,N_12299);
nand U15612 (N_15612,N_13950,N_13747);
and U15613 (N_15613,N_13696,N_12777);
or U15614 (N_15614,N_13815,N_12968);
nand U15615 (N_15615,N_13299,N_13382);
or U15616 (N_15616,N_13881,N_13816);
and U15617 (N_15617,N_12189,N_13136);
and U15618 (N_15618,N_13617,N_13402);
and U15619 (N_15619,N_12954,N_13033);
nor U15620 (N_15620,N_13608,N_13052);
or U15621 (N_15621,N_12946,N_13342);
nand U15622 (N_15622,N_12083,N_13549);
nand U15623 (N_15623,N_13152,N_12152);
nand U15624 (N_15624,N_12126,N_12039);
xnor U15625 (N_15625,N_12956,N_12999);
xnor U15626 (N_15626,N_12401,N_13764);
or U15627 (N_15627,N_13431,N_12171);
or U15628 (N_15628,N_12030,N_13894);
or U15629 (N_15629,N_12232,N_13278);
xnor U15630 (N_15630,N_13554,N_12457);
or U15631 (N_15631,N_12867,N_12640);
or U15632 (N_15632,N_13414,N_12477);
and U15633 (N_15633,N_12484,N_12703);
or U15634 (N_15634,N_13641,N_13601);
xor U15635 (N_15635,N_13794,N_13413);
and U15636 (N_15636,N_12811,N_13109);
and U15637 (N_15637,N_12200,N_12490);
and U15638 (N_15638,N_12752,N_13491);
nand U15639 (N_15639,N_13712,N_12052);
and U15640 (N_15640,N_12832,N_13226);
or U15641 (N_15641,N_13976,N_12154);
or U15642 (N_15642,N_13903,N_12770);
nor U15643 (N_15643,N_13124,N_12835);
xnor U15644 (N_15644,N_13595,N_12138);
and U15645 (N_15645,N_12181,N_13552);
and U15646 (N_15646,N_12545,N_12388);
and U15647 (N_15647,N_13031,N_12452);
nand U15648 (N_15648,N_13188,N_12009);
xnor U15649 (N_15649,N_13389,N_13743);
and U15650 (N_15650,N_12747,N_12843);
and U15651 (N_15651,N_12814,N_12824);
nor U15652 (N_15652,N_12985,N_12660);
nand U15653 (N_15653,N_13279,N_13443);
or U15654 (N_15654,N_13884,N_13939);
or U15655 (N_15655,N_13342,N_13283);
and U15656 (N_15656,N_13549,N_12640);
nor U15657 (N_15657,N_12747,N_12892);
nor U15658 (N_15658,N_13278,N_13272);
or U15659 (N_15659,N_13176,N_13501);
or U15660 (N_15660,N_13132,N_13534);
nand U15661 (N_15661,N_12125,N_12327);
and U15662 (N_15662,N_13249,N_13730);
xnor U15663 (N_15663,N_12596,N_12512);
and U15664 (N_15664,N_13008,N_13194);
and U15665 (N_15665,N_13120,N_12643);
xnor U15666 (N_15666,N_12270,N_12851);
nand U15667 (N_15667,N_12643,N_13853);
nor U15668 (N_15668,N_13720,N_13093);
and U15669 (N_15669,N_13868,N_12059);
nor U15670 (N_15670,N_13957,N_12283);
xor U15671 (N_15671,N_13323,N_12109);
and U15672 (N_15672,N_13303,N_12163);
and U15673 (N_15673,N_13109,N_12064);
and U15674 (N_15674,N_12805,N_12068);
or U15675 (N_15675,N_12833,N_12177);
nor U15676 (N_15676,N_12252,N_12996);
nand U15677 (N_15677,N_12309,N_13817);
and U15678 (N_15678,N_12196,N_12615);
nand U15679 (N_15679,N_13955,N_12040);
xnor U15680 (N_15680,N_13009,N_12961);
and U15681 (N_15681,N_12405,N_13826);
and U15682 (N_15682,N_13358,N_12846);
or U15683 (N_15683,N_13580,N_13509);
nand U15684 (N_15684,N_12237,N_12337);
and U15685 (N_15685,N_12437,N_12854);
nor U15686 (N_15686,N_12312,N_13205);
or U15687 (N_15687,N_13699,N_13034);
and U15688 (N_15688,N_12743,N_12338);
xnor U15689 (N_15689,N_12235,N_13876);
nand U15690 (N_15690,N_13323,N_13952);
nand U15691 (N_15691,N_13000,N_13051);
xor U15692 (N_15692,N_13988,N_13409);
nor U15693 (N_15693,N_12403,N_12940);
nand U15694 (N_15694,N_13174,N_13243);
nand U15695 (N_15695,N_13467,N_13892);
nand U15696 (N_15696,N_12108,N_13895);
or U15697 (N_15697,N_12534,N_13139);
or U15698 (N_15698,N_12489,N_12884);
or U15699 (N_15699,N_12785,N_13223);
nor U15700 (N_15700,N_13795,N_13191);
xor U15701 (N_15701,N_13487,N_12639);
or U15702 (N_15702,N_13614,N_12992);
and U15703 (N_15703,N_12052,N_13677);
xnor U15704 (N_15704,N_12281,N_13945);
nand U15705 (N_15705,N_12149,N_12432);
nand U15706 (N_15706,N_12739,N_13289);
nand U15707 (N_15707,N_12860,N_13851);
or U15708 (N_15708,N_12910,N_13019);
xnor U15709 (N_15709,N_12576,N_13963);
or U15710 (N_15710,N_12471,N_12749);
nor U15711 (N_15711,N_13886,N_13956);
nand U15712 (N_15712,N_12880,N_12931);
or U15713 (N_15713,N_12023,N_12634);
nand U15714 (N_15714,N_13371,N_13413);
nand U15715 (N_15715,N_12431,N_13399);
nand U15716 (N_15716,N_12413,N_13690);
nand U15717 (N_15717,N_12991,N_12813);
nor U15718 (N_15718,N_13109,N_12487);
nor U15719 (N_15719,N_13746,N_12784);
and U15720 (N_15720,N_12252,N_12757);
and U15721 (N_15721,N_12543,N_12339);
nor U15722 (N_15722,N_12894,N_12067);
or U15723 (N_15723,N_13228,N_13639);
nor U15724 (N_15724,N_13540,N_13337);
nor U15725 (N_15725,N_13883,N_12781);
or U15726 (N_15726,N_12853,N_13228);
and U15727 (N_15727,N_13537,N_13182);
or U15728 (N_15728,N_13658,N_12372);
nand U15729 (N_15729,N_12760,N_13329);
nor U15730 (N_15730,N_13222,N_13670);
nand U15731 (N_15731,N_13259,N_12727);
xnor U15732 (N_15732,N_12917,N_13504);
and U15733 (N_15733,N_13920,N_12928);
and U15734 (N_15734,N_12368,N_12768);
nor U15735 (N_15735,N_13793,N_13419);
xnor U15736 (N_15736,N_13077,N_12691);
nand U15737 (N_15737,N_12140,N_13495);
and U15738 (N_15738,N_13822,N_13142);
and U15739 (N_15739,N_12110,N_13538);
nor U15740 (N_15740,N_13018,N_13320);
and U15741 (N_15741,N_13403,N_12206);
xor U15742 (N_15742,N_13957,N_12967);
xnor U15743 (N_15743,N_12701,N_13617);
or U15744 (N_15744,N_13330,N_12351);
nand U15745 (N_15745,N_13973,N_12435);
nor U15746 (N_15746,N_13697,N_13959);
xnor U15747 (N_15747,N_12458,N_13150);
xnor U15748 (N_15748,N_12674,N_13392);
and U15749 (N_15749,N_12085,N_13547);
xnor U15750 (N_15750,N_12349,N_13413);
xnor U15751 (N_15751,N_13069,N_13963);
and U15752 (N_15752,N_13412,N_13190);
xor U15753 (N_15753,N_13872,N_12712);
or U15754 (N_15754,N_13647,N_12231);
nand U15755 (N_15755,N_12548,N_12590);
nor U15756 (N_15756,N_12426,N_12441);
or U15757 (N_15757,N_13670,N_12665);
nor U15758 (N_15758,N_13163,N_12396);
nand U15759 (N_15759,N_12002,N_12582);
nor U15760 (N_15760,N_13892,N_12034);
nand U15761 (N_15761,N_13712,N_12909);
nor U15762 (N_15762,N_13105,N_12657);
and U15763 (N_15763,N_12158,N_13204);
xor U15764 (N_15764,N_12378,N_13145);
nand U15765 (N_15765,N_13468,N_12157);
xnor U15766 (N_15766,N_13347,N_13611);
or U15767 (N_15767,N_12610,N_12114);
and U15768 (N_15768,N_12850,N_12061);
xnor U15769 (N_15769,N_12478,N_13104);
and U15770 (N_15770,N_13629,N_12182);
nor U15771 (N_15771,N_13188,N_12915);
or U15772 (N_15772,N_12986,N_13817);
nor U15773 (N_15773,N_13670,N_12377);
nand U15774 (N_15774,N_12132,N_13854);
and U15775 (N_15775,N_12181,N_13053);
xor U15776 (N_15776,N_12656,N_12671);
or U15777 (N_15777,N_12002,N_12779);
nand U15778 (N_15778,N_12603,N_13522);
and U15779 (N_15779,N_12281,N_13638);
or U15780 (N_15780,N_13387,N_12782);
and U15781 (N_15781,N_13925,N_12602);
xor U15782 (N_15782,N_13131,N_13850);
or U15783 (N_15783,N_12225,N_12187);
or U15784 (N_15784,N_12040,N_13030);
or U15785 (N_15785,N_12072,N_12796);
xor U15786 (N_15786,N_13329,N_13497);
or U15787 (N_15787,N_12479,N_12177);
nand U15788 (N_15788,N_12520,N_13408);
nand U15789 (N_15789,N_12848,N_13472);
and U15790 (N_15790,N_13703,N_12864);
nor U15791 (N_15791,N_12793,N_13970);
and U15792 (N_15792,N_12897,N_12892);
xor U15793 (N_15793,N_12517,N_13886);
xor U15794 (N_15794,N_13457,N_12432);
xor U15795 (N_15795,N_12284,N_13688);
nand U15796 (N_15796,N_13168,N_12927);
and U15797 (N_15797,N_13764,N_12112);
xnor U15798 (N_15798,N_13118,N_12960);
and U15799 (N_15799,N_12373,N_12998);
and U15800 (N_15800,N_12074,N_13267);
and U15801 (N_15801,N_12435,N_13658);
nand U15802 (N_15802,N_13652,N_12693);
xnor U15803 (N_15803,N_13145,N_12676);
and U15804 (N_15804,N_13116,N_12966);
nand U15805 (N_15805,N_13884,N_13110);
nor U15806 (N_15806,N_13442,N_12604);
nand U15807 (N_15807,N_12650,N_13677);
or U15808 (N_15808,N_13791,N_13180);
nand U15809 (N_15809,N_13170,N_13756);
or U15810 (N_15810,N_13394,N_13762);
nor U15811 (N_15811,N_13051,N_13948);
nor U15812 (N_15812,N_13224,N_12806);
nand U15813 (N_15813,N_13979,N_12819);
and U15814 (N_15814,N_12168,N_12346);
or U15815 (N_15815,N_12122,N_13074);
and U15816 (N_15816,N_13947,N_12323);
or U15817 (N_15817,N_12181,N_13579);
and U15818 (N_15818,N_13301,N_13322);
xnor U15819 (N_15819,N_13043,N_13142);
xnor U15820 (N_15820,N_13118,N_13207);
or U15821 (N_15821,N_12585,N_12329);
nor U15822 (N_15822,N_12820,N_13004);
and U15823 (N_15823,N_13228,N_13010);
nand U15824 (N_15824,N_12756,N_12351);
nand U15825 (N_15825,N_12317,N_12388);
and U15826 (N_15826,N_12801,N_13824);
xor U15827 (N_15827,N_13890,N_12319);
xor U15828 (N_15828,N_12098,N_12514);
or U15829 (N_15829,N_13595,N_13201);
nor U15830 (N_15830,N_13101,N_13450);
xor U15831 (N_15831,N_12866,N_13474);
and U15832 (N_15832,N_13654,N_13166);
nand U15833 (N_15833,N_13006,N_13371);
or U15834 (N_15834,N_13680,N_13489);
or U15835 (N_15835,N_13881,N_13932);
nand U15836 (N_15836,N_13424,N_12089);
nand U15837 (N_15837,N_13747,N_13860);
nor U15838 (N_15838,N_12829,N_12640);
xor U15839 (N_15839,N_13672,N_13452);
or U15840 (N_15840,N_13173,N_13642);
or U15841 (N_15841,N_12342,N_13052);
nor U15842 (N_15842,N_12878,N_12003);
xor U15843 (N_15843,N_13023,N_13768);
nand U15844 (N_15844,N_12844,N_13089);
xnor U15845 (N_15845,N_13325,N_12943);
nand U15846 (N_15846,N_12043,N_13167);
or U15847 (N_15847,N_13418,N_12464);
or U15848 (N_15848,N_13755,N_12483);
and U15849 (N_15849,N_12027,N_13851);
nor U15850 (N_15850,N_12716,N_13718);
or U15851 (N_15851,N_12342,N_12860);
nor U15852 (N_15852,N_13290,N_12668);
or U15853 (N_15853,N_12782,N_13475);
nand U15854 (N_15854,N_12529,N_13568);
xnor U15855 (N_15855,N_13067,N_13168);
and U15856 (N_15856,N_12618,N_12946);
and U15857 (N_15857,N_12330,N_13582);
nand U15858 (N_15858,N_13954,N_12911);
nor U15859 (N_15859,N_12204,N_13044);
nor U15860 (N_15860,N_12705,N_12228);
nor U15861 (N_15861,N_13765,N_13057);
and U15862 (N_15862,N_13805,N_13299);
nand U15863 (N_15863,N_13706,N_13408);
xor U15864 (N_15864,N_12646,N_12077);
nand U15865 (N_15865,N_12656,N_12191);
nand U15866 (N_15866,N_12919,N_12707);
xor U15867 (N_15867,N_12540,N_12299);
xor U15868 (N_15868,N_13835,N_12054);
and U15869 (N_15869,N_12884,N_13736);
and U15870 (N_15870,N_13660,N_12256);
nor U15871 (N_15871,N_13998,N_13094);
nand U15872 (N_15872,N_12905,N_12333);
and U15873 (N_15873,N_12233,N_13347);
xor U15874 (N_15874,N_13379,N_12817);
xor U15875 (N_15875,N_12670,N_13587);
nor U15876 (N_15876,N_13441,N_12670);
xor U15877 (N_15877,N_12703,N_12285);
and U15878 (N_15878,N_13366,N_12984);
or U15879 (N_15879,N_13200,N_12492);
nor U15880 (N_15880,N_13564,N_12149);
nand U15881 (N_15881,N_13738,N_13429);
or U15882 (N_15882,N_13786,N_13333);
xnor U15883 (N_15883,N_12035,N_12634);
xor U15884 (N_15884,N_13314,N_13858);
xor U15885 (N_15885,N_12679,N_13353);
xnor U15886 (N_15886,N_12553,N_13712);
nor U15887 (N_15887,N_13305,N_13109);
and U15888 (N_15888,N_13196,N_13455);
nor U15889 (N_15889,N_13455,N_12810);
xnor U15890 (N_15890,N_12560,N_12366);
and U15891 (N_15891,N_12275,N_13871);
and U15892 (N_15892,N_12526,N_13888);
and U15893 (N_15893,N_13859,N_13845);
nor U15894 (N_15894,N_13093,N_13541);
nor U15895 (N_15895,N_12525,N_12997);
xor U15896 (N_15896,N_13987,N_13966);
or U15897 (N_15897,N_13020,N_13861);
nand U15898 (N_15898,N_12453,N_12256);
nor U15899 (N_15899,N_12914,N_12169);
and U15900 (N_15900,N_13863,N_13078);
and U15901 (N_15901,N_12616,N_13088);
or U15902 (N_15902,N_13154,N_12830);
or U15903 (N_15903,N_13521,N_12216);
or U15904 (N_15904,N_13101,N_12382);
xor U15905 (N_15905,N_12363,N_12715);
xnor U15906 (N_15906,N_13376,N_13016);
and U15907 (N_15907,N_12151,N_13874);
or U15908 (N_15908,N_13706,N_12108);
nand U15909 (N_15909,N_13340,N_13513);
xnor U15910 (N_15910,N_12023,N_13378);
and U15911 (N_15911,N_13693,N_13080);
xor U15912 (N_15912,N_13299,N_12239);
nor U15913 (N_15913,N_13641,N_12146);
or U15914 (N_15914,N_13555,N_13140);
xor U15915 (N_15915,N_13540,N_12033);
xor U15916 (N_15916,N_12673,N_13227);
nand U15917 (N_15917,N_13312,N_12013);
or U15918 (N_15918,N_12376,N_13504);
nand U15919 (N_15919,N_13231,N_13865);
nor U15920 (N_15920,N_12217,N_13678);
nand U15921 (N_15921,N_13245,N_13102);
or U15922 (N_15922,N_13161,N_12955);
nor U15923 (N_15923,N_13873,N_13036);
nor U15924 (N_15924,N_13495,N_12283);
nand U15925 (N_15925,N_12210,N_12083);
xnor U15926 (N_15926,N_12275,N_12646);
nor U15927 (N_15927,N_12306,N_12361);
or U15928 (N_15928,N_13400,N_13891);
and U15929 (N_15929,N_13407,N_12321);
nor U15930 (N_15930,N_13629,N_13391);
or U15931 (N_15931,N_13308,N_12716);
or U15932 (N_15932,N_12870,N_12369);
nand U15933 (N_15933,N_12163,N_12970);
xor U15934 (N_15934,N_13664,N_13781);
and U15935 (N_15935,N_12207,N_13732);
and U15936 (N_15936,N_13308,N_12450);
nor U15937 (N_15937,N_13643,N_13436);
nand U15938 (N_15938,N_12796,N_13491);
xor U15939 (N_15939,N_13135,N_12561);
and U15940 (N_15940,N_13948,N_13012);
or U15941 (N_15941,N_12132,N_13749);
nor U15942 (N_15942,N_13255,N_13167);
xor U15943 (N_15943,N_13395,N_12090);
nand U15944 (N_15944,N_12196,N_13015);
nand U15945 (N_15945,N_13043,N_13452);
nor U15946 (N_15946,N_13407,N_12481);
or U15947 (N_15947,N_13919,N_13412);
nor U15948 (N_15948,N_13058,N_12828);
xor U15949 (N_15949,N_13241,N_13907);
and U15950 (N_15950,N_13327,N_12871);
and U15951 (N_15951,N_13977,N_12238);
and U15952 (N_15952,N_12609,N_13045);
xnor U15953 (N_15953,N_12581,N_12245);
nand U15954 (N_15954,N_13339,N_13301);
xnor U15955 (N_15955,N_12733,N_12586);
and U15956 (N_15956,N_12073,N_12737);
and U15957 (N_15957,N_12281,N_12392);
nor U15958 (N_15958,N_12572,N_13404);
or U15959 (N_15959,N_12076,N_13586);
nand U15960 (N_15960,N_13298,N_13982);
and U15961 (N_15961,N_12294,N_12292);
nor U15962 (N_15962,N_13393,N_13089);
nor U15963 (N_15963,N_12366,N_12030);
or U15964 (N_15964,N_12628,N_13469);
or U15965 (N_15965,N_13956,N_12134);
xnor U15966 (N_15966,N_13031,N_13035);
nand U15967 (N_15967,N_12533,N_12226);
xnor U15968 (N_15968,N_13082,N_13726);
nand U15969 (N_15969,N_13866,N_12126);
and U15970 (N_15970,N_13094,N_13735);
and U15971 (N_15971,N_13367,N_12872);
and U15972 (N_15972,N_13352,N_12835);
nand U15973 (N_15973,N_12987,N_13755);
xor U15974 (N_15974,N_13894,N_13944);
or U15975 (N_15975,N_13873,N_12374);
nor U15976 (N_15976,N_13881,N_12759);
and U15977 (N_15977,N_12735,N_12488);
or U15978 (N_15978,N_13680,N_13557);
nand U15979 (N_15979,N_13743,N_13520);
or U15980 (N_15980,N_13827,N_12499);
or U15981 (N_15981,N_13686,N_12795);
xor U15982 (N_15982,N_13925,N_12647);
xnor U15983 (N_15983,N_12900,N_12178);
and U15984 (N_15984,N_12266,N_12564);
xor U15985 (N_15985,N_13378,N_12131);
or U15986 (N_15986,N_12893,N_13445);
nor U15987 (N_15987,N_13890,N_12717);
nand U15988 (N_15988,N_13722,N_13145);
or U15989 (N_15989,N_12995,N_13820);
and U15990 (N_15990,N_13805,N_12971);
and U15991 (N_15991,N_12426,N_13911);
xnor U15992 (N_15992,N_12432,N_12465);
and U15993 (N_15993,N_12681,N_12750);
nand U15994 (N_15994,N_13378,N_13856);
nand U15995 (N_15995,N_12846,N_12606);
and U15996 (N_15996,N_12977,N_12113);
xor U15997 (N_15997,N_12896,N_12557);
nand U15998 (N_15998,N_12001,N_12537);
and U15999 (N_15999,N_12898,N_12762);
xor U16000 (N_16000,N_14623,N_15550);
or U16001 (N_16001,N_14521,N_14838);
or U16002 (N_16002,N_14015,N_14556);
or U16003 (N_16003,N_14708,N_15791);
and U16004 (N_16004,N_14898,N_15307);
or U16005 (N_16005,N_15914,N_14505);
xnor U16006 (N_16006,N_15235,N_14850);
xnor U16007 (N_16007,N_15176,N_14735);
nor U16008 (N_16008,N_14224,N_15023);
and U16009 (N_16009,N_15941,N_14226);
nor U16010 (N_16010,N_15872,N_14084);
and U16011 (N_16011,N_15196,N_14785);
or U16012 (N_16012,N_15219,N_15802);
and U16013 (N_16013,N_15835,N_15597);
or U16014 (N_16014,N_15614,N_15027);
nand U16015 (N_16015,N_15447,N_15549);
nor U16016 (N_16016,N_14570,N_15841);
nor U16017 (N_16017,N_14789,N_14345);
and U16018 (N_16018,N_15243,N_14208);
and U16019 (N_16019,N_14327,N_15092);
or U16020 (N_16020,N_15789,N_15364);
xor U16021 (N_16021,N_15168,N_14925);
nor U16022 (N_16022,N_15800,N_14494);
xnor U16023 (N_16023,N_15359,N_14605);
nor U16024 (N_16024,N_15014,N_14949);
nand U16025 (N_16025,N_15151,N_15683);
or U16026 (N_16026,N_14389,N_15652);
nor U16027 (N_16027,N_14752,N_14739);
or U16028 (N_16028,N_15001,N_14315);
or U16029 (N_16029,N_14852,N_14006);
nand U16030 (N_16030,N_15996,N_15101);
or U16031 (N_16031,N_15177,N_14042);
xnor U16032 (N_16032,N_15838,N_15230);
or U16033 (N_16033,N_14741,N_14927);
or U16034 (N_16034,N_14929,N_14894);
nor U16035 (N_16035,N_14507,N_14943);
nand U16036 (N_16036,N_14397,N_14981);
and U16037 (N_16037,N_14629,N_14816);
xor U16038 (N_16038,N_15118,N_14294);
nand U16039 (N_16039,N_14278,N_14732);
and U16040 (N_16040,N_14303,N_15312);
nor U16041 (N_16041,N_14583,N_14827);
xnor U16042 (N_16042,N_15329,N_15391);
and U16043 (N_16043,N_14447,N_14098);
xnor U16044 (N_16044,N_14300,N_15668);
nor U16045 (N_16045,N_14237,N_14119);
xor U16046 (N_16046,N_15541,N_14384);
and U16047 (N_16047,N_14870,N_15911);
or U16048 (N_16048,N_15333,N_14390);
and U16049 (N_16049,N_15191,N_14823);
nor U16050 (N_16050,N_15565,N_14259);
nor U16051 (N_16051,N_14691,N_15755);
and U16052 (N_16052,N_15165,N_15068);
and U16053 (N_16053,N_15041,N_14211);
xnor U16054 (N_16054,N_14436,N_15891);
or U16055 (N_16055,N_14087,N_14256);
or U16056 (N_16056,N_15639,N_14736);
and U16057 (N_16057,N_15873,N_14808);
or U16058 (N_16058,N_14292,N_15904);
or U16059 (N_16059,N_15558,N_15090);
or U16060 (N_16060,N_15782,N_14562);
xor U16061 (N_16061,N_14887,N_15519);
and U16062 (N_16062,N_14698,N_14148);
or U16063 (N_16063,N_15610,N_14221);
and U16064 (N_16064,N_14320,N_14817);
or U16065 (N_16065,N_15984,N_14670);
or U16066 (N_16066,N_15384,N_15464);
and U16067 (N_16067,N_14968,N_15407);
nand U16068 (N_16068,N_14257,N_15170);
xnor U16069 (N_16069,N_14932,N_14241);
xor U16070 (N_16070,N_14486,N_14339);
xnor U16071 (N_16071,N_15578,N_15819);
and U16072 (N_16072,N_14988,N_14767);
and U16073 (N_16073,N_15640,N_14975);
and U16074 (N_16074,N_15035,N_15267);
xnor U16075 (N_16075,N_14888,N_15255);
or U16076 (N_16076,N_15822,N_14859);
or U16077 (N_16077,N_14040,N_15404);
or U16078 (N_16078,N_14642,N_14343);
and U16079 (N_16079,N_15448,N_15069);
xor U16080 (N_16080,N_15964,N_14409);
xnor U16081 (N_16081,N_14464,N_14810);
or U16082 (N_16082,N_15415,N_14719);
and U16083 (N_16083,N_14703,N_15539);
nor U16084 (N_16084,N_15326,N_15145);
or U16085 (N_16085,N_15479,N_15829);
or U16086 (N_16086,N_14172,N_14529);
or U16087 (N_16087,N_14867,N_14000);
nor U16088 (N_16088,N_14655,N_15757);
xor U16089 (N_16089,N_14854,N_15394);
nand U16090 (N_16090,N_14373,N_15222);
or U16091 (N_16091,N_15074,N_15022);
or U16092 (N_16092,N_14588,N_15313);
and U16093 (N_16093,N_14560,N_15294);
xor U16094 (N_16094,N_14701,N_15544);
nand U16095 (N_16095,N_14768,N_15306);
xnor U16096 (N_16096,N_15225,N_15982);
xnor U16097 (N_16097,N_15923,N_15559);
xor U16098 (N_16098,N_15005,N_14531);
and U16099 (N_16099,N_14990,N_14095);
nor U16100 (N_16100,N_14037,N_15143);
or U16101 (N_16101,N_15778,N_15402);
and U16102 (N_16102,N_14206,N_15707);
and U16103 (N_16103,N_14500,N_14950);
xnor U16104 (N_16104,N_14820,N_15908);
nor U16105 (N_16105,N_14019,N_14763);
and U16106 (N_16106,N_15254,N_15481);
nor U16107 (N_16107,N_15477,N_15528);
and U16108 (N_16108,N_14902,N_15799);
and U16109 (N_16109,N_15180,N_15855);
xor U16110 (N_16110,N_14731,N_15038);
xor U16111 (N_16111,N_14794,N_14082);
nand U16112 (N_16112,N_14075,N_15399);
nor U16113 (N_16113,N_14566,N_15651);
or U16114 (N_16114,N_15928,N_14967);
xnor U16115 (N_16115,N_14352,N_15379);
and U16116 (N_16116,N_14871,N_15521);
nand U16117 (N_16117,N_15042,N_14607);
or U16118 (N_16118,N_14126,N_15874);
nand U16119 (N_16119,N_14836,N_15737);
xnor U16120 (N_16120,N_15787,N_14393);
nor U16121 (N_16121,N_15728,N_15796);
xor U16122 (N_16122,N_15317,N_14717);
nor U16123 (N_16123,N_15451,N_14745);
nor U16124 (N_16124,N_14355,N_14506);
and U16125 (N_16125,N_15825,N_14749);
nor U16126 (N_16126,N_14465,N_15608);
or U16127 (N_16127,N_15513,N_15190);
nand U16128 (N_16128,N_15771,N_15609);
and U16129 (N_16129,N_14460,N_15797);
nor U16130 (N_16130,N_15248,N_15357);
nor U16131 (N_16131,N_14142,N_14830);
and U16132 (N_16132,N_14041,N_14919);
or U16133 (N_16133,N_14485,N_15476);
xnor U16134 (N_16134,N_15950,N_15435);
nor U16135 (N_16135,N_14323,N_15154);
or U16136 (N_16136,N_15163,N_15779);
xor U16137 (N_16137,N_15089,N_14157);
nor U16138 (N_16138,N_14534,N_14600);
or U16139 (N_16139,N_14127,N_15434);
and U16140 (N_16140,N_15518,N_15221);
nor U16141 (N_16141,N_14565,N_15161);
nand U16142 (N_16142,N_14350,N_14723);
xnor U16143 (N_16143,N_14262,N_15381);
nor U16144 (N_16144,N_14603,N_15334);
and U16145 (N_16145,N_15512,N_15113);
and U16146 (N_16146,N_14367,N_15320);
xnor U16147 (N_16147,N_14601,N_15625);
and U16148 (N_16148,N_15656,N_15722);
nor U16149 (N_16149,N_14059,N_14673);
nand U16150 (N_16150,N_14772,N_14503);
and U16151 (N_16151,N_14400,N_15700);
nor U16152 (N_16152,N_15929,N_14223);
nand U16153 (N_16153,N_15805,N_15785);
nand U16154 (N_16154,N_14415,N_15783);
nand U16155 (N_16155,N_14689,N_15413);
xor U16156 (N_16156,N_15837,N_15875);
and U16157 (N_16157,N_15818,N_14989);
nor U16158 (N_16158,N_15416,N_15523);
nand U16159 (N_16159,N_14276,N_14387);
nand U16160 (N_16160,N_14564,N_14143);
and U16161 (N_16161,N_15581,N_14614);
and U16162 (N_16162,N_14769,N_14942);
xnor U16163 (N_16163,N_14751,N_14840);
xnor U16164 (N_16164,N_15252,N_15378);
or U16165 (N_16165,N_15985,N_14442);
or U16166 (N_16166,N_14302,N_15446);
or U16167 (N_16167,N_14742,N_15946);
and U16168 (N_16168,N_15004,N_15637);
and U16169 (N_16169,N_14044,N_14755);
and U16170 (N_16170,N_14330,N_15450);
nand U16171 (N_16171,N_14429,N_15099);
nand U16172 (N_16172,N_15775,N_15536);
nand U16173 (N_16173,N_14790,N_14250);
or U16174 (N_16174,N_15650,N_15573);
xnor U16175 (N_16175,N_14192,N_15696);
nor U16176 (N_16176,N_14579,N_15355);
or U16177 (N_16177,N_14010,N_15529);
nor U16178 (N_16178,N_14586,N_15987);
xnor U16179 (N_16179,N_14504,N_15495);
nor U16180 (N_16180,N_14585,N_15804);
xor U16181 (N_16181,N_14449,N_15178);
xor U16182 (N_16182,N_14285,N_15265);
nor U16183 (N_16183,N_15406,N_14002);
and U16184 (N_16184,N_14648,N_15286);
and U16185 (N_16185,N_15957,N_15989);
or U16186 (N_16186,N_14162,N_15643);
and U16187 (N_16187,N_15365,N_14283);
and U16188 (N_16188,N_15932,N_14592);
or U16189 (N_16189,N_15842,N_15944);
and U16190 (N_16190,N_14083,N_14552);
and U16191 (N_16191,N_14108,N_14619);
or U16192 (N_16192,N_14471,N_15232);
or U16193 (N_16193,N_14166,N_14379);
nor U16194 (N_16194,N_15462,N_15882);
or U16195 (N_16195,N_14631,N_15098);
or U16196 (N_16196,N_14261,N_14185);
or U16197 (N_16197,N_15997,N_15492);
xor U16198 (N_16198,N_15863,N_15955);
or U16199 (N_16199,N_14814,N_15893);
and U16200 (N_16200,N_14864,N_14092);
xnor U16201 (N_16201,N_14284,N_15183);
or U16202 (N_16202,N_14225,N_15515);
nor U16203 (N_16203,N_14425,N_14604);
and U16204 (N_16204,N_15621,N_15999);
nor U16205 (N_16205,N_15684,N_15403);
or U16206 (N_16206,N_15272,N_15965);
xor U16207 (N_16207,N_15150,N_14744);
or U16208 (N_16208,N_15345,N_15776);
nor U16209 (N_16209,N_14011,N_14457);
nand U16210 (N_16210,N_14883,N_14826);
nor U16211 (N_16211,N_15292,N_14641);
nand U16212 (N_16212,N_14740,N_14258);
or U16213 (N_16213,N_14331,N_14365);
nor U16214 (N_16214,N_14175,N_14363);
or U16215 (N_16215,N_15121,N_15681);
nor U16216 (N_16216,N_15120,N_14117);
nand U16217 (N_16217,N_14154,N_15769);
and U16218 (N_16218,N_15352,N_14813);
nor U16219 (N_16219,N_14617,N_15314);
or U16220 (N_16220,N_14882,N_15566);
and U16221 (N_16221,N_14061,N_14178);
or U16222 (N_16222,N_15386,N_15777);
nor U16223 (N_16223,N_14984,N_14351);
xor U16224 (N_16224,N_15302,N_15432);
nor U16225 (N_16225,N_14128,N_14892);
nand U16226 (N_16226,N_15046,N_14626);
or U16227 (N_16227,N_15241,N_14359);
xor U16228 (N_16228,N_15820,N_15714);
nor U16229 (N_16229,N_14797,N_14637);
nand U16230 (N_16230,N_14780,N_14891);
xor U16231 (N_16231,N_15052,N_15043);
nand U16232 (N_16232,N_14347,N_15290);
xnor U16233 (N_16233,N_15361,N_15615);
nand U16234 (N_16234,N_15439,N_14134);
xnor U16235 (N_16235,N_15546,N_14805);
and U16236 (N_16236,N_14133,N_14665);
nand U16237 (N_16237,N_14299,N_14458);
nor U16238 (N_16238,N_14841,N_14640);
and U16239 (N_16239,N_14973,N_15613);
nor U16240 (N_16240,N_14383,N_14498);
xor U16241 (N_16241,N_15367,N_15634);
or U16242 (N_16242,N_15438,N_14115);
nand U16243 (N_16243,N_15973,N_14992);
xor U16244 (N_16244,N_14634,N_15542);
and U16245 (N_16245,N_15327,N_15057);
nand U16246 (N_16246,N_15605,N_14706);
nor U16247 (N_16247,N_14649,N_15720);
nor U16248 (N_16248,N_15694,N_15452);
and U16249 (N_16249,N_14856,N_15134);
and U16250 (N_16250,N_14636,N_14957);
xnor U16251 (N_16251,N_15482,N_14606);
nand U16252 (N_16252,N_15516,N_14497);
nor U16253 (N_16253,N_14169,N_14613);
or U16254 (N_16254,N_15470,N_15461);
or U16255 (N_16255,N_15736,N_15358);
nand U16256 (N_16256,N_15039,N_14100);
and U16257 (N_16257,N_15580,N_15507);
nor U16258 (N_16258,N_15260,N_14775);
nand U16259 (N_16259,N_15018,N_15500);
nor U16260 (N_16260,N_14356,N_14110);
or U16261 (N_16261,N_15490,N_14954);
or U16262 (N_16262,N_15952,N_15902);
xor U16263 (N_16263,N_14269,N_14150);
xnor U16264 (N_16264,N_15679,N_14478);
nand U16265 (N_16265,N_14322,N_15008);
or U16266 (N_16266,N_14496,N_14035);
nand U16267 (N_16267,N_14987,N_14252);
and U16268 (N_16268,N_14516,N_15733);
and U16269 (N_16269,N_14274,N_14783);
or U16270 (N_16270,N_15037,N_14155);
and U16271 (N_16271,N_14316,N_15295);
nor U16272 (N_16272,N_15934,N_14120);
nand U16273 (N_16273,N_14526,N_14822);
nand U16274 (N_16274,N_15075,N_15132);
or U16275 (N_16275,N_14027,N_14419);
and U16276 (N_16276,N_15535,N_14054);
nor U16277 (N_16277,N_15383,N_14366);
and U16278 (N_16278,N_15199,N_15278);
nand U16279 (N_16279,N_15554,N_14369);
and U16280 (N_16280,N_14554,N_15641);
nor U16281 (N_16281,N_15764,N_15044);
nor U16282 (N_16282,N_14832,N_14595);
and U16283 (N_16283,N_14156,N_15473);
or U16284 (N_16284,N_15362,N_14525);
or U16285 (N_16285,N_14624,N_14945);
nor U16286 (N_16286,N_14561,N_15200);
nor U16287 (N_16287,N_15620,N_14053);
or U16288 (N_16288,N_15724,N_14812);
or U16289 (N_16289,N_14212,N_15187);
or U16290 (N_16290,N_15878,N_15856);
or U16291 (N_16291,N_14238,N_15095);
nand U16292 (N_16292,N_14833,N_15892);
nor U16293 (N_16293,N_15685,N_15316);
xor U16294 (N_16294,N_15033,N_15382);
nor U16295 (N_16295,N_15017,N_15747);
xor U16296 (N_16296,N_14646,N_14482);
and U16297 (N_16297,N_14946,N_14334);
nor U16298 (N_16298,N_14545,N_14970);
nand U16299 (N_16299,N_15305,N_15116);
and U16300 (N_16300,N_15472,N_14675);
xnor U16301 (N_16301,N_14375,N_15560);
or U16302 (N_16302,N_14268,N_14845);
xor U16303 (N_16303,N_15171,N_14936);
nand U16304 (N_16304,N_15644,N_15029);
xnor U16305 (N_16305,N_15138,N_14983);
xor U16306 (N_16306,N_14718,N_15971);
xor U16307 (N_16307,N_15746,N_15576);
nand U16308 (N_16308,N_14911,N_15377);
nor U16309 (N_16309,N_15545,N_14802);
and U16310 (N_16310,N_14978,N_15555);
nand U16311 (N_16311,N_15096,N_14074);
and U16312 (N_16312,N_14272,N_15082);
nor U16313 (N_16313,N_15725,N_14112);
nand U16314 (N_16314,N_14743,N_15489);
or U16315 (N_16315,N_15649,N_15488);
and U16316 (N_16316,N_15890,N_14851);
or U16317 (N_16317,N_14240,N_15175);
nand U16318 (N_16318,N_14395,N_15976);
or U16319 (N_16319,N_14441,N_14884);
xor U16320 (N_16320,N_15795,N_15711);
or U16321 (N_16321,N_15400,N_15259);
nand U16322 (N_16322,N_15673,N_15061);
nor U16323 (N_16323,N_14063,N_15894);
and U16324 (N_16324,N_14265,N_15678);
and U16325 (N_16325,N_14874,N_14993);
and U16326 (N_16326,N_15296,N_15013);
xnor U16327 (N_16327,N_15790,N_14941);
xor U16328 (N_16328,N_15215,N_15126);
nand U16329 (N_16329,N_15596,N_14944);
nor U16330 (N_16330,N_15885,N_15048);
nand U16331 (N_16331,N_14553,N_14530);
nor U16332 (N_16332,N_14182,N_15066);
nor U16333 (N_16333,N_15072,N_14523);
or U16334 (N_16334,N_15859,N_15318);
nor U16335 (N_16335,N_15496,N_14349);
nand U16336 (N_16336,N_14492,N_15664);
or U16337 (N_16337,N_14860,N_14293);
xor U16338 (N_16338,N_15223,N_14620);
or U16339 (N_16339,N_15677,N_15209);
xor U16340 (N_16340,N_14408,N_15194);
nand U16341 (N_16341,N_14979,N_14661);
xor U16342 (N_16342,N_15437,N_14446);
nor U16343 (N_16343,N_15374,N_14920);
nor U16344 (N_16344,N_15823,N_15718);
or U16345 (N_16345,N_15672,N_14414);
xnor U16346 (N_16346,N_14904,N_15988);
or U16347 (N_16347,N_15245,N_15030);
xor U16348 (N_16348,N_14519,N_14760);
nand U16349 (N_16349,N_14167,N_15360);
and U16350 (N_16350,N_15181,N_14628);
xor U16351 (N_16351,N_15195,N_15508);
nor U16352 (N_16352,N_14179,N_14536);
and U16353 (N_16353,N_15563,N_14829);
or U16354 (N_16354,N_14145,N_15285);
or U16355 (N_16355,N_14109,N_15784);
nand U16356 (N_16356,N_14219,N_15561);
xor U16357 (N_16357,N_15593,N_15173);
or U16358 (N_16358,N_14779,N_14372);
and U16359 (N_16359,N_15993,N_14914);
nor U16360 (N_16360,N_14287,N_15808);
or U16361 (N_16361,N_15397,N_14078);
xnor U16362 (N_16362,N_15655,N_14499);
or U16363 (N_16363,N_15275,N_15137);
xor U16364 (N_16364,N_15063,N_15433);
and U16365 (N_16365,N_15671,N_14513);
and U16366 (N_16366,N_15021,N_14515);
nor U16367 (N_16367,N_14958,N_14404);
nor U16368 (N_16368,N_15310,N_15938);
or U16369 (N_16369,N_15412,N_14924);
xnor U16370 (N_16370,N_15207,N_15642);
xor U16371 (N_16371,N_14277,N_14643);
nor U16372 (N_16372,N_15411,N_15526);
nor U16373 (N_16373,N_14216,N_15564);
xor U16374 (N_16374,N_14026,N_15141);
nand U16375 (N_16375,N_15760,N_15459);
xor U16376 (N_16376,N_15011,N_15826);
nor U16377 (N_16377,N_15401,N_14454);
xor U16378 (N_16378,N_14558,N_15761);
or U16379 (N_16379,N_14312,N_14342);
or U16380 (N_16380,N_14424,N_15675);
xor U16381 (N_16381,N_14213,N_14985);
nor U16382 (N_16382,N_14125,N_14897);
nor U16383 (N_16383,N_15570,N_14451);
xor U16384 (N_16384,N_14076,N_14638);
nand U16385 (N_16385,N_15497,N_15547);
nand U16386 (N_16386,N_15309,N_14848);
xnor U16387 (N_16387,N_15587,N_15436);
or U16388 (N_16388,N_14239,N_15060);
and U16389 (N_16389,N_15786,N_14472);
nand U16390 (N_16390,N_15870,N_14587);
nand U16391 (N_16391,N_15522,N_15801);
xor U16392 (N_16392,N_14774,N_14430);
nor U16393 (N_16393,N_15636,N_14090);
nor U16394 (N_16394,N_14459,N_14444);
nand U16395 (N_16395,N_14996,N_14544);
and U16396 (N_16396,N_14378,N_14502);
xor U16397 (N_16397,N_15686,N_14060);
or U16398 (N_16398,N_14227,N_15741);
nand U16399 (N_16399,N_14580,N_14008);
nor U16400 (N_16400,N_15167,N_14466);
or U16401 (N_16401,N_15336,N_14692);
xnor U16402 (N_16402,N_15136,N_14876);
and U16403 (N_16403,N_15595,N_15107);
nand U16404 (N_16404,N_15097,N_15146);
nand U16405 (N_16405,N_15626,N_14190);
nor U16406 (N_16406,N_14467,N_15380);
nand U16407 (N_16407,N_15426,N_15453);
nor U16408 (N_16408,N_15884,N_15117);
nand U16409 (N_16409,N_14361,N_14462);
and U16410 (N_16410,N_14686,N_14886);
and U16411 (N_16411,N_15592,N_14056);
and U16412 (N_16412,N_14693,N_14140);
nor U16413 (N_16413,N_15846,N_14475);
xnor U16414 (N_16414,N_15140,N_14955);
and U16415 (N_16415,N_14687,N_15727);
xor U16416 (N_16416,N_15688,N_15133);
nor U16417 (N_16417,N_14030,N_14057);
xor U16418 (N_16418,N_15674,N_14308);
and U16419 (N_16419,N_15645,N_14158);
and U16420 (N_16420,N_14807,N_15659);
or U16421 (N_16421,N_14131,N_14847);
nand U16422 (N_16422,N_14715,N_15748);
or U16423 (N_16423,N_15111,N_15833);
nand U16424 (N_16424,N_15551,N_14517);
and U16425 (N_16425,N_14382,N_14088);
or U16426 (N_16426,N_14737,N_15667);
or U16427 (N_16427,N_14371,N_14524);
and U16428 (N_16428,N_15611,N_14291);
xor U16429 (N_16429,N_14136,N_15653);
nand U16430 (N_16430,N_15000,N_14537);
nor U16431 (N_16431,N_14249,N_15735);
xnor U16432 (N_16432,N_14263,N_15331);
and U16433 (N_16433,N_15851,N_15858);
xor U16434 (N_16434,N_14652,N_14994);
and U16435 (N_16435,N_15393,N_15291);
and U16436 (N_16436,N_14193,N_15032);
xor U16437 (N_16437,N_14555,N_15930);
nor U16438 (N_16438,N_15420,N_14803);
or U16439 (N_16439,N_14039,N_15257);
xor U16440 (N_16440,N_15569,N_14234);
or U16441 (N_16441,N_15375,N_15575);
nand U16442 (N_16442,N_14275,N_15509);
xnor U16443 (N_16443,N_15019,N_14905);
nand U16444 (N_16444,N_15240,N_14702);
nor U16445 (N_16445,N_14581,N_14426);
nor U16446 (N_16446,N_15654,N_15629);
nand U16447 (N_16447,N_15886,N_15354);
nor U16448 (N_16448,N_14591,N_14385);
nand U16449 (N_16449,N_14325,N_14358);
nand U16450 (N_16450,N_14445,N_15734);
and U16451 (N_16451,N_15504,N_15498);
xor U16452 (N_16452,N_14934,N_15937);
xnor U16453 (N_16453,N_15591,N_15369);
nand U16454 (N_16454,N_14963,N_14217);
or U16455 (N_16455,N_14654,N_15015);
nand U16456 (N_16456,N_15197,N_15752);
or U16457 (N_16457,N_15236,N_14681);
and U16458 (N_16458,N_14705,N_14357);
or U16459 (N_16459,N_15088,N_14021);
nor U16460 (N_16460,N_15185,N_15622);
or U16461 (N_16461,N_15319,N_15288);
nor U16462 (N_16462,N_15942,N_14089);
xnor U16463 (N_16463,N_15662,N_14046);
nor U16464 (N_16464,N_14309,N_14574);
nand U16465 (N_16465,N_15189,N_15648);
xor U16466 (N_16466,N_14846,N_14288);
xnor U16467 (N_16467,N_15814,N_15774);
or U16468 (N_16468,N_14512,N_15332);
nand U16469 (N_16469,N_14551,N_14657);
nor U16470 (N_16470,N_15898,N_14427);
nand U16471 (N_16471,N_15441,N_14599);
and U16472 (N_16472,N_14313,N_14535);
or U16473 (N_16473,N_15690,N_14939);
and U16474 (N_16474,N_15348,N_14889);
or U16475 (N_16475,N_14036,N_15910);
or U16476 (N_16476,N_14048,N_15160);
or U16477 (N_16477,N_15765,N_14656);
nor U16478 (N_16478,N_15297,N_15865);
and U16479 (N_16479,N_15062,N_15912);
and U16480 (N_16480,N_15612,N_15773);
xor U16481 (N_16481,N_14571,N_15740);
nor U16482 (N_16482,N_14197,N_15351);
xnor U16483 (N_16483,N_14340,N_15281);
or U16484 (N_16484,N_15469,N_14766);
or U16485 (N_16485,N_14877,N_14144);
or U16486 (N_16486,N_15182,N_14184);
xor U16487 (N_16487,N_14509,N_15457);
nand U16488 (N_16488,N_14577,N_15896);
xnor U16489 (N_16489,N_14953,N_15442);
nor U16490 (N_16490,N_15918,N_14243);
or U16491 (N_16491,N_14784,N_14612);
and U16492 (N_16492,N_14633,N_15958);
or U16493 (N_16493,N_15227,N_15342);
nor U16494 (N_16494,N_14203,N_15335);
xor U16495 (N_16495,N_15903,N_14764);
nand U16496 (N_16496,N_14049,N_15205);
nand U16497 (N_16497,N_14793,N_14246);
nand U16498 (N_16498,N_15951,N_15139);
and U16499 (N_16499,N_15466,N_14218);
nand U16500 (N_16500,N_14796,N_14280);
and U16501 (N_16501,N_15478,N_14456);
or U16502 (N_16502,N_15078,N_14786);
or U16503 (N_16503,N_14388,N_14149);
nand U16504 (N_16504,N_14065,N_15485);
nand U16505 (N_16505,N_14443,N_14549);
nor U16506 (N_16506,N_14964,N_15834);
or U16507 (N_16507,N_14123,N_14900);
nand U16508 (N_16508,N_15753,N_14111);
and U16509 (N_16509,N_15864,N_14220);
and U16510 (N_16510,N_15166,N_15330);
or U16511 (N_16511,N_15986,N_14428);
xor U16512 (N_16512,N_15056,N_15689);
xor U16513 (N_16513,N_14672,N_15020);
nand U16514 (N_16514,N_15794,N_14489);
nand U16515 (N_16515,N_14837,N_15172);
and U16516 (N_16516,N_15244,N_15184);
nand U16517 (N_16517,N_14559,N_14189);
nand U16518 (N_16518,N_14396,N_14399);
and U16519 (N_16519,N_15809,N_14912);
or U16520 (N_16520,N_15224,N_15503);
nand U16521 (N_16521,N_15229,N_15991);
and U16522 (N_16522,N_15906,N_14286);
xnor U16523 (N_16523,N_15520,N_15271);
nor U16524 (N_16524,N_14016,N_15607);
or U16525 (N_16525,N_14129,N_14279);
nor U16526 (N_16526,N_14440,N_15743);
and U16527 (N_16527,N_15850,N_15721);
nand U16528 (N_16528,N_15449,N_15340);
and U16529 (N_16529,N_14022,N_15263);
and U16530 (N_16530,N_14940,N_14625);
nor U16531 (N_16531,N_15584,N_14938);
or U16532 (N_16532,N_15103,N_15155);
or U16533 (N_16533,N_14228,N_15623);
nand U16534 (N_16534,N_14077,N_14677);
xor U16535 (N_16535,N_15658,N_15218);
xor U16536 (N_16536,N_15660,N_15630);
nand U16537 (N_16537,N_14033,N_14319);
or U16538 (N_16538,N_14105,N_15206);
xnor U16539 (N_16539,N_14392,N_15738);
xor U16540 (N_16540,N_14873,N_15368);
or U16541 (N_16541,N_14282,N_15739);
nand U16542 (N_16542,N_14974,N_15980);
nor U16543 (N_16543,N_15862,N_15372);
nand U16544 (N_16544,N_14377,N_14194);
or U16545 (N_16545,N_14073,N_14405);
and U16546 (N_16546,N_14508,N_15483);
nand U16547 (N_16547,N_15843,N_14959);
or U16548 (N_16548,N_14907,N_14122);
nand U16549 (N_16549,N_14844,N_14421);
or U16550 (N_16550,N_14488,N_15149);
or U16551 (N_16551,N_14720,N_15025);
and U16552 (N_16552,N_14163,N_15421);
nor U16553 (N_16553,N_15242,N_14610);
and U16554 (N_16554,N_14106,N_14281);
xor U16555 (N_16555,N_14017,N_14542);
nor U16556 (N_16556,N_15772,N_15055);
xor U16557 (N_16557,N_14200,N_15983);
and U16558 (N_16558,N_14251,N_15646);
or U16559 (N_16559,N_15484,N_15213);
nor U16560 (N_16560,N_14187,N_15635);
nor U16561 (N_16561,N_14976,N_14962);
nand U16562 (N_16562,N_15967,N_15553);
or U16563 (N_16563,N_15759,N_15128);
xnor U16564 (N_16564,N_15010,N_14403);
and U16565 (N_16565,N_15444,N_15148);
or U16566 (N_16566,N_14307,N_15692);
nor U16567 (N_16567,N_15931,N_14951);
nand U16568 (N_16568,N_15754,N_14757);
nor U16569 (N_16569,N_15631,N_15493);
nand U16570 (N_16570,N_15174,N_15424);
or U16571 (N_16571,N_14432,N_14792);
and U16572 (N_16572,N_14653,N_15251);
nor U16573 (N_16573,N_14013,N_14198);
nand U16574 (N_16574,N_15328,N_15460);
or U16575 (N_16575,N_14437,N_15119);
and U16576 (N_16576,N_15114,N_14748);
and U16577 (N_16577,N_14930,N_14028);
nand U16578 (N_16578,N_14401,N_15666);
nand U16579 (N_16579,N_15792,N_15705);
or U16580 (N_16580,N_14434,N_15346);
nand U16581 (N_16581,N_15045,N_14031);
nor U16582 (N_16582,N_14977,N_14791);
and U16583 (N_16583,N_14153,N_14247);
xor U16584 (N_16584,N_14009,N_15943);
nor U16585 (N_16585,N_15505,N_15687);
and U16586 (N_16586,N_14899,N_15638);
nor U16587 (N_16587,N_14242,N_14861);
and U16588 (N_16588,N_14402,N_14045);
nand U16589 (N_16589,N_14146,N_14248);
xor U16590 (N_16590,N_15086,N_14104);
nor U16591 (N_16591,N_15186,N_14913);
or U16592 (N_16592,N_15990,N_15419);
or U16593 (N_16593,N_15936,N_15543);
or U16594 (N_16594,N_15344,N_14295);
nand U16595 (N_16595,N_15531,N_14326);
xor U16596 (N_16596,N_14147,N_14582);
or U16597 (N_16597,N_15719,N_14114);
nor U16598 (N_16598,N_14541,N_15959);
and U16599 (N_16599,N_14094,N_15350);
or U16600 (N_16600,N_15385,N_15708);
nor U16601 (N_16601,N_14699,N_15203);
or U16602 (N_16602,N_15266,N_15866);
xnor U16603 (N_16603,N_15373,N_14232);
and U16604 (N_16604,N_15836,N_15371);
nand U16605 (N_16605,N_15927,N_14164);
nor U16606 (N_16606,N_14584,N_14159);
nor U16607 (N_16607,N_15710,N_15815);
or U16608 (N_16608,N_14615,N_14650);
or U16609 (N_16609,N_15234,N_14096);
xnor U16610 (N_16610,N_14778,N_14885);
and U16611 (N_16611,N_15909,N_14066);
or U16612 (N_16612,N_14341,N_15279);
or U16613 (N_16613,N_15854,N_15703);
nor U16614 (N_16614,N_15940,N_15284);
and U16615 (N_16615,N_14091,N_14866);
nand U16616 (N_16616,N_15210,N_14346);
and U16617 (N_16617,N_14353,N_14483);
and U16618 (N_16618,N_14107,N_14647);
nor U16619 (N_16619,N_14991,N_15907);
and U16620 (N_16620,N_14102,N_15803);
or U16621 (N_16621,N_15729,N_15028);
and U16622 (N_16622,N_15860,N_15122);
xor U16623 (N_16623,N_14233,N_14514);
nor U16624 (N_16624,N_15123,N_15768);
xor U16625 (N_16625,N_14215,N_14290);
nor U16626 (N_16626,N_14335,N_15388);
xor U16627 (N_16627,N_14669,N_15530);
nor U16628 (N_16628,N_15009,N_15273);
and U16629 (N_16629,N_14880,N_15916);
and U16630 (N_16630,N_14253,N_14696);
or U16631 (N_16631,N_14546,N_14770);
or U16632 (N_16632,N_15070,N_15961);
xor U16633 (N_16633,N_15156,N_14097);
and U16634 (N_16634,N_15852,N_15353);
nor U16635 (N_16635,N_14865,N_14306);
nand U16636 (N_16636,N_14130,N_14025);
or U16637 (N_16637,N_15162,N_14165);
nand U16638 (N_16638,N_15876,N_14132);
and U16639 (N_16639,N_14527,N_14999);
nor U16640 (N_16640,N_14543,N_15763);
and U16641 (N_16641,N_15398,N_15995);
nand U16642 (N_16642,N_15300,N_14690);
or U16643 (N_16643,N_15202,N_15169);
or U16644 (N_16644,N_15661,N_14995);
nor U16645 (N_16645,N_15280,N_14923);
nor U16646 (N_16646,N_15974,N_15465);
nand U16647 (N_16647,N_15467,N_14759);
nand U16648 (N_16648,N_14332,N_14207);
nand U16649 (N_16649,N_14819,N_15065);
xnor U16650 (N_16650,N_14093,N_14713);
or U16651 (N_16651,N_14244,N_15704);
nand U16652 (N_16652,N_15208,N_15304);
nor U16653 (N_16653,N_14590,N_14070);
nand U16654 (N_16654,N_15387,N_14199);
or U16655 (N_16655,N_15053,N_15619);
xnor U16656 (N_16656,N_15723,N_14298);
nor U16657 (N_16657,N_15839,N_15083);
nand U16658 (N_16658,N_14362,N_14501);
and U16659 (N_16659,N_15253,N_15389);
nor U16660 (N_16660,N_15730,N_14881);
nor U16661 (N_16661,N_14666,N_15770);
nand U16662 (N_16662,N_14103,N_14398);
nor U16663 (N_16663,N_15480,N_15193);
nor U16664 (N_16664,N_15579,N_15036);
and U16665 (N_16665,N_14455,N_14329);
xor U16666 (N_16666,N_14801,N_14338);
nor U16667 (N_16667,N_15347,N_14782);
nand U16668 (N_16668,N_15603,N_15844);
or U16669 (N_16669,N_14124,N_15925);
nand U16670 (N_16670,N_15939,N_14597);
and U16671 (N_16671,N_14289,N_14236);
xnor U16672 (N_16672,N_15054,N_14842);
and U16673 (N_16673,N_15109,N_15978);
nor U16674 (N_16674,N_15751,N_15425);
and U16675 (N_16675,N_15917,N_15897);
or U16676 (N_16676,N_15102,N_14738);
nor U16677 (N_16677,N_15237,N_14917);
or U16678 (N_16678,N_15217,N_15857);
or U16679 (N_16679,N_14317,N_14645);
nor U16680 (N_16680,N_14849,N_15443);
xnor U16681 (N_16681,N_14573,N_14180);
and U16682 (N_16682,N_14071,N_14495);
or U16683 (N_16683,N_14952,N_15418);
and U16684 (N_16684,N_15682,N_14660);
xnor U16685 (N_16685,N_15556,N_14064);
nand U16686 (N_16686,N_15192,N_14410);
and U16687 (N_16687,N_15486,N_14260);
nor U16688 (N_16688,N_15806,N_15298);
and U16689 (N_16689,N_14001,N_15502);
nor U16690 (N_16690,N_14214,N_15606);
or U16691 (N_16691,N_15695,N_15693);
nand U16692 (N_16692,N_15158,N_15067);
and U16693 (N_16693,N_15888,N_15762);
xor U16694 (N_16694,N_15676,N_15968);
nand U16695 (N_16695,N_15970,N_14118);
and U16696 (N_16696,N_14452,N_14024);
nor U16697 (N_16697,N_15848,N_14622);
xor U16698 (N_16698,N_15617,N_15463);
xor U16699 (N_16699,N_15913,N_15270);
and U16700 (N_16700,N_14141,N_14032);
nand U16701 (N_16701,N_15562,N_14520);
nand U16702 (N_16702,N_15106,N_14980);
xor U16703 (N_16703,N_15824,N_14728);
nand U16704 (N_16704,N_15899,N_15571);
or U16705 (N_16705,N_14918,N_15474);
nor U16706 (N_16706,N_14678,N_14890);
nor U16707 (N_16707,N_14853,N_14101);
nand U16708 (N_16708,N_14477,N_15742);
nor U16709 (N_16709,N_14697,N_15709);
nor U16710 (N_16710,N_14230,N_15458);
or U16711 (N_16711,N_14616,N_14522);
or U16712 (N_16712,N_15915,N_14863);
nor U16713 (N_16713,N_15201,N_15491);
nor U16714 (N_16714,N_15475,N_14231);
or U16715 (N_16715,N_15124,N_14539);
xnor U16716 (N_16716,N_14376,N_15159);
nor U16717 (N_16717,N_15325,N_14632);
or U16718 (N_16718,N_14576,N_14018);
or U16719 (N_16719,N_15157,N_15430);
and U16720 (N_16720,N_14479,N_14879);
and U16721 (N_16721,N_15577,N_15258);
and U16722 (N_16722,N_15599,N_15992);
nand U16723 (N_16723,N_14602,N_14971);
nand U16724 (N_16724,N_15905,N_14858);
nor U16725 (N_16725,N_15525,N_14412);
and U16726 (N_16726,N_14762,N_14765);
or U16727 (N_16727,N_15766,N_14468);
and U16728 (N_16728,N_14435,N_15956);
nand U16729 (N_16729,N_14305,N_15071);
and U16730 (N_16730,N_15663,N_15287);
xnor U16731 (N_16731,N_14799,N_14080);
nor U16732 (N_16732,N_14191,N_14965);
or U16733 (N_16733,N_14005,N_14270);
and U16734 (N_16734,N_15699,N_14725);
xnor U16735 (N_16735,N_14547,N_14928);
nand U16736 (N_16736,N_14611,N_15428);
nor U16737 (N_16737,N_15264,N_15816);
xnor U16738 (N_16738,N_15975,N_14644);
nor U16739 (N_16739,N_14659,N_15105);
or U16740 (N_16740,N_14413,N_15147);
xnor U16741 (N_16741,N_14055,N_14202);
nor U16742 (N_16742,N_15301,N_14463);
xor U16743 (N_16743,N_15582,N_14273);
and U16744 (N_16744,N_14380,N_14896);
and U16745 (N_16745,N_14997,N_15131);
nor U16746 (N_16746,N_14982,N_14205);
xnor U16747 (N_16747,N_14235,N_14116);
nor U16748 (N_16748,N_14364,N_14609);
and U16749 (N_16749,N_15744,N_14310);
nand U16750 (N_16750,N_15414,N_15510);
nand U16751 (N_16751,N_14658,N_14915);
or U16752 (N_16752,N_15431,N_15588);
or U16753 (N_16753,N_15142,N_15869);
or U16754 (N_16754,N_14050,N_14787);
xor U16755 (N_16755,N_15262,N_15810);
and U16756 (N_16756,N_14909,N_15047);
and U16757 (N_16757,N_15293,N_15600);
and U16758 (N_16758,N_14344,N_15871);
and U16759 (N_16759,N_15706,N_14043);
nand U16760 (N_16760,N_15152,N_15003);
xnor U16761 (N_16761,N_14007,N_15948);
xnor U16762 (N_16762,N_14533,N_15007);
or U16763 (N_16763,N_15583,N_14381);
xnor U16764 (N_16764,N_15994,N_15188);
nor U16765 (N_16765,N_14160,N_15828);
or U16766 (N_16766,N_15880,N_14003);
nor U16767 (N_16767,N_15557,N_15572);
or U16768 (N_16768,N_15269,N_15511);
or U16769 (N_16769,N_15422,N_15051);
nand U16770 (N_16770,N_15471,N_14360);
nor U16771 (N_16771,N_15283,N_14598);
nand U16772 (N_16772,N_15574,N_14047);
nand U16773 (N_16773,N_15050,N_15501);
or U16774 (N_16774,N_15356,N_14473);
xor U16775 (N_16775,N_14411,N_14795);
xnor U16776 (N_16776,N_15895,N_14688);
nor U16777 (N_16777,N_15049,N_14948);
nor U16778 (N_16778,N_14085,N_14121);
nand U16779 (N_16779,N_14174,N_15323);
or U16780 (N_16780,N_14773,N_15514);
or U16781 (N_16781,N_15016,N_15887);
nand U16782 (N_16782,N_14862,N_14834);
and U16783 (N_16783,N_15408,N_14806);
and U16784 (N_16784,N_15455,N_15130);
or U16785 (N_16785,N_15780,N_14875);
and U16786 (N_16786,N_15534,N_14781);
or U16787 (N_16787,N_15665,N_14694);
and U16788 (N_16788,N_14406,N_14222);
and U16789 (N_16789,N_14267,N_15840);
and U16790 (N_16790,N_15532,N_15084);
nor U16791 (N_16791,N_14548,N_14271);
xor U16792 (N_16792,N_15499,N_14969);
and U16793 (N_16793,N_15376,N_15506);
nand U16794 (N_16794,N_15979,N_14135);
xor U16795 (N_16795,N_15034,N_14771);
nand U16796 (N_16796,N_15081,N_14750);
xor U16797 (N_16797,N_15040,N_15093);
nor U16798 (N_16798,N_15094,N_14474);
or U16799 (N_16799,N_14800,N_14439);
or U16800 (N_16800,N_15691,N_15552);
nand U16801 (N_16801,N_14391,N_14297);
nand U16802 (N_16802,N_15924,N_14314);
nor U16803 (N_16803,N_14416,N_15756);
xor U16804 (N_16804,N_14181,N_15311);
nor U16805 (N_16805,N_15793,N_14868);
xnor U16806 (N_16806,N_15601,N_15085);
or U16807 (N_16807,N_14304,N_14753);
and U16808 (N_16808,N_15715,N_14578);
xnor U16809 (N_16809,N_14469,N_14621);
or U16810 (N_16810,N_15405,N_14168);
nor U16811 (N_16811,N_14855,N_15981);
and U16812 (N_16812,N_15487,N_14433);
xnor U16813 (N_16813,N_14821,N_14538);
nand U16814 (N_16814,N_15079,N_14386);
or U16815 (N_16815,N_14324,N_15632);
nand U16816 (N_16816,N_15827,N_15239);
nor U16817 (N_16817,N_15745,N_15628);
nand U16818 (N_16818,N_15627,N_14777);
xnor U16819 (N_16819,N_15633,N_15618);
xor U16820 (N_16820,N_15922,N_14589);
xor U16821 (N_16821,N_15299,N_14724);
xor U16822 (N_16822,N_15540,N_14910);
xor U16823 (N_16823,N_14714,N_15669);
nand U16824 (N_16824,N_15115,N_15900);
xnor U16825 (N_16825,N_15445,N_15830);
or U16826 (N_16826,N_14333,N_15657);
nand U16827 (N_16827,N_15390,N_14072);
nand U16828 (N_16828,N_15216,N_14895);
xor U16829 (N_16829,N_14476,N_14746);
nor U16830 (N_16830,N_14418,N_14255);
nand U16831 (N_16831,N_15125,N_14461);
nand U16832 (N_16832,N_15256,N_14682);
xor U16833 (N_16833,N_14081,N_15527);
or U16834 (N_16834,N_14528,N_14062);
xor U16835 (N_16835,N_14099,N_14630);
xnor U16836 (N_16836,N_15494,N_14843);
and U16837 (N_16837,N_14788,N_14662);
or U16838 (N_16838,N_14722,N_14704);
nor U16839 (N_16839,N_15716,N_14068);
xnor U16840 (N_16840,N_14683,N_15228);
nor U16841 (N_16841,N_15135,N_14532);
and U16842 (N_16842,N_15919,N_14711);
nor U16843 (N_16843,N_14438,N_14998);
nor U16844 (N_16844,N_15594,N_14901);
nor U16845 (N_16845,N_15568,N_14761);
xor U16846 (N_16846,N_14935,N_15006);
nor U16847 (N_16847,N_14857,N_15524);
or U16848 (N_16848,N_15108,N_15849);
and U16849 (N_16849,N_14758,N_14204);
or U16850 (N_16850,N_14020,N_15953);
xnor U16851 (N_16851,N_14422,N_15315);
xor U16852 (N_16852,N_14679,N_15726);
and U16853 (N_16853,N_14960,N_14872);
nand U16854 (N_16854,N_14137,N_14337);
or U16855 (N_16855,N_14921,N_14138);
xnor U16856 (N_16856,N_15998,N_15417);
nor U16857 (N_16857,N_15921,N_14450);
and U16858 (N_16858,N_15781,N_14947);
xnor U16859 (N_16859,N_15586,N_15058);
xor U16860 (N_16860,N_15901,N_14575);
nor U16861 (N_16861,N_14511,N_14493);
or U16862 (N_16862,N_15831,N_15962);
nor U16863 (N_16863,N_15226,N_14839);
nand U16864 (N_16864,N_15077,N_14370);
or U16865 (N_16865,N_15247,N_14139);
xor U16866 (N_16866,N_14926,N_15024);
nor U16867 (N_16867,N_15713,N_15616);
nor U16868 (N_16868,N_15749,N_15410);
xor U16869 (N_16869,N_15602,N_15680);
nand U16870 (N_16870,N_14937,N_14721);
nand U16871 (N_16871,N_14869,N_14594);
nor U16872 (N_16872,N_14726,N_14710);
xnor U16873 (N_16873,N_14563,N_15701);
and U16874 (N_16874,N_14804,N_15268);
nor U16875 (N_16875,N_15324,N_14014);
and U16876 (N_16876,N_15338,N_15767);
nand U16877 (N_16877,N_14368,N_15712);
xor U16878 (N_16878,N_14733,N_15960);
xor U16879 (N_16879,N_15026,N_15321);
and U16880 (N_16880,N_15002,N_15104);
xnor U16881 (N_16881,N_15059,N_15881);
xnor U16882 (N_16882,N_14680,N_14933);
and U16883 (N_16883,N_15702,N_15889);
nand U16884 (N_16884,N_14034,N_15129);
nand U16885 (N_16885,N_15468,N_15949);
or U16886 (N_16886,N_14052,N_15073);
xor U16887 (N_16887,N_15211,N_15788);
nand U16888 (N_16888,N_15867,N_14151);
nor U16889 (N_16889,N_15598,N_15590);
nor U16890 (N_16890,N_14328,N_15144);
nor U16891 (N_16891,N_14956,N_15349);
and U16892 (N_16892,N_15538,N_15087);
xnor U16893 (N_16893,N_14627,N_14818);
and U16894 (N_16894,N_14798,N_14161);
nand U16895 (N_16895,N_14023,N_14903);
or U16896 (N_16896,N_15112,N_15972);
nand U16897 (N_16897,N_14825,N_14170);
and U16898 (N_16898,N_14481,N_15926);
nand U16899 (N_16899,N_15647,N_14173);
nand U16900 (N_16900,N_15935,N_14490);
or U16901 (N_16901,N_14051,N_15604);
nor U16902 (N_16902,N_15807,N_14550);
xnor U16903 (N_16903,N_14651,N_14747);
nor U16904 (N_16904,N_15697,N_15214);
nor U16905 (N_16905,N_15879,N_14707);
nand U16906 (N_16906,N_14712,N_15883);
and U16907 (N_16907,N_14815,N_15969);
or U16908 (N_16908,N_14674,N_14754);
and U16909 (N_16909,N_15396,N_14069);
and U16910 (N_16910,N_15758,N_14195);
nor U16911 (N_16911,N_14729,N_14453);
xor U16912 (N_16912,N_14916,N_15731);
xor U16913 (N_16913,N_15813,N_14264);
xor U16914 (N_16914,N_14635,N_15031);
nand U16915 (N_16915,N_14596,N_14177);
xnor U16916 (N_16916,N_15339,N_15456);
and U16917 (N_16917,N_14668,N_14510);
and U16918 (N_16918,N_14196,N_14296);
nor U16919 (N_16919,N_14906,N_14354);
nand U16920 (N_16920,N_14663,N_14431);
or U16921 (N_16921,N_14188,N_15517);
and U16922 (N_16922,N_14664,N_15337);
or U16923 (N_16923,N_14986,N_15164);
or U16924 (N_16924,N_15427,N_14374);
and U16925 (N_16925,N_14301,N_15100);
xor U16926 (N_16926,N_14593,N_14407);
nor U16927 (N_16927,N_14186,N_15429);
xnor U16928 (N_16928,N_14776,N_15395);
and U16929 (N_16929,N_14311,N_14824);
nand U16930 (N_16930,N_15817,N_14423);
and U16931 (N_16931,N_15845,N_15861);
nor U16932 (N_16932,N_14671,N_14608);
xor U16933 (N_16933,N_14029,N_14639);
nor U16934 (N_16934,N_15548,N_15249);
nor U16935 (N_16935,N_15812,N_14756);
or U16936 (N_16936,N_14321,N_14448);
or U16937 (N_16937,N_15276,N_14245);
or U16938 (N_16938,N_14183,N_15847);
and U16939 (N_16939,N_15933,N_14676);
nand U16940 (N_16940,N_14727,N_15440);
xor U16941 (N_16941,N_15732,N_15585);
and U16942 (N_16942,N_15212,N_14058);
xor U16943 (N_16943,N_15308,N_15204);
nor U16944 (N_16944,N_15080,N_15153);
nand U16945 (N_16945,N_15261,N_14908);
xor U16946 (N_16946,N_14420,N_15282);
and U16947 (N_16947,N_14079,N_14567);
xnor U16948 (N_16948,N_14491,N_15717);
xnor U16949 (N_16949,N_15920,N_15366);
nor U16950 (N_16950,N_14667,N_15220);
or U16951 (N_16951,N_14318,N_14734);
nand U16952 (N_16952,N_14557,N_14540);
nor U16953 (N_16953,N_15977,N_14684);
xnor U16954 (N_16954,N_15064,N_14113);
or U16955 (N_16955,N_15798,N_15091);
xor U16956 (N_16956,N_14266,N_15392);
and U16957 (N_16957,N_14210,N_14394);
or U16958 (N_16958,N_15963,N_14700);
xnor U16959 (N_16959,N_14336,N_14709);
nand U16960 (N_16960,N_14470,N_15341);
nor U16961 (N_16961,N_14484,N_15370);
nand U16962 (N_16962,N_15012,N_15537);
nor U16963 (N_16963,N_15954,N_14004);
xnor U16964 (N_16964,N_15832,N_15277);
or U16965 (N_16965,N_15868,N_15811);
nand U16966 (N_16966,N_14966,N_15409);
nor U16967 (N_16967,N_15698,N_15624);
nand U16968 (N_16968,N_15363,N_14695);
nand U16969 (N_16969,N_14716,N_14229);
nor U16970 (N_16970,N_15322,N_15966);
and U16971 (N_16971,N_14209,N_14086);
nor U16972 (N_16972,N_14038,N_15947);
and U16973 (N_16973,N_15198,N_15127);
xor U16974 (N_16974,N_15423,N_14618);
nand U16975 (N_16975,N_14809,N_14961);
and U16976 (N_16976,N_15246,N_15567);
xor U16977 (N_16977,N_15076,N_14568);
and U16978 (N_16978,N_15821,N_14348);
and U16979 (N_16979,N_14171,N_15238);
xnor U16980 (N_16980,N_15274,N_15289);
or U16981 (N_16981,N_15877,N_14480);
and U16982 (N_16982,N_15750,N_14152);
xor U16983 (N_16983,N_15179,N_14878);
nor U16984 (N_16984,N_14685,N_14487);
nand U16985 (N_16985,N_14176,N_14254);
nand U16986 (N_16986,N_15110,N_14012);
nor U16987 (N_16987,N_14922,N_14067);
or U16988 (N_16988,N_14569,N_14730);
and U16989 (N_16989,N_14835,N_14572);
nor U16990 (N_16990,N_14931,N_14972);
nor U16991 (N_16991,N_15533,N_15231);
and U16992 (N_16992,N_15233,N_15853);
or U16993 (N_16993,N_14201,N_15589);
nor U16994 (N_16994,N_14828,N_15250);
and U16995 (N_16995,N_14831,N_15303);
nor U16996 (N_16996,N_15343,N_14811);
or U16997 (N_16997,N_14518,N_14417);
nor U16998 (N_16998,N_15454,N_15945);
xnor U16999 (N_16999,N_15670,N_14893);
or U17000 (N_17000,N_15996,N_14072);
or U17001 (N_17001,N_15381,N_14024);
nor U17002 (N_17002,N_15991,N_14720);
and U17003 (N_17003,N_15509,N_15384);
nand U17004 (N_17004,N_14321,N_15746);
nand U17005 (N_17005,N_14965,N_15130);
and U17006 (N_17006,N_15890,N_15450);
nor U17007 (N_17007,N_15771,N_14787);
nor U17008 (N_17008,N_15934,N_14568);
and U17009 (N_17009,N_14236,N_14076);
and U17010 (N_17010,N_15910,N_14986);
nor U17011 (N_17011,N_15998,N_14943);
nor U17012 (N_17012,N_15600,N_15553);
or U17013 (N_17013,N_14352,N_15262);
nand U17014 (N_17014,N_14065,N_15944);
or U17015 (N_17015,N_15668,N_15593);
or U17016 (N_17016,N_14709,N_14702);
xor U17017 (N_17017,N_14931,N_15225);
nor U17018 (N_17018,N_14173,N_15038);
or U17019 (N_17019,N_15389,N_15056);
nand U17020 (N_17020,N_15327,N_15961);
and U17021 (N_17021,N_14390,N_15206);
or U17022 (N_17022,N_14815,N_15172);
xor U17023 (N_17023,N_14872,N_15740);
or U17024 (N_17024,N_15996,N_14494);
and U17025 (N_17025,N_15850,N_14772);
or U17026 (N_17026,N_14310,N_15023);
and U17027 (N_17027,N_14011,N_15872);
xnor U17028 (N_17028,N_15928,N_15868);
or U17029 (N_17029,N_14088,N_15916);
xnor U17030 (N_17030,N_15130,N_14389);
or U17031 (N_17031,N_15398,N_14661);
nand U17032 (N_17032,N_14970,N_15000);
or U17033 (N_17033,N_15721,N_14733);
nor U17034 (N_17034,N_15639,N_14923);
nor U17035 (N_17035,N_14595,N_14319);
and U17036 (N_17036,N_14448,N_15298);
nand U17037 (N_17037,N_15943,N_14763);
xnor U17038 (N_17038,N_14430,N_15742);
xor U17039 (N_17039,N_15378,N_14916);
xor U17040 (N_17040,N_14832,N_15731);
and U17041 (N_17041,N_14708,N_15799);
nor U17042 (N_17042,N_15219,N_15402);
and U17043 (N_17043,N_15469,N_14364);
and U17044 (N_17044,N_14285,N_14954);
nand U17045 (N_17045,N_14026,N_14529);
nand U17046 (N_17046,N_14204,N_14181);
and U17047 (N_17047,N_15286,N_14766);
or U17048 (N_17048,N_14033,N_15197);
nand U17049 (N_17049,N_15252,N_15460);
xnor U17050 (N_17050,N_15195,N_14465);
or U17051 (N_17051,N_14401,N_14314);
and U17052 (N_17052,N_14160,N_15315);
or U17053 (N_17053,N_14123,N_15718);
xnor U17054 (N_17054,N_15427,N_15579);
and U17055 (N_17055,N_15452,N_15903);
nor U17056 (N_17056,N_15098,N_15529);
xor U17057 (N_17057,N_14736,N_14672);
or U17058 (N_17058,N_14229,N_15772);
and U17059 (N_17059,N_14292,N_15498);
xnor U17060 (N_17060,N_14474,N_14938);
and U17061 (N_17061,N_14219,N_14550);
nor U17062 (N_17062,N_14785,N_14642);
nand U17063 (N_17063,N_15590,N_15359);
xnor U17064 (N_17064,N_15508,N_15485);
or U17065 (N_17065,N_14806,N_15377);
nor U17066 (N_17066,N_14435,N_14563);
or U17067 (N_17067,N_14904,N_15766);
xnor U17068 (N_17068,N_14920,N_14873);
nand U17069 (N_17069,N_14583,N_14406);
or U17070 (N_17070,N_15227,N_14889);
and U17071 (N_17071,N_15717,N_14970);
or U17072 (N_17072,N_15336,N_14183);
nor U17073 (N_17073,N_14125,N_14638);
xnor U17074 (N_17074,N_14120,N_14596);
nor U17075 (N_17075,N_15175,N_14692);
or U17076 (N_17076,N_15283,N_14708);
and U17077 (N_17077,N_14309,N_14592);
nor U17078 (N_17078,N_15846,N_15238);
and U17079 (N_17079,N_15951,N_14976);
nand U17080 (N_17080,N_15049,N_15358);
and U17081 (N_17081,N_15843,N_15076);
xnor U17082 (N_17082,N_14143,N_15594);
and U17083 (N_17083,N_14131,N_14708);
or U17084 (N_17084,N_15482,N_15805);
or U17085 (N_17085,N_15570,N_15559);
or U17086 (N_17086,N_15076,N_14463);
nor U17087 (N_17087,N_14657,N_15455);
and U17088 (N_17088,N_15357,N_14092);
nand U17089 (N_17089,N_14736,N_14292);
and U17090 (N_17090,N_14053,N_15988);
and U17091 (N_17091,N_15851,N_14845);
or U17092 (N_17092,N_15358,N_15387);
and U17093 (N_17093,N_15198,N_14208);
or U17094 (N_17094,N_14194,N_15461);
nor U17095 (N_17095,N_14172,N_14286);
and U17096 (N_17096,N_15697,N_15281);
nand U17097 (N_17097,N_15412,N_14592);
nand U17098 (N_17098,N_14995,N_14560);
nand U17099 (N_17099,N_14330,N_14595);
nor U17100 (N_17100,N_14606,N_15397);
or U17101 (N_17101,N_14736,N_14173);
nor U17102 (N_17102,N_14526,N_14511);
and U17103 (N_17103,N_15654,N_15747);
and U17104 (N_17104,N_14298,N_14271);
and U17105 (N_17105,N_14100,N_15189);
nand U17106 (N_17106,N_14249,N_15846);
nand U17107 (N_17107,N_14582,N_14345);
or U17108 (N_17108,N_14045,N_14779);
nand U17109 (N_17109,N_15313,N_15588);
nor U17110 (N_17110,N_14239,N_14793);
and U17111 (N_17111,N_14920,N_15833);
and U17112 (N_17112,N_14650,N_15426);
and U17113 (N_17113,N_15303,N_14815);
xnor U17114 (N_17114,N_14351,N_14270);
xnor U17115 (N_17115,N_15224,N_14950);
nand U17116 (N_17116,N_15197,N_15532);
nand U17117 (N_17117,N_15667,N_15353);
nand U17118 (N_17118,N_15929,N_14863);
nor U17119 (N_17119,N_15117,N_15937);
and U17120 (N_17120,N_15480,N_15766);
nor U17121 (N_17121,N_14088,N_14747);
or U17122 (N_17122,N_14127,N_15072);
and U17123 (N_17123,N_15958,N_15899);
nor U17124 (N_17124,N_14438,N_15360);
nor U17125 (N_17125,N_14285,N_15296);
nand U17126 (N_17126,N_14248,N_14102);
xor U17127 (N_17127,N_15534,N_14205);
nand U17128 (N_17128,N_15979,N_15649);
nand U17129 (N_17129,N_15986,N_15039);
or U17130 (N_17130,N_15448,N_14619);
nor U17131 (N_17131,N_15620,N_15859);
or U17132 (N_17132,N_14632,N_14892);
or U17133 (N_17133,N_15110,N_14871);
xor U17134 (N_17134,N_15100,N_15815);
nor U17135 (N_17135,N_14427,N_14358);
or U17136 (N_17136,N_14766,N_14676);
nand U17137 (N_17137,N_15448,N_15098);
or U17138 (N_17138,N_15552,N_14528);
nand U17139 (N_17139,N_14198,N_15592);
and U17140 (N_17140,N_15139,N_15222);
nor U17141 (N_17141,N_15299,N_15507);
nand U17142 (N_17142,N_15239,N_14873);
nand U17143 (N_17143,N_14672,N_15604);
and U17144 (N_17144,N_14646,N_14773);
and U17145 (N_17145,N_15785,N_15514);
and U17146 (N_17146,N_15352,N_15712);
nand U17147 (N_17147,N_15505,N_15111);
nand U17148 (N_17148,N_14905,N_14097);
or U17149 (N_17149,N_15923,N_15272);
nand U17150 (N_17150,N_15453,N_15070);
nor U17151 (N_17151,N_14663,N_15075);
nand U17152 (N_17152,N_15748,N_15604);
nand U17153 (N_17153,N_15618,N_14417);
and U17154 (N_17154,N_15043,N_14045);
or U17155 (N_17155,N_15453,N_15820);
xnor U17156 (N_17156,N_14498,N_14721);
or U17157 (N_17157,N_14963,N_14391);
and U17158 (N_17158,N_15452,N_15510);
and U17159 (N_17159,N_15583,N_14943);
nor U17160 (N_17160,N_14101,N_14750);
nand U17161 (N_17161,N_14737,N_15958);
nor U17162 (N_17162,N_14658,N_15867);
nor U17163 (N_17163,N_14704,N_14069);
nor U17164 (N_17164,N_15716,N_14950);
nand U17165 (N_17165,N_15365,N_15916);
xor U17166 (N_17166,N_15878,N_14871);
and U17167 (N_17167,N_14121,N_14735);
nor U17168 (N_17168,N_15109,N_15840);
or U17169 (N_17169,N_14422,N_14857);
nor U17170 (N_17170,N_15200,N_14051);
nor U17171 (N_17171,N_14008,N_14457);
or U17172 (N_17172,N_15173,N_14255);
xnor U17173 (N_17173,N_14393,N_15577);
or U17174 (N_17174,N_14081,N_15882);
and U17175 (N_17175,N_14974,N_15618);
and U17176 (N_17176,N_14471,N_15884);
or U17177 (N_17177,N_14868,N_14973);
or U17178 (N_17178,N_15149,N_15577);
xnor U17179 (N_17179,N_15697,N_15775);
nand U17180 (N_17180,N_14157,N_14319);
nand U17181 (N_17181,N_15622,N_14187);
or U17182 (N_17182,N_14637,N_15568);
nor U17183 (N_17183,N_15312,N_14185);
or U17184 (N_17184,N_14175,N_15351);
or U17185 (N_17185,N_14943,N_15111);
and U17186 (N_17186,N_15848,N_15628);
nand U17187 (N_17187,N_15117,N_15931);
and U17188 (N_17188,N_15484,N_14587);
or U17189 (N_17189,N_15530,N_14867);
or U17190 (N_17190,N_14235,N_15647);
xnor U17191 (N_17191,N_15513,N_15114);
nor U17192 (N_17192,N_15846,N_14611);
nor U17193 (N_17193,N_14792,N_14569);
or U17194 (N_17194,N_14829,N_15848);
xor U17195 (N_17195,N_15693,N_14855);
nor U17196 (N_17196,N_14602,N_14725);
and U17197 (N_17197,N_15801,N_15838);
or U17198 (N_17198,N_15202,N_14709);
or U17199 (N_17199,N_14265,N_15576);
and U17200 (N_17200,N_15586,N_14790);
xnor U17201 (N_17201,N_14589,N_14877);
nand U17202 (N_17202,N_14533,N_14011);
xor U17203 (N_17203,N_14133,N_15653);
xor U17204 (N_17204,N_15971,N_14630);
and U17205 (N_17205,N_14836,N_15053);
xor U17206 (N_17206,N_15744,N_15499);
nand U17207 (N_17207,N_15806,N_14285);
and U17208 (N_17208,N_15586,N_14966);
xor U17209 (N_17209,N_14023,N_14938);
xor U17210 (N_17210,N_14642,N_14197);
nand U17211 (N_17211,N_14013,N_14248);
and U17212 (N_17212,N_15145,N_15911);
xor U17213 (N_17213,N_15065,N_15657);
nor U17214 (N_17214,N_15996,N_15015);
nor U17215 (N_17215,N_15895,N_15981);
or U17216 (N_17216,N_15211,N_15725);
xor U17217 (N_17217,N_15116,N_14429);
or U17218 (N_17218,N_14864,N_14615);
xnor U17219 (N_17219,N_15288,N_14168);
nor U17220 (N_17220,N_15020,N_15659);
nand U17221 (N_17221,N_15003,N_15698);
or U17222 (N_17222,N_15353,N_14643);
nor U17223 (N_17223,N_14446,N_14675);
and U17224 (N_17224,N_15831,N_14727);
nor U17225 (N_17225,N_14311,N_15743);
and U17226 (N_17226,N_14333,N_15007);
and U17227 (N_17227,N_14417,N_14287);
or U17228 (N_17228,N_14289,N_14407);
nand U17229 (N_17229,N_14037,N_14605);
xnor U17230 (N_17230,N_15157,N_15410);
or U17231 (N_17231,N_15370,N_15673);
xnor U17232 (N_17232,N_14775,N_14680);
nor U17233 (N_17233,N_15116,N_15357);
or U17234 (N_17234,N_14412,N_14468);
xor U17235 (N_17235,N_14881,N_14172);
or U17236 (N_17236,N_14352,N_15573);
or U17237 (N_17237,N_14444,N_14141);
or U17238 (N_17238,N_14607,N_14498);
nand U17239 (N_17239,N_15752,N_15890);
xnor U17240 (N_17240,N_14342,N_14880);
nor U17241 (N_17241,N_14835,N_15009);
xnor U17242 (N_17242,N_14222,N_14970);
nor U17243 (N_17243,N_14863,N_15067);
and U17244 (N_17244,N_14864,N_15060);
and U17245 (N_17245,N_14293,N_14085);
nor U17246 (N_17246,N_15477,N_15060);
nor U17247 (N_17247,N_15696,N_14041);
nor U17248 (N_17248,N_14294,N_14099);
or U17249 (N_17249,N_15201,N_14805);
xor U17250 (N_17250,N_14415,N_15175);
xor U17251 (N_17251,N_15819,N_15478);
nor U17252 (N_17252,N_14458,N_14661);
or U17253 (N_17253,N_15666,N_15807);
and U17254 (N_17254,N_14840,N_15667);
or U17255 (N_17255,N_15923,N_14823);
xnor U17256 (N_17256,N_15473,N_14140);
and U17257 (N_17257,N_14089,N_15257);
and U17258 (N_17258,N_15014,N_15161);
xnor U17259 (N_17259,N_14598,N_14214);
or U17260 (N_17260,N_14097,N_14774);
and U17261 (N_17261,N_15358,N_14934);
or U17262 (N_17262,N_15510,N_14901);
xnor U17263 (N_17263,N_15253,N_14424);
nand U17264 (N_17264,N_14316,N_15159);
nor U17265 (N_17265,N_15973,N_14275);
nand U17266 (N_17266,N_15414,N_15925);
nor U17267 (N_17267,N_15159,N_14878);
or U17268 (N_17268,N_14096,N_14713);
nor U17269 (N_17269,N_15012,N_14679);
and U17270 (N_17270,N_15134,N_14143);
nor U17271 (N_17271,N_15876,N_14489);
xnor U17272 (N_17272,N_15744,N_14608);
or U17273 (N_17273,N_15734,N_14759);
xnor U17274 (N_17274,N_14683,N_14571);
or U17275 (N_17275,N_14132,N_14998);
nor U17276 (N_17276,N_15162,N_15933);
nor U17277 (N_17277,N_15318,N_14049);
nor U17278 (N_17278,N_14999,N_14415);
and U17279 (N_17279,N_15982,N_15913);
xor U17280 (N_17280,N_15848,N_14929);
nand U17281 (N_17281,N_14435,N_14075);
and U17282 (N_17282,N_14376,N_14031);
nor U17283 (N_17283,N_14187,N_14479);
and U17284 (N_17284,N_14352,N_14690);
nand U17285 (N_17285,N_15104,N_14308);
and U17286 (N_17286,N_15573,N_15029);
nor U17287 (N_17287,N_14149,N_15101);
nor U17288 (N_17288,N_15567,N_14444);
xnor U17289 (N_17289,N_15377,N_14018);
xor U17290 (N_17290,N_14716,N_15642);
nor U17291 (N_17291,N_14714,N_15216);
xor U17292 (N_17292,N_15340,N_14823);
or U17293 (N_17293,N_14437,N_14338);
nand U17294 (N_17294,N_14125,N_14533);
nand U17295 (N_17295,N_15831,N_15066);
xor U17296 (N_17296,N_14568,N_14086);
or U17297 (N_17297,N_15492,N_14487);
nor U17298 (N_17298,N_14162,N_14983);
xor U17299 (N_17299,N_14010,N_14583);
and U17300 (N_17300,N_14119,N_14055);
nand U17301 (N_17301,N_14907,N_14029);
nor U17302 (N_17302,N_15702,N_14486);
and U17303 (N_17303,N_15487,N_15859);
nor U17304 (N_17304,N_15327,N_14022);
or U17305 (N_17305,N_14924,N_15151);
nand U17306 (N_17306,N_14408,N_14045);
or U17307 (N_17307,N_15131,N_14906);
nand U17308 (N_17308,N_15751,N_15181);
nor U17309 (N_17309,N_15963,N_14368);
nand U17310 (N_17310,N_14545,N_14662);
nand U17311 (N_17311,N_14077,N_14107);
nor U17312 (N_17312,N_14091,N_14272);
xor U17313 (N_17313,N_15854,N_15626);
or U17314 (N_17314,N_14198,N_15415);
nor U17315 (N_17315,N_14265,N_14130);
xnor U17316 (N_17316,N_14098,N_15619);
xnor U17317 (N_17317,N_14331,N_15961);
or U17318 (N_17318,N_14978,N_15272);
and U17319 (N_17319,N_15014,N_15938);
nor U17320 (N_17320,N_15149,N_14403);
and U17321 (N_17321,N_15555,N_15751);
nor U17322 (N_17322,N_15876,N_15566);
nand U17323 (N_17323,N_14234,N_15416);
or U17324 (N_17324,N_15563,N_15324);
xnor U17325 (N_17325,N_14744,N_15016);
nand U17326 (N_17326,N_15172,N_14436);
and U17327 (N_17327,N_15089,N_14266);
nand U17328 (N_17328,N_15325,N_15438);
nor U17329 (N_17329,N_14939,N_14186);
nand U17330 (N_17330,N_15747,N_15358);
xor U17331 (N_17331,N_14778,N_15057);
nor U17332 (N_17332,N_15280,N_15461);
nand U17333 (N_17333,N_15382,N_15146);
nor U17334 (N_17334,N_14830,N_15181);
or U17335 (N_17335,N_14719,N_15212);
xor U17336 (N_17336,N_15094,N_14445);
nand U17337 (N_17337,N_14879,N_14579);
nor U17338 (N_17338,N_14947,N_14365);
nand U17339 (N_17339,N_14620,N_14615);
xnor U17340 (N_17340,N_15157,N_15052);
nand U17341 (N_17341,N_14266,N_14515);
or U17342 (N_17342,N_14781,N_15571);
nand U17343 (N_17343,N_15569,N_14618);
or U17344 (N_17344,N_15323,N_14782);
nor U17345 (N_17345,N_14301,N_14082);
nand U17346 (N_17346,N_14359,N_14387);
and U17347 (N_17347,N_14303,N_14185);
or U17348 (N_17348,N_15858,N_15900);
nand U17349 (N_17349,N_14413,N_14751);
xor U17350 (N_17350,N_15442,N_15957);
nand U17351 (N_17351,N_14923,N_14955);
and U17352 (N_17352,N_15384,N_15723);
and U17353 (N_17353,N_14833,N_15182);
and U17354 (N_17354,N_14601,N_14458);
xnor U17355 (N_17355,N_15585,N_15975);
nor U17356 (N_17356,N_15145,N_15966);
nor U17357 (N_17357,N_14320,N_14008);
xnor U17358 (N_17358,N_14140,N_14324);
xor U17359 (N_17359,N_14010,N_15916);
nand U17360 (N_17360,N_15502,N_15395);
and U17361 (N_17361,N_14198,N_15419);
nand U17362 (N_17362,N_14416,N_15589);
xnor U17363 (N_17363,N_14360,N_15850);
nand U17364 (N_17364,N_14449,N_14720);
and U17365 (N_17365,N_15980,N_14574);
or U17366 (N_17366,N_14404,N_15478);
xnor U17367 (N_17367,N_15767,N_14030);
or U17368 (N_17368,N_15663,N_14993);
xor U17369 (N_17369,N_15795,N_15555);
xnor U17370 (N_17370,N_15735,N_15059);
and U17371 (N_17371,N_14321,N_14745);
xor U17372 (N_17372,N_14858,N_14948);
nor U17373 (N_17373,N_15281,N_14191);
nand U17374 (N_17374,N_14011,N_14294);
or U17375 (N_17375,N_15180,N_14142);
nand U17376 (N_17376,N_14849,N_15908);
and U17377 (N_17377,N_15849,N_15989);
and U17378 (N_17378,N_15785,N_14016);
and U17379 (N_17379,N_15520,N_14555);
nor U17380 (N_17380,N_15997,N_14097);
xnor U17381 (N_17381,N_14183,N_14359);
nand U17382 (N_17382,N_15406,N_14176);
nor U17383 (N_17383,N_15902,N_14785);
or U17384 (N_17384,N_15801,N_14580);
nand U17385 (N_17385,N_14225,N_14277);
nand U17386 (N_17386,N_14727,N_15219);
nand U17387 (N_17387,N_15528,N_14829);
nor U17388 (N_17388,N_14309,N_14423);
and U17389 (N_17389,N_14083,N_15407);
and U17390 (N_17390,N_15703,N_15698);
xnor U17391 (N_17391,N_15782,N_14055);
xor U17392 (N_17392,N_15639,N_14387);
nand U17393 (N_17393,N_15929,N_14517);
and U17394 (N_17394,N_15257,N_15429);
and U17395 (N_17395,N_15257,N_15720);
nand U17396 (N_17396,N_14683,N_15211);
xnor U17397 (N_17397,N_14748,N_15278);
xor U17398 (N_17398,N_14233,N_15633);
or U17399 (N_17399,N_15016,N_14927);
or U17400 (N_17400,N_15985,N_14800);
and U17401 (N_17401,N_14102,N_14808);
nand U17402 (N_17402,N_15582,N_15751);
and U17403 (N_17403,N_14837,N_14967);
or U17404 (N_17404,N_14583,N_14611);
nand U17405 (N_17405,N_15143,N_14326);
or U17406 (N_17406,N_15376,N_14880);
nand U17407 (N_17407,N_14621,N_15408);
xor U17408 (N_17408,N_14906,N_15661);
or U17409 (N_17409,N_15055,N_15647);
nand U17410 (N_17410,N_15086,N_15807);
and U17411 (N_17411,N_15249,N_15276);
and U17412 (N_17412,N_14681,N_15653);
and U17413 (N_17413,N_14000,N_14967);
and U17414 (N_17414,N_15149,N_14063);
nor U17415 (N_17415,N_15522,N_15644);
and U17416 (N_17416,N_14577,N_15224);
nand U17417 (N_17417,N_15084,N_15284);
or U17418 (N_17418,N_15398,N_14037);
or U17419 (N_17419,N_15844,N_15666);
nand U17420 (N_17420,N_14371,N_15454);
nor U17421 (N_17421,N_15548,N_14757);
xor U17422 (N_17422,N_14497,N_15261);
and U17423 (N_17423,N_15663,N_15265);
xor U17424 (N_17424,N_14459,N_14298);
nand U17425 (N_17425,N_14125,N_15336);
xor U17426 (N_17426,N_14425,N_14085);
nor U17427 (N_17427,N_14492,N_15784);
or U17428 (N_17428,N_15290,N_14589);
and U17429 (N_17429,N_14992,N_14599);
and U17430 (N_17430,N_14840,N_15985);
and U17431 (N_17431,N_14197,N_15977);
nand U17432 (N_17432,N_14206,N_14476);
xnor U17433 (N_17433,N_15755,N_14611);
or U17434 (N_17434,N_14523,N_14775);
and U17435 (N_17435,N_15193,N_14003);
and U17436 (N_17436,N_14961,N_14550);
and U17437 (N_17437,N_15984,N_14759);
and U17438 (N_17438,N_14754,N_15899);
nor U17439 (N_17439,N_14436,N_15344);
nor U17440 (N_17440,N_15603,N_14671);
nor U17441 (N_17441,N_14356,N_15135);
nor U17442 (N_17442,N_15488,N_15417);
nor U17443 (N_17443,N_14218,N_14016);
and U17444 (N_17444,N_15868,N_14393);
nand U17445 (N_17445,N_14189,N_14376);
xnor U17446 (N_17446,N_15166,N_14180);
nand U17447 (N_17447,N_15323,N_14502);
nor U17448 (N_17448,N_14704,N_14733);
or U17449 (N_17449,N_14653,N_14820);
xnor U17450 (N_17450,N_15250,N_14944);
nand U17451 (N_17451,N_15179,N_14409);
xor U17452 (N_17452,N_15883,N_15007);
nand U17453 (N_17453,N_15104,N_15755);
nor U17454 (N_17454,N_14973,N_14031);
and U17455 (N_17455,N_15086,N_15198);
and U17456 (N_17456,N_14685,N_15749);
or U17457 (N_17457,N_14039,N_14520);
nand U17458 (N_17458,N_14245,N_15626);
and U17459 (N_17459,N_15677,N_14694);
xor U17460 (N_17460,N_15362,N_14983);
or U17461 (N_17461,N_14260,N_15960);
and U17462 (N_17462,N_14836,N_14816);
nand U17463 (N_17463,N_15673,N_14675);
nand U17464 (N_17464,N_14175,N_14562);
or U17465 (N_17465,N_15236,N_14765);
xnor U17466 (N_17466,N_14482,N_14942);
xnor U17467 (N_17467,N_14538,N_14197);
nand U17468 (N_17468,N_15771,N_14418);
xnor U17469 (N_17469,N_14020,N_15309);
xnor U17470 (N_17470,N_14390,N_15353);
nand U17471 (N_17471,N_15166,N_15019);
nor U17472 (N_17472,N_14994,N_15013);
or U17473 (N_17473,N_14266,N_15506);
xor U17474 (N_17474,N_15741,N_14276);
nor U17475 (N_17475,N_15832,N_15368);
nor U17476 (N_17476,N_14728,N_14513);
xnor U17477 (N_17477,N_14813,N_15529);
nand U17478 (N_17478,N_15618,N_15263);
and U17479 (N_17479,N_15051,N_15873);
nor U17480 (N_17480,N_14644,N_14250);
or U17481 (N_17481,N_14350,N_15999);
xor U17482 (N_17482,N_15422,N_14330);
xor U17483 (N_17483,N_15980,N_15612);
nand U17484 (N_17484,N_14933,N_15624);
or U17485 (N_17485,N_15538,N_15197);
xnor U17486 (N_17486,N_14947,N_15185);
nand U17487 (N_17487,N_15042,N_14783);
nand U17488 (N_17488,N_15176,N_14182);
xor U17489 (N_17489,N_15263,N_14336);
or U17490 (N_17490,N_14482,N_14010);
xor U17491 (N_17491,N_15729,N_14050);
nand U17492 (N_17492,N_15290,N_15695);
and U17493 (N_17493,N_15390,N_14264);
nand U17494 (N_17494,N_14531,N_14424);
and U17495 (N_17495,N_15147,N_15023);
and U17496 (N_17496,N_15321,N_15504);
nand U17497 (N_17497,N_14441,N_14086);
or U17498 (N_17498,N_15032,N_14926);
or U17499 (N_17499,N_14883,N_14858);
xor U17500 (N_17500,N_15711,N_14468);
nor U17501 (N_17501,N_15296,N_14467);
nor U17502 (N_17502,N_14128,N_15863);
xor U17503 (N_17503,N_15059,N_15824);
xor U17504 (N_17504,N_15999,N_15280);
xor U17505 (N_17505,N_15508,N_15216);
and U17506 (N_17506,N_15916,N_15829);
nand U17507 (N_17507,N_15626,N_15016);
or U17508 (N_17508,N_14175,N_15983);
or U17509 (N_17509,N_15668,N_15011);
or U17510 (N_17510,N_15304,N_15152);
nand U17511 (N_17511,N_14671,N_14529);
nand U17512 (N_17512,N_15030,N_15695);
or U17513 (N_17513,N_14509,N_15839);
nor U17514 (N_17514,N_14027,N_14422);
nor U17515 (N_17515,N_14718,N_15626);
nor U17516 (N_17516,N_14841,N_15594);
xnor U17517 (N_17517,N_15543,N_15200);
nor U17518 (N_17518,N_14867,N_14221);
nand U17519 (N_17519,N_15265,N_14686);
or U17520 (N_17520,N_14360,N_14509);
and U17521 (N_17521,N_15521,N_14377);
or U17522 (N_17522,N_15380,N_15652);
and U17523 (N_17523,N_14507,N_14122);
nor U17524 (N_17524,N_14595,N_14998);
xor U17525 (N_17525,N_14775,N_14669);
nand U17526 (N_17526,N_15190,N_15778);
xnor U17527 (N_17527,N_15940,N_15963);
nor U17528 (N_17528,N_14303,N_15229);
nor U17529 (N_17529,N_14586,N_15438);
xor U17530 (N_17530,N_14093,N_15163);
nand U17531 (N_17531,N_14316,N_15739);
and U17532 (N_17532,N_14457,N_15940);
xor U17533 (N_17533,N_14650,N_14150);
and U17534 (N_17534,N_15165,N_15245);
or U17535 (N_17535,N_14174,N_14347);
nor U17536 (N_17536,N_15654,N_14682);
nor U17537 (N_17537,N_14492,N_14664);
nand U17538 (N_17538,N_14635,N_15134);
and U17539 (N_17539,N_15579,N_14390);
nand U17540 (N_17540,N_15487,N_14349);
xor U17541 (N_17541,N_15774,N_14485);
and U17542 (N_17542,N_15923,N_14143);
or U17543 (N_17543,N_15018,N_14009);
xnor U17544 (N_17544,N_15068,N_14333);
or U17545 (N_17545,N_14893,N_15038);
nand U17546 (N_17546,N_15639,N_14043);
nor U17547 (N_17547,N_14271,N_14223);
nand U17548 (N_17548,N_15460,N_15427);
nand U17549 (N_17549,N_14197,N_15865);
nor U17550 (N_17550,N_15469,N_15898);
or U17551 (N_17551,N_15195,N_14904);
or U17552 (N_17552,N_14202,N_15816);
nand U17553 (N_17553,N_15097,N_15339);
xnor U17554 (N_17554,N_14294,N_14096);
or U17555 (N_17555,N_14024,N_15544);
and U17556 (N_17556,N_14545,N_14333);
and U17557 (N_17557,N_14298,N_14578);
xnor U17558 (N_17558,N_14015,N_14179);
and U17559 (N_17559,N_15487,N_14627);
or U17560 (N_17560,N_15819,N_14591);
nor U17561 (N_17561,N_15343,N_15538);
or U17562 (N_17562,N_14150,N_15210);
and U17563 (N_17563,N_14426,N_14919);
xnor U17564 (N_17564,N_15299,N_15198);
and U17565 (N_17565,N_15346,N_15062);
and U17566 (N_17566,N_15579,N_14581);
nor U17567 (N_17567,N_14500,N_14446);
xor U17568 (N_17568,N_14978,N_15193);
and U17569 (N_17569,N_15231,N_14499);
or U17570 (N_17570,N_14393,N_15122);
nor U17571 (N_17571,N_15211,N_15218);
nor U17572 (N_17572,N_14568,N_15343);
and U17573 (N_17573,N_15015,N_15055);
or U17574 (N_17574,N_15815,N_15128);
xnor U17575 (N_17575,N_15126,N_14730);
nand U17576 (N_17576,N_14524,N_14312);
nand U17577 (N_17577,N_14443,N_14524);
and U17578 (N_17578,N_15016,N_14961);
or U17579 (N_17579,N_14962,N_15681);
and U17580 (N_17580,N_14742,N_15851);
and U17581 (N_17581,N_14414,N_14393);
xnor U17582 (N_17582,N_15758,N_14872);
nor U17583 (N_17583,N_14095,N_15668);
or U17584 (N_17584,N_15403,N_15492);
nor U17585 (N_17585,N_14596,N_14487);
or U17586 (N_17586,N_15960,N_15848);
nand U17587 (N_17587,N_15191,N_14053);
xnor U17588 (N_17588,N_14219,N_14916);
and U17589 (N_17589,N_14100,N_14866);
or U17590 (N_17590,N_15004,N_14216);
and U17591 (N_17591,N_15208,N_14724);
xnor U17592 (N_17592,N_15861,N_15315);
xor U17593 (N_17593,N_14593,N_14557);
xnor U17594 (N_17594,N_15880,N_15522);
or U17595 (N_17595,N_14256,N_14357);
or U17596 (N_17596,N_14477,N_15693);
and U17597 (N_17597,N_14670,N_15652);
and U17598 (N_17598,N_14997,N_14482);
nor U17599 (N_17599,N_15659,N_14032);
and U17600 (N_17600,N_14592,N_14535);
xnor U17601 (N_17601,N_14300,N_14154);
nor U17602 (N_17602,N_15663,N_15235);
xnor U17603 (N_17603,N_14009,N_14089);
or U17604 (N_17604,N_14173,N_15829);
xnor U17605 (N_17605,N_15093,N_15507);
nor U17606 (N_17606,N_15116,N_15604);
xnor U17607 (N_17607,N_14273,N_14681);
or U17608 (N_17608,N_14700,N_15514);
or U17609 (N_17609,N_14724,N_15527);
nor U17610 (N_17610,N_14783,N_14706);
and U17611 (N_17611,N_15693,N_15384);
nor U17612 (N_17612,N_15033,N_15868);
nand U17613 (N_17613,N_14119,N_14542);
and U17614 (N_17614,N_15711,N_14246);
nand U17615 (N_17615,N_15382,N_14388);
xnor U17616 (N_17616,N_14208,N_15639);
nand U17617 (N_17617,N_14566,N_14803);
or U17618 (N_17618,N_15601,N_14460);
and U17619 (N_17619,N_14758,N_14459);
nor U17620 (N_17620,N_14489,N_14392);
xnor U17621 (N_17621,N_15055,N_15862);
or U17622 (N_17622,N_14197,N_15598);
nand U17623 (N_17623,N_15014,N_14634);
nor U17624 (N_17624,N_15057,N_15373);
or U17625 (N_17625,N_14492,N_15212);
or U17626 (N_17626,N_14145,N_14762);
nor U17627 (N_17627,N_14342,N_15654);
or U17628 (N_17628,N_15836,N_15625);
and U17629 (N_17629,N_15707,N_15069);
xor U17630 (N_17630,N_14515,N_15278);
or U17631 (N_17631,N_15303,N_14714);
and U17632 (N_17632,N_14806,N_15866);
or U17633 (N_17633,N_14268,N_15402);
xnor U17634 (N_17634,N_15390,N_14526);
nand U17635 (N_17635,N_14873,N_15713);
or U17636 (N_17636,N_15599,N_14415);
or U17637 (N_17637,N_15120,N_15682);
nand U17638 (N_17638,N_15969,N_14393);
nand U17639 (N_17639,N_14194,N_15589);
or U17640 (N_17640,N_14558,N_14095);
or U17641 (N_17641,N_14034,N_15976);
or U17642 (N_17642,N_15345,N_15594);
and U17643 (N_17643,N_14218,N_15989);
xor U17644 (N_17644,N_15115,N_15937);
and U17645 (N_17645,N_14139,N_15347);
and U17646 (N_17646,N_15846,N_14462);
xor U17647 (N_17647,N_15890,N_15879);
or U17648 (N_17648,N_15633,N_15729);
nand U17649 (N_17649,N_15138,N_14129);
nand U17650 (N_17650,N_15187,N_14046);
and U17651 (N_17651,N_14702,N_14130);
or U17652 (N_17652,N_15087,N_14189);
or U17653 (N_17653,N_14926,N_14354);
nor U17654 (N_17654,N_14284,N_15628);
nand U17655 (N_17655,N_14990,N_14777);
nand U17656 (N_17656,N_14723,N_14151);
xor U17657 (N_17657,N_14807,N_14144);
nand U17658 (N_17658,N_14588,N_14465);
and U17659 (N_17659,N_14371,N_14287);
and U17660 (N_17660,N_14656,N_15325);
and U17661 (N_17661,N_15139,N_14441);
nor U17662 (N_17662,N_15646,N_14149);
and U17663 (N_17663,N_14170,N_15151);
and U17664 (N_17664,N_14738,N_14388);
or U17665 (N_17665,N_14662,N_15156);
xor U17666 (N_17666,N_14412,N_15069);
xor U17667 (N_17667,N_14904,N_14038);
and U17668 (N_17668,N_15622,N_14779);
and U17669 (N_17669,N_14452,N_14347);
and U17670 (N_17670,N_14398,N_15021);
xnor U17671 (N_17671,N_15004,N_14930);
or U17672 (N_17672,N_14042,N_15060);
xor U17673 (N_17673,N_15691,N_15939);
or U17674 (N_17674,N_14108,N_15742);
xor U17675 (N_17675,N_14307,N_14142);
and U17676 (N_17676,N_14630,N_15134);
or U17677 (N_17677,N_15703,N_14616);
nand U17678 (N_17678,N_14077,N_14835);
nand U17679 (N_17679,N_15562,N_14522);
nor U17680 (N_17680,N_14115,N_14018);
or U17681 (N_17681,N_14491,N_14461);
nor U17682 (N_17682,N_14713,N_14630);
nor U17683 (N_17683,N_14004,N_15699);
nand U17684 (N_17684,N_14378,N_15783);
xnor U17685 (N_17685,N_14434,N_15171);
xnor U17686 (N_17686,N_14838,N_15738);
xnor U17687 (N_17687,N_14281,N_14600);
xor U17688 (N_17688,N_14897,N_15690);
nor U17689 (N_17689,N_15479,N_14013);
nand U17690 (N_17690,N_14255,N_15253);
nor U17691 (N_17691,N_14850,N_14150);
or U17692 (N_17692,N_14585,N_15238);
and U17693 (N_17693,N_14697,N_15797);
xnor U17694 (N_17694,N_14307,N_15915);
xnor U17695 (N_17695,N_14175,N_15249);
nand U17696 (N_17696,N_14220,N_15703);
xnor U17697 (N_17697,N_14588,N_14287);
nand U17698 (N_17698,N_15570,N_14341);
xor U17699 (N_17699,N_14562,N_14969);
and U17700 (N_17700,N_14017,N_15914);
nand U17701 (N_17701,N_14968,N_14411);
or U17702 (N_17702,N_15001,N_15280);
or U17703 (N_17703,N_14053,N_14472);
nand U17704 (N_17704,N_14875,N_14140);
xor U17705 (N_17705,N_14310,N_14099);
and U17706 (N_17706,N_14590,N_15220);
xor U17707 (N_17707,N_15422,N_14299);
nor U17708 (N_17708,N_14844,N_14542);
nand U17709 (N_17709,N_14096,N_14547);
nand U17710 (N_17710,N_14226,N_15637);
or U17711 (N_17711,N_15670,N_15833);
or U17712 (N_17712,N_14244,N_15244);
and U17713 (N_17713,N_15965,N_14343);
and U17714 (N_17714,N_14010,N_14713);
nor U17715 (N_17715,N_14633,N_14750);
nand U17716 (N_17716,N_15732,N_14808);
and U17717 (N_17717,N_15424,N_14439);
xnor U17718 (N_17718,N_14562,N_15924);
nand U17719 (N_17719,N_14291,N_14319);
and U17720 (N_17720,N_15973,N_14202);
xnor U17721 (N_17721,N_14291,N_14643);
xnor U17722 (N_17722,N_15017,N_15777);
and U17723 (N_17723,N_14226,N_14035);
xnor U17724 (N_17724,N_15023,N_15478);
or U17725 (N_17725,N_15358,N_15134);
and U17726 (N_17726,N_14374,N_15063);
and U17727 (N_17727,N_15589,N_15041);
nor U17728 (N_17728,N_15359,N_14301);
or U17729 (N_17729,N_15514,N_15328);
or U17730 (N_17730,N_14320,N_14951);
and U17731 (N_17731,N_15476,N_14589);
and U17732 (N_17732,N_15769,N_14170);
nor U17733 (N_17733,N_15079,N_15067);
or U17734 (N_17734,N_14649,N_15869);
or U17735 (N_17735,N_15831,N_15714);
and U17736 (N_17736,N_14712,N_14300);
xnor U17737 (N_17737,N_14063,N_15092);
and U17738 (N_17738,N_15578,N_15098);
nor U17739 (N_17739,N_14466,N_15424);
nor U17740 (N_17740,N_15092,N_14020);
xor U17741 (N_17741,N_15365,N_15485);
or U17742 (N_17742,N_15410,N_15548);
and U17743 (N_17743,N_15664,N_14827);
nor U17744 (N_17744,N_14103,N_14059);
xor U17745 (N_17745,N_15617,N_14940);
or U17746 (N_17746,N_15457,N_14927);
and U17747 (N_17747,N_15501,N_14647);
nand U17748 (N_17748,N_14101,N_14015);
nand U17749 (N_17749,N_15908,N_14664);
nand U17750 (N_17750,N_15130,N_15156);
or U17751 (N_17751,N_14143,N_15142);
and U17752 (N_17752,N_14148,N_15968);
xor U17753 (N_17753,N_15429,N_14378);
nor U17754 (N_17754,N_14295,N_15578);
nor U17755 (N_17755,N_15972,N_15169);
nand U17756 (N_17756,N_14867,N_15397);
xor U17757 (N_17757,N_14405,N_15025);
xor U17758 (N_17758,N_15319,N_14274);
nand U17759 (N_17759,N_15556,N_15068);
and U17760 (N_17760,N_14959,N_15580);
nor U17761 (N_17761,N_14749,N_14085);
nand U17762 (N_17762,N_14946,N_15751);
nor U17763 (N_17763,N_15455,N_15840);
or U17764 (N_17764,N_14706,N_15206);
nand U17765 (N_17765,N_15805,N_15986);
nand U17766 (N_17766,N_14917,N_14642);
nand U17767 (N_17767,N_14338,N_15390);
nand U17768 (N_17768,N_15600,N_15500);
xor U17769 (N_17769,N_15061,N_15161);
nor U17770 (N_17770,N_14156,N_14321);
xnor U17771 (N_17771,N_15165,N_15905);
or U17772 (N_17772,N_15408,N_14215);
or U17773 (N_17773,N_14009,N_14805);
xnor U17774 (N_17774,N_15820,N_15981);
nand U17775 (N_17775,N_14842,N_14099);
xnor U17776 (N_17776,N_15301,N_14304);
xnor U17777 (N_17777,N_15224,N_15164);
xnor U17778 (N_17778,N_14258,N_15717);
xor U17779 (N_17779,N_15184,N_14009);
nand U17780 (N_17780,N_15465,N_15805);
nor U17781 (N_17781,N_15160,N_15513);
nand U17782 (N_17782,N_15689,N_14786);
or U17783 (N_17783,N_14355,N_14320);
or U17784 (N_17784,N_14709,N_14233);
xnor U17785 (N_17785,N_15373,N_14002);
nand U17786 (N_17786,N_15413,N_14773);
nor U17787 (N_17787,N_14586,N_14715);
and U17788 (N_17788,N_14938,N_15344);
nand U17789 (N_17789,N_15284,N_14143);
nand U17790 (N_17790,N_15449,N_15208);
xor U17791 (N_17791,N_14978,N_14709);
and U17792 (N_17792,N_14459,N_14173);
nor U17793 (N_17793,N_14904,N_14507);
xnor U17794 (N_17794,N_15132,N_15077);
and U17795 (N_17795,N_15151,N_15607);
xnor U17796 (N_17796,N_15464,N_14636);
and U17797 (N_17797,N_15301,N_14741);
nor U17798 (N_17798,N_15969,N_15434);
nand U17799 (N_17799,N_15573,N_14696);
nor U17800 (N_17800,N_14008,N_14764);
nand U17801 (N_17801,N_15465,N_15506);
and U17802 (N_17802,N_14325,N_14476);
and U17803 (N_17803,N_15980,N_15066);
and U17804 (N_17804,N_15699,N_15355);
nand U17805 (N_17805,N_14798,N_14905);
and U17806 (N_17806,N_14045,N_14625);
nor U17807 (N_17807,N_14429,N_14456);
nand U17808 (N_17808,N_14505,N_15336);
or U17809 (N_17809,N_14315,N_14997);
nor U17810 (N_17810,N_15350,N_14794);
or U17811 (N_17811,N_14315,N_14968);
and U17812 (N_17812,N_14339,N_14455);
and U17813 (N_17813,N_14185,N_15538);
nor U17814 (N_17814,N_15779,N_14072);
xnor U17815 (N_17815,N_14225,N_14014);
nor U17816 (N_17816,N_14363,N_15485);
nand U17817 (N_17817,N_15378,N_15742);
nand U17818 (N_17818,N_14289,N_15233);
and U17819 (N_17819,N_14507,N_14949);
nand U17820 (N_17820,N_14202,N_15488);
nand U17821 (N_17821,N_15387,N_14171);
xor U17822 (N_17822,N_14731,N_15597);
or U17823 (N_17823,N_15272,N_14703);
nand U17824 (N_17824,N_15796,N_14550);
nand U17825 (N_17825,N_14237,N_14969);
xor U17826 (N_17826,N_14748,N_14990);
nand U17827 (N_17827,N_15753,N_15113);
or U17828 (N_17828,N_15497,N_15376);
nor U17829 (N_17829,N_14712,N_14796);
nor U17830 (N_17830,N_14602,N_14691);
nand U17831 (N_17831,N_14562,N_14706);
or U17832 (N_17832,N_14118,N_15745);
xor U17833 (N_17833,N_15022,N_15342);
nand U17834 (N_17834,N_15700,N_15365);
and U17835 (N_17835,N_14250,N_14398);
xor U17836 (N_17836,N_14848,N_15312);
xnor U17837 (N_17837,N_14213,N_15150);
or U17838 (N_17838,N_15276,N_14892);
xor U17839 (N_17839,N_15400,N_15128);
or U17840 (N_17840,N_15113,N_14829);
and U17841 (N_17841,N_15168,N_14604);
xor U17842 (N_17842,N_14495,N_14110);
nand U17843 (N_17843,N_15820,N_14190);
nor U17844 (N_17844,N_14044,N_15809);
and U17845 (N_17845,N_14850,N_15915);
or U17846 (N_17846,N_15684,N_15915);
and U17847 (N_17847,N_14826,N_15517);
xor U17848 (N_17848,N_14367,N_15262);
or U17849 (N_17849,N_14045,N_14666);
or U17850 (N_17850,N_15215,N_14399);
or U17851 (N_17851,N_14551,N_14444);
nand U17852 (N_17852,N_14971,N_14779);
nor U17853 (N_17853,N_14310,N_15665);
xor U17854 (N_17854,N_14084,N_14602);
and U17855 (N_17855,N_15405,N_15237);
nor U17856 (N_17856,N_14047,N_14416);
or U17857 (N_17857,N_14567,N_15751);
and U17858 (N_17858,N_15071,N_15980);
nand U17859 (N_17859,N_15908,N_14835);
nor U17860 (N_17860,N_14091,N_15439);
nand U17861 (N_17861,N_14820,N_15184);
nor U17862 (N_17862,N_15359,N_14885);
and U17863 (N_17863,N_15371,N_14926);
nor U17864 (N_17864,N_15425,N_15433);
xor U17865 (N_17865,N_15457,N_14940);
nor U17866 (N_17866,N_14569,N_15698);
and U17867 (N_17867,N_15011,N_14346);
xor U17868 (N_17868,N_14905,N_15189);
nand U17869 (N_17869,N_15281,N_14756);
and U17870 (N_17870,N_15045,N_15337);
and U17871 (N_17871,N_15690,N_15636);
or U17872 (N_17872,N_14026,N_14311);
xor U17873 (N_17873,N_14066,N_14763);
nor U17874 (N_17874,N_15332,N_14566);
or U17875 (N_17875,N_14221,N_15299);
nand U17876 (N_17876,N_14678,N_14957);
nor U17877 (N_17877,N_15368,N_15443);
or U17878 (N_17878,N_15871,N_14606);
and U17879 (N_17879,N_14548,N_14747);
xnor U17880 (N_17880,N_15001,N_14211);
or U17881 (N_17881,N_15953,N_14104);
or U17882 (N_17882,N_14894,N_14843);
nand U17883 (N_17883,N_14483,N_15387);
or U17884 (N_17884,N_14684,N_14369);
nand U17885 (N_17885,N_14441,N_14482);
xnor U17886 (N_17886,N_15345,N_15446);
nor U17887 (N_17887,N_14888,N_15847);
or U17888 (N_17888,N_15503,N_15373);
xor U17889 (N_17889,N_14909,N_14636);
or U17890 (N_17890,N_14691,N_15080);
nand U17891 (N_17891,N_14323,N_14585);
xnor U17892 (N_17892,N_14529,N_15033);
and U17893 (N_17893,N_15835,N_14440);
nand U17894 (N_17894,N_14379,N_14510);
nor U17895 (N_17895,N_14020,N_15243);
nor U17896 (N_17896,N_15682,N_15152);
and U17897 (N_17897,N_14759,N_15833);
nor U17898 (N_17898,N_15977,N_15620);
or U17899 (N_17899,N_15192,N_14041);
nand U17900 (N_17900,N_15143,N_15329);
nand U17901 (N_17901,N_15899,N_15703);
nand U17902 (N_17902,N_15135,N_14995);
nor U17903 (N_17903,N_15640,N_15351);
or U17904 (N_17904,N_15778,N_15079);
xnor U17905 (N_17905,N_15099,N_14935);
or U17906 (N_17906,N_14326,N_15423);
nand U17907 (N_17907,N_15612,N_14952);
and U17908 (N_17908,N_15084,N_14892);
nor U17909 (N_17909,N_15945,N_15343);
nor U17910 (N_17910,N_14684,N_14249);
and U17911 (N_17911,N_15149,N_15706);
or U17912 (N_17912,N_15987,N_15269);
nor U17913 (N_17913,N_14865,N_14547);
xor U17914 (N_17914,N_15450,N_14935);
nand U17915 (N_17915,N_15644,N_15517);
nor U17916 (N_17916,N_15733,N_15535);
or U17917 (N_17917,N_15739,N_14435);
or U17918 (N_17918,N_15205,N_15109);
and U17919 (N_17919,N_15597,N_15717);
and U17920 (N_17920,N_14965,N_14553);
nor U17921 (N_17921,N_14560,N_15166);
nor U17922 (N_17922,N_14281,N_14551);
and U17923 (N_17923,N_15163,N_15368);
xnor U17924 (N_17924,N_15262,N_14676);
or U17925 (N_17925,N_14576,N_14418);
nor U17926 (N_17926,N_15747,N_14694);
nor U17927 (N_17927,N_15218,N_14624);
nor U17928 (N_17928,N_15655,N_14288);
and U17929 (N_17929,N_15837,N_14538);
nand U17930 (N_17930,N_14635,N_15799);
xnor U17931 (N_17931,N_14519,N_15000);
nand U17932 (N_17932,N_15367,N_15352);
nor U17933 (N_17933,N_15364,N_14413);
nor U17934 (N_17934,N_14640,N_15411);
or U17935 (N_17935,N_15157,N_15022);
or U17936 (N_17936,N_15242,N_15992);
or U17937 (N_17937,N_15470,N_15918);
nand U17938 (N_17938,N_14022,N_15528);
nand U17939 (N_17939,N_14285,N_14394);
xnor U17940 (N_17940,N_14150,N_15403);
and U17941 (N_17941,N_15280,N_15902);
nand U17942 (N_17942,N_15870,N_14448);
and U17943 (N_17943,N_15196,N_14598);
nor U17944 (N_17944,N_14158,N_14409);
xor U17945 (N_17945,N_15216,N_15511);
nor U17946 (N_17946,N_14954,N_15662);
and U17947 (N_17947,N_14934,N_14074);
xor U17948 (N_17948,N_15479,N_15367);
xor U17949 (N_17949,N_15867,N_15035);
xor U17950 (N_17950,N_14893,N_14753);
or U17951 (N_17951,N_15620,N_14180);
nand U17952 (N_17952,N_14130,N_14712);
nor U17953 (N_17953,N_15546,N_15600);
nand U17954 (N_17954,N_14737,N_14493);
nor U17955 (N_17955,N_14793,N_14459);
nand U17956 (N_17956,N_14238,N_14904);
nand U17957 (N_17957,N_15679,N_15609);
and U17958 (N_17958,N_14854,N_15786);
xnor U17959 (N_17959,N_15457,N_14332);
xnor U17960 (N_17960,N_15883,N_15142);
and U17961 (N_17961,N_15079,N_15326);
nand U17962 (N_17962,N_15205,N_15719);
xnor U17963 (N_17963,N_15932,N_15737);
nand U17964 (N_17964,N_14006,N_14338);
or U17965 (N_17965,N_14015,N_14242);
xor U17966 (N_17966,N_15274,N_14955);
or U17967 (N_17967,N_14386,N_14762);
or U17968 (N_17968,N_14747,N_15689);
xnor U17969 (N_17969,N_14858,N_14760);
nand U17970 (N_17970,N_15936,N_14118);
and U17971 (N_17971,N_15735,N_15111);
nand U17972 (N_17972,N_15686,N_15896);
and U17973 (N_17973,N_14419,N_14114);
xor U17974 (N_17974,N_15250,N_14671);
xor U17975 (N_17975,N_14767,N_14474);
xor U17976 (N_17976,N_15983,N_14345);
nor U17977 (N_17977,N_15259,N_14479);
nor U17978 (N_17978,N_14815,N_14665);
or U17979 (N_17979,N_14782,N_15326);
and U17980 (N_17980,N_15599,N_15935);
nor U17981 (N_17981,N_14901,N_14380);
or U17982 (N_17982,N_15488,N_14861);
and U17983 (N_17983,N_14359,N_14785);
xnor U17984 (N_17984,N_14129,N_14940);
xnor U17985 (N_17985,N_14349,N_15207);
nand U17986 (N_17986,N_14615,N_14720);
and U17987 (N_17987,N_15996,N_15783);
xnor U17988 (N_17988,N_15902,N_14557);
nor U17989 (N_17989,N_15951,N_14681);
or U17990 (N_17990,N_14689,N_14302);
or U17991 (N_17991,N_15357,N_14005);
xnor U17992 (N_17992,N_15078,N_14359);
or U17993 (N_17993,N_15790,N_14305);
nand U17994 (N_17994,N_15280,N_15881);
nor U17995 (N_17995,N_14989,N_15865);
nor U17996 (N_17996,N_14352,N_14144);
nor U17997 (N_17997,N_15468,N_15289);
nor U17998 (N_17998,N_15707,N_15351);
nor U17999 (N_17999,N_15026,N_15162);
xnor U18000 (N_18000,N_16595,N_17142);
or U18001 (N_18001,N_17128,N_17503);
and U18002 (N_18002,N_16184,N_17667);
or U18003 (N_18003,N_16265,N_16285);
nand U18004 (N_18004,N_16131,N_16896);
nor U18005 (N_18005,N_16474,N_16255);
xnor U18006 (N_18006,N_17624,N_16885);
nor U18007 (N_18007,N_17760,N_16149);
nand U18008 (N_18008,N_16738,N_16725);
nand U18009 (N_18009,N_17119,N_16127);
xnor U18010 (N_18010,N_16205,N_17860);
xor U18011 (N_18011,N_17429,N_16855);
and U18012 (N_18012,N_17514,N_16552);
nand U18013 (N_18013,N_16578,N_17446);
xor U18014 (N_18014,N_17932,N_16848);
nand U18015 (N_18015,N_17013,N_17647);
nor U18016 (N_18016,N_16555,N_16367);
xnor U18017 (N_18017,N_16527,N_16816);
and U18018 (N_18018,N_17071,N_16806);
and U18019 (N_18019,N_17536,N_16753);
xor U18020 (N_18020,N_16280,N_16424);
nor U18021 (N_18021,N_17234,N_16965);
nor U18022 (N_18022,N_16530,N_17072);
or U18023 (N_18023,N_17088,N_17131);
nor U18024 (N_18024,N_17347,N_16465);
and U18025 (N_18025,N_17442,N_16640);
and U18026 (N_18026,N_16650,N_16894);
nand U18027 (N_18027,N_17901,N_17517);
or U18028 (N_18028,N_17688,N_16204);
nand U18029 (N_18029,N_17036,N_17921);
xnor U18030 (N_18030,N_16931,N_17318);
nor U18031 (N_18031,N_17525,N_17368);
and U18032 (N_18032,N_17462,N_17965);
and U18033 (N_18033,N_16416,N_17610);
and U18034 (N_18034,N_16408,N_17654);
xnor U18035 (N_18035,N_17835,N_17244);
nand U18036 (N_18036,N_17821,N_17376);
nor U18037 (N_18037,N_17896,N_16322);
and U18038 (N_18038,N_17478,N_16443);
nand U18039 (N_18039,N_17951,N_16203);
nor U18040 (N_18040,N_16202,N_16976);
nand U18041 (N_18041,N_17053,N_16063);
xnor U18042 (N_18042,N_16318,N_16981);
nand U18043 (N_18043,N_16395,N_16256);
xnor U18044 (N_18044,N_16351,N_16475);
or U18045 (N_18045,N_16073,N_17355);
xor U18046 (N_18046,N_17962,N_17634);
or U18047 (N_18047,N_17162,N_17192);
nor U18048 (N_18048,N_16244,N_16150);
nand U18049 (N_18049,N_17201,N_17778);
and U18050 (N_18050,N_17764,N_17326);
and U18051 (N_18051,N_16748,N_17532);
nand U18052 (N_18052,N_16226,N_17285);
or U18053 (N_18053,N_16636,N_17560);
xor U18054 (N_18054,N_16476,N_16959);
and U18055 (N_18055,N_17362,N_17475);
xor U18056 (N_18056,N_17351,N_16009);
nand U18057 (N_18057,N_17570,N_17078);
and U18058 (N_18058,N_17676,N_16145);
and U18059 (N_18059,N_16752,N_17440);
xnor U18060 (N_18060,N_17000,N_17976);
and U18061 (N_18061,N_16935,N_16167);
nor U18062 (N_18062,N_17884,N_16209);
or U18063 (N_18063,N_17613,N_17887);
xnor U18064 (N_18064,N_16000,N_16100);
nand U18065 (N_18065,N_17695,N_16524);
nor U18066 (N_18066,N_16308,N_16215);
nor U18067 (N_18067,N_16767,N_16891);
or U18068 (N_18068,N_16470,N_16034);
nand U18069 (N_18069,N_17450,N_16397);
nand U18070 (N_18070,N_17200,N_17196);
and U18071 (N_18071,N_17328,N_17158);
xnor U18072 (N_18072,N_16220,N_17199);
nor U18073 (N_18073,N_17081,N_16511);
xnor U18074 (N_18074,N_17419,N_17424);
nor U18075 (N_18075,N_17639,N_16197);
nand U18076 (N_18076,N_16594,N_17674);
and U18077 (N_18077,N_17578,N_17390);
xor U18078 (N_18078,N_17495,N_17793);
nand U18079 (N_18079,N_17227,N_17294);
nor U18080 (N_18080,N_17255,N_17640);
or U18081 (N_18081,N_16386,N_16573);
and U18082 (N_18082,N_17319,N_16104);
and U18083 (N_18083,N_16022,N_17261);
xnor U18084 (N_18084,N_16579,N_16762);
xnor U18085 (N_18085,N_17470,N_16529);
nor U18086 (N_18086,N_16460,N_16320);
xnor U18087 (N_18087,N_16082,N_16996);
or U18088 (N_18088,N_17927,N_16638);
xor U18089 (N_18089,N_16958,N_16795);
nand U18090 (N_18090,N_16512,N_16764);
xor U18091 (N_18091,N_17739,N_16080);
and U18092 (N_18092,N_16301,N_16381);
nand U18093 (N_18093,N_17248,N_17744);
xor U18094 (N_18094,N_16742,N_17147);
nand U18095 (N_18095,N_16405,N_17477);
nand U18096 (N_18096,N_16309,N_16939);
xnor U18097 (N_18097,N_16757,N_17980);
nand U18098 (N_18098,N_17191,N_17480);
nand U18099 (N_18099,N_17689,N_16562);
xor U18100 (N_18100,N_16102,N_16334);
nor U18101 (N_18101,N_16542,N_16263);
xnor U18102 (N_18102,N_17183,N_16355);
and U18103 (N_18103,N_16856,N_17505);
and U18104 (N_18104,N_16012,N_16124);
or U18105 (N_18105,N_16923,N_16081);
or U18106 (N_18106,N_17970,N_17742);
nand U18107 (N_18107,N_16766,N_17839);
nor U18108 (N_18108,N_17543,N_17338);
xor U18109 (N_18109,N_16600,N_17583);
xnor U18110 (N_18110,N_17703,N_16982);
nor U18111 (N_18111,N_16793,N_16175);
nor U18112 (N_18112,N_17267,N_16791);
nand U18113 (N_18113,N_17940,N_17037);
and U18114 (N_18114,N_16781,N_16566);
nand U18115 (N_18115,N_17637,N_17763);
xnor U18116 (N_18116,N_17912,N_17762);
and U18117 (N_18117,N_17611,N_17410);
or U18118 (N_18118,N_17116,N_17311);
or U18119 (N_18119,N_17367,N_17207);
or U18120 (N_18120,N_17213,N_16754);
nor U18121 (N_18121,N_16664,N_16517);
nor U18122 (N_18122,N_17862,N_17672);
nand U18123 (N_18123,N_16974,N_17723);
or U18124 (N_18124,N_16143,N_16484);
xor U18125 (N_18125,N_16788,N_17915);
and U18126 (N_18126,N_17365,N_16444);
xor U18127 (N_18127,N_16151,N_16042);
nand U18128 (N_18128,N_17902,N_16735);
xnor U18129 (N_18129,N_17516,N_17945);
nor U18130 (N_18130,N_16006,N_16553);
nor U18131 (N_18131,N_17774,N_17299);
nor U18132 (N_18132,N_16048,N_17504);
and U18133 (N_18133,N_16087,N_17799);
nor U18134 (N_18134,N_17729,N_17321);
xnor U18135 (N_18135,N_17603,N_16119);
nand U18136 (N_18136,N_17057,N_17794);
and U18137 (N_18137,N_16538,N_16148);
nand U18138 (N_18138,N_17435,N_16704);
nand U18139 (N_18139,N_17087,N_17469);
nand U18140 (N_18140,N_16654,N_16147);
xnor U18141 (N_18141,N_16350,N_16930);
nor U18142 (N_18142,N_17448,N_16259);
nor U18143 (N_18143,N_17911,N_17892);
or U18144 (N_18144,N_16967,N_17768);
or U18145 (N_18145,N_16125,N_17609);
nand U18146 (N_18146,N_17079,N_17974);
xnor U18147 (N_18147,N_16095,N_16239);
nand U18148 (N_18148,N_16294,N_17206);
nand U18149 (N_18149,N_16633,N_17716);
and U18150 (N_18150,N_16266,N_16647);
or U18151 (N_18151,N_16665,N_17378);
nand U18152 (N_18152,N_16356,N_16372);
nand U18153 (N_18153,N_17230,N_17264);
and U18154 (N_18154,N_16845,N_17414);
nor U18155 (N_18155,N_16477,N_17222);
or U18156 (N_18156,N_17956,N_17101);
and U18157 (N_18157,N_16488,N_17841);
and U18158 (N_18158,N_16260,N_17784);
xor U18159 (N_18159,N_16419,N_16662);
xor U18160 (N_18160,N_16839,N_16606);
and U18161 (N_18161,N_16236,N_17738);
or U18162 (N_18162,N_17132,N_17562);
nand U18163 (N_18163,N_17075,N_17698);
xor U18164 (N_18164,N_16522,N_16815);
nor U18165 (N_18165,N_16956,N_17858);
and U18166 (N_18166,N_17095,N_16655);
xnor U18167 (N_18167,N_16669,N_17882);
and U18168 (N_18168,N_16780,N_16380);
and U18169 (N_18169,N_16980,N_16347);
nand U18170 (N_18170,N_17052,N_16067);
or U18171 (N_18171,N_17467,N_17438);
xor U18172 (N_18172,N_17541,N_16937);
and U18173 (N_18173,N_17046,N_17530);
nand U18174 (N_18174,N_17117,N_17850);
and U18175 (N_18175,N_17341,N_17907);
and U18176 (N_18176,N_17169,N_16548);
xnor U18177 (N_18177,N_16534,N_17812);
nor U18178 (N_18178,N_17682,N_16375);
or U18179 (N_18179,N_17418,N_17312);
xnor U18180 (N_18180,N_16758,N_16680);
and U18181 (N_18181,N_16195,N_16106);
nand U18182 (N_18182,N_16770,N_17831);
and U18183 (N_18183,N_17937,N_17398);
nor U18184 (N_18184,N_17310,N_17969);
nor U18185 (N_18185,N_17822,N_17387);
and U18186 (N_18186,N_17651,N_16139);
nand U18187 (N_18187,N_17944,N_17662);
and U18188 (N_18188,N_17186,N_16394);
nand U18189 (N_18189,N_17967,N_16952);
xnor U18190 (N_18190,N_17681,N_17174);
or U18191 (N_18191,N_16545,N_17084);
xnor U18192 (N_18192,N_16450,N_17515);
nand U18193 (N_18193,N_16805,N_16178);
and U18194 (N_18194,N_17719,N_16155);
or U18195 (N_18195,N_17995,N_17224);
and U18196 (N_18196,N_16506,N_17718);
xor U18197 (N_18197,N_17500,N_17752);
and U18198 (N_18198,N_17332,N_16036);
nand U18199 (N_18199,N_16218,N_17291);
xor U18200 (N_18200,N_16064,N_16298);
nand U18201 (N_18201,N_17041,N_17823);
nor U18202 (N_18202,N_17648,N_16154);
nand U18203 (N_18203,N_17804,N_16532);
or U18204 (N_18204,N_16072,N_16508);
nand U18205 (N_18205,N_17371,N_16363);
xor U18206 (N_18206,N_17109,N_17876);
or U18207 (N_18207,N_17096,N_16843);
xnor U18208 (N_18208,N_16188,N_16132);
nand U18209 (N_18209,N_17272,N_16570);
xor U18210 (N_18210,N_17628,N_16249);
nor U18211 (N_18211,N_16688,N_17342);
or U18212 (N_18212,N_16797,N_16851);
xor U18213 (N_18213,N_17148,N_17796);
nand U18214 (N_18214,N_16040,N_16702);
nand U18215 (N_18215,N_17614,N_16520);
or U18216 (N_18216,N_16467,N_17406);
and U18217 (N_18217,N_17528,N_16645);
and U18218 (N_18218,N_16019,N_17849);
or U18219 (N_18219,N_16163,N_17020);
xnor U18220 (N_18220,N_16317,N_16238);
nor U18221 (N_18221,N_17030,N_17021);
and U18222 (N_18222,N_16964,N_17577);
or U18223 (N_18223,N_17687,N_17430);
nor U18224 (N_18224,N_16761,N_16993);
and U18225 (N_18225,N_17722,N_17670);
nor U18226 (N_18226,N_16228,N_16369);
or U18227 (N_18227,N_16101,N_16945);
nor U18228 (N_18228,N_16133,N_16246);
xor U18229 (N_18229,N_16326,N_16768);
and U18230 (N_18230,N_17409,N_16316);
xnor U18231 (N_18231,N_17236,N_16804);
nand U18232 (N_18232,N_17708,N_17276);
xor U18233 (N_18233,N_17444,N_17391);
nand U18234 (N_18234,N_16707,N_17114);
and U18235 (N_18235,N_17608,N_16635);
nor U18236 (N_18236,N_17431,N_17066);
or U18237 (N_18237,N_17950,N_16021);
or U18238 (N_18238,N_17226,N_16617);
and U18239 (N_18239,N_16271,N_16303);
and U18240 (N_18240,N_17059,N_16389);
nor U18241 (N_18241,N_17568,N_17173);
nand U18242 (N_18242,N_16750,N_17949);
nand U18243 (N_18243,N_16359,N_16947);
nor U18244 (N_18244,N_16050,N_17298);
and U18245 (N_18245,N_16212,N_17212);
nand U18246 (N_18246,N_16927,N_17994);
or U18247 (N_18247,N_17238,N_17049);
nand U18248 (N_18248,N_17315,N_17552);
or U18249 (N_18249,N_16733,N_16737);
nand U18250 (N_18250,N_17653,N_17243);
or U18251 (N_18251,N_17463,N_16897);
and U18252 (N_18252,N_16504,N_17566);
and U18253 (N_18253,N_16300,N_17171);
and U18254 (N_18254,N_17385,N_17141);
nand U18255 (N_18255,N_17352,N_17237);
and U18256 (N_18256,N_16018,N_17874);
and U18257 (N_18257,N_16189,N_16975);
xor U18258 (N_18258,N_16144,N_17537);
xnor U18259 (N_18259,N_17957,N_17220);
or U18260 (N_18260,N_17554,N_17880);
or U18261 (N_18261,N_16518,N_17557);
nor U18262 (N_18262,N_17485,N_16473);
xnor U18263 (N_18263,N_17677,N_16599);
nor U18264 (N_18264,N_16321,N_16091);
xor U18265 (N_18265,N_16948,N_16810);
xor U18266 (N_18266,N_17824,N_16920);
and U18267 (N_18267,N_17612,N_17643);
nor U18268 (N_18268,N_16113,N_16516);
or U18269 (N_18269,N_16463,N_16830);
xnor U18270 (N_18270,N_16686,N_17425);
or U18271 (N_18271,N_16963,N_16028);
nand U18272 (N_18272,N_17520,N_17591);
and U18273 (N_18273,N_17073,N_16284);
or U18274 (N_18274,N_17426,N_17999);
and U18275 (N_18275,N_16961,N_17184);
xor U18276 (N_18276,N_17179,N_17403);
or U18277 (N_18277,N_16162,N_16052);
and U18278 (N_18278,N_17713,N_16016);
or U18279 (N_18279,N_16357,N_16418);
xor U18280 (N_18280,N_16201,N_16344);
nor U18281 (N_18281,N_17094,N_16245);
nand U18282 (N_18282,N_16934,N_16279);
nor U18283 (N_18283,N_16850,N_16017);
and U18284 (N_18284,N_17534,N_17345);
nand U18285 (N_18285,N_16916,N_16437);
xor U18286 (N_18286,N_17407,N_16602);
nand U18287 (N_18287,N_16786,N_17788);
xnor U18288 (N_18288,N_17456,N_17211);
xnor U18289 (N_18289,N_17655,N_16448);
nor U18290 (N_18290,N_16105,N_17535);
nand U18291 (N_18291,N_16242,N_17549);
or U18292 (N_18292,N_16728,N_16718);
or U18293 (N_18293,N_16183,N_16071);
nor U18294 (N_18294,N_17010,N_16924);
or U18295 (N_18295,N_16865,N_16581);
or U18296 (N_18296,N_16402,N_17806);
xor U18297 (N_18297,N_16660,N_17130);
or U18298 (N_18298,N_17394,N_17574);
xor U18299 (N_18299,N_16466,N_16953);
and U18300 (N_18300,N_16248,N_17437);
xnor U18301 (N_18301,N_17558,N_16898);
xnor U18302 (N_18302,N_17089,N_16694);
nor U18303 (N_18303,N_16940,N_16565);
and U18304 (N_18304,N_16293,N_17451);
nand U18305 (N_18305,N_16447,N_17496);
nor U18306 (N_18306,N_16421,N_16099);
or U18307 (N_18307,N_17547,N_16888);
or U18308 (N_18308,N_17623,N_16333);
and U18309 (N_18309,N_16656,N_16305);
and U18310 (N_18310,N_16751,N_17218);
and U18311 (N_18311,N_17068,N_16783);
nand U18312 (N_18312,N_17331,N_16563);
nor U18313 (N_18313,N_17984,N_17472);
or U18314 (N_18314,N_16904,N_16486);
nand U18315 (N_18315,N_17313,N_17616);
and U18316 (N_18316,N_17193,N_17922);
xnor U18317 (N_18317,N_16663,N_16746);
and U18318 (N_18318,N_17559,N_17930);
or U18319 (N_18319,N_16169,N_16391);
or U18320 (N_18320,N_16196,N_17625);
or U18321 (N_18321,N_17097,N_17959);
and U18322 (N_18322,N_16313,N_17303);
nand U18323 (N_18323,N_16023,N_17777);
or U18324 (N_18324,N_17971,N_16564);
and U18325 (N_18325,N_16682,N_16229);
or U18326 (N_18326,N_16921,N_16110);
or U18327 (N_18327,N_17513,N_16960);
xnor U18328 (N_18328,N_16270,N_16510);
xnor U18329 (N_18329,N_16800,N_17697);
or U18330 (N_18330,N_17601,N_17293);
xnor U18331 (N_18331,N_16612,N_16059);
xor U18332 (N_18332,N_16053,N_17527);
or U18333 (N_18333,N_17942,N_17404);
nand U18334 (N_18334,N_16560,N_17575);
xnor U18335 (N_18335,N_17917,N_16706);
xnor U18336 (N_18336,N_16319,N_16708);
or U18337 (N_18337,N_17208,N_17960);
xnor U18338 (N_18338,N_17282,N_16991);
xor U18339 (N_18339,N_17675,N_17747);
nand U18340 (N_18340,N_17666,N_17910);
and U18341 (N_18341,N_16684,N_17275);
xnor U18342 (N_18342,N_17510,N_16900);
nand U18343 (N_18343,N_17709,N_16451);
nor U18344 (N_18344,N_17808,N_16464);
nand U18345 (N_18345,N_17606,N_16601);
nor U18346 (N_18346,N_16299,N_17065);
nor U18347 (N_18347,N_17811,N_17900);
nor U18348 (N_18348,N_17617,N_16013);
or U18349 (N_18349,N_17359,N_17242);
nand U18350 (N_18350,N_16526,N_17443);
or U18351 (N_18351,N_17402,N_16364);
xor U18352 (N_18352,N_17754,N_17413);
nor U18353 (N_18353,N_16371,N_16138);
or U18354 (N_18354,N_17644,N_17353);
and U18355 (N_18355,N_16247,N_17361);
nand U18356 (N_18356,N_16613,N_16509);
nor U18357 (N_18357,N_17767,N_17098);
nand U18358 (N_18358,N_17863,N_17813);
or U18359 (N_18359,N_16373,N_16908);
xnor U18360 (N_18360,N_17724,N_16035);
and U18361 (N_18361,N_17953,N_17107);
nand U18362 (N_18362,N_17987,N_16586);
nor U18363 (N_18363,N_17092,N_16061);
xnor U18364 (N_18364,N_16076,N_17473);
or U18365 (N_18365,N_16918,N_16871);
xor U18366 (N_18366,N_16692,N_16241);
or U18367 (N_18367,N_17569,N_17167);
nor U18368 (N_18368,N_16648,N_17388);
or U18369 (N_18369,N_16584,N_16025);
nor U18370 (N_18370,N_16734,N_16157);
nand U18371 (N_18371,N_16668,N_17320);
and U18372 (N_18372,N_17453,N_17110);
xor U18373 (N_18373,N_17205,N_17787);
nor U18374 (N_18374,N_17460,N_17792);
or U18375 (N_18375,N_16041,N_16938);
xor U18376 (N_18376,N_16409,N_16576);
or U18377 (N_18377,N_16610,N_17306);
nor U18378 (N_18378,N_17899,N_17112);
xor U18379 (N_18379,N_17363,N_16130);
and U18380 (N_18380,N_16785,N_16010);
or U18381 (N_18381,N_16630,N_17017);
and U18382 (N_18382,N_16075,N_17025);
or U18383 (N_18383,N_17690,N_17300);
and U18384 (N_18384,N_17563,N_17157);
nor U18385 (N_18385,N_16114,N_16970);
xnor U18386 (N_18386,N_16875,N_17152);
and U18387 (N_18387,N_17122,N_16158);
nor U18388 (N_18388,N_17358,N_16026);
and U18389 (N_18389,N_16343,N_17731);
xnor U18390 (N_18390,N_16365,N_17176);
nor U18391 (N_18391,N_16066,N_17405);
or U18392 (N_18392,N_17124,N_16252);
nor U18393 (N_18393,N_17604,N_17581);
xnor U18394 (N_18394,N_17859,N_17125);
xor U18395 (N_18395,N_17877,N_16643);
xor U18396 (N_18396,N_17062,N_17786);
xnor U18397 (N_18397,N_16603,N_16760);
nand U18398 (N_18398,N_17836,N_16911);
and U18399 (N_18399,N_16759,N_17782);
or U18400 (N_18400,N_16291,N_17271);
nor U18401 (N_18401,N_17684,N_16136);
xor U18402 (N_18402,N_17228,N_17343);
nand U18403 (N_18403,N_17187,N_16596);
xor U18404 (N_18404,N_16146,N_17870);
nor U18405 (N_18405,N_17381,N_17465);
and U18406 (N_18406,N_16598,N_17329);
nand U18407 (N_18407,N_17985,N_17780);
xor U18408 (N_18408,N_17364,N_16813);
xnor U18409 (N_18409,N_17177,N_16919);
xnor U18410 (N_18410,N_17621,N_16834);
nand U18411 (N_18411,N_16832,N_17597);
or U18412 (N_18412,N_16176,N_16628);
nor U18413 (N_18413,N_16634,N_17016);
and U18414 (N_18414,N_16847,N_17254);
nor U18415 (N_18415,N_17233,N_17753);
or U18416 (N_18416,N_17576,N_16886);
nand U18417 (N_18417,N_17502,N_16452);
xnor U18418 (N_18418,N_17375,N_16112);
xor U18419 (N_18419,N_17416,N_16852);
and U18420 (N_18420,N_17216,N_16393);
or U18421 (N_18421,N_16696,N_17531);
xnor U18422 (N_18422,N_17631,N_16868);
xor U18423 (N_18423,N_16749,N_16282);
xor U18424 (N_18424,N_17638,N_17867);
xor U18425 (N_18425,N_16987,N_16056);
and U18426 (N_18426,N_17123,N_16887);
nand U18427 (N_18427,N_16253,N_16156);
or U18428 (N_18428,N_16121,N_16722);
xor U18429 (N_18429,N_17323,N_16362);
xor U18430 (N_18430,N_16611,N_16949);
xor U18431 (N_18431,N_17166,N_16128);
nor U18432 (N_18432,N_17652,N_16547);
nor U18433 (N_18433,N_17428,N_17120);
or U18434 (N_18434,N_16739,N_17251);
and U18435 (N_18435,N_16942,N_16328);
and U18436 (N_18436,N_17727,N_17290);
nor U18437 (N_18437,N_16103,N_16926);
xnor U18438 (N_18438,N_17449,N_16336);
nor U18439 (N_18439,N_16011,N_17197);
and U18440 (N_18440,N_17512,N_16427);
xnor U18441 (N_18441,N_16337,N_16191);
or U18442 (N_18442,N_16497,N_17439);
xor U18443 (N_18443,N_16626,N_16455);
or U18444 (N_18444,N_16901,N_16062);
nand U18445 (N_18445,N_16377,N_16186);
and U18446 (N_18446,N_17397,N_16962);
or U18447 (N_18447,N_16556,N_16994);
nor U18448 (N_18448,N_16107,N_17399);
xnor U18449 (N_18449,N_16194,N_17339);
nand U18450 (N_18450,N_16666,N_16462);
xnor U18451 (N_18451,N_17873,N_17573);
nand U18452 (N_18452,N_16430,N_16999);
or U18453 (N_18453,N_17524,N_17668);
nor U18454 (N_18454,N_17814,N_17348);
and U18455 (N_18455,N_17153,N_16230);
and U18456 (N_18456,N_16514,N_17337);
nor U18457 (N_18457,N_16479,N_16237);
or U18458 (N_18458,N_16142,N_17033);
nand U18459 (N_18459,N_17801,N_17189);
nor U18460 (N_18460,N_17529,N_17746);
xnor U18461 (N_18461,N_17400,N_17269);
nor U18462 (N_18462,N_17393,N_16033);
xnor U18463 (N_18463,N_16232,N_16172);
xor U18464 (N_18464,N_17471,N_17802);
or U18465 (N_18465,N_17305,N_16801);
nor U18466 (N_18466,N_17113,N_16833);
nor U18467 (N_18467,N_16401,N_17544);
xnor U18468 (N_18468,N_17834,N_16480);
or U18469 (N_18469,N_16472,N_16727);
and U18470 (N_18470,N_17245,N_16597);
nor U18471 (N_18471,N_16623,N_16705);
xnor U18472 (N_18472,N_16436,N_16903);
or U18473 (N_18473,N_17050,N_16446);
or U18474 (N_18474,N_16489,N_16312);
nand U18475 (N_18475,N_16039,N_17249);
and U18476 (N_18476,N_17977,N_17629);
nand U18477 (N_18477,N_16568,N_16854);
nor U18478 (N_18478,N_16681,N_16951);
nand U18479 (N_18479,N_17572,N_17004);
or U18480 (N_18480,N_16348,N_16358);
and U18481 (N_18481,N_16881,N_17856);
nand U18482 (N_18482,N_17993,N_16429);
nand U18483 (N_18483,N_16030,N_17555);
nand U18484 (N_18484,N_17454,N_17307);
xor U18485 (N_18485,N_16928,N_16907);
or U18486 (N_18486,N_16714,N_16159);
nor U18487 (N_18487,N_17182,N_17235);
xnor U18488 (N_18488,N_16792,N_16413);
nor U18489 (N_18489,N_16917,N_17587);
and U18490 (N_18490,N_17487,N_17539);
nand U18491 (N_18491,N_16292,N_17165);
and U18492 (N_18492,N_17024,N_17015);
and U18493 (N_18493,N_17292,N_17336);
or U18494 (N_18494,N_17240,N_16272);
nand U18495 (N_18495,N_17659,N_17002);
nor U18496 (N_18496,N_16483,N_16278);
or U18497 (N_18497,N_17086,N_16281);
xnor U18498 (N_18498,N_16307,N_16659);
or U18499 (N_18499,N_17284,N_16608);
and U18500 (N_18500,N_17357,N_16857);
and U18501 (N_18501,N_17370,N_17898);
xor U18502 (N_18502,N_17714,N_17889);
nor U18503 (N_18503,N_17408,N_16382);
nor U18504 (N_18504,N_17934,N_17933);
xor U18505 (N_18505,N_17210,N_16554);
nor U18506 (N_18506,N_17734,N_16240);
xor U18507 (N_18507,N_17458,N_17476);
nor U18508 (N_18508,N_16997,N_17180);
or U18509 (N_18509,N_17966,N_17209);
nand U18510 (N_18510,N_16743,N_17006);
nor U18511 (N_18511,N_16153,N_17441);
nand U18512 (N_18512,N_17720,N_17302);
nand U18513 (N_18513,N_17296,N_17461);
and U18514 (N_18514,N_17947,N_16674);
xnor U18515 (N_18515,N_16763,N_16933);
xnor U18516 (N_18516,N_17711,N_17997);
nor U18517 (N_18517,N_17257,N_16955);
xor U18518 (N_18518,N_17975,N_16615);
nor U18519 (N_18519,N_17386,N_16880);
xor U18520 (N_18520,N_16863,N_16721);
nor U18521 (N_18521,N_17871,N_16093);
nor U18522 (N_18522,N_16097,N_16528);
and U18523 (N_18523,N_17260,N_17149);
and U18524 (N_18524,N_17526,N_17875);
xnor U18525 (N_18525,N_16929,N_16495);
xnor U18526 (N_18526,N_16619,N_16164);
nand U18527 (N_18527,N_17241,N_17145);
and U18528 (N_18528,N_16776,N_16315);
and U18529 (N_18529,N_17693,N_17519);
and U18530 (N_18530,N_17935,N_17826);
nand U18531 (N_18531,N_16211,N_16989);
nor U18532 (N_18532,N_17853,N_17288);
nand U18533 (N_18533,N_17038,N_17350);
and U18534 (N_18534,N_17795,N_17333);
xnor U18535 (N_18535,N_17783,N_16435);
xnor U18536 (N_18536,N_17736,N_17061);
and U18537 (N_18537,N_16841,N_16689);
and U18538 (N_18538,N_17175,N_17383);
nor U18539 (N_18539,N_16616,N_17929);
or U18540 (N_18540,N_17595,N_16001);
nand U18541 (N_18541,N_17818,N_17973);
xnor U18542 (N_18542,N_17080,N_16914);
nand U18543 (N_18543,N_16620,N_17815);
nor U18544 (N_18544,N_16789,N_16837);
xor U18545 (N_18545,N_16227,N_17263);
and U18546 (N_18546,N_17646,N_17048);
or U18547 (N_18547,N_16677,N_17567);
or U18548 (N_18548,N_17830,N_16539);
and U18549 (N_18549,N_16079,N_16494);
and U18550 (N_18550,N_16944,N_17384);
or U18551 (N_18551,N_16507,N_16049);
nor U18552 (N_18552,N_17770,N_17256);
nand U18553 (N_18553,N_17489,N_17420);
nand U18554 (N_18554,N_17982,N_17214);
or U18555 (N_18555,N_16353,N_17215);
or U18556 (N_18556,N_16166,N_17981);
xor U18557 (N_18557,N_16206,N_17642);
nand U18558 (N_18558,N_16161,N_17138);
nand U18559 (N_18559,N_16014,N_17908);
nand U18560 (N_18560,N_16607,N_17317);
xnor U18561 (N_18561,N_16913,N_17219);
or U18562 (N_18562,N_16137,N_17968);
nor U18563 (N_18563,N_16024,N_17588);
or U18564 (N_18564,N_17630,N_17584);
xnor U18565 (N_18565,N_16029,N_16740);
nor U18566 (N_18566,N_16192,N_17492);
nor U18567 (N_18567,N_17895,N_17809);
and U18568 (N_18568,N_17730,N_16811);
nor U18569 (N_18569,N_16331,N_17955);
nor U18570 (N_18570,N_17304,N_16314);
nand U18571 (N_18571,N_17106,N_16712);
nand U18572 (N_18572,N_17958,N_16902);
and U18573 (N_18573,N_17607,N_17926);
nor U18574 (N_18574,N_17599,N_16442);
or U18575 (N_18575,N_16765,N_17064);
nand U18576 (N_18576,N_16417,N_16275);
nand U18577 (N_18577,N_17551,N_17700);
xnor U18578 (N_18578,N_16519,N_16869);
nand U18579 (N_18579,N_17807,N_16972);
or U18580 (N_18580,N_17952,N_16219);
nor U18581 (N_18581,N_16412,N_16879);
or U18582 (N_18582,N_16771,N_16569);
and U18583 (N_18583,N_16724,N_17848);
xor U18584 (N_18584,N_17810,N_17923);
and U18585 (N_18585,N_16814,N_17027);
xnor U18586 (N_18586,N_17301,N_17636);
nor U18587 (N_18587,N_16392,N_16878);
and U18588 (N_18588,N_17832,N_17622);
xor U18589 (N_18589,N_17790,N_16135);
nand U18590 (N_18590,N_16329,N_16370);
xor U18591 (N_18591,N_16731,N_16349);
nor U18592 (N_18592,N_16779,N_16558);
xnor U18593 (N_18593,N_16716,N_17797);
and U18594 (N_18594,N_16941,N_16820);
nand U18595 (N_18595,N_16234,N_16045);
nor U18596 (N_18596,N_16836,N_16973);
and U18597 (N_18597,N_16604,N_16605);
nand U18598 (N_18598,N_16591,N_16629);
or U18599 (N_18599,N_16730,N_16872);
xnor U18600 (N_18600,N_17773,N_17499);
nor U18601 (N_18601,N_17042,N_16003);
nor U18602 (N_18602,N_17671,N_16084);
nor U18603 (N_18603,N_17396,N_17129);
nor U18604 (N_18604,N_17289,N_16637);
nor U18605 (N_18605,N_16168,N_17377);
or U18606 (N_18606,N_17865,N_16502);
nor U18607 (N_18607,N_17619,N_17266);
nor U18608 (N_18608,N_17372,N_17732);
nor U18609 (N_18609,N_17344,N_16819);
nor U18610 (N_18610,N_17885,N_17281);
or U18611 (N_18611,N_17028,N_17829);
or U18612 (N_18612,N_16438,N_17586);
nor U18613 (N_18613,N_17270,N_16667);
or U18614 (N_18614,N_16756,N_16031);
xor U18615 (N_18615,N_16687,N_17434);
nor U18616 (N_18616,N_16008,N_16261);
or U18617 (N_18617,N_16126,N_17888);
nor U18618 (N_18618,N_17308,N_16078);
nand U18619 (N_18619,N_17704,N_17857);
nand U18620 (N_18620,N_16283,N_17992);
or U18621 (N_18621,N_16171,N_16561);
nor U18622 (N_18622,N_17661,N_16523);
or U18623 (N_18623,N_17602,N_16876);
or U18624 (N_18624,N_17433,N_16807);
or U18625 (N_18625,N_16589,N_17548);
and U18626 (N_18626,N_17509,N_16866);
nand U18627 (N_18627,N_17474,N_17247);
or U18628 (N_18628,N_17229,N_17737);
nor U18629 (N_18629,N_17274,N_17820);
xnor U18630 (N_18630,N_16910,N_17771);
xnor U18631 (N_18631,N_16971,N_16257);
nand U18632 (N_18632,N_16658,N_17897);
and U18633 (N_18633,N_17571,N_17605);
and U18634 (N_18634,N_17268,N_16890);
nand U18635 (N_18635,N_16327,N_17745);
and U18636 (N_18636,N_16932,N_16808);
xnor U18637 (N_18637,N_16777,N_17279);
nor U18638 (N_18638,N_16818,N_17144);
or U18639 (N_18639,N_16440,N_17855);
and U18640 (N_18640,N_16835,N_16396);
xnor U18641 (N_18641,N_16366,N_17481);
or U18642 (N_18642,N_16860,N_17582);
and U18643 (N_18643,N_16368,N_17972);
xnor U18644 (N_18644,N_17758,N_17497);
or U18645 (N_18645,N_17259,N_17633);
nand U18646 (N_18646,N_17991,N_16533);
xor U18647 (N_18647,N_16468,N_17914);
or U18648 (N_18648,N_17273,N_17203);
xnor U18649 (N_18649,N_16276,N_16210);
nor U18650 (N_18650,N_17800,N_17983);
and U18651 (N_18651,N_17185,N_17447);
and U18652 (N_18652,N_16699,N_17354);
nand U18653 (N_18653,N_16893,N_16057);
or U18654 (N_18654,N_16311,N_16683);
nor U18655 (N_18655,N_16407,N_17085);
or U18656 (N_18656,N_17421,N_17003);
or U18657 (N_18657,N_16096,N_17904);
nand U18658 (N_18658,N_17093,N_17803);
nor U18659 (N_18659,N_16492,N_16490);
nor U18660 (N_18660,N_16361,N_17369);
nand U18661 (N_18661,N_16840,N_16269);
or U18662 (N_18662,N_17842,N_16642);
or U18663 (N_18663,N_17894,N_16173);
and U18664 (N_18664,N_17253,N_17872);
and U18665 (N_18665,N_17936,N_16709);
and U18666 (N_18666,N_16134,N_17840);
nor U18667 (N_18667,N_17135,N_16826);
or U18668 (N_18668,N_16160,N_16221);
or U18669 (N_18669,N_16775,N_17295);
nand U18670 (N_18670,N_17978,N_17658);
xor U18671 (N_18671,N_16700,N_17594);
nor U18672 (N_18672,N_16549,N_16713);
nand U18673 (N_18673,N_17265,N_17852);
or U18674 (N_18674,N_16445,N_16092);
nor U18675 (N_18675,N_16109,N_17150);
or U18676 (N_18676,N_16264,N_16592);
xor U18677 (N_18677,N_17005,N_16574);
nand U18678 (N_18678,N_16849,N_16354);
nor U18679 (N_18679,N_16360,N_16388);
xor U18680 (N_18680,N_17466,N_16572);
or U18681 (N_18681,N_17702,N_17436);
or U18682 (N_18682,N_16411,N_17232);
nor U18683 (N_18683,N_16732,N_16899);
nand U18684 (N_18684,N_16691,N_16288);
xnor U18685 (N_18685,N_17725,N_17349);
xor U18686 (N_18686,N_17422,N_17838);
and U18687 (N_18687,N_17798,N_17710);
xor U18688 (N_18688,N_16129,N_17726);
nor U18689 (N_18689,N_16652,N_16338);
and U18690 (N_18690,N_17928,N_17772);
nand U18691 (N_18691,N_16794,N_16977);
nor U18692 (N_18692,N_17156,N_17360);
nor U18693 (N_18693,N_16222,N_16831);
nor U18694 (N_18694,N_17590,N_17665);
xor U18695 (N_18695,N_16335,N_16180);
and U18696 (N_18696,N_16685,N_17507);
nor U18697 (N_18697,N_17925,N_16624);
or U18698 (N_18698,N_17067,N_17696);
or U18699 (N_18699,N_16404,N_16641);
or U18700 (N_18700,N_17001,N_17715);
and U18701 (N_18701,N_17151,N_17161);
nand U18702 (N_18702,N_16745,N_16043);
and U18703 (N_18703,N_17680,N_16827);
and U18704 (N_18704,N_16649,N_16456);
xor U18705 (N_18705,N_17750,N_16593);
or U18706 (N_18706,N_17488,N_17632);
and U18707 (N_18707,N_16676,N_16822);
nand U18708 (N_18708,N_17789,N_17412);
or U18709 (N_18709,N_16339,N_17008);
or U18710 (N_18710,N_16697,N_16859);
xnor U18711 (N_18711,N_16174,N_17890);
nand U18712 (N_18712,N_16790,N_17776);
or U18713 (N_18713,N_16123,N_16342);
or U18714 (N_18714,N_17924,N_17140);
nand U18715 (N_18715,N_16296,N_16858);
xor U18716 (N_18716,N_17262,N_17751);
xnor U18717 (N_18717,N_17854,N_17379);
or U18718 (N_18718,N_16796,N_17076);
or U18719 (N_18719,N_17881,N_17920);
nor U18720 (N_18720,N_16541,N_16531);
xnor U18721 (N_18721,N_17019,N_16821);
nand U18722 (N_18722,N_16302,N_16609);
nand U18723 (N_18723,N_17479,N_16906);
xor U18724 (N_18724,N_17740,N_17277);
xor U18725 (N_18725,N_16625,N_16387);
xor U18726 (N_18726,N_16179,N_16423);
nor U18727 (N_18727,N_17506,N_16233);
xnor U18728 (N_18728,N_17861,N_16673);
or U18729 (N_18729,N_17432,N_17334);
nand U18730 (N_18730,N_16117,N_17694);
nor U18731 (N_18731,N_16825,N_16829);
or U18732 (N_18732,N_16824,N_16864);
nand U18733 (N_18733,N_17864,N_17755);
nand U18734 (N_18734,N_16310,N_16672);
xnor U18735 (N_18735,N_17483,N_16711);
or U18736 (N_18736,N_16406,N_16671);
or U18737 (N_18737,N_17931,N_16984);
and U18738 (N_18738,N_17592,N_17194);
nor U18739 (N_18739,N_17998,N_17741);
nor U18740 (N_18740,N_16415,N_16414);
xor U18741 (N_18741,N_17190,N_16098);
nand U18742 (N_18742,N_16698,N_16032);
nand U18743 (N_18743,N_17121,N_17058);
nand U18744 (N_18744,N_17160,N_17650);
xor U18745 (N_18745,N_17553,N_16346);
xor U18746 (N_18746,N_16715,N_17728);
or U18747 (N_18747,N_16439,N_16089);
nand U18748 (N_18748,N_17395,N_17717);
or U18749 (N_18749,N_16870,N_17879);
or U18750 (N_18750,N_17663,N_16122);
xor U18751 (N_18751,N_16216,N_16877);
xnor U18752 (N_18752,N_16557,N_16223);
nor U18753 (N_18753,N_17380,N_16703);
nor U18754 (N_18754,N_16111,N_17615);
or U18755 (N_18755,N_16295,N_17287);
or U18756 (N_18756,N_17979,N_16037);
and U18757 (N_18757,N_17511,N_17221);
xnor U18758 (N_18758,N_16500,N_17325);
xnor U18759 (N_18759,N_17986,N_16892);
nand U18760 (N_18760,N_17819,N_16559);
or U18761 (N_18761,N_17007,N_16583);
nor U18762 (N_18762,N_17996,N_17545);
or U18763 (N_18763,N_17490,N_17133);
nand U18764 (N_18764,N_17673,N_17225);
nor U18765 (N_18765,N_16498,N_17735);
xnor U18766 (N_18766,N_17686,N_17706);
xnor U18767 (N_18767,N_17837,N_17766);
xnor U18768 (N_18768,N_16181,N_17104);
and U18769 (N_18769,N_16587,N_17330);
nand U18770 (N_18770,N_16225,N_17580);
xor U18771 (N_18771,N_17401,N_17283);
xor U18772 (N_18772,N_16828,N_17692);
or U18773 (N_18773,N_17593,N_16842);
xor U18774 (N_18774,N_16459,N_16690);
or U18775 (N_18775,N_16646,N_17635);
nand U18776 (N_18776,N_16345,N_17163);
nand U18777 (N_18777,N_16736,N_16817);
nor U18778 (N_18778,N_16544,N_17188);
and U18779 (N_18779,N_17869,N_17946);
nor U18780 (N_18780,N_17948,N_17366);
and U18781 (N_18781,N_17664,N_16653);
nand U18782 (N_18782,N_16874,N_16496);
or U18783 (N_18783,N_17679,N_17833);
nand U18784 (N_18784,N_17195,N_16844);
nor U18785 (N_18785,N_16614,N_16995);
xor U18786 (N_18786,N_16047,N_17641);
and U18787 (N_18787,N_17961,N_16546);
or U18788 (N_18788,N_16912,N_16376);
xor U18789 (N_18789,N_16883,N_16379);
or U18790 (N_18790,N_17701,N_16182);
or U18791 (N_18791,N_17721,N_17851);
and U18792 (N_18792,N_16585,N_16140);
or U18793 (N_18793,N_17546,N_16231);
nand U18794 (N_18794,N_16478,N_16978);
or U18795 (N_18795,N_16501,N_17082);
or U18796 (N_18796,N_17054,N_16540);
nor U18797 (N_18797,N_17749,N_16434);
and U18798 (N_18798,N_16784,N_17943);
or U18799 (N_18799,N_17493,N_16701);
nand U18800 (N_18800,N_17828,N_16200);
or U18801 (N_18801,N_17645,N_17678);
nor U18802 (N_18802,N_17217,N_16809);
or U18803 (N_18803,N_17805,N_16274);
and U18804 (N_18804,N_16661,N_17501);
xor U18805 (N_18805,N_16772,N_16431);
and U18806 (N_18806,N_17105,N_17022);
and U18807 (N_18807,N_16950,N_17111);
nand U18808 (N_18808,N_17040,N_17316);
nand U18809 (N_18809,N_17906,N_16118);
xor U18810 (N_18810,N_17585,N_16755);
xor U18811 (N_18811,N_16267,N_16846);
nor U18812 (N_18812,N_17779,N_16324);
or U18813 (N_18813,N_16513,N_17707);
nand U18814 (N_18814,N_17047,N_16088);
nand U18815 (N_18815,N_17126,N_16262);
and U18816 (N_18816,N_17115,N_16207);
or U18817 (N_18817,N_17009,N_17374);
or U18818 (N_18818,N_16895,N_17521);
and U18819 (N_18819,N_16943,N_17491);
or U18820 (N_18820,N_16503,N_16720);
or U18821 (N_18821,N_17452,N_16873);
or U18822 (N_18822,N_17246,N_17415);
xnor U18823 (N_18823,N_16969,N_17712);
and U18824 (N_18824,N_17314,N_17649);
or U18825 (N_18825,N_17324,N_16812);
nor U18826 (N_18826,N_17032,N_16051);
nor U18827 (N_18827,N_16332,N_17155);
or U18828 (N_18828,N_16352,N_16618);
xor U18829 (N_18829,N_16190,N_17769);
xnor U18830 (N_18830,N_16915,N_17775);
nor U18831 (N_18831,N_17523,N_17035);
and U18832 (N_18832,N_16243,N_16384);
xnor U18833 (N_18833,N_16773,N_16487);
and U18834 (N_18834,N_16575,N_17846);
nand U18835 (N_18835,N_17533,N_16979);
nand U18836 (N_18836,N_16287,N_16485);
xor U18837 (N_18837,N_17044,N_17411);
nand U18838 (N_18838,N_17029,N_17143);
nor U18839 (N_18839,N_16710,N_17280);
nand U18840 (N_18840,N_16719,N_17963);
and U18841 (N_18841,N_16968,N_17159);
or U18842 (N_18842,N_16251,N_16670);
nor U18843 (N_18843,N_17231,N_16505);
and U18844 (N_18844,N_17757,N_16853);
and U18845 (N_18845,N_16070,N_16988);
and U18846 (N_18846,N_17893,N_17913);
nor U18847 (N_18847,N_17459,N_17699);
xor U18848 (N_18848,N_17018,N_16966);
or U18849 (N_18849,N_17102,N_16020);
and U18850 (N_18850,N_17100,N_16170);
nand U18851 (N_18851,N_16065,N_16069);
nor U18852 (N_18852,N_17045,N_16422);
nor U18853 (N_18853,N_17626,N_16799);
and U18854 (N_18854,N_16550,N_17445);
or U18855 (N_18855,N_17518,N_16208);
nor U18856 (N_18856,N_17561,N_16453);
nand U18857 (N_18857,N_17919,N_16420);
and U18858 (N_18858,N_16454,N_16651);
nor U18859 (N_18859,N_17181,N_16060);
nor U18860 (N_18860,N_17204,N_17542);
nand U18861 (N_18861,N_17620,N_17556);
nand U18862 (N_18862,N_16383,N_16769);
and U18863 (N_18863,N_16723,N_16803);
xnor U18864 (N_18864,N_16861,N_17382);
nand U18865 (N_18865,N_17988,N_17905);
xnor U18866 (N_18866,N_17034,N_17565);
nand U18867 (N_18867,N_17761,N_17618);
nand U18868 (N_18868,N_16838,N_16588);
and U18869 (N_18869,N_17012,N_17154);
and U18870 (N_18870,N_17866,N_17198);
xor U18871 (N_18871,N_16323,N_16068);
nand U18872 (N_18872,N_16922,N_16774);
or U18873 (N_18873,N_17990,N_16449);
or U18874 (N_18874,N_16297,N_17579);
nor U18875 (N_18875,N_16426,N_17356);
and U18876 (N_18876,N_16695,N_16521);
and U18877 (N_18877,N_17168,N_17868);
or U18878 (N_18878,N_17083,N_17989);
xor U18879 (N_18879,N_17258,N_17278);
or U18880 (N_18880,N_16120,N_17791);
or U18881 (N_18881,N_16054,N_17055);
nor U18882 (N_18882,N_16499,N_17843);
and U18883 (N_18883,N_17014,N_16905);
nand U18884 (N_18884,N_16432,N_17417);
nand U18885 (N_18885,N_16235,N_16213);
nor U18886 (N_18886,N_16007,N_17118);
nand U18887 (N_18887,N_17756,N_16177);
nor U18888 (N_18888,N_16410,N_17023);
or U18889 (N_18889,N_17389,N_16290);
xnor U18890 (N_18890,N_16224,N_16403);
xnor U18891 (N_18891,N_17494,N_17964);
or U18892 (N_18892,N_16679,N_16535);
xor U18893 (N_18893,N_17077,N_17108);
xor U18894 (N_18894,N_16152,N_16055);
nand U18895 (N_18895,N_16425,N_16086);
xor U18896 (N_18896,N_16867,N_16002);
nand U18897 (N_18897,N_17891,N_16567);
or U18898 (N_18898,N_16108,N_16627);
and U18899 (N_18899,N_17043,N_17139);
nand U18900 (N_18900,N_17596,N_16525);
nor U18901 (N_18901,N_17134,N_17486);
xnor U18902 (N_18902,N_17878,N_16693);
nor U18903 (N_18903,N_16782,N_16741);
xor U18904 (N_18904,N_16015,N_16577);
xor U18905 (N_18905,N_17137,N_17845);
nand U18906 (N_18906,N_16992,N_16185);
or U18907 (N_18907,N_16038,N_16571);
or U18908 (N_18908,N_17598,N_16141);
or U18909 (N_18909,N_17508,N_17457);
nor U18910 (N_18910,N_17941,N_16090);
xnor U18911 (N_18911,N_16374,N_16491);
or U18912 (N_18912,N_16481,N_17844);
xor U18913 (N_18913,N_16340,N_17589);
nor U18914 (N_18914,N_16925,N_16537);
nor U18915 (N_18915,N_16747,N_17322);
xnor U18916 (N_18916,N_16325,N_17427);
xnor U18917 (N_18917,N_17056,N_16077);
or U18918 (N_18918,N_16622,N_16273);
and U18919 (N_18919,N_16957,N_16289);
xnor U18920 (N_18920,N_17223,N_17026);
xnor U18921 (N_18921,N_16254,N_17916);
xor U18922 (N_18922,N_17091,N_17090);
xnor U18923 (N_18923,N_16936,N_16399);
nand U18924 (N_18924,N_16778,N_16580);
nor U18925 (N_18925,N_16787,N_16717);
nand U18926 (N_18926,N_16983,N_17392);
xor U18927 (N_18927,N_16457,N_17060);
nor U18928 (N_18928,N_16005,N_16433);
xnor U18929 (N_18929,N_17051,N_17886);
or U18930 (N_18930,N_17309,N_17286);
xor U18931 (N_18931,N_16985,N_17748);
nor U18932 (N_18932,N_16882,N_17733);
xor U18933 (N_18933,N_16862,N_17816);
nand U18934 (N_18934,N_16058,N_17468);
nor U18935 (N_18935,N_16744,N_16536);
and U18936 (N_18936,N_16004,N_17522);
or U18937 (N_18937,N_17170,N_17939);
nand U18938 (N_18938,N_16990,N_17938);
nand U18939 (N_18939,N_16027,N_17743);
nor U18940 (N_18940,N_17759,N_16644);
or U18941 (N_18941,N_17127,N_17039);
nor U18942 (N_18942,N_16286,N_16657);
xnor U18943 (N_18943,N_17464,N_17781);
nand U18944 (N_18944,N_17250,N_16085);
and U18945 (N_18945,N_16458,N_17070);
and U18946 (N_18946,N_16306,N_16304);
or U18947 (N_18947,N_17564,N_16074);
nor U18948 (N_18948,N_16187,N_16884);
nor U18949 (N_18949,N_16889,N_16193);
nand U18950 (N_18950,N_16675,N_16998);
xnor U18951 (N_18951,N_16046,N_16199);
nand U18952 (N_18952,N_16515,N_16044);
xnor U18953 (N_18953,N_17883,N_17327);
or U18954 (N_18954,N_16469,N_16582);
nand U18955 (N_18955,N_17099,N_16398);
nor U18956 (N_18956,N_17669,N_16823);
nand U18957 (N_18957,N_16639,N_17627);
or U18958 (N_18958,N_17164,N_17335);
or U18959 (N_18959,N_16986,N_17909);
nand U18960 (N_18960,N_16909,N_17817);
nand U18961 (N_18961,N_17297,N_17600);
and U18962 (N_18962,N_17954,N_16165);
nand U18963 (N_18963,N_16590,N_17455);
nand U18964 (N_18964,N_16083,N_17069);
nor U18965 (N_18965,N_17482,N_16441);
and U18966 (N_18966,N_17785,N_17011);
nand U18967 (N_18967,N_16250,N_16493);
and U18968 (N_18968,N_17903,N_17691);
xor U18969 (N_18969,N_16330,N_16115);
or U18970 (N_18970,N_16632,N_17172);
nand U18971 (N_18971,N_16551,N_17178);
or U18972 (N_18972,N_16954,N_17146);
nor U18973 (N_18973,N_17918,N_16471);
or U18974 (N_18974,N_16094,N_17657);
and U18975 (N_18975,N_16621,N_17340);
or U18976 (N_18976,N_16217,N_17423);
nor U18977 (N_18977,N_17685,N_16258);
nand U18978 (N_18978,N_16946,N_17063);
nor U18979 (N_18979,N_16631,N_16482);
nand U18980 (N_18980,N_17827,N_17498);
or U18981 (N_18981,N_16400,N_16277);
nand U18982 (N_18982,N_16116,N_17252);
and U18983 (N_18983,N_16729,N_17550);
nand U18984 (N_18984,N_16341,N_17373);
xnor U18985 (N_18985,N_16678,N_16390);
xor U18986 (N_18986,N_17660,N_17705);
nor U18987 (N_18987,N_17239,N_17540);
or U18988 (N_18988,N_17136,N_16428);
or U18989 (N_18989,N_17683,N_17538);
xnor U18990 (N_18990,N_16268,N_16378);
xnor U18991 (N_18991,N_17484,N_16385);
and U18992 (N_18992,N_17825,N_17346);
nor U18993 (N_18993,N_17074,N_17202);
or U18994 (N_18994,N_17656,N_17765);
xor U18995 (N_18995,N_17031,N_16726);
or U18996 (N_18996,N_16198,N_16798);
or U18997 (N_18997,N_16461,N_17847);
nor U18998 (N_18998,N_16802,N_17103);
nand U18999 (N_18999,N_16543,N_16214);
or U19000 (N_19000,N_17526,N_17319);
and U19001 (N_19001,N_16637,N_17903);
nor U19002 (N_19002,N_17439,N_16033);
xor U19003 (N_19003,N_17919,N_17128);
nand U19004 (N_19004,N_17240,N_17137);
nor U19005 (N_19005,N_16009,N_16483);
and U19006 (N_19006,N_17526,N_16116);
nor U19007 (N_19007,N_17243,N_17857);
or U19008 (N_19008,N_17514,N_16130);
or U19009 (N_19009,N_16701,N_17707);
and U19010 (N_19010,N_17236,N_17645);
xor U19011 (N_19011,N_16404,N_17280);
nand U19012 (N_19012,N_16242,N_17370);
nor U19013 (N_19013,N_17452,N_16267);
nor U19014 (N_19014,N_16335,N_17828);
nor U19015 (N_19015,N_16227,N_17628);
nor U19016 (N_19016,N_17430,N_16261);
nand U19017 (N_19017,N_17933,N_17980);
or U19018 (N_19018,N_17861,N_16858);
nand U19019 (N_19019,N_16442,N_17213);
and U19020 (N_19020,N_17889,N_16054);
nor U19021 (N_19021,N_17897,N_16309);
and U19022 (N_19022,N_16468,N_16366);
xor U19023 (N_19023,N_17152,N_16978);
and U19024 (N_19024,N_17389,N_16148);
nor U19025 (N_19025,N_16952,N_17940);
nand U19026 (N_19026,N_16497,N_16237);
nand U19027 (N_19027,N_17353,N_16195);
and U19028 (N_19028,N_16830,N_16898);
nand U19029 (N_19029,N_17515,N_17576);
xnor U19030 (N_19030,N_17677,N_17343);
nor U19031 (N_19031,N_16421,N_16870);
or U19032 (N_19032,N_16311,N_17717);
nor U19033 (N_19033,N_17558,N_16035);
or U19034 (N_19034,N_16119,N_17060);
xnor U19035 (N_19035,N_17027,N_17530);
nor U19036 (N_19036,N_17643,N_16051);
or U19037 (N_19037,N_16688,N_17914);
nand U19038 (N_19038,N_16025,N_17187);
nand U19039 (N_19039,N_16843,N_16704);
xnor U19040 (N_19040,N_17653,N_16325);
xnor U19041 (N_19041,N_17504,N_16863);
nor U19042 (N_19042,N_16473,N_17033);
nand U19043 (N_19043,N_17287,N_17093);
and U19044 (N_19044,N_17769,N_16148);
xor U19045 (N_19045,N_17081,N_16685);
nor U19046 (N_19046,N_16044,N_16612);
or U19047 (N_19047,N_17907,N_17994);
nand U19048 (N_19048,N_17056,N_17562);
and U19049 (N_19049,N_17753,N_16918);
or U19050 (N_19050,N_17909,N_16178);
xor U19051 (N_19051,N_17489,N_17252);
and U19052 (N_19052,N_17243,N_16262);
or U19053 (N_19053,N_16618,N_16644);
or U19054 (N_19054,N_17651,N_17134);
nor U19055 (N_19055,N_17732,N_17569);
xnor U19056 (N_19056,N_16244,N_16897);
nand U19057 (N_19057,N_17495,N_16432);
xnor U19058 (N_19058,N_16342,N_17694);
and U19059 (N_19059,N_16759,N_17803);
and U19060 (N_19060,N_17118,N_17849);
nor U19061 (N_19061,N_16697,N_17138);
or U19062 (N_19062,N_17232,N_16659);
xor U19063 (N_19063,N_16743,N_17749);
xnor U19064 (N_19064,N_17637,N_17780);
xor U19065 (N_19065,N_17640,N_17469);
or U19066 (N_19066,N_17304,N_17425);
nand U19067 (N_19067,N_17363,N_16766);
xor U19068 (N_19068,N_17033,N_16959);
and U19069 (N_19069,N_17725,N_16265);
nand U19070 (N_19070,N_17913,N_17709);
nand U19071 (N_19071,N_16825,N_16046);
nand U19072 (N_19072,N_17321,N_16363);
and U19073 (N_19073,N_17874,N_16342);
nand U19074 (N_19074,N_16122,N_17560);
or U19075 (N_19075,N_16168,N_17160);
nand U19076 (N_19076,N_17053,N_17529);
nor U19077 (N_19077,N_17365,N_17092);
and U19078 (N_19078,N_17122,N_16518);
or U19079 (N_19079,N_16943,N_16287);
xnor U19080 (N_19080,N_16497,N_16174);
and U19081 (N_19081,N_17078,N_17353);
nand U19082 (N_19082,N_16021,N_16826);
nand U19083 (N_19083,N_16226,N_16448);
xor U19084 (N_19084,N_17228,N_16500);
xnor U19085 (N_19085,N_17815,N_16977);
and U19086 (N_19086,N_17751,N_16677);
nor U19087 (N_19087,N_16746,N_17852);
or U19088 (N_19088,N_17291,N_17513);
nor U19089 (N_19089,N_17734,N_17331);
or U19090 (N_19090,N_17829,N_16836);
nor U19091 (N_19091,N_17506,N_17815);
and U19092 (N_19092,N_17871,N_17565);
and U19093 (N_19093,N_17722,N_16041);
xnor U19094 (N_19094,N_17681,N_17981);
xnor U19095 (N_19095,N_17279,N_17484);
nand U19096 (N_19096,N_16943,N_16096);
and U19097 (N_19097,N_16413,N_16937);
nor U19098 (N_19098,N_17860,N_17870);
and U19099 (N_19099,N_17890,N_17126);
xor U19100 (N_19100,N_16608,N_17412);
xor U19101 (N_19101,N_16309,N_17917);
xnor U19102 (N_19102,N_17277,N_16775);
or U19103 (N_19103,N_16249,N_16667);
nand U19104 (N_19104,N_17126,N_16271);
nand U19105 (N_19105,N_17267,N_16303);
nor U19106 (N_19106,N_17256,N_17847);
nand U19107 (N_19107,N_16133,N_17803);
or U19108 (N_19108,N_17881,N_16998);
and U19109 (N_19109,N_16847,N_16353);
nand U19110 (N_19110,N_16452,N_17473);
nand U19111 (N_19111,N_16644,N_16452);
xnor U19112 (N_19112,N_17120,N_17983);
or U19113 (N_19113,N_16510,N_17244);
xnor U19114 (N_19114,N_17467,N_16337);
and U19115 (N_19115,N_17802,N_16367);
and U19116 (N_19116,N_16023,N_17502);
nand U19117 (N_19117,N_16140,N_16501);
nor U19118 (N_19118,N_17896,N_16311);
and U19119 (N_19119,N_17100,N_16701);
and U19120 (N_19120,N_17837,N_17221);
and U19121 (N_19121,N_16006,N_16109);
and U19122 (N_19122,N_16969,N_17666);
or U19123 (N_19123,N_17726,N_17735);
nor U19124 (N_19124,N_16919,N_17715);
nor U19125 (N_19125,N_17835,N_17940);
xor U19126 (N_19126,N_16755,N_16917);
xnor U19127 (N_19127,N_16216,N_17695);
xnor U19128 (N_19128,N_16173,N_17082);
and U19129 (N_19129,N_17342,N_17073);
xor U19130 (N_19130,N_16851,N_16065);
nor U19131 (N_19131,N_17151,N_16556);
nand U19132 (N_19132,N_17623,N_16592);
nor U19133 (N_19133,N_16855,N_16816);
or U19134 (N_19134,N_17494,N_17048);
xnor U19135 (N_19135,N_17680,N_16004);
nand U19136 (N_19136,N_16758,N_16266);
xnor U19137 (N_19137,N_17683,N_16951);
xor U19138 (N_19138,N_17681,N_16447);
or U19139 (N_19139,N_17529,N_16480);
nor U19140 (N_19140,N_17835,N_17246);
nand U19141 (N_19141,N_16116,N_17113);
or U19142 (N_19142,N_17368,N_17932);
nor U19143 (N_19143,N_17277,N_16972);
and U19144 (N_19144,N_16748,N_17731);
and U19145 (N_19145,N_17209,N_16609);
xnor U19146 (N_19146,N_16218,N_16504);
nor U19147 (N_19147,N_16282,N_17463);
nand U19148 (N_19148,N_16036,N_17180);
xnor U19149 (N_19149,N_16918,N_17068);
and U19150 (N_19150,N_16866,N_16085);
nor U19151 (N_19151,N_16972,N_16796);
and U19152 (N_19152,N_16013,N_17412);
xor U19153 (N_19153,N_17771,N_17493);
nand U19154 (N_19154,N_16936,N_16773);
xnor U19155 (N_19155,N_17155,N_16696);
or U19156 (N_19156,N_16045,N_17779);
nor U19157 (N_19157,N_16587,N_16298);
or U19158 (N_19158,N_17352,N_16125);
xor U19159 (N_19159,N_16061,N_16074);
xor U19160 (N_19160,N_17224,N_16826);
and U19161 (N_19161,N_16131,N_17428);
and U19162 (N_19162,N_17925,N_16262);
xor U19163 (N_19163,N_17854,N_17972);
nor U19164 (N_19164,N_16398,N_16859);
or U19165 (N_19165,N_16966,N_16313);
or U19166 (N_19166,N_16723,N_17537);
nand U19167 (N_19167,N_17476,N_16061);
nand U19168 (N_19168,N_17943,N_16214);
xnor U19169 (N_19169,N_17410,N_17099);
nor U19170 (N_19170,N_16377,N_16133);
xnor U19171 (N_19171,N_17835,N_16619);
or U19172 (N_19172,N_17028,N_16102);
nor U19173 (N_19173,N_17786,N_16357);
xor U19174 (N_19174,N_17302,N_16034);
and U19175 (N_19175,N_17268,N_16690);
and U19176 (N_19176,N_16224,N_17231);
nand U19177 (N_19177,N_16625,N_17746);
and U19178 (N_19178,N_17842,N_16711);
or U19179 (N_19179,N_17966,N_17271);
nand U19180 (N_19180,N_16985,N_17137);
xnor U19181 (N_19181,N_17971,N_16881);
nand U19182 (N_19182,N_17935,N_16469);
nand U19183 (N_19183,N_16848,N_17698);
xnor U19184 (N_19184,N_16740,N_16596);
nand U19185 (N_19185,N_16672,N_16424);
or U19186 (N_19186,N_16176,N_17639);
or U19187 (N_19187,N_16975,N_16874);
nand U19188 (N_19188,N_17143,N_17223);
and U19189 (N_19189,N_16505,N_17916);
nand U19190 (N_19190,N_17646,N_17449);
nand U19191 (N_19191,N_17589,N_16241);
xnor U19192 (N_19192,N_17171,N_16431);
and U19193 (N_19193,N_16873,N_17909);
nor U19194 (N_19194,N_17770,N_17879);
nor U19195 (N_19195,N_16223,N_16231);
and U19196 (N_19196,N_16803,N_17306);
and U19197 (N_19197,N_16718,N_17721);
and U19198 (N_19198,N_16417,N_16835);
nand U19199 (N_19199,N_17422,N_16306);
xnor U19200 (N_19200,N_17294,N_16705);
and U19201 (N_19201,N_16095,N_16382);
and U19202 (N_19202,N_17479,N_16665);
nand U19203 (N_19203,N_16199,N_17664);
or U19204 (N_19204,N_17939,N_17131);
and U19205 (N_19205,N_17902,N_16493);
and U19206 (N_19206,N_16891,N_17464);
xor U19207 (N_19207,N_16381,N_17038);
or U19208 (N_19208,N_17275,N_16594);
nand U19209 (N_19209,N_17289,N_16759);
nand U19210 (N_19210,N_16899,N_17254);
xor U19211 (N_19211,N_16492,N_17721);
xor U19212 (N_19212,N_16640,N_17432);
and U19213 (N_19213,N_17089,N_16574);
or U19214 (N_19214,N_16402,N_16493);
nand U19215 (N_19215,N_16853,N_17632);
nand U19216 (N_19216,N_17766,N_16177);
or U19217 (N_19217,N_16312,N_17212);
nor U19218 (N_19218,N_16594,N_16649);
xor U19219 (N_19219,N_16742,N_17453);
xnor U19220 (N_19220,N_17989,N_16385);
and U19221 (N_19221,N_16512,N_16656);
xnor U19222 (N_19222,N_17028,N_17092);
and U19223 (N_19223,N_16753,N_16549);
or U19224 (N_19224,N_17910,N_17408);
or U19225 (N_19225,N_17164,N_17605);
and U19226 (N_19226,N_17148,N_16398);
and U19227 (N_19227,N_17472,N_16065);
or U19228 (N_19228,N_17930,N_17500);
xnor U19229 (N_19229,N_17645,N_16399);
xnor U19230 (N_19230,N_16286,N_17238);
nor U19231 (N_19231,N_17877,N_16532);
or U19232 (N_19232,N_16962,N_17558);
nor U19233 (N_19233,N_16334,N_16555);
nand U19234 (N_19234,N_17045,N_17351);
nor U19235 (N_19235,N_17087,N_17148);
nand U19236 (N_19236,N_16456,N_17420);
nand U19237 (N_19237,N_16176,N_17788);
or U19238 (N_19238,N_17972,N_17621);
nor U19239 (N_19239,N_16359,N_16328);
nor U19240 (N_19240,N_17054,N_16388);
nand U19241 (N_19241,N_17013,N_16514);
nand U19242 (N_19242,N_16926,N_16451);
or U19243 (N_19243,N_16541,N_16733);
nand U19244 (N_19244,N_16486,N_17289);
xor U19245 (N_19245,N_16500,N_17391);
nand U19246 (N_19246,N_17742,N_16739);
nand U19247 (N_19247,N_16015,N_17214);
nor U19248 (N_19248,N_17257,N_17504);
xor U19249 (N_19249,N_16751,N_16476);
and U19250 (N_19250,N_16279,N_16545);
and U19251 (N_19251,N_16447,N_17432);
xnor U19252 (N_19252,N_17832,N_17101);
nor U19253 (N_19253,N_16663,N_17859);
nand U19254 (N_19254,N_17300,N_17098);
nor U19255 (N_19255,N_16106,N_17495);
nand U19256 (N_19256,N_16003,N_16238);
xnor U19257 (N_19257,N_16754,N_17530);
and U19258 (N_19258,N_16385,N_16230);
xor U19259 (N_19259,N_16146,N_17210);
nand U19260 (N_19260,N_16106,N_16895);
or U19261 (N_19261,N_17418,N_17625);
nand U19262 (N_19262,N_17681,N_17381);
xnor U19263 (N_19263,N_16202,N_17459);
nor U19264 (N_19264,N_17762,N_17332);
and U19265 (N_19265,N_16057,N_16770);
or U19266 (N_19266,N_17961,N_17298);
or U19267 (N_19267,N_17944,N_17020);
and U19268 (N_19268,N_16582,N_17141);
and U19269 (N_19269,N_17926,N_17318);
nand U19270 (N_19270,N_16735,N_17393);
xnor U19271 (N_19271,N_17543,N_17043);
xnor U19272 (N_19272,N_17186,N_16200);
nor U19273 (N_19273,N_17868,N_17055);
nand U19274 (N_19274,N_17441,N_17954);
xnor U19275 (N_19275,N_17794,N_17490);
xnor U19276 (N_19276,N_16681,N_16648);
nor U19277 (N_19277,N_17560,N_16178);
xor U19278 (N_19278,N_16264,N_17018);
and U19279 (N_19279,N_16131,N_17654);
nand U19280 (N_19280,N_16995,N_16798);
and U19281 (N_19281,N_17992,N_16308);
nor U19282 (N_19282,N_17092,N_16631);
nor U19283 (N_19283,N_17233,N_17987);
nor U19284 (N_19284,N_16092,N_16310);
nand U19285 (N_19285,N_17676,N_16723);
nor U19286 (N_19286,N_16042,N_16318);
xor U19287 (N_19287,N_16596,N_16277);
and U19288 (N_19288,N_17704,N_17131);
nor U19289 (N_19289,N_16356,N_16450);
nor U19290 (N_19290,N_16005,N_17223);
xor U19291 (N_19291,N_17358,N_16946);
nor U19292 (N_19292,N_17408,N_16423);
xor U19293 (N_19293,N_16796,N_17182);
nand U19294 (N_19294,N_17892,N_16894);
nor U19295 (N_19295,N_17004,N_17389);
and U19296 (N_19296,N_17088,N_17587);
nor U19297 (N_19297,N_16558,N_16746);
nand U19298 (N_19298,N_17911,N_17168);
and U19299 (N_19299,N_17930,N_16152);
or U19300 (N_19300,N_16328,N_16868);
and U19301 (N_19301,N_17243,N_17615);
nor U19302 (N_19302,N_16314,N_17751);
or U19303 (N_19303,N_17661,N_16886);
or U19304 (N_19304,N_17081,N_16785);
nand U19305 (N_19305,N_16720,N_17109);
xor U19306 (N_19306,N_17735,N_16509);
xor U19307 (N_19307,N_16390,N_16302);
and U19308 (N_19308,N_17741,N_16447);
nor U19309 (N_19309,N_17220,N_16514);
nand U19310 (N_19310,N_16175,N_16970);
and U19311 (N_19311,N_16078,N_17896);
xor U19312 (N_19312,N_17140,N_16478);
and U19313 (N_19313,N_17201,N_16123);
nand U19314 (N_19314,N_16499,N_16708);
nor U19315 (N_19315,N_16997,N_16651);
nor U19316 (N_19316,N_16729,N_17189);
or U19317 (N_19317,N_17284,N_17403);
nand U19318 (N_19318,N_16788,N_17418);
and U19319 (N_19319,N_16807,N_16449);
or U19320 (N_19320,N_16341,N_16661);
or U19321 (N_19321,N_16540,N_17619);
nor U19322 (N_19322,N_17989,N_16108);
nor U19323 (N_19323,N_17684,N_16494);
nor U19324 (N_19324,N_16758,N_16062);
nor U19325 (N_19325,N_16339,N_16624);
and U19326 (N_19326,N_16268,N_17328);
nand U19327 (N_19327,N_16767,N_17989);
or U19328 (N_19328,N_17969,N_17426);
nor U19329 (N_19329,N_16532,N_16864);
nor U19330 (N_19330,N_17375,N_16098);
xor U19331 (N_19331,N_17437,N_17008);
xor U19332 (N_19332,N_16965,N_16812);
xnor U19333 (N_19333,N_16464,N_16331);
or U19334 (N_19334,N_17648,N_16122);
xor U19335 (N_19335,N_16443,N_16414);
or U19336 (N_19336,N_16629,N_17318);
xnor U19337 (N_19337,N_17854,N_17047);
xor U19338 (N_19338,N_17276,N_16068);
or U19339 (N_19339,N_17536,N_16619);
nand U19340 (N_19340,N_17770,N_16148);
xor U19341 (N_19341,N_17998,N_16836);
xor U19342 (N_19342,N_16855,N_16250);
or U19343 (N_19343,N_16328,N_16143);
xor U19344 (N_19344,N_17303,N_17264);
nor U19345 (N_19345,N_16415,N_16145);
and U19346 (N_19346,N_17720,N_17647);
or U19347 (N_19347,N_17722,N_17427);
or U19348 (N_19348,N_17864,N_17909);
nand U19349 (N_19349,N_17798,N_17963);
xnor U19350 (N_19350,N_16509,N_17989);
nand U19351 (N_19351,N_16430,N_17878);
nor U19352 (N_19352,N_16160,N_16074);
xor U19353 (N_19353,N_16928,N_17615);
and U19354 (N_19354,N_16313,N_16425);
and U19355 (N_19355,N_17730,N_17601);
and U19356 (N_19356,N_16381,N_16240);
and U19357 (N_19357,N_16506,N_17050);
and U19358 (N_19358,N_16344,N_16082);
xnor U19359 (N_19359,N_17562,N_16139);
and U19360 (N_19360,N_16798,N_17004);
xor U19361 (N_19361,N_16198,N_16060);
nand U19362 (N_19362,N_16196,N_16497);
and U19363 (N_19363,N_17377,N_16803);
nand U19364 (N_19364,N_16543,N_16791);
xor U19365 (N_19365,N_16582,N_16437);
nand U19366 (N_19366,N_16028,N_16665);
nand U19367 (N_19367,N_17934,N_17511);
nor U19368 (N_19368,N_16246,N_16118);
and U19369 (N_19369,N_17305,N_17193);
nor U19370 (N_19370,N_17809,N_16936);
nand U19371 (N_19371,N_17666,N_17276);
nor U19372 (N_19372,N_17278,N_17123);
xnor U19373 (N_19373,N_16099,N_16664);
nand U19374 (N_19374,N_17128,N_16749);
and U19375 (N_19375,N_17075,N_17889);
or U19376 (N_19376,N_16182,N_16988);
nor U19377 (N_19377,N_17666,N_16983);
xnor U19378 (N_19378,N_16059,N_16307);
nand U19379 (N_19379,N_16519,N_17569);
nor U19380 (N_19380,N_16483,N_16335);
xor U19381 (N_19381,N_17378,N_17422);
or U19382 (N_19382,N_17552,N_16521);
xor U19383 (N_19383,N_17065,N_16093);
or U19384 (N_19384,N_16280,N_17749);
nand U19385 (N_19385,N_17838,N_16976);
nor U19386 (N_19386,N_16370,N_17023);
and U19387 (N_19387,N_16753,N_17765);
nand U19388 (N_19388,N_17309,N_17072);
xor U19389 (N_19389,N_17860,N_17723);
nand U19390 (N_19390,N_16659,N_17122);
and U19391 (N_19391,N_16909,N_17856);
xor U19392 (N_19392,N_17294,N_16537);
or U19393 (N_19393,N_17722,N_17521);
nor U19394 (N_19394,N_16076,N_16988);
and U19395 (N_19395,N_17498,N_17491);
nand U19396 (N_19396,N_16470,N_17673);
nand U19397 (N_19397,N_17469,N_16463);
xnor U19398 (N_19398,N_17356,N_17586);
nand U19399 (N_19399,N_16376,N_17893);
nor U19400 (N_19400,N_16650,N_16484);
or U19401 (N_19401,N_16205,N_17023);
nand U19402 (N_19402,N_17325,N_17909);
nor U19403 (N_19403,N_17432,N_16618);
nand U19404 (N_19404,N_17762,N_17439);
nor U19405 (N_19405,N_16884,N_17562);
nand U19406 (N_19406,N_16243,N_16005);
nor U19407 (N_19407,N_16293,N_17600);
nand U19408 (N_19408,N_17235,N_17841);
or U19409 (N_19409,N_17970,N_16442);
and U19410 (N_19410,N_17541,N_17337);
nand U19411 (N_19411,N_16307,N_17473);
nand U19412 (N_19412,N_17256,N_17356);
nand U19413 (N_19413,N_16391,N_16064);
nand U19414 (N_19414,N_16755,N_16856);
and U19415 (N_19415,N_17505,N_17846);
nand U19416 (N_19416,N_16048,N_17992);
or U19417 (N_19417,N_16724,N_17398);
and U19418 (N_19418,N_16668,N_17523);
xor U19419 (N_19419,N_16888,N_16249);
xor U19420 (N_19420,N_17202,N_17967);
nand U19421 (N_19421,N_16994,N_17931);
nor U19422 (N_19422,N_17636,N_17453);
or U19423 (N_19423,N_17240,N_16812);
and U19424 (N_19424,N_17531,N_16862);
xor U19425 (N_19425,N_16562,N_17644);
nand U19426 (N_19426,N_16908,N_17996);
and U19427 (N_19427,N_17314,N_16673);
nand U19428 (N_19428,N_17860,N_17750);
or U19429 (N_19429,N_16436,N_16914);
nor U19430 (N_19430,N_16920,N_17248);
or U19431 (N_19431,N_17229,N_16644);
and U19432 (N_19432,N_16417,N_16528);
xor U19433 (N_19433,N_16069,N_17647);
or U19434 (N_19434,N_17508,N_16946);
nor U19435 (N_19435,N_16163,N_17369);
nor U19436 (N_19436,N_17609,N_16160);
nor U19437 (N_19437,N_17582,N_16043);
and U19438 (N_19438,N_17751,N_17714);
nand U19439 (N_19439,N_17370,N_16398);
nand U19440 (N_19440,N_16323,N_16261);
nand U19441 (N_19441,N_17390,N_17179);
nor U19442 (N_19442,N_17229,N_16446);
nand U19443 (N_19443,N_17069,N_16548);
or U19444 (N_19444,N_16481,N_16072);
nor U19445 (N_19445,N_17021,N_17222);
or U19446 (N_19446,N_17567,N_17195);
or U19447 (N_19447,N_16020,N_16457);
nor U19448 (N_19448,N_17292,N_16110);
or U19449 (N_19449,N_16156,N_16576);
or U19450 (N_19450,N_17086,N_17541);
or U19451 (N_19451,N_16472,N_17587);
nand U19452 (N_19452,N_17302,N_17950);
nor U19453 (N_19453,N_16889,N_16835);
nor U19454 (N_19454,N_16812,N_17592);
nand U19455 (N_19455,N_16985,N_16170);
nor U19456 (N_19456,N_16342,N_16305);
nor U19457 (N_19457,N_17791,N_16018);
and U19458 (N_19458,N_17536,N_16320);
or U19459 (N_19459,N_16577,N_17220);
and U19460 (N_19460,N_17958,N_16083);
xnor U19461 (N_19461,N_17627,N_16072);
nand U19462 (N_19462,N_17779,N_16783);
nor U19463 (N_19463,N_17943,N_16101);
or U19464 (N_19464,N_17527,N_16046);
nand U19465 (N_19465,N_16382,N_17912);
nor U19466 (N_19466,N_16599,N_16958);
xor U19467 (N_19467,N_16065,N_17234);
xnor U19468 (N_19468,N_16232,N_16889);
and U19469 (N_19469,N_16140,N_17129);
nand U19470 (N_19470,N_16966,N_17032);
nor U19471 (N_19471,N_16901,N_16094);
xor U19472 (N_19472,N_16221,N_17063);
xnor U19473 (N_19473,N_16528,N_17761);
or U19474 (N_19474,N_17876,N_16253);
nand U19475 (N_19475,N_17297,N_17419);
and U19476 (N_19476,N_17629,N_16308);
nand U19477 (N_19477,N_16990,N_16247);
nand U19478 (N_19478,N_16795,N_17686);
nor U19479 (N_19479,N_17691,N_17922);
and U19480 (N_19480,N_16183,N_16651);
and U19481 (N_19481,N_17127,N_17681);
nand U19482 (N_19482,N_17708,N_16529);
nor U19483 (N_19483,N_17535,N_16440);
or U19484 (N_19484,N_16512,N_16401);
or U19485 (N_19485,N_16383,N_16323);
or U19486 (N_19486,N_17052,N_16909);
nand U19487 (N_19487,N_16595,N_17547);
nand U19488 (N_19488,N_17550,N_17491);
xor U19489 (N_19489,N_16742,N_17165);
nand U19490 (N_19490,N_16274,N_17330);
nor U19491 (N_19491,N_17688,N_16488);
nand U19492 (N_19492,N_16967,N_16537);
and U19493 (N_19493,N_16229,N_17693);
and U19494 (N_19494,N_17245,N_16125);
nor U19495 (N_19495,N_17030,N_16946);
and U19496 (N_19496,N_17266,N_16001);
and U19497 (N_19497,N_16462,N_16456);
and U19498 (N_19498,N_16229,N_17163);
nand U19499 (N_19499,N_17396,N_16826);
and U19500 (N_19500,N_16916,N_16241);
nor U19501 (N_19501,N_16909,N_17901);
xor U19502 (N_19502,N_17359,N_16745);
or U19503 (N_19503,N_17331,N_17805);
and U19504 (N_19504,N_17076,N_17051);
and U19505 (N_19505,N_16246,N_17886);
xnor U19506 (N_19506,N_16946,N_17787);
and U19507 (N_19507,N_17693,N_16550);
and U19508 (N_19508,N_16962,N_17669);
or U19509 (N_19509,N_17056,N_16882);
and U19510 (N_19510,N_17267,N_17172);
and U19511 (N_19511,N_16456,N_17854);
nand U19512 (N_19512,N_16294,N_16851);
nor U19513 (N_19513,N_16247,N_16868);
and U19514 (N_19514,N_17896,N_17785);
nor U19515 (N_19515,N_17059,N_16945);
xnor U19516 (N_19516,N_16485,N_17621);
xnor U19517 (N_19517,N_17766,N_16191);
nor U19518 (N_19518,N_17307,N_17031);
and U19519 (N_19519,N_17357,N_16206);
and U19520 (N_19520,N_16864,N_16379);
or U19521 (N_19521,N_17902,N_17151);
or U19522 (N_19522,N_16635,N_17120);
nor U19523 (N_19523,N_17790,N_17381);
xnor U19524 (N_19524,N_16661,N_17522);
and U19525 (N_19525,N_16155,N_16531);
nor U19526 (N_19526,N_17956,N_17099);
xor U19527 (N_19527,N_17383,N_17230);
or U19528 (N_19528,N_16943,N_17054);
or U19529 (N_19529,N_17408,N_16780);
xor U19530 (N_19530,N_17964,N_16892);
and U19531 (N_19531,N_17867,N_17204);
nand U19532 (N_19532,N_16777,N_17624);
or U19533 (N_19533,N_16171,N_16039);
and U19534 (N_19534,N_16948,N_16545);
xor U19535 (N_19535,N_16582,N_17522);
nand U19536 (N_19536,N_16834,N_17433);
xor U19537 (N_19537,N_16881,N_17650);
xor U19538 (N_19538,N_17392,N_17340);
and U19539 (N_19539,N_17278,N_17589);
nor U19540 (N_19540,N_16969,N_17668);
or U19541 (N_19541,N_16074,N_17850);
xor U19542 (N_19542,N_17511,N_16148);
xnor U19543 (N_19543,N_17249,N_16786);
xnor U19544 (N_19544,N_17115,N_16985);
or U19545 (N_19545,N_16150,N_16763);
nor U19546 (N_19546,N_16008,N_17641);
nand U19547 (N_19547,N_17183,N_16185);
or U19548 (N_19548,N_16202,N_16363);
nor U19549 (N_19549,N_17270,N_17108);
nor U19550 (N_19550,N_17502,N_16574);
nor U19551 (N_19551,N_17830,N_17691);
or U19552 (N_19552,N_16297,N_17573);
or U19553 (N_19553,N_16353,N_17728);
and U19554 (N_19554,N_17710,N_16097);
and U19555 (N_19555,N_16108,N_17330);
and U19556 (N_19556,N_17380,N_16163);
xnor U19557 (N_19557,N_16032,N_16764);
and U19558 (N_19558,N_17398,N_16051);
xnor U19559 (N_19559,N_16164,N_16509);
xor U19560 (N_19560,N_17258,N_16616);
nor U19561 (N_19561,N_16104,N_16189);
and U19562 (N_19562,N_17731,N_16757);
nand U19563 (N_19563,N_17636,N_17784);
and U19564 (N_19564,N_16206,N_17024);
or U19565 (N_19565,N_16175,N_17990);
xor U19566 (N_19566,N_16378,N_16361);
or U19567 (N_19567,N_17045,N_16129);
or U19568 (N_19568,N_16136,N_16612);
nor U19569 (N_19569,N_16793,N_16295);
xnor U19570 (N_19570,N_16479,N_16281);
nand U19571 (N_19571,N_17406,N_16725);
and U19572 (N_19572,N_17311,N_17938);
and U19573 (N_19573,N_17974,N_16270);
or U19574 (N_19574,N_16242,N_17675);
xor U19575 (N_19575,N_16135,N_17721);
or U19576 (N_19576,N_16222,N_16679);
or U19577 (N_19577,N_16101,N_16972);
nand U19578 (N_19578,N_17570,N_17067);
nor U19579 (N_19579,N_17075,N_16772);
or U19580 (N_19580,N_16059,N_16920);
nor U19581 (N_19581,N_17160,N_16045);
and U19582 (N_19582,N_16688,N_16814);
xnor U19583 (N_19583,N_16974,N_16387);
or U19584 (N_19584,N_16847,N_17014);
and U19585 (N_19585,N_17570,N_16676);
or U19586 (N_19586,N_17011,N_16319);
nor U19587 (N_19587,N_16097,N_17025);
and U19588 (N_19588,N_16991,N_17016);
or U19589 (N_19589,N_16086,N_17192);
nor U19590 (N_19590,N_17378,N_17878);
nand U19591 (N_19591,N_17950,N_16307);
xor U19592 (N_19592,N_17838,N_16763);
xor U19593 (N_19593,N_17274,N_17339);
nor U19594 (N_19594,N_16417,N_17814);
or U19595 (N_19595,N_16521,N_17571);
and U19596 (N_19596,N_16327,N_17278);
xnor U19597 (N_19597,N_16702,N_17440);
xor U19598 (N_19598,N_16416,N_16665);
nand U19599 (N_19599,N_16660,N_16146);
or U19600 (N_19600,N_17014,N_17388);
and U19601 (N_19601,N_16825,N_17169);
and U19602 (N_19602,N_17352,N_17792);
nand U19603 (N_19603,N_16229,N_16631);
nor U19604 (N_19604,N_17792,N_17501);
nor U19605 (N_19605,N_17531,N_17752);
nand U19606 (N_19606,N_16180,N_16880);
and U19607 (N_19607,N_17823,N_17382);
or U19608 (N_19608,N_16940,N_17405);
and U19609 (N_19609,N_17371,N_17492);
xnor U19610 (N_19610,N_17529,N_16959);
and U19611 (N_19611,N_16273,N_16111);
nand U19612 (N_19612,N_17565,N_16356);
and U19613 (N_19613,N_17230,N_17458);
nand U19614 (N_19614,N_16277,N_16819);
and U19615 (N_19615,N_17402,N_16598);
nand U19616 (N_19616,N_17957,N_16363);
and U19617 (N_19617,N_16079,N_16120);
and U19618 (N_19618,N_16086,N_17878);
nor U19619 (N_19619,N_17495,N_16912);
nand U19620 (N_19620,N_16236,N_16859);
xor U19621 (N_19621,N_16604,N_17152);
nand U19622 (N_19622,N_17920,N_16198);
and U19623 (N_19623,N_17635,N_17087);
and U19624 (N_19624,N_16072,N_17055);
or U19625 (N_19625,N_17446,N_16028);
nor U19626 (N_19626,N_17436,N_17921);
nand U19627 (N_19627,N_17763,N_16311);
nand U19628 (N_19628,N_16446,N_16008);
xnor U19629 (N_19629,N_16126,N_17427);
or U19630 (N_19630,N_16565,N_16490);
nand U19631 (N_19631,N_17962,N_17759);
nand U19632 (N_19632,N_17892,N_17754);
xnor U19633 (N_19633,N_16927,N_17357);
nand U19634 (N_19634,N_17254,N_16951);
and U19635 (N_19635,N_17763,N_16361);
or U19636 (N_19636,N_17725,N_16400);
or U19637 (N_19637,N_16809,N_16570);
nand U19638 (N_19638,N_16006,N_16560);
xor U19639 (N_19639,N_16724,N_16753);
or U19640 (N_19640,N_16776,N_16501);
xnor U19641 (N_19641,N_17700,N_16042);
nand U19642 (N_19642,N_17596,N_16230);
and U19643 (N_19643,N_16355,N_17310);
and U19644 (N_19644,N_17549,N_17855);
xor U19645 (N_19645,N_16640,N_17418);
xnor U19646 (N_19646,N_17695,N_16024);
nor U19647 (N_19647,N_17207,N_17285);
and U19648 (N_19648,N_17498,N_16993);
or U19649 (N_19649,N_16934,N_16234);
xor U19650 (N_19650,N_17808,N_17034);
nor U19651 (N_19651,N_17503,N_16289);
or U19652 (N_19652,N_17444,N_17046);
xnor U19653 (N_19653,N_17544,N_17145);
xnor U19654 (N_19654,N_17256,N_16611);
xnor U19655 (N_19655,N_16960,N_16627);
xor U19656 (N_19656,N_16586,N_16181);
xnor U19657 (N_19657,N_16625,N_17378);
or U19658 (N_19658,N_16877,N_17889);
or U19659 (N_19659,N_16031,N_17208);
nor U19660 (N_19660,N_16929,N_17408);
xor U19661 (N_19661,N_17508,N_17210);
xor U19662 (N_19662,N_16240,N_16438);
xnor U19663 (N_19663,N_17916,N_17811);
nand U19664 (N_19664,N_16289,N_16463);
and U19665 (N_19665,N_17225,N_17281);
and U19666 (N_19666,N_17914,N_17096);
nor U19667 (N_19667,N_17914,N_17166);
nor U19668 (N_19668,N_17913,N_16210);
xnor U19669 (N_19669,N_16593,N_17185);
or U19670 (N_19670,N_16304,N_17276);
or U19671 (N_19671,N_16166,N_16357);
or U19672 (N_19672,N_17150,N_16590);
nand U19673 (N_19673,N_17862,N_17298);
or U19674 (N_19674,N_17719,N_16819);
or U19675 (N_19675,N_16199,N_17153);
and U19676 (N_19676,N_17805,N_16023);
nor U19677 (N_19677,N_17667,N_17949);
and U19678 (N_19678,N_16925,N_17318);
nand U19679 (N_19679,N_16754,N_17319);
nand U19680 (N_19680,N_17979,N_17334);
or U19681 (N_19681,N_16086,N_16130);
xor U19682 (N_19682,N_17329,N_16229);
nor U19683 (N_19683,N_16387,N_16410);
nand U19684 (N_19684,N_17378,N_16272);
nand U19685 (N_19685,N_17292,N_16388);
nor U19686 (N_19686,N_17031,N_16102);
or U19687 (N_19687,N_17703,N_16638);
nor U19688 (N_19688,N_17765,N_16264);
xor U19689 (N_19689,N_16766,N_17346);
xnor U19690 (N_19690,N_16690,N_17933);
nor U19691 (N_19691,N_17711,N_17502);
nand U19692 (N_19692,N_16919,N_16353);
or U19693 (N_19693,N_16411,N_16857);
nand U19694 (N_19694,N_16524,N_17879);
xor U19695 (N_19695,N_17118,N_17909);
xnor U19696 (N_19696,N_17454,N_16771);
and U19697 (N_19697,N_16758,N_16167);
nand U19698 (N_19698,N_16778,N_16596);
xnor U19699 (N_19699,N_16737,N_17554);
nand U19700 (N_19700,N_17947,N_17404);
xnor U19701 (N_19701,N_17544,N_17833);
nand U19702 (N_19702,N_16093,N_17967);
and U19703 (N_19703,N_16255,N_17943);
and U19704 (N_19704,N_17964,N_17585);
nor U19705 (N_19705,N_16377,N_16818);
nor U19706 (N_19706,N_16297,N_17953);
and U19707 (N_19707,N_17432,N_17504);
xor U19708 (N_19708,N_17809,N_16375);
or U19709 (N_19709,N_16236,N_16166);
or U19710 (N_19710,N_17449,N_16542);
xor U19711 (N_19711,N_17916,N_17045);
nor U19712 (N_19712,N_16479,N_17422);
nor U19713 (N_19713,N_16203,N_17198);
nand U19714 (N_19714,N_17514,N_16279);
nand U19715 (N_19715,N_17055,N_17512);
nor U19716 (N_19716,N_16306,N_16936);
nor U19717 (N_19717,N_17133,N_16701);
nand U19718 (N_19718,N_17666,N_17131);
or U19719 (N_19719,N_16570,N_17333);
nor U19720 (N_19720,N_16405,N_16481);
nand U19721 (N_19721,N_16144,N_16986);
or U19722 (N_19722,N_17727,N_17192);
nand U19723 (N_19723,N_17898,N_17991);
nand U19724 (N_19724,N_16492,N_16459);
nor U19725 (N_19725,N_17372,N_17439);
nand U19726 (N_19726,N_16631,N_16886);
nor U19727 (N_19727,N_16077,N_16233);
or U19728 (N_19728,N_16536,N_16131);
nand U19729 (N_19729,N_16933,N_17868);
and U19730 (N_19730,N_16124,N_17170);
xor U19731 (N_19731,N_17120,N_16515);
and U19732 (N_19732,N_17236,N_17286);
and U19733 (N_19733,N_16493,N_17447);
or U19734 (N_19734,N_16156,N_17626);
xnor U19735 (N_19735,N_17242,N_17976);
and U19736 (N_19736,N_17821,N_16495);
and U19737 (N_19737,N_16872,N_17600);
xor U19738 (N_19738,N_16130,N_16361);
and U19739 (N_19739,N_17312,N_16973);
nor U19740 (N_19740,N_17982,N_16189);
nor U19741 (N_19741,N_17706,N_17092);
nor U19742 (N_19742,N_16014,N_17053);
xor U19743 (N_19743,N_16356,N_17113);
or U19744 (N_19744,N_17588,N_17360);
nand U19745 (N_19745,N_17023,N_17384);
nor U19746 (N_19746,N_16985,N_16119);
and U19747 (N_19747,N_16793,N_16807);
or U19748 (N_19748,N_16974,N_17464);
nand U19749 (N_19749,N_17094,N_17584);
xor U19750 (N_19750,N_16315,N_17706);
xnor U19751 (N_19751,N_17501,N_17789);
nand U19752 (N_19752,N_17669,N_17060);
nand U19753 (N_19753,N_17110,N_17456);
and U19754 (N_19754,N_16313,N_17406);
nand U19755 (N_19755,N_17001,N_17788);
nor U19756 (N_19756,N_16571,N_17173);
and U19757 (N_19757,N_16909,N_17908);
xor U19758 (N_19758,N_17301,N_16730);
or U19759 (N_19759,N_16240,N_17816);
nand U19760 (N_19760,N_16655,N_17512);
nand U19761 (N_19761,N_16276,N_16907);
xnor U19762 (N_19762,N_16085,N_17895);
or U19763 (N_19763,N_17166,N_16811);
and U19764 (N_19764,N_17302,N_17061);
nand U19765 (N_19765,N_16321,N_17544);
or U19766 (N_19766,N_16308,N_17880);
and U19767 (N_19767,N_16344,N_17947);
nor U19768 (N_19768,N_16040,N_16892);
and U19769 (N_19769,N_17932,N_17815);
xor U19770 (N_19770,N_17825,N_17795);
xor U19771 (N_19771,N_16340,N_17874);
xor U19772 (N_19772,N_16132,N_17822);
nand U19773 (N_19773,N_16973,N_17983);
xnor U19774 (N_19774,N_17259,N_17150);
or U19775 (N_19775,N_16190,N_16480);
xnor U19776 (N_19776,N_17902,N_16903);
nor U19777 (N_19777,N_16078,N_17229);
nand U19778 (N_19778,N_17286,N_16479);
and U19779 (N_19779,N_17273,N_16609);
xor U19780 (N_19780,N_17546,N_16322);
nor U19781 (N_19781,N_17450,N_17169);
or U19782 (N_19782,N_17937,N_16564);
and U19783 (N_19783,N_17661,N_17365);
nor U19784 (N_19784,N_17290,N_16195);
xor U19785 (N_19785,N_16329,N_17327);
nand U19786 (N_19786,N_16291,N_16679);
nand U19787 (N_19787,N_17113,N_17928);
xor U19788 (N_19788,N_16898,N_16368);
nand U19789 (N_19789,N_16192,N_16731);
xnor U19790 (N_19790,N_17232,N_17201);
nand U19791 (N_19791,N_16139,N_16150);
or U19792 (N_19792,N_16572,N_16909);
or U19793 (N_19793,N_17675,N_17114);
or U19794 (N_19794,N_17567,N_16635);
and U19795 (N_19795,N_16462,N_16998);
nor U19796 (N_19796,N_16611,N_16463);
xor U19797 (N_19797,N_17361,N_17907);
nor U19798 (N_19798,N_17761,N_16801);
nand U19799 (N_19799,N_17063,N_16608);
nor U19800 (N_19800,N_16731,N_16269);
or U19801 (N_19801,N_17585,N_17813);
or U19802 (N_19802,N_17068,N_16271);
nor U19803 (N_19803,N_16145,N_16822);
or U19804 (N_19804,N_16553,N_17344);
and U19805 (N_19805,N_16986,N_16830);
xor U19806 (N_19806,N_16201,N_17586);
or U19807 (N_19807,N_17963,N_16666);
and U19808 (N_19808,N_17411,N_17046);
xor U19809 (N_19809,N_17548,N_17201);
nor U19810 (N_19810,N_16526,N_16784);
nand U19811 (N_19811,N_16832,N_16261);
and U19812 (N_19812,N_17473,N_16692);
nand U19813 (N_19813,N_16605,N_17089);
nor U19814 (N_19814,N_16886,N_17212);
nand U19815 (N_19815,N_17943,N_17328);
or U19816 (N_19816,N_17546,N_16939);
or U19817 (N_19817,N_17880,N_16230);
nor U19818 (N_19818,N_17096,N_17078);
and U19819 (N_19819,N_16397,N_16169);
or U19820 (N_19820,N_16695,N_16603);
nand U19821 (N_19821,N_16403,N_17062);
and U19822 (N_19822,N_17868,N_17437);
nand U19823 (N_19823,N_17847,N_17027);
nor U19824 (N_19824,N_16364,N_16433);
xor U19825 (N_19825,N_17610,N_17120);
xor U19826 (N_19826,N_16224,N_17361);
nor U19827 (N_19827,N_16585,N_17684);
or U19828 (N_19828,N_16069,N_16925);
and U19829 (N_19829,N_16536,N_16270);
and U19830 (N_19830,N_17530,N_16447);
and U19831 (N_19831,N_17834,N_17549);
or U19832 (N_19832,N_17575,N_16714);
xnor U19833 (N_19833,N_16196,N_16037);
nor U19834 (N_19834,N_17865,N_17629);
xor U19835 (N_19835,N_16450,N_17411);
xor U19836 (N_19836,N_17929,N_16299);
and U19837 (N_19837,N_16720,N_16136);
or U19838 (N_19838,N_16588,N_16085);
or U19839 (N_19839,N_17861,N_17240);
nand U19840 (N_19840,N_17582,N_16408);
nor U19841 (N_19841,N_17873,N_17969);
nand U19842 (N_19842,N_16537,N_17284);
nand U19843 (N_19843,N_17833,N_17714);
xnor U19844 (N_19844,N_16171,N_17156);
and U19845 (N_19845,N_17194,N_16154);
xnor U19846 (N_19846,N_16381,N_17861);
and U19847 (N_19847,N_16302,N_17136);
nand U19848 (N_19848,N_16066,N_17923);
nor U19849 (N_19849,N_16285,N_17593);
and U19850 (N_19850,N_16014,N_17325);
xor U19851 (N_19851,N_17922,N_17312);
nand U19852 (N_19852,N_17609,N_16803);
and U19853 (N_19853,N_16450,N_17257);
nand U19854 (N_19854,N_16524,N_16452);
and U19855 (N_19855,N_17152,N_16666);
nand U19856 (N_19856,N_17292,N_16637);
nor U19857 (N_19857,N_17596,N_16416);
nand U19858 (N_19858,N_17019,N_17559);
nor U19859 (N_19859,N_17045,N_17308);
and U19860 (N_19860,N_17592,N_17681);
or U19861 (N_19861,N_16820,N_17833);
nor U19862 (N_19862,N_17831,N_16014);
and U19863 (N_19863,N_17927,N_16928);
nor U19864 (N_19864,N_17927,N_17916);
nor U19865 (N_19865,N_17659,N_17074);
or U19866 (N_19866,N_16449,N_17715);
xor U19867 (N_19867,N_17717,N_17126);
and U19868 (N_19868,N_16336,N_16138);
nor U19869 (N_19869,N_17205,N_16384);
or U19870 (N_19870,N_17856,N_16510);
nor U19871 (N_19871,N_17467,N_16726);
nor U19872 (N_19872,N_16788,N_17473);
nor U19873 (N_19873,N_17460,N_17384);
and U19874 (N_19874,N_16089,N_17127);
nor U19875 (N_19875,N_16303,N_17750);
or U19876 (N_19876,N_17881,N_16732);
nor U19877 (N_19877,N_16330,N_17915);
nand U19878 (N_19878,N_17696,N_17095);
xnor U19879 (N_19879,N_16620,N_17338);
nor U19880 (N_19880,N_16661,N_16756);
and U19881 (N_19881,N_16603,N_17966);
xnor U19882 (N_19882,N_16181,N_17523);
nor U19883 (N_19883,N_16295,N_17353);
and U19884 (N_19884,N_17296,N_17395);
nor U19885 (N_19885,N_16944,N_17336);
nor U19886 (N_19886,N_16824,N_16530);
nor U19887 (N_19887,N_17076,N_17823);
nand U19888 (N_19888,N_16486,N_17780);
or U19889 (N_19889,N_17110,N_17950);
nand U19890 (N_19890,N_16699,N_16724);
and U19891 (N_19891,N_17332,N_17282);
and U19892 (N_19892,N_17226,N_16466);
nor U19893 (N_19893,N_17741,N_16674);
xnor U19894 (N_19894,N_17073,N_16308);
xor U19895 (N_19895,N_17453,N_16184);
and U19896 (N_19896,N_17649,N_16696);
and U19897 (N_19897,N_17537,N_16288);
nand U19898 (N_19898,N_17730,N_17827);
nor U19899 (N_19899,N_17563,N_16346);
xor U19900 (N_19900,N_16282,N_17161);
xnor U19901 (N_19901,N_16943,N_17503);
nand U19902 (N_19902,N_17318,N_16732);
nand U19903 (N_19903,N_16545,N_17114);
and U19904 (N_19904,N_17603,N_17620);
or U19905 (N_19905,N_16523,N_17991);
nor U19906 (N_19906,N_16209,N_16900);
nand U19907 (N_19907,N_16213,N_17888);
and U19908 (N_19908,N_16266,N_16574);
nand U19909 (N_19909,N_17484,N_16749);
xnor U19910 (N_19910,N_16399,N_17115);
and U19911 (N_19911,N_16222,N_16281);
and U19912 (N_19912,N_17803,N_17967);
or U19913 (N_19913,N_17445,N_17453);
nor U19914 (N_19914,N_17335,N_16000);
nand U19915 (N_19915,N_16405,N_16157);
and U19916 (N_19916,N_16554,N_16359);
nor U19917 (N_19917,N_16193,N_16535);
xor U19918 (N_19918,N_16400,N_17936);
nor U19919 (N_19919,N_16887,N_16208);
xnor U19920 (N_19920,N_17357,N_16858);
or U19921 (N_19921,N_16418,N_17095);
or U19922 (N_19922,N_17880,N_16284);
nor U19923 (N_19923,N_16349,N_16772);
nor U19924 (N_19924,N_17337,N_17667);
or U19925 (N_19925,N_17265,N_17683);
xnor U19926 (N_19926,N_17573,N_16802);
and U19927 (N_19927,N_17449,N_17847);
nand U19928 (N_19928,N_17701,N_17184);
or U19929 (N_19929,N_16387,N_17314);
nor U19930 (N_19930,N_16768,N_16219);
or U19931 (N_19931,N_16820,N_17670);
xnor U19932 (N_19932,N_16199,N_16362);
or U19933 (N_19933,N_16076,N_17144);
nand U19934 (N_19934,N_16281,N_17797);
nand U19935 (N_19935,N_17825,N_16543);
nand U19936 (N_19936,N_17435,N_17058);
nor U19937 (N_19937,N_17461,N_17153);
and U19938 (N_19938,N_16703,N_16756);
nor U19939 (N_19939,N_17586,N_17947);
nand U19940 (N_19940,N_16109,N_16537);
nand U19941 (N_19941,N_16443,N_17425);
nand U19942 (N_19942,N_17284,N_17130);
nor U19943 (N_19943,N_16071,N_16451);
and U19944 (N_19944,N_16405,N_16508);
and U19945 (N_19945,N_17092,N_17842);
nor U19946 (N_19946,N_17257,N_16805);
or U19947 (N_19947,N_16240,N_16674);
and U19948 (N_19948,N_16463,N_16989);
nor U19949 (N_19949,N_16048,N_17972);
and U19950 (N_19950,N_16571,N_16766);
and U19951 (N_19951,N_17097,N_16715);
nor U19952 (N_19952,N_16126,N_17477);
nand U19953 (N_19953,N_16849,N_16793);
nor U19954 (N_19954,N_16895,N_17365);
xor U19955 (N_19955,N_17059,N_17022);
xnor U19956 (N_19956,N_16640,N_16260);
xnor U19957 (N_19957,N_17546,N_17882);
and U19958 (N_19958,N_17445,N_16901);
and U19959 (N_19959,N_17847,N_17162);
xor U19960 (N_19960,N_17916,N_16337);
xnor U19961 (N_19961,N_17549,N_17978);
nor U19962 (N_19962,N_17745,N_16488);
nand U19963 (N_19963,N_16592,N_16550);
xor U19964 (N_19964,N_17620,N_16533);
nand U19965 (N_19965,N_17982,N_17794);
xor U19966 (N_19966,N_17066,N_16729);
nor U19967 (N_19967,N_17602,N_17162);
or U19968 (N_19968,N_16850,N_17813);
nand U19969 (N_19969,N_16788,N_17271);
nand U19970 (N_19970,N_16716,N_17458);
or U19971 (N_19971,N_16696,N_17898);
xnor U19972 (N_19972,N_17212,N_17441);
and U19973 (N_19973,N_16131,N_17077);
nand U19974 (N_19974,N_17305,N_17432);
nor U19975 (N_19975,N_17500,N_17001);
nor U19976 (N_19976,N_16169,N_17437);
and U19977 (N_19977,N_17725,N_16464);
nand U19978 (N_19978,N_16666,N_16230);
nand U19979 (N_19979,N_16814,N_17426);
nor U19980 (N_19980,N_16435,N_16723);
or U19981 (N_19981,N_16228,N_17523);
nor U19982 (N_19982,N_17518,N_16129);
nand U19983 (N_19983,N_17129,N_16125);
or U19984 (N_19984,N_17441,N_17667);
nor U19985 (N_19985,N_17099,N_17226);
and U19986 (N_19986,N_16380,N_17231);
nor U19987 (N_19987,N_17457,N_16211);
or U19988 (N_19988,N_17215,N_17522);
nor U19989 (N_19989,N_16516,N_16281);
or U19990 (N_19990,N_16564,N_17436);
and U19991 (N_19991,N_17917,N_16929);
xnor U19992 (N_19992,N_16951,N_16484);
or U19993 (N_19993,N_17603,N_17510);
nor U19994 (N_19994,N_16450,N_17275);
nor U19995 (N_19995,N_16052,N_16370);
nor U19996 (N_19996,N_17857,N_17984);
nor U19997 (N_19997,N_16602,N_17923);
nand U19998 (N_19998,N_16107,N_17486);
and U19999 (N_19999,N_16373,N_16578);
xnor U20000 (N_20000,N_18062,N_19051);
xnor U20001 (N_20001,N_18731,N_18971);
xnor U20002 (N_20002,N_19953,N_18986);
nor U20003 (N_20003,N_19490,N_18614);
or U20004 (N_20004,N_19140,N_19338);
xor U20005 (N_20005,N_18835,N_19088);
nand U20006 (N_20006,N_18354,N_19450);
and U20007 (N_20007,N_19472,N_19565);
nor U20008 (N_20008,N_18815,N_19353);
and U20009 (N_20009,N_19530,N_19112);
nor U20010 (N_20010,N_19972,N_18647);
xor U20011 (N_20011,N_18782,N_19185);
nand U20012 (N_20012,N_18116,N_18444);
or U20013 (N_20013,N_18576,N_18405);
or U20014 (N_20014,N_18061,N_19485);
and U20015 (N_20015,N_18644,N_19725);
xor U20016 (N_20016,N_19383,N_18247);
and U20017 (N_20017,N_18013,N_19645);
or U20018 (N_20018,N_18775,N_19853);
or U20019 (N_20019,N_18708,N_18492);
nor U20020 (N_20020,N_19003,N_19376);
xor U20021 (N_20021,N_18888,N_19845);
xor U20022 (N_20022,N_19087,N_18338);
nand U20023 (N_20023,N_18886,N_18317);
nor U20024 (N_20024,N_19979,N_19504);
or U20025 (N_20025,N_18240,N_19539);
or U20026 (N_20026,N_18617,N_19055);
xor U20027 (N_20027,N_19021,N_19555);
nand U20028 (N_20028,N_19017,N_19924);
nand U20029 (N_20029,N_19095,N_18859);
xnor U20030 (N_20030,N_18352,N_19451);
nor U20031 (N_20031,N_19691,N_19908);
nand U20032 (N_20032,N_19946,N_19011);
or U20033 (N_20033,N_19998,N_18229);
xnor U20034 (N_20034,N_18372,N_19640);
xor U20035 (N_20035,N_19697,N_18106);
nand U20036 (N_20036,N_19287,N_19015);
and U20037 (N_20037,N_19390,N_18786);
and U20038 (N_20038,N_18509,N_18831);
xor U20039 (N_20039,N_18760,N_18908);
nor U20040 (N_20040,N_18281,N_18422);
and U20041 (N_20041,N_18494,N_19005);
nor U20042 (N_20042,N_18022,N_18525);
or U20043 (N_20043,N_18611,N_18928);
xor U20044 (N_20044,N_18342,N_18858);
xnor U20045 (N_20045,N_19121,N_18333);
nand U20046 (N_20046,N_19856,N_19909);
or U20047 (N_20047,N_19732,N_19476);
or U20048 (N_20048,N_18748,N_18954);
xnor U20049 (N_20049,N_19742,N_19984);
or U20050 (N_20050,N_18181,N_18121);
or U20051 (N_20051,N_18452,N_18083);
xor U20052 (N_20052,N_19409,N_18995);
or U20053 (N_20053,N_18699,N_19335);
nor U20054 (N_20054,N_19291,N_18103);
and U20055 (N_20055,N_18978,N_19801);
and U20056 (N_20056,N_19181,N_19010);
xnor U20057 (N_20057,N_19913,N_19880);
nand U20058 (N_20058,N_19760,N_18958);
xnor U20059 (N_20059,N_18302,N_19431);
nor U20060 (N_20060,N_19144,N_18718);
nor U20061 (N_20061,N_18001,N_18358);
or U20062 (N_20062,N_19631,N_19001);
or U20063 (N_20063,N_19955,N_19411);
xor U20064 (N_20064,N_19986,N_18568);
or U20065 (N_20065,N_18111,N_18047);
xor U20066 (N_20066,N_18015,N_19568);
nand U20067 (N_20067,N_19625,N_18987);
nor U20068 (N_20068,N_19414,N_19574);
xor U20069 (N_20069,N_19728,N_18080);
and U20070 (N_20070,N_18843,N_19292);
xnor U20071 (N_20071,N_18875,N_18553);
and U20072 (N_20072,N_18988,N_18286);
nand U20073 (N_20073,N_19293,N_18517);
nor U20074 (N_20074,N_18341,N_18176);
or U20075 (N_20075,N_18648,N_19024);
xor U20076 (N_20076,N_19107,N_19586);
nand U20077 (N_20077,N_19670,N_19580);
nand U20078 (N_20078,N_18051,N_19309);
nand U20079 (N_20079,N_19723,N_18747);
nand U20080 (N_20080,N_19378,N_19491);
nand U20081 (N_20081,N_18736,N_18825);
nand U20082 (N_20082,N_18994,N_18897);
nor U20083 (N_20083,N_18998,N_19030);
or U20084 (N_20084,N_18232,N_19759);
or U20085 (N_20085,N_18651,N_19859);
and U20086 (N_20086,N_19086,N_19848);
xnor U20087 (N_20087,N_18893,N_18441);
or U20088 (N_20088,N_18909,N_19989);
nand U20089 (N_20089,N_18299,N_19246);
xnor U20090 (N_20090,N_19754,N_19791);
and U20091 (N_20091,N_19306,N_18347);
or U20092 (N_20092,N_18570,N_18841);
or U20093 (N_20093,N_18857,N_18134);
nand U20094 (N_20094,N_18283,N_19199);
xnor U20095 (N_20095,N_19193,N_19289);
xor U20096 (N_20096,N_18887,N_19183);
xor U20097 (N_20097,N_18109,N_19660);
and U20098 (N_20098,N_18690,N_19581);
and U20099 (N_20099,N_18534,N_18707);
xor U20100 (N_20100,N_18619,N_19419);
and U20101 (N_20101,N_18860,N_18253);
nor U20102 (N_20102,N_18011,N_19659);
and U20103 (N_20103,N_18276,N_18749);
and U20104 (N_20104,N_18673,N_18429);
nand U20105 (N_20105,N_18810,N_19943);
xor U20106 (N_20106,N_18615,N_18064);
or U20107 (N_20107,N_18365,N_18221);
nor U20108 (N_20108,N_19970,N_18059);
nor U20109 (N_20109,N_19620,N_18379);
xor U20110 (N_20110,N_19784,N_19263);
nor U20111 (N_20111,N_18472,N_18003);
nor U20112 (N_20112,N_18495,N_18682);
xor U20113 (N_20113,N_19212,N_18091);
xnor U20114 (N_20114,N_19394,N_19014);
nand U20115 (N_20115,N_19059,N_18496);
and U20116 (N_20116,N_19142,N_19458);
or U20117 (N_20117,N_19919,N_19375);
or U20118 (N_20118,N_19103,N_19060);
nor U20119 (N_20119,N_18703,N_19813);
xnor U20120 (N_20120,N_19843,N_18331);
nand U20121 (N_20121,N_18827,N_19531);
and U20122 (N_20122,N_18766,N_18204);
nand U20123 (N_20123,N_19905,N_18095);
xnor U20124 (N_20124,N_18222,N_19439);
nand U20125 (N_20125,N_19332,N_18813);
or U20126 (N_20126,N_19280,N_18520);
nor U20127 (N_20127,N_18265,N_19285);
nor U20128 (N_20128,N_19435,N_18845);
xnor U20129 (N_20129,N_19511,N_19399);
nor U20130 (N_20130,N_19552,N_19178);
xnor U20131 (N_20131,N_19713,N_19622);
nand U20132 (N_20132,N_18772,N_18260);
nand U20133 (N_20133,N_19255,N_19778);
nor U20134 (N_20134,N_18144,N_19575);
nand U20135 (N_20135,N_19223,N_19685);
nor U20136 (N_20136,N_19453,N_18256);
nor U20137 (N_20137,N_19669,N_18921);
or U20138 (N_20138,N_18547,N_19388);
and U20139 (N_20139,N_19166,N_18211);
nor U20140 (N_20140,N_18814,N_19649);
nand U20141 (N_20141,N_18744,N_18851);
and U20142 (N_20142,N_19612,N_19683);
nor U20143 (N_20143,N_18044,N_18470);
nor U20144 (N_20144,N_18196,N_19762);
or U20145 (N_20145,N_19259,N_18239);
nor U20146 (N_20146,N_18562,N_18397);
nor U20147 (N_20147,N_18582,N_18032);
xor U20148 (N_20148,N_19392,N_19161);
nand U20149 (N_20149,N_19308,N_19823);
xnor U20150 (N_20150,N_18267,N_19885);
or U20151 (N_20151,N_19057,N_18459);
xnor U20152 (N_20152,N_19701,N_18714);
xor U20153 (N_20153,N_18237,N_19344);
or U20154 (N_20154,N_19237,N_19933);
and U20155 (N_20155,N_19960,N_19500);
xor U20156 (N_20156,N_19747,N_18764);
and U20157 (N_20157,N_19047,N_19693);
nor U20158 (N_20158,N_19618,N_18923);
nor U20159 (N_20159,N_18861,N_19863);
nand U20160 (N_20160,N_19895,N_19652);
nand U20161 (N_20161,N_18991,N_18193);
or U20162 (N_20162,N_18770,N_18242);
or U20163 (N_20163,N_18440,N_19318);
and U20164 (N_20164,N_19882,N_18901);
xnor U20165 (N_20165,N_19427,N_19825);
and U20166 (N_20166,N_18637,N_18633);
or U20167 (N_20167,N_19042,N_18321);
xor U20168 (N_20168,N_19039,N_19331);
nor U20169 (N_20169,N_19727,N_18305);
xnor U20170 (N_20170,N_19113,N_19459);
xor U20171 (N_20171,N_19938,N_18937);
or U20172 (N_20172,N_19780,N_19231);
nor U20173 (N_20173,N_18866,N_18005);
and U20174 (N_20174,N_18498,N_19815);
xnor U20175 (N_20175,N_18178,N_19334);
nand U20176 (N_20176,N_18235,N_19322);
xnor U20177 (N_20177,N_19311,N_19248);
and U20178 (N_20178,N_18752,N_18674);
nand U20179 (N_20179,N_19177,N_19266);
nand U20180 (N_20180,N_19934,N_19542);
xnor U20181 (N_20181,N_18130,N_18241);
nand U20182 (N_20182,N_18628,N_19134);
and U20183 (N_20183,N_18603,N_19797);
and U20184 (N_20184,N_19785,N_18107);
nor U20185 (N_20185,N_18082,N_18715);
nor U20186 (N_20186,N_19601,N_18497);
xor U20187 (N_20187,N_18504,N_18078);
nand U20188 (N_20188,N_19241,N_18550);
xor U20189 (N_20189,N_19428,N_19209);
nor U20190 (N_20190,N_19092,N_19692);
and U20191 (N_20191,N_18934,N_19886);
or U20192 (N_20192,N_19977,N_19589);
nand U20193 (N_20193,N_19556,N_18931);
or U20194 (N_20194,N_19483,N_19076);
or U20195 (N_20195,N_18746,N_18230);
nand U20196 (N_20196,N_19499,N_19070);
nand U20197 (N_20197,N_18713,N_19916);
xor U20198 (N_20198,N_18566,N_19571);
and U20199 (N_20199,N_18359,N_19745);
and U20200 (N_20200,N_18410,N_19284);
or U20201 (N_20201,N_18910,N_19341);
xor U20202 (N_20202,N_19270,N_19438);
and U20203 (N_20203,N_18869,N_18643);
nor U20204 (N_20204,N_18724,N_18785);
nand U20205 (N_20205,N_18669,N_19858);
or U20206 (N_20206,N_18090,N_18412);
xnor U20207 (N_20207,N_18318,N_18362);
nand U20208 (N_20208,N_18623,N_19603);
nand U20209 (N_20209,N_19085,N_19487);
or U20210 (N_20210,N_18695,N_19247);
and U20211 (N_20211,N_18946,N_19407);
nor U20212 (N_20212,N_19605,N_19983);
and U20213 (N_20213,N_18650,N_19031);
nand U20214 (N_20214,N_19604,N_19307);
nand U20215 (N_20215,N_18882,N_18108);
nor U20216 (N_20216,N_19911,N_19035);
nor U20217 (N_20217,N_19303,N_18035);
nor U20218 (N_20218,N_19523,N_19936);
nand U20219 (N_20219,N_19243,N_19668);
or U20220 (N_20220,N_18712,N_18126);
nand U20221 (N_20221,N_18640,N_19041);
nor U20222 (N_20222,N_19746,N_18533);
or U20223 (N_20223,N_18645,N_18700);
and U20224 (N_20224,N_18335,N_19213);
nor U20225 (N_20225,N_19221,N_18368);
nand U20226 (N_20226,N_19371,N_19739);
xor U20227 (N_20227,N_18828,N_18544);
nor U20228 (N_20228,N_19091,N_18480);
nand U20229 (N_20229,N_19698,N_19633);
nand U20230 (N_20230,N_18630,N_18549);
xnor U20231 (N_20231,N_19374,N_19448);
and U20232 (N_20232,N_19796,N_19950);
xnor U20233 (N_20233,N_18250,N_19721);
and U20234 (N_20234,N_18300,N_18967);
and U20235 (N_20235,N_19412,N_18689);
nor U20236 (N_20236,N_19834,N_18491);
or U20237 (N_20237,N_18164,N_19675);
and U20238 (N_20238,N_18052,N_19029);
or U20239 (N_20239,N_19462,N_18865);
and U20240 (N_20240,N_19071,N_18826);
xor U20241 (N_20241,N_18873,N_18990);
nor U20242 (N_20242,N_19521,N_19912);
xnor U20243 (N_20243,N_18408,N_18275);
xnor U20244 (N_20244,N_19551,N_18583);
nor U20245 (N_20245,N_19657,N_19838);
or U20246 (N_20246,N_19861,N_18319);
or U20247 (N_20247,N_18529,N_19854);
nand U20248 (N_20248,N_18442,N_18200);
xor U20249 (N_20249,N_18058,N_19951);
or U20250 (N_20250,N_19585,N_18536);
nor U20251 (N_20251,N_18042,N_18666);
nor U20252 (N_20252,N_19962,N_18320);
and U20253 (N_20253,N_19360,N_19626);
nand U20254 (N_20254,N_19461,N_19227);
xnor U20255 (N_20255,N_19937,N_18601);
or U20256 (N_20256,N_19094,N_19764);
xor U20257 (N_20257,N_18883,N_18487);
nand U20258 (N_20258,N_19628,N_19106);
and U20259 (N_20259,N_19321,N_18343);
xnor U20260 (N_20260,N_18684,N_18187);
nand U20261 (N_20261,N_19803,N_19545);
or U20262 (N_20262,N_19592,N_18661);
and U20263 (N_20263,N_19982,N_19547);
nand U20264 (N_20264,N_18754,N_19268);
nor U20265 (N_20265,N_19023,N_18626);
nand U20266 (N_20266,N_19369,N_19105);
and U20267 (N_20267,N_19794,N_19229);
nor U20268 (N_20268,N_18165,N_19567);
or U20269 (N_20269,N_18539,N_19114);
and U20270 (N_20270,N_19154,N_19874);
nor U20271 (N_20271,N_19295,N_18556);
xnor U20272 (N_20272,N_19968,N_18149);
nand U20273 (N_20273,N_19599,N_19365);
or U20274 (N_20274,N_19839,N_18722);
and U20275 (N_20275,N_18298,N_19034);
and U20276 (N_20276,N_18559,N_19281);
and U20277 (N_20277,N_19948,N_18905);
nor U20278 (N_20278,N_19703,N_18890);
or U20279 (N_20279,N_19143,N_19492);
nand U20280 (N_20280,N_19329,N_18273);
xor U20281 (N_20281,N_18019,N_18632);
nand U20282 (N_20282,N_19829,N_19686);
nand U20283 (N_20283,N_19918,N_19061);
or U20284 (N_20284,N_19827,N_19347);
nor U20285 (N_20285,N_18739,N_18171);
or U20286 (N_20286,N_19751,N_19920);
and U20287 (N_20287,N_19277,N_18488);
and U20288 (N_20288,N_19674,N_19340);
and U20289 (N_20289,N_18756,N_19323);
nand U20290 (N_20290,N_18657,N_19783);
and U20291 (N_20291,N_18952,N_19124);
and U20292 (N_20292,N_19137,N_18705);
nor U20293 (N_20293,N_19852,N_18425);
or U20294 (N_20294,N_19484,N_18027);
and U20295 (N_20295,N_19647,N_19196);
nor U20296 (N_20296,N_18796,N_19345);
nor U20297 (N_20297,N_18146,N_18411);
or U20298 (N_20298,N_19102,N_19546);
xnor U20299 (N_20299,N_19509,N_18268);
nand U20300 (N_20300,N_18112,N_18166);
and U20301 (N_20301,N_18940,N_18367);
or U20302 (N_20302,N_18293,N_18043);
nand U20303 (N_20303,N_19127,N_18501);
nor U20304 (N_20304,N_18092,N_18351);
nor U20305 (N_20305,N_18409,N_19187);
xor U20306 (N_20306,N_19389,N_18117);
xor U20307 (N_20307,N_18919,N_18711);
nand U20308 (N_20308,N_19866,N_19179);
xnor U20309 (N_20309,N_18432,N_18622);
nor U20310 (N_20310,N_19282,N_19973);
xnor U20311 (N_20311,N_18132,N_18194);
or U20312 (N_20312,N_19468,N_19969);
and U20313 (N_20313,N_19735,N_18765);
and U20314 (N_20314,N_18589,N_19877);
nand U20315 (N_20315,N_18399,N_18269);
nand U20316 (N_20316,N_19274,N_19890);
and U20317 (N_20317,N_18198,N_19704);
xor U20318 (N_20318,N_19678,N_18096);
xor U20319 (N_20319,N_19405,N_19457);
or U20320 (N_20320,N_19715,N_18717);
nor U20321 (N_20321,N_18607,N_19129);
and U20322 (N_20322,N_19145,N_19415);
nand U20323 (N_20323,N_19639,N_19296);
and U20324 (N_20324,N_19447,N_19860);
xor U20325 (N_20325,N_19025,N_19352);
xor U20326 (N_20326,N_19477,N_18789);
xnor U20327 (N_20327,N_18244,N_19812);
or U20328 (N_20328,N_18602,N_18590);
nand U20329 (N_20329,N_19520,N_18340);
and U20330 (N_20330,N_19297,N_19327);
and U20331 (N_20331,N_18920,N_18304);
or U20332 (N_20332,N_18140,N_19190);
nor U20333 (N_20333,N_18124,N_19109);
xor U20334 (N_20334,N_18207,N_19755);
or U20335 (N_20335,N_19370,N_19786);
nor U20336 (N_20336,N_18678,N_18093);
or U20337 (N_20337,N_18864,N_18687);
xnor U20338 (N_20338,N_19522,N_18474);
or U20339 (N_20339,N_18862,N_19188);
or U20340 (N_20340,N_19907,N_19654);
or U20341 (N_20341,N_19426,N_18025);
nor U20342 (N_20342,N_19065,N_18026);
nor U20343 (N_20343,N_18469,N_19108);
nor U20344 (N_20344,N_18757,N_18809);
nor U20345 (N_20345,N_19771,N_19312);
and U20346 (N_20346,N_18729,N_18515);
nor U20347 (N_20347,N_19207,N_18447);
and U20348 (N_20348,N_18677,N_19804);
or U20349 (N_20349,N_18264,N_18021);
nor U20350 (N_20350,N_19578,N_19743);
xnor U20351 (N_20351,N_18899,N_19596);
and U20352 (N_20352,N_18720,N_19182);
or U20353 (N_20353,N_18569,N_18113);
xor U20354 (N_20354,N_19623,N_18353);
or U20355 (N_20355,N_19146,N_19806);
and U20356 (N_20356,N_18926,N_19326);
nand U20357 (N_20357,N_18068,N_19929);
or U20358 (N_20358,N_18932,N_18324);
and U20359 (N_20359,N_18339,N_19769);
xor U20360 (N_20360,N_18933,N_18427);
or U20361 (N_20361,N_19254,N_18219);
xor U20362 (N_20362,N_19090,N_18822);
nand U20363 (N_20363,N_18629,N_18031);
and U20364 (N_20364,N_18389,N_18050);
nor U20365 (N_20365,N_18803,N_18778);
or U20366 (N_20366,N_19644,N_19372);
nor U20367 (N_20367,N_18769,N_19342);
and U20368 (N_20368,N_18385,N_18101);
nor U20369 (N_20369,N_18552,N_18592);
or U20370 (N_20370,N_19481,N_18783);
xor U20371 (N_20371,N_19766,N_19009);
nand U20372 (N_20372,N_19115,N_18581);
nor U20373 (N_20373,N_18072,N_19077);
and U20374 (N_20374,N_18332,N_18055);
or U20375 (N_20375,N_18842,N_18139);
nor U20376 (N_20376,N_19452,N_19662);
nor U20377 (N_20377,N_19767,N_19162);
nor U20378 (N_20378,N_19891,N_19563);
xor U20379 (N_20379,N_18685,N_18605);
nand U20380 (N_20380,N_18274,N_19286);
xor U20381 (N_20381,N_19663,N_19423);
xor U20382 (N_20382,N_18099,N_19512);
nand U20383 (N_20383,N_18541,N_18018);
nor U20384 (N_20384,N_18400,N_18968);
and U20385 (N_20385,N_18161,N_19135);
and U20386 (N_20386,N_19044,N_19097);
nor U20387 (N_20387,N_18431,N_19757);
or U20388 (N_20388,N_18356,N_18464);
or U20389 (N_20389,N_18401,N_18449);
nor U20390 (N_20390,N_18780,N_18852);
nand U20391 (N_20391,N_19733,N_18642);
nand U20392 (N_20392,N_18471,N_19359);
nor U20393 (N_20393,N_19434,N_19401);
and U20394 (N_20394,N_18191,N_19294);
nand U20395 (N_20395,N_18020,N_19573);
nand U20396 (N_20396,N_18925,N_18475);
nand U20397 (N_20397,N_18192,N_18426);
nand U20398 (N_20398,N_18964,N_18531);
nand U20399 (N_20399,N_18949,N_18584);
or U20400 (N_20400,N_18070,N_19595);
or U20401 (N_20401,N_19174,N_19089);
or U20402 (N_20402,N_19446,N_18554);
and U20403 (N_20403,N_19337,N_19054);
nand U20404 (N_20404,N_19387,N_19781);
nor U20405 (N_20405,N_18565,N_19258);
or U20406 (N_20406,N_18836,N_18818);
and U20407 (N_20407,N_18246,N_19965);
or U20408 (N_20408,N_18378,N_18532);
or U20409 (N_20409,N_19851,N_18430);
nand U20410 (N_20410,N_18580,N_18781);
or U20411 (N_20411,N_18519,N_19798);
or U20412 (N_20412,N_19471,N_18036);
nand U20413 (N_20413,N_18310,N_19238);
nor U20414 (N_20414,N_19032,N_19515);
xor U20415 (N_20415,N_18002,N_18428);
nand U20416 (N_20416,N_18621,N_18732);
xnor U20417 (N_20417,N_18418,N_19598);
and U20418 (N_20418,N_18199,N_18454);
or U20419 (N_20419,N_18077,N_19328);
nor U20420 (N_20420,N_18545,N_18252);
nor U20421 (N_20421,N_19516,N_18792);
nor U20422 (N_20422,N_19175,N_19104);
and U20423 (N_20423,N_18692,N_18327);
xor U20424 (N_20424,N_19607,N_19153);
xor U20425 (N_20425,N_18201,N_19699);
nor U20426 (N_20426,N_18750,N_19538);
or U20427 (N_20427,N_19430,N_18799);
nor U20428 (N_20428,N_18227,N_19753);
xor U20429 (N_20429,N_19433,N_18423);
nand U20430 (N_20430,N_18524,N_19824);
and U20431 (N_20431,N_18087,N_19894);
and U20432 (N_20432,N_19688,N_19192);
nor U20433 (N_20433,N_18942,N_19206);
nor U20434 (N_20434,N_19718,N_18505);
and U20435 (N_20435,N_19330,N_19579);
nor U20436 (N_20436,N_18955,N_18326);
nor U20437 (N_20437,N_19493,N_19963);
xnor U20438 (N_20438,N_19385,N_18228);
nand U20439 (N_20439,N_18179,N_18900);
or U20440 (N_20440,N_19810,N_18506);
and U20441 (N_20441,N_19404,N_19532);
xor U20442 (N_20442,N_18261,N_19535);
xnor U20443 (N_20443,N_18450,N_18213);
nor U20444 (N_20444,N_19475,N_19410);
nand U20445 (N_20445,N_18725,N_18877);
xnor U20446 (N_20446,N_18694,N_18402);
and U20447 (N_20447,N_19952,N_19807);
xnor U20448 (N_20448,N_19792,N_18177);
and U20449 (N_20449,N_19141,N_18175);
nand U20450 (N_20450,N_18793,N_18127);
nand U20451 (N_20451,N_19587,N_18763);
xor U20452 (N_20452,N_19036,N_19418);
nor U20453 (N_20453,N_19325,N_18133);
and U20454 (N_20454,N_18325,N_18163);
xnor U20455 (N_20455,N_19793,N_19597);
or U20456 (N_20456,N_19830,N_19478);
nor U20457 (N_20457,N_19865,N_18948);
nand U20458 (N_20458,N_19550,N_19437);
and U20459 (N_20459,N_19068,N_18413);
or U20460 (N_20460,N_19903,N_18638);
xnor U20461 (N_20461,N_18985,N_18184);
or U20462 (N_20462,N_18587,N_19988);
and U20463 (N_20463,N_19445,N_18599);
or U20464 (N_20464,N_18652,N_18114);
nor U20465 (N_20465,N_19777,N_19226);
or U20466 (N_20466,N_19975,N_18217);
xor U20467 (N_20467,N_19901,N_19120);
xor U20468 (N_20468,N_18710,N_19682);
and U20469 (N_20469,N_18243,N_18701);
nor U20470 (N_20470,N_19696,N_19165);
or U20471 (N_20471,N_18484,N_19987);
nor U20472 (N_20472,N_19653,N_19078);
and U20473 (N_20473,N_19313,N_19038);
xor U20474 (N_20474,N_18616,N_19033);
nor U20475 (N_20475,N_18723,N_19186);
nand U20476 (N_20476,N_18680,N_18074);
nor U20477 (N_20477,N_19250,N_18263);
nor U20478 (N_20478,N_19636,N_18188);
and U20479 (N_20479,N_18936,N_18169);
and U20480 (N_20480,N_18593,N_18557);
nand U20481 (N_20481,N_19529,N_18041);
nor U20482 (N_20482,N_19847,N_19716);
xnor U20483 (N_20483,N_18456,N_19170);
nor U20484 (N_20484,N_19350,N_18182);
nand U20485 (N_20485,N_19508,N_18500);
xnor U20486 (N_20486,N_18636,N_18371);
nor U20487 (N_20487,N_18151,N_19621);
and U20488 (N_20488,N_18595,N_19261);
xor U20489 (N_20489,N_18336,N_19930);
and U20490 (N_20490,N_18688,N_18473);
or U20491 (N_20491,N_18510,N_19466);
nand U20492 (N_20492,N_18067,N_18066);
nand U20493 (N_20493,N_19533,N_18386);
or U20494 (N_20494,N_19230,N_18137);
or U20495 (N_20495,N_19004,N_18311);
nor U20496 (N_20496,N_18821,N_18328);
nor U20497 (N_20497,N_18322,N_18730);
nand U20498 (N_20498,N_19463,N_19406);
nand U20499 (N_20499,N_19220,N_18168);
and U20500 (N_20500,N_18435,N_18131);
or U20501 (N_20501,N_18817,N_19299);
nor U20502 (N_20502,N_18697,N_18664);
xor U20503 (N_20503,N_18445,N_19518);
or U20504 (N_20504,N_18896,N_18308);
and U20505 (N_20505,N_18214,N_18384);
nor U20506 (N_20506,N_19302,N_18158);
and U20507 (N_20507,N_18639,N_18075);
nand U20508 (N_20508,N_19677,N_19782);
nand U20509 (N_20509,N_19158,N_18125);
or U20510 (N_20510,N_18996,N_18906);
xnor U20511 (N_20511,N_19204,N_19173);
nor U20512 (N_20512,N_18060,N_19191);
and U20513 (N_20513,N_19687,N_18794);
or U20514 (N_20514,N_19027,N_18223);
nor U20515 (N_20515,N_19658,N_19208);
and U20516 (N_20516,N_18254,N_18844);
xor U20517 (N_20517,N_18608,N_18220);
and U20518 (N_20518,N_19400,N_18790);
and U20519 (N_20519,N_19393,N_19641);
nand U20520 (N_20520,N_19235,N_19734);
or U20521 (N_20521,N_18759,N_18610);
nor U20522 (N_20522,N_18884,N_19464);
and U20523 (N_20523,N_18693,N_18951);
nor U20524 (N_20524,N_18935,N_18577);
and U20525 (N_20525,N_18558,N_19744);
nand U20526 (N_20526,N_19333,N_19849);
nor U20527 (N_20527,N_19577,N_19432);
nor U20528 (N_20528,N_18800,N_19954);
xnor U20529 (N_20529,N_18037,N_19123);
or U20530 (N_20530,N_18895,N_19961);
xnor U20531 (N_20531,N_18993,N_18160);
nor U20532 (N_20532,N_18627,N_19482);
xnor U20533 (N_20533,N_19283,N_19528);
xor U20534 (N_20534,N_19775,N_18820);
nand U20535 (N_20535,N_18743,N_19981);
and U20536 (N_20536,N_18672,N_18811);
nand U20537 (N_20537,N_19809,N_19811);
nor U20538 (N_20538,N_19857,N_19288);
and U20539 (N_20539,N_19850,N_18259);
or U20540 (N_20540,N_19712,N_19897);
and U20541 (N_20541,N_18784,N_18604);
and U20542 (N_20542,N_18433,N_18773);
or U20543 (N_20543,N_19867,N_18676);
or U20544 (N_20544,N_18395,N_18788);
xor U20545 (N_20545,N_19560,N_18088);
xor U20546 (N_20546,N_18742,N_19656);
or U20547 (N_20547,N_18634,N_19197);
nor U20548 (N_20548,N_18138,N_18834);
nor U20549 (N_20549,N_18056,N_19841);
nand U20550 (N_20550,N_19202,N_19486);
and U20551 (N_20551,N_18309,N_18465);
or U20552 (N_20552,N_19480,N_18655);
nand U20553 (N_20553,N_18316,N_18249);
nand U20554 (N_20554,N_18514,N_19148);
or U20555 (N_20555,N_18658,N_19256);
xor U20556 (N_20556,N_19242,N_18089);
and U20557 (N_20557,N_19772,N_18804);
or U20558 (N_20558,N_19667,N_18406);
and U20559 (N_20559,N_18073,N_19736);
or U20560 (N_20560,N_19872,N_18902);
nand U20561 (N_20561,N_18017,N_19902);
xnor U20562 (N_20562,N_18383,N_18363);
or U20563 (N_20563,N_19357,N_18904);
or U20564 (N_20564,N_18618,N_18596);
and U20565 (N_20565,N_18120,N_19949);
nand U20566 (N_20566,N_18812,N_19210);
xor U20567 (N_20567,N_18856,N_19099);
xor U20568 (N_20568,N_19671,N_19172);
nor U20569 (N_20569,N_18659,N_18446);
and U20570 (N_20570,N_19875,N_19756);
xor U20571 (N_20571,N_18045,N_18189);
nor U20572 (N_20572,N_18962,N_18195);
xnor U20573 (N_20573,N_19386,N_19217);
nand U20574 (N_20574,N_19133,N_18758);
xnor U20575 (N_20575,N_18334,N_19132);
xor U20576 (N_20576,N_19494,N_18997);
and U20577 (N_20577,N_18704,N_19828);
xor U20578 (N_20578,N_18361,N_18816);
and U20579 (N_20579,N_18210,N_19768);
and U20580 (N_20580,N_19497,N_19893);
nor U20581 (N_20581,N_18663,N_19642);
nor U20582 (N_20582,N_19548,N_19046);
xor U20583 (N_20583,N_19672,N_18838);
nand U20584 (N_20584,N_19634,N_18156);
xnor U20585 (N_20585,N_19527,N_18624);
xor U20586 (N_20586,N_18040,N_19900);
xor U20587 (N_20587,N_19167,N_18289);
or U20588 (N_20588,N_19496,N_18301);
nor U20589 (N_20589,N_19422,N_19429);
xor U20590 (N_20590,N_18668,N_18231);
nand U20591 (N_20591,N_18355,N_18466);
xor U20592 (N_20592,N_19351,N_18038);
and U20593 (N_20593,N_18315,N_19996);
or U20594 (N_20594,N_18600,N_18548);
nor U20595 (N_20595,N_18918,N_19966);
and U20596 (N_20596,N_19022,N_19540);
nor U20597 (N_20597,N_19377,N_19100);
and U20598 (N_20598,N_18963,N_18251);
xor U20599 (N_20599,N_19084,N_18512);
nand U20600 (N_20600,N_18499,N_18924);
xnor U20601 (N_20601,N_19402,N_19562);
xnor U20602 (N_20602,N_18914,N_19366);
or U20603 (N_20603,N_18233,N_19876);
xor U20604 (N_20604,N_18609,N_18404);
nand U20605 (N_20605,N_18523,N_19232);
and U20606 (N_20606,N_18771,N_18294);
nand U20607 (N_20607,N_19278,N_18588);
and U20608 (N_20608,N_18155,N_19610);
nand U20609 (N_20609,N_18129,N_19638);
xnor U20610 (N_20610,N_19368,N_19064);
nor U20611 (N_20611,N_19110,N_18185);
xor U20612 (N_20612,N_18572,N_18513);
nand U20613 (N_20613,N_19380,N_18502);
xnor U20614 (N_20614,N_18303,N_18482);
or U20615 (N_20615,N_18881,N_19842);
or U20616 (N_20616,N_18009,N_18727);
nor U20617 (N_20617,N_18453,N_18313);
or U20618 (N_20618,N_18944,N_19364);
xnor U20619 (N_20619,N_19684,N_19750);
or U20620 (N_20620,N_18797,N_19171);
nand U20621 (N_20621,N_18917,N_19939);
or U20622 (N_20622,N_19524,N_19262);
nand U20623 (N_20623,N_18024,N_19469);
and U20624 (N_20624,N_18039,N_19835);
nor U20625 (N_20625,N_19082,N_18257);
or U20626 (N_20626,N_19637,N_18180);
and U20627 (N_20627,N_18903,N_19264);
and U20628 (N_20628,N_18392,N_18876);
xor U20629 (N_20629,N_19506,N_19053);
and U20630 (N_20630,N_18119,N_19514);
xor U20631 (N_20631,N_19239,N_19219);
xor U20632 (N_20632,N_19976,N_18393);
or U20633 (N_20633,N_18916,N_18135);
nand U20634 (N_20634,N_18521,N_18270);
nor U20635 (N_20635,N_19519,N_18455);
or U20636 (N_20636,N_18414,N_19320);
and U20637 (N_20637,N_18437,N_18415);
nand U20638 (N_20638,N_18049,N_19788);
nand U20639 (N_20639,N_18665,N_18733);
and U20640 (N_20640,N_18443,N_19730);
xnor U20641 (N_20641,N_18183,N_19228);
or U20642 (N_20642,N_19898,N_18329);
nand U20643 (N_20643,N_18010,N_19617);
nor U20644 (N_20644,N_18461,N_19971);
xor U20645 (N_20645,N_19705,N_19600);
nor U20646 (N_20646,N_18462,N_18943);
xor U20647 (N_20647,N_18776,N_18102);
nand U20648 (N_20648,N_19474,N_18612);
and U20649 (N_20649,N_18398,N_18777);
and U20650 (N_20650,N_19343,N_19310);
nor U20651 (N_20651,N_18128,N_18973);
and U20652 (N_20652,N_18063,N_18660);
nand U20653 (N_20653,N_18065,N_18885);
nor U20654 (N_20654,N_19074,N_19758);
or U20655 (N_20655,N_19444,N_18306);
and U20656 (N_20656,N_19436,N_18868);
and U20657 (N_20657,N_18008,N_19348);
or U20658 (N_20658,N_18613,N_19941);
or U20659 (N_20659,N_19576,N_19553);
nand U20660 (N_20660,N_18795,N_19218);
nor U20661 (N_20661,N_18915,N_18396);
xnor U20662 (N_20662,N_19517,N_18737);
nand U20663 (N_20663,N_19304,N_19695);
nand U20664 (N_20664,N_19056,N_18974);
xnor U20665 (N_20665,N_18071,N_18203);
or U20666 (N_20666,N_19870,N_18085);
xor U20667 (N_20667,N_18848,N_19666);
xnor U20668 (N_20668,N_18671,N_19449);
and U20669 (N_20669,N_18706,N_19502);
nand U20670 (N_20670,N_18563,N_18476);
nor U20671 (N_20671,N_19507,N_19871);
xnor U20672 (N_20672,N_18551,N_19417);
xnor U20673 (N_20673,N_18798,N_19591);
nor U20674 (N_20674,N_19346,N_19584);
or U20675 (N_20675,N_19467,N_19837);
or U20676 (N_20676,N_19566,N_19151);
or U20677 (N_20677,N_18202,N_19862);
and U20678 (N_20678,N_18805,N_18929);
nand U20679 (N_20679,N_18947,N_18215);
nand U20680 (N_20680,N_18631,N_18238);
nor U20681 (N_20681,N_18808,N_18573);
xnor U20682 (N_20682,N_18755,N_18649);
xor U20683 (N_20683,N_18898,N_18598);
nand U20684 (N_20684,N_18762,N_18277);
or U20685 (N_20685,N_18807,N_19680);
nor U20686 (N_20686,N_19316,N_18779);
nor U20687 (N_20687,N_19111,N_18537);
nand U20688 (N_20688,N_18285,N_19000);
and U20689 (N_20689,N_18162,N_18486);
nand U20690 (N_20690,N_19822,N_19673);
and U20691 (N_20691,N_19441,N_18076);
and U20692 (N_20692,N_18702,N_18438);
nor U20693 (N_20693,N_19510,N_18457);
nor U20694 (N_20694,N_19252,N_18448);
nand U20695 (N_20695,N_18147,N_19367);
xor U20696 (N_20696,N_19999,N_19763);
xnor U20697 (N_20697,N_18419,N_19016);
xor U20698 (N_20698,N_18197,N_19873);
or U20699 (N_20699,N_19225,N_19883);
xnor U20700 (N_20700,N_18745,N_19363);
or U20701 (N_20701,N_19265,N_19201);
nor U20702 (N_20702,N_19928,N_19921);
xnor U20703 (N_20703,N_18508,N_18291);
xor U20704 (N_20704,N_19572,N_19917);
or U20705 (N_20705,N_18097,N_18597);
or U20706 (N_20706,N_18375,N_18170);
nor U20707 (N_20707,N_19081,N_18258);
xnor U20708 (N_20708,N_18255,N_19470);
xor U20709 (N_20709,N_19062,N_19544);
or U20710 (N_20710,N_19269,N_18046);
xor U20711 (N_20711,N_19855,N_19910);
xor U20712 (N_20712,N_19152,N_18979);
or U20713 (N_20713,N_18094,N_19679);
nand U20714 (N_20714,N_18625,N_18791);
nand U20715 (N_20715,N_19790,N_19608);
nand U20716 (N_20716,N_18683,N_18982);
nand U20717 (N_20717,N_19040,N_19189);
nand U20718 (N_20718,N_19706,N_18594);
nor U20719 (N_20719,N_18679,N_19012);
nor U20720 (N_20720,N_18840,N_19028);
and U20721 (N_20721,N_19101,N_18287);
xor U20722 (N_20722,N_19125,N_18478);
nor U20723 (N_20723,N_18959,N_19761);
nand U20724 (N_20724,N_19534,N_19722);
xnor U20725 (N_20725,N_18266,N_18945);
xor U20726 (N_20726,N_18574,N_19319);
xor U20727 (N_20727,N_19495,N_18738);
nor U20728 (N_20728,N_18387,N_19537);
xnor U20729 (N_20729,N_18989,N_18892);
and U20730 (N_20730,N_18479,N_18976);
nor U20731 (N_20731,N_19942,N_18292);
nand U20732 (N_20732,N_18575,N_19465);
nor U20733 (N_20733,N_18123,N_19787);
xor U20734 (N_20734,N_19800,N_19935);
nor U20735 (N_20735,N_19833,N_19892);
or U20736 (N_20736,N_19072,N_19130);
nand U20737 (N_20737,N_19726,N_19974);
and U20738 (N_20738,N_19947,N_18346);
and U20739 (N_20739,N_18248,N_19315);
xnor U20740 (N_20740,N_18416,N_19398);
nand U20741 (N_20741,N_18670,N_18110);
xnor U20742 (N_20742,N_18878,N_19702);
nor U20743 (N_20743,N_18434,N_19049);
nor U20744 (N_20744,N_18118,N_19992);
nor U20745 (N_20745,N_19932,N_18726);
xor U20746 (N_20746,N_18960,N_19802);
nand U20747 (N_20747,N_18728,N_19301);
or U20748 (N_20748,N_19997,N_18307);
nand U20749 (N_20749,N_18157,N_19558);
xor U20750 (N_20750,N_19554,N_19779);
and U20751 (N_20751,N_18740,N_18561);
xor U20752 (N_20752,N_18774,N_19440);
xnor U20753 (N_20753,N_18350,N_19194);
or U20754 (N_20754,N_18209,N_18586);
or U20755 (N_20755,N_18084,N_18829);
nor U20756 (N_20756,N_19149,N_19249);
nand U20757 (N_20757,N_19564,N_19632);
and U20758 (N_20758,N_18801,N_19339);
nand U20759 (N_20759,N_19007,N_18208);
xor U20760 (N_20760,N_19655,N_19700);
or U20761 (N_20761,N_18212,N_19817);
nand U20762 (N_20762,N_18330,N_19362);
nand U20763 (N_20763,N_19222,N_19831);
nand U20764 (N_20764,N_19244,N_19118);
or U20765 (N_20765,N_18141,N_19720);
nand U20766 (N_20766,N_19080,N_19358);
and U20767 (N_20767,N_19690,N_19045);
nor U20768 (N_20768,N_19570,N_18992);
and U20769 (N_20769,N_19795,N_18567);
nor U20770 (N_20770,N_18543,N_19711);
nand U20771 (N_20771,N_19155,N_18691);
and U20772 (N_20772,N_18234,N_19373);
nand U20773 (N_20773,N_19018,N_18262);
or U20774 (N_20774,N_19940,N_19416);
or U20775 (N_20775,N_18390,N_18850);
and U20776 (N_20776,N_18768,N_18407);
xnor U20777 (N_20777,N_19846,N_19138);
xnor U20778 (N_20778,N_19075,N_18662);
or U20779 (N_20779,N_18369,N_19543);
nand U20780 (N_20780,N_19993,N_18719);
and U20781 (N_20781,N_18079,N_19557);
nor U20782 (N_20782,N_18104,N_18606);
xnor U20783 (N_20783,N_19245,N_18518);
nand U20784 (N_20784,N_18014,N_19126);
nor U20785 (N_20785,N_18635,N_18337);
or U20786 (N_20786,N_18709,N_19501);
or U20787 (N_20787,N_18527,N_18016);
xor U20788 (N_20788,N_19272,N_19594);
xnor U20789 (N_20789,N_19273,N_19216);
nand U20790 (N_20790,N_18535,N_18086);
or U20791 (N_20791,N_19391,N_19931);
and U20792 (N_20792,N_19995,N_18839);
nor U20793 (N_20793,N_18830,N_18880);
xor U20794 (N_20794,N_19887,N_19994);
xor U20795 (N_20795,N_18507,N_19240);
and U20796 (N_20796,N_18054,N_18981);
and U20797 (N_20797,N_19408,N_19819);
xnor U20798 (N_20798,N_18373,N_19160);
nor U20799 (N_20799,N_18734,N_18528);
nor U20800 (N_20800,N_19665,N_19630);
and U20801 (N_20801,N_19324,N_18142);
nand U20802 (N_20802,N_18172,N_19455);
xnor U20803 (N_20803,N_19019,N_18468);
nand U20804 (N_20804,N_18394,N_18891);
or U20805 (N_20805,N_18853,N_19180);
nand U20806 (N_20806,N_18436,N_18364);
nand U20807 (N_20807,N_19253,N_18028);
nor U20808 (N_20808,N_19505,N_19421);
xor U20809 (N_20809,N_19460,N_19168);
nor U20810 (N_20810,N_19498,N_19602);
xnor U20811 (N_20811,N_18245,N_19864);
or U20812 (N_20812,N_19058,N_19714);
and U20813 (N_20813,N_19629,N_19719);
or U20814 (N_20814,N_19279,N_19741);
or U20815 (N_20815,N_18922,N_19305);
nand U20816 (N_20816,N_18190,N_19395);
nand U20817 (N_20817,N_19063,N_19648);
and U20818 (N_20818,N_19832,N_19879);
xnor U20819 (N_20819,N_18100,N_19776);
xnor U20820 (N_20820,N_19878,N_19957);
or U20821 (N_20821,N_19425,N_18530);
xor U20822 (N_20822,N_18912,N_18483);
and U20823 (N_20823,N_18391,N_18837);
xnor U20824 (N_20824,N_19650,N_19396);
or U20825 (N_20825,N_18295,N_18961);
nand U20826 (N_20826,N_19043,N_19150);
nand U20827 (N_20827,N_19814,N_19117);
and U20828 (N_20828,N_19098,N_18280);
xor U20829 (N_20829,N_18023,N_18004);
nand U20830 (N_20830,N_18366,N_19748);
or U20831 (N_20831,N_19914,N_18956);
nand U20832 (N_20832,N_19899,N_19413);
nor U20833 (N_20833,N_19356,N_19156);
or U20834 (N_20834,N_18721,N_18620);
xor U20835 (N_20835,N_18136,N_18823);
nor U20836 (N_20836,N_18894,N_19073);
xor U20837 (N_20837,N_19868,N_19915);
or U20838 (N_20838,N_19616,N_19361);
or U20839 (N_20839,N_18216,N_18143);
and U20840 (N_20840,N_18975,N_18578);
nor U20841 (N_20841,N_18485,N_19224);
nor U20842 (N_20842,N_18186,N_18122);
nand U20843 (N_20843,N_18641,N_18927);
or U20844 (N_20844,N_19131,N_19869);
nand U20845 (N_20845,N_18941,N_19922);
xnor U20846 (N_20846,N_19765,N_19959);
or U20847 (N_20847,N_19752,N_19176);
nand U20848 (N_20848,N_18686,N_18957);
nand U20849 (N_20849,N_19379,N_18867);
nand U20850 (N_20850,N_19048,N_18115);
nor U20851 (N_20851,N_19773,N_19008);
or U20852 (N_20852,N_19275,N_18716);
and U20853 (N_20853,N_18105,N_19881);
and U20854 (N_20854,N_19980,N_18481);
xor U20855 (N_20855,N_18874,N_19945);
nand U20856 (N_20856,N_18284,N_19163);
and U20857 (N_20857,N_18950,N_19083);
or U20858 (N_20858,N_18591,N_19643);
and U20859 (N_20859,N_18493,N_18154);
and U20860 (N_20860,N_18271,N_19298);
nand U20861 (N_20861,N_18819,N_19985);
nand U20862 (N_20862,N_19805,N_19317);
nand U20863 (N_20863,N_19205,N_18272);
nor U20864 (N_20864,N_18205,N_19456);
nor U20865 (N_20865,N_19789,N_19355);
nand U20866 (N_20866,N_19067,N_19906);
and U20867 (N_20867,N_18698,N_18226);
nand U20868 (N_20868,N_19694,N_18420);
nand U20869 (N_20869,N_19770,N_19403);
and U20870 (N_20870,N_18889,N_19276);
nand U20871 (N_20871,N_18297,N_18439);
or U20872 (N_20872,N_18218,N_18938);
xor U20873 (N_20873,N_18735,N_18224);
and U20874 (N_20874,N_19606,N_18490);
nor U20875 (N_20875,N_18053,N_18048);
xor U20876 (N_20876,N_19676,N_19958);
xor U20877 (N_20877,N_19200,N_19525);
nor U20878 (N_20878,N_19991,N_18977);
nor U20879 (N_20879,N_18012,N_18787);
xor U20880 (N_20880,N_18999,N_18806);
and U20881 (N_20881,N_18279,N_18225);
xor U20882 (N_20882,N_18761,N_18458);
nand U20883 (N_20883,N_19384,N_18345);
or U20884 (N_20884,N_19164,N_18388);
or U20885 (N_20885,N_19503,N_19904);
or U20886 (N_20886,N_18753,N_18542);
xor U20887 (N_20887,N_18953,N_18546);
nand U20888 (N_20888,N_19611,N_19541);
and U20889 (N_20889,N_19836,N_19710);
nor U20890 (N_20890,N_19889,N_19840);
nand U20891 (N_20891,N_19944,N_18370);
nand U20892 (N_20892,N_18000,N_18278);
and U20893 (N_20893,N_19271,N_19198);
or U20894 (N_20894,N_18516,N_19473);
xor U20895 (N_20895,N_19927,N_19002);
nor U20896 (N_20896,N_18854,N_19233);
xnor U20897 (N_20897,N_19314,N_19651);
and U20898 (N_20898,N_19749,N_19203);
nor U20899 (N_20899,N_19096,N_18846);
nand U20900 (N_20900,N_18847,N_19443);
xnor U20901 (N_20901,N_19821,N_19526);
or U20902 (N_20902,N_19006,N_18296);
nor U20903 (N_20903,N_19052,N_18571);
and U20904 (N_20904,N_19026,N_19050);
nand U20905 (N_20905,N_19808,N_18477);
xnor U20906 (N_20906,N_19707,N_19967);
and U20907 (N_20907,N_19615,N_18646);
xor U20908 (N_20908,N_19635,N_19737);
xor U20909 (N_20909,N_18832,N_18489);
nor U20910 (N_20910,N_19820,N_19420);
xnor U20911 (N_20911,N_19619,N_18538);
nand U20912 (N_20912,N_18939,N_19559);
and U20913 (N_20913,N_18872,N_19119);
nand U20914 (N_20914,N_19382,N_18029);
or U20915 (N_20915,N_18526,N_19627);
and U20916 (N_20916,N_19990,N_18503);
nand U20917 (N_20917,N_18377,N_19122);
or U20918 (N_20918,N_18057,N_18511);
and U20919 (N_20919,N_19336,N_19593);
or U20920 (N_20920,N_19664,N_18344);
xnor U20921 (N_20921,N_18206,N_18767);
nor U20922 (N_20922,N_18376,N_18870);
and U20923 (N_20923,N_19424,N_19442);
nor U20924 (N_20924,N_19349,N_19454);
nand U20925 (N_20925,N_18236,N_18145);
or U20926 (N_20926,N_18751,N_19844);
or U20927 (N_20927,N_19799,N_19724);
xnor U20928 (N_20928,N_18824,N_19136);
nand U20929 (N_20929,N_19020,N_18540);
and U20930 (N_20930,N_18357,N_19609);
xnor U20931 (N_20931,N_19956,N_18451);
nor U20932 (N_20932,N_19738,N_18965);
nand U20933 (N_20933,N_19590,N_19290);
or U20934 (N_20934,N_18033,N_18148);
nand U20935 (N_20935,N_19717,N_18863);
nand U20936 (N_20936,N_18911,N_19925);
nand U20937 (N_20937,N_18555,N_18380);
nor U20938 (N_20938,N_18460,N_19729);
or U20939 (N_20939,N_19826,N_18006);
or U20940 (N_20940,N_19588,N_19037);
and U20941 (N_20941,N_18007,N_18833);
nor U20942 (N_20942,N_19066,N_19116);
and U20943 (N_20943,N_18173,N_18656);
nand U20944 (N_20944,N_18969,N_19488);
xnor U20945 (N_20945,N_19184,N_18681);
and U20946 (N_20946,N_18098,N_19689);
or U20947 (N_20947,N_18966,N_18382);
and U20948 (N_20948,N_18424,N_18913);
nor U20949 (N_20949,N_18467,N_19964);
nand U20950 (N_20950,N_18871,N_18314);
and U20951 (N_20951,N_18348,N_19614);
or U20952 (N_20952,N_19569,N_19978);
nand U20953 (N_20953,N_18696,N_18653);
xor U20954 (N_20954,N_19926,N_18879);
or U20955 (N_20955,N_18984,N_18349);
nor U20956 (N_20956,N_18153,N_19381);
xor U20957 (N_20957,N_19251,N_18290);
nand U20958 (N_20958,N_18970,N_19646);
nand U20959 (N_20959,N_18855,N_18907);
and U20960 (N_20960,N_18654,N_18667);
nand U20961 (N_20961,N_19128,N_18374);
and U20962 (N_20962,N_19582,N_18360);
and U20963 (N_20963,N_19139,N_19147);
or U20964 (N_20964,N_18849,N_18034);
nand U20965 (N_20965,N_18381,N_19300);
or U20966 (N_20966,N_18980,N_18972);
xor U20967 (N_20967,N_19079,N_18675);
nand U20968 (N_20968,N_18417,N_18403);
nand U20969 (N_20969,N_19536,N_19159);
xor U20970 (N_20970,N_19013,N_19169);
xnor U20971 (N_20971,N_19740,N_19397);
nor U20972 (N_20972,N_18069,N_19234);
nor U20973 (N_20973,N_18152,N_19236);
xnor U20974 (N_20974,N_18030,N_18983);
nor U20975 (N_20975,N_19708,N_19093);
xor U20976 (N_20976,N_18560,N_18741);
and U20977 (N_20977,N_18323,N_19709);
nor U20978 (N_20978,N_19884,N_19731);
or U20979 (N_20979,N_19774,N_18282);
nor U20980 (N_20980,N_19896,N_19624);
xor U20981 (N_20981,N_19195,N_19214);
nor U20982 (N_20982,N_19513,N_19818);
xnor U20983 (N_20983,N_19613,N_19069);
and U20984 (N_20984,N_18579,N_18081);
or U20985 (N_20985,N_19260,N_18930);
nor U20986 (N_20986,N_19479,N_19489);
and U20987 (N_20987,N_19354,N_18159);
or U20988 (N_20988,N_18174,N_19681);
or U20989 (N_20989,N_18167,N_18522);
nor U20990 (N_20990,N_18463,N_18421);
or U20991 (N_20991,N_19583,N_19923);
or U20992 (N_20992,N_18150,N_19549);
nor U20993 (N_20993,N_19661,N_19888);
and U20994 (N_20994,N_18288,N_19157);
nor U20995 (N_20995,N_18312,N_18585);
and U20996 (N_20996,N_19267,N_19215);
and U20997 (N_20997,N_18564,N_19561);
nand U20998 (N_20998,N_18802,N_19816);
xor U20999 (N_20999,N_19257,N_19211);
xnor U21000 (N_21000,N_18712,N_19381);
nand U21001 (N_21001,N_19315,N_18752);
nand U21002 (N_21002,N_18531,N_18097);
or U21003 (N_21003,N_19025,N_18430);
nand U21004 (N_21004,N_18287,N_19203);
or U21005 (N_21005,N_18375,N_18336);
or U21006 (N_21006,N_19889,N_19317);
or U21007 (N_21007,N_19223,N_18588);
nor U21008 (N_21008,N_18798,N_19250);
or U21009 (N_21009,N_18978,N_18363);
or U21010 (N_21010,N_18494,N_18375);
and U21011 (N_21011,N_19389,N_18827);
nor U21012 (N_21012,N_18485,N_18706);
or U21013 (N_21013,N_19684,N_19103);
nor U21014 (N_21014,N_18077,N_18831);
or U21015 (N_21015,N_19168,N_19090);
xnor U21016 (N_21016,N_19275,N_19403);
and U21017 (N_21017,N_19327,N_19935);
xnor U21018 (N_21018,N_18164,N_19285);
nor U21019 (N_21019,N_18478,N_18239);
xor U21020 (N_21020,N_19486,N_18993);
nand U21021 (N_21021,N_19068,N_18827);
and U21022 (N_21022,N_19821,N_19642);
nor U21023 (N_21023,N_19011,N_18179);
xor U21024 (N_21024,N_19659,N_18490);
or U21025 (N_21025,N_18003,N_18774);
nand U21026 (N_21026,N_19429,N_19341);
and U21027 (N_21027,N_18487,N_18459);
or U21028 (N_21028,N_19878,N_19374);
and U21029 (N_21029,N_19066,N_18012);
and U21030 (N_21030,N_19278,N_18942);
nor U21031 (N_21031,N_18898,N_19806);
xnor U21032 (N_21032,N_18173,N_19513);
xor U21033 (N_21033,N_18034,N_19415);
xnor U21034 (N_21034,N_19993,N_19587);
or U21035 (N_21035,N_18814,N_19272);
xor U21036 (N_21036,N_18233,N_19867);
nor U21037 (N_21037,N_19441,N_19861);
and U21038 (N_21038,N_19771,N_19245);
and U21039 (N_21039,N_19364,N_19840);
nand U21040 (N_21040,N_18965,N_18867);
xnor U21041 (N_21041,N_18398,N_19773);
xnor U21042 (N_21042,N_19552,N_18014);
xnor U21043 (N_21043,N_19936,N_19915);
nor U21044 (N_21044,N_18262,N_19705);
xor U21045 (N_21045,N_19779,N_19627);
xor U21046 (N_21046,N_19425,N_18509);
or U21047 (N_21047,N_19496,N_19838);
nor U21048 (N_21048,N_19075,N_19271);
nand U21049 (N_21049,N_18310,N_18878);
and U21050 (N_21050,N_18537,N_18612);
nand U21051 (N_21051,N_19922,N_19174);
nand U21052 (N_21052,N_19494,N_19098);
or U21053 (N_21053,N_18051,N_19704);
nand U21054 (N_21054,N_18600,N_18324);
or U21055 (N_21055,N_19658,N_19797);
xor U21056 (N_21056,N_18960,N_18145);
and U21057 (N_21057,N_18803,N_18371);
xor U21058 (N_21058,N_18869,N_19360);
or U21059 (N_21059,N_18869,N_18905);
nand U21060 (N_21060,N_18302,N_18911);
and U21061 (N_21061,N_19582,N_18070);
and U21062 (N_21062,N_18261,N_18979);
nand U21063 (N_21063,N_19992,N_19180);
or U21064 (N_21064,N_18944,N_19791);
nor U21065 (N_21065,N_19464,N_18464);
xnor U21066 (N_21066,N_18416,N_18242);
nand U21067 (N_21067,N_18570,N_19700);
and U21068 (N_21068,N_19702,N_19643);
and U21069 (N_21069,N_19590,N_18078);
and U21070 (N_21070,N_19108,N_19755);
or U21071 (N_21071,N_18259,N_19042);
and U21072 (N_21072,N_18293,N_19529);
and U21073 (N_21073,N_18084,N_19390);
nand U21074 (N_21074,N_18779,N_18362);
xnor U21075 (N_21075,N_19743,N_18025);
nand U21076 (N_21076,N_19655,N_18770);
nor U21077 (N_21077,N_19780,N_18041);
or U21078 (N_21078,N_18203,N_18164);
nand U21079 (N_21079,N_19947,N_18646);
xor U21080 (N_21080,N_18636,N_18704);
and U21081 (N_21081,N_19449,N_18287);
nand U21082 (N_21082,N_18296,N_19482);
nor U21083 (N_21083,N_19698,N_19512);
or U21084 (N_21084,N_18806,N_19001);
xnor U21085 (N_21085,N_18079,N_19825);
nand U21086 (N_21086,N_18219,N_19159);
nor U21087 (N_21087,N_18900,N_19088);
nand U21088 (N_21088,N_19107,N_19337);
or U21089 (N_21089,N_19747,N_19945);
nor U21090 (N_21090,N_19705,N_18483);
nand U21091 (N_21091,N_19662,N_19362);
and U21092 (N_21092,N_19582,N_18590);
nand U21093 (N_21093,N_19415,N_19806);
xnor U21094 (N_21094,N_19681,N_18393);
or U21095 (N_21095,N_19451,N_18257);
nor U21096 (N_21096,N_19768,N_18085);
nor U21097 (N_21097,N_19615,N_19690);
xor U21098 (N_21098,N_18878,N_19169);
nand U21099 (N_21099,N_19658,N_19914);
nand U21100 (N_21100,N_19493,N_19152);
and U21101 (N_21101,N_19325,N_19833);
nor U21102 (N_21102,N_18911,N_19952);
xor U21103 (N_21103,N_18034,N_18858);
nor U21104 (N_21104,N_18135,N_19006);
xor U21105 (N_21105,N_18567,N_18524);
nand U21106 (N_21106,N_19045,N_19250);
nor U21107 (N_21107,N_19981,N_19196);
nand U21108 (N_21108,N_19208,N_18661);
and U21109 (N_21109,N_19782,N_18131);
nand U21110 (N_21110,N_18060,N_19588);
xor U21111 (N_21111,N_18061,N_18456);
or U21112 (N_21112,N_18075,N_19883);
xnor U21113 (N_21113,N_18671,N_19415);
and U21114 (N_21114,N_18720,N_19283);
nand U21115 (N_21115,N_18413,N_18426);
nand U21116 (N_21116,N_19653,N_19655);
nor U21117 (N_21117,N_19556,N_18543);
nor U21118 (N_21118,N_18196,N_18681);
nor U21119 (N_21119,N_18401,N_19861);
and U21120 (N_21120,N_19221,N_18083);
or U21121 (N_21121,N_18222,N_18560);
and U21122 (N_21122,N_19128,N_18936);
and U21123 (N_21123,N_18269,N_19270);
nor U21124 (N_21124,N_19506,N_18099);
nand U21125 (N_21125,N_19861,N_19339);
or U21126 (N_21126,N_19046,N_19797);
and U21127 (N_21127,N_19667,N_18648);
xnor U21128 (N_21128,N_19095,N_19900);
and U21129 (N_21129,N_18742,N_19191);
or U21130 (N_21130,N_19563,N_19238);
and U21131 (N_21131,N_19020,N_18463);
or U21132 (N_21132,N_19191,N_19565);
and U21133 (N_21133,N_18525,N_19461);
and U21134 (N_21134,N_19661,N_18392);
nand U21135 (N_21135,N_18870,N_18488);
nand U21136 (N_21136,N_18712,N_19788);
and U21137 (N_21137,N_19244,N_19890);
nand U21138 (N_21138,N_18807,N_18769);
and U21139 (N_21139,N_19058,N_19528);
and U21140 (N_21140,N_18076,N_18908);
or U21141 (N_21141,N_18411,N_18170);
and U21142 (N_21142,N_18258,N_18594);
xnor U21143 (N_21143,N_18897,N_19119);
nand U21144 (N_21144,N_19321,N_18889);
xor U21145 (N_21145,N_19022,N_18984);
nand U21146 (N_21146,N_19371,N_18670);
xnor U21147 (N_21147,N_19997,N_19014);
and U21148 (N_21148,N_18824,N_18126);
nor U21149 (N_21149,N_19877,N_18471);
and U21150 (N_21150,N_19626,N_18075);
or U21151 (N_21151,N_18692,N_19412);
nor U21152 (N_21152,N_18854,N_18641);
and U21153 (N_21153,N_19437,N_19480);
xor U21154 (N_21154,N_19960,N_18143);
or U21155 (N_21155,N_19491,N_18384);
and U21156 (N_21156,N_19478,N_19319);
nor U21157 (N_21157,N_19542,N_19693);
nor U21158 (N_21158,N_18627,N_19033);
nand U21159 (N_21159,N_18058,N_18724);
nand U21160 (N_21160,N_18886,N_18147);
and U21161 (N_21161,N_18229,N_19488);
or U21162 (N_21162,N_18123,N_19337);
and U21163 (N_21163,N_18974,N_19269);
xnor U21164 (N_21164,N_19076,N_19751);
nand U21165 (N_21165,N_18676,N_19199);
nor U21166 (N_21166,N_19281,N_19688);
and U21167 (N_21167,N_19348,N_18050);
or U21168 (N_21168,N_19007,N_19260);
nand U21169 (N_21169,N_18749,N_19026);
nand U21170 (N_21170,N_19284,N_18195);
and U21171 (N_21171,N_19068,N_18035);
or U21172 (N_21172,N_19735,N_19227);
and U21173 (N_21173,N_19992,N_18547);
or U21174 (N_21174,N_19318,N_18346);
nor U21175 (N_21175,N_18875,N_18923);
nand U21176 (N_21176,N_18960,N_19726);
or U21177 (N_21177,N_19750,N_19038);
xnor U21178 (N_21178,N_19938,N_18013);
or U21179 (N_21179,N_18625,N_19397);
nor U21180 (N_21180,N_19289,N_18903);
and U21181 (N_21181,N_19025,N_18060);
xor U21182 (N_21182,N_18985,N_18109);
and U21183 (N_21183,N_18878,N_19767);
nor U21184 (N_21184,N_19123,N_18946);
nand U21185 (N_21185,N_19174,N_18888);
nor U21186 (N_21186,N_18852,N_19825);
and U21187 (N_21187,N_18271,N_19531);
or U21188 (N_21188,N_19273,N_18731);
xor U21189 (N_21189,N_19514,N_19265);
xor U21190 (N_21190,N_19035,N_18637);
and U21191 (N_21191,N_18647,N_18167);
nor U21192 (N_21192,N_18436,N_19487);
or U21193 (N_21193,N_18211,N_18274);
xnor U21194 (N_21194,N_19226,N_18276);
nand U21195 (N_21195,N_19039,N_18457);
and U21196 (N_21196,N_19394,N_18814);
nor U21197 (N_21197,N_18327,N_18502);
xor U21198 (N_21198,N_19855,N_19566);
nand U21199 (N_21199,N_18424,N_18196);
nor U21200 (N_21200,N_19627,N_18071);
and U21201 (N_21201,N_18096,N_19858);
nor U21202 (N_21202,N_18526,N_19192);
nand U21203 (N_21203,N_18204,N_19803);
nor U21204 (N_21204,N_19960,N_19315);
xnor U21205 (N_21205,N_18453,N_18259);
nand U21206 (N_21206,N_19522,N_19057);
nand U21207 (N_21207,N_18155,N_19762);
xnor U21208 (N_21208,N_18975,N_19060);
nand U21209 (N_21209,N_18506,N_18624);
nor U21210 (N_21210,N_18534,N_19740);
or U21211 (N_21211,N_18817,N_19246);
xnor U21212 (N_21212,N_19435,N_18234);
xor U21213 (N_21213,N_18446,N_19400);
or U21214 (N_21214,N_18133,N_19303);
xor U21215 (N_21215,N_19660,N_18346);
xnor U21216 (N_21216,N_18693,N_18948);
xnor U21217 (N_21217,N_19940,N_19374);
nor U21218 (N_21218,N_19049,N_19980);
nor U21219 (N_21219,N_19947,N_19988);
nor U21220 (N_21220,N_18352,N_18543);
or U21221 (N_21221,N_18162,N_18881);
nand U21222 (N_21222,N_18002,N_18988);
nand U21223 (N_21223,N_18587,N_18890);
and U21224 (N_21224,N_18826,N_18534);
or U21225 (N_21225,N_19291,N_18642);
or U21226 (N_21226,N_19624,N_19876);
xnor U21227 (N_21227,N_19160,N_19937);
nand U21228 (N_21228,N_18986,N_19293);
xnor U21229 (N_21229,N_19180,N_19868);
nor U21230 (N_21230,N_19722,N_19379);
and U21231 (N_21231,N_19643,N_19880);
and U21232 (N_21232,N_18468,N_18812);
and U21233 (N_21233,N_19796,N_18079);
and U21234 (N_21234,N_19507,N_19191);
and U21235 (N_21235,N_18370,N_18529);
nor U21236 (N_21236,N_19535,N_19463);
and U21237 (N_21237,N_19467,N_19333);
or U21238 (N_21238,N_19239,N_19421);
xnor U21239 (N_21239,N_18968,N_19929);
or U21240 (N_21240,N_18717,N_19597);
and U21241 (N_21241,N_18069,N_18623);
and U21242 (N_21242,N_18401,N_18426);
nand U21243 (N_21243,N_19336,N_18770);
or U21244 (N_21244,N_19443,N_18069);
xnor U21245 (N_21245,N_18361,N_18701);
nand U21246 (N_21246,N_19164,N_18247);
nand U21247 (N_21247,N_19889,N_19418);
nand U21248 (N_21248,N_18749,N_19574);
nand U21249 (N_21249,N_19490,N_19994);
and U21250 (N_21250,N_18276,N_18146);
nor U21251 (N_21251,N_19121,N_18560);
nor U21252 (N_21252,N_19679,N_18323);
xor U21253 (N_21253,N_18323,N_18541);
nor U21254 (N_21254,N_19781,N_19528);
nor U21255 (N_21255,N_19761,N_19104);
xnor U21256 (N_21256,N_19902,N_19780);
xnor U21257 (N_21257,N_19266,N_18334);
or U21258 (N_21258,N_18293,N_19178);
and U21259 (N_21259,N_18949,N_18722);
xnor U21260 (N_21260,N_19904,N_19125);
nand U21261 (N_21261,N_19680,N_19700);
nand U21262 (N_21262,N_18672,N_18071);
or U21263 (N_21263,N_19072,N_18463);
nor U21264 (N_21264,N_18463,N_19165);
or U21265 (N_21265,N_19938,N_19251);
and U21266 (N_21266,N_18836,N_19555);
and U21267 (N_21267,N_19104,N_18025);
xor U21268 (N_21268,N_18553,N_19078);
xor U21269 (N_21269,N_18512,N_19869);
nor U21270 (N_21270,N_19558,N_19597);
or U21271 (N_21271,N_19830,N_18393);
and U21272 (N_21272,N_19620,N_19656);
nand U21273 (N_21273,N_18361,N_18805);
nand U21274 (N_21274,N_19957,N_18531);
nor U21275 (N_21275,N_18295,N_18538);
xor U21276 (N_21276,N_18090,N_19283);
or U21277 (N_21277,N_19922,N_18963);
nand U21278 (N_21278,N_18395,N_18235);
and U21279 (N_21279,N_19294,N_19740);
or U21280 (N_21280,N_19042,N_19912);
and U21281 (N_21281,N_19486,N_18630);
or U21282 (N_21282,N_19732,N_19729);
and U21283 (N_21283,N_19144,N_19360);
xor U21284 (N_21284,N_19125,N_18688);
nor U21285 (N_21285,N_18557,N_18896);
or U21286 (N_21286,N_18175,N_19229);
nand U21287 (N_21287,N_19070,N_18920);
xnor U21288 (N_21288,N_18395,N_19761);
nor U21289 (N_21289,N_18170,N_18963);
and U21290 (N_21290,N_19490,N_19378);
or U21291 (N_21291,N_19284,N_19904);
nor U21292 (N_21292,N_19341,N_18765);
nor U21293 (N_21293,N_18127,N_19121);
or U21294 (N_21294,N_18244,N_18523);
nand U21295 (N_21295,N_18328,N_19811);
and U21296 (N_21296,N_19943,N_19120);
nand U21297 (N_21297,N_19963,N_18157);
nor U21298 (N_21298,N_19818,N_18527);
xor U21299 (N_21299,N_18688,N_18394);
nand U21300 (N_21300,N_19563,N_18536);
xnor U21301 (N_21301,N_18580,N_19824);
xor U21302 (N_21302,N_18768,N_19525);
and U21303 (N_21303,N_18654,N_18908);
or U21304 (N_21304,N_18530,N_19343);
and U21305 (N_21305,N_18169,N_19280);
nor U21306 (N_21306,N_18450,N_19172);
nand U21307 (N_21307,N_19541,N_19432);
nand U21308 (N_21308,N_18717,N_19666);
nor U21309 (N_21309,N_19816,N_19291);
xor U21310 (N_21310,N_18107,N_18730);
and U21311 (N_21311,N_19310,N_19378);
xnor U21312 (N_21312,N_18279,N_19381);
or U21313 (N_21313,N_18212,N_18464);
nand U21314 (N_21314,N_18175,N_19464);
xnor U21315 (N_21315,N_18999,N_18196);
or U21316 (N_21316,N_18968,N_18802);
or U21317 (N_21317,N_19878,N_18031);
and U21318 (N_21318,N_18636,N_18703);
nand U21319 (N_21319,N_19981,N_19992);
and U21320 (N_21320,N_18382,N_18659);
and U21321 (N_21321,N_18027,N_18924);
nand U21322 (N_21322,N_19999,N_19853);
nand U21323 (N_21323,N_19375,N_19125);
nand U21324 (N_21324,N_19910,N_18339);
nand U21325 (N_21325,N_18598,N_18584);
or U21326 (N_21326,N_19235,N_19250);
nor U21327 (N_21327,N_19635,N_19768);
xnor U21328 (N_21328,N_18981,N_18120);
xor U21329 (N_21329,N_19400,N_18870);
and U21330 (N_21330,N_18614,N_18302);
and U21331 (N_21331,N_18089,N_18832);
xnor U21332 (N_21332,N_19542,N_19928);
xor U21333 (N_21333,N_19073,N_18526);
xnor U21334 (N_21334,N_18031,N_18330);
and U21335 (N_21335,N_18853,N_18400);
or U21336 (N_21336,N_18508,N_18295);
nor U21337 (N_21337,N_18049,N_18959);
nor U21338 (N_21338,N_19173,N_18238);
or U21339 (N_21339,N_19797,N_18906);
nand U21340 (N_21340,N_19141,N_19079);
or U21341 (N_21341,N_19623,N_18216);
or U21342 (N_21342,N_19754,N_18287);
xor U21343 (N_21343,N_18361,N_19766);
nand U21344 (N_21344,N_19548,N_18740);
nand U21345 (N_21345,N_19924,N_19364);
xor U21346 (N_21346,N_19199,N_19001);
or U21347 (N_21347,N_19786,N_18475);
and U21348 (N_21348,N_18069,N_19168);
xnor U21349 (N_21349,N_18915,N_19764);
or U21350 (N_21350,N_19001,N_19395);
nor U21351 (N_21351,N_19741,N_18987);
nand U21352 (N_21352,N_18460,N_18097);
nor U21353 (N_21353,N_18511,N_19534);
or U21354 (N_21354,N_19467,N_18322);
nand U21355 (N_21355,N_18399,N_18549);
nand U21356 (N_21356,N_19791,N_18521);
or U21357 (N_21357,N_18162,N_18018);
nand U21358 (N_21358,N_19460,N_18907);
xor U21359 (N_21359,N_18601,N_19782);
nor U21360 (N_21360,N_18624,N_18269);
or U21361 (N_21361,N_19432,N_19478);
nand U21362 (N_21362,N_18675,N_18075);
xor U21363 (N_21363,N_18794,N_19925);
or U21364 (N_21364,N_18890,N_18115);
nand U21365 (N_21365,N_18811,N_18596);
nor U21366 (N_21366,N_18873,N_18039);
xor U21367 (N_21367,N_18897,N_18658);
nor U21368 (N_21368,N_19995,N_18865);
nand U21369 (N_21369,N_19557,N_19954);
nand U21370 (N_21370,N_19566,N_19042);
xor U21371 (N_21371,N_18877,N_19781);
nor U21372 (N_21372,N_18791,N_18518);
or U21373 (N_21373,N_19916,N_19004);
or U21374 (N_21374,N_18690,N_18692);
xnor U21375 (N_21375,N_18450,N_19822);
xor U21376 (N_21376,N_19747,N_18012);
or U21377 (N_21377,N_18479,N_19101);
or U21378 (N_21378,N_19141,N_18717);
nand U21379 (N_21379,N_18574,N_19478);
nor U21380 (N_21380,N_19616,N_18001);
or U21381 (N_21381,N_18865,N_18401);
or U21382 (N_21382,N_18202,N_18521);
or U21383 (N_21383,N_18844,N_19647);
and U21384 (N_21384,N_19363,N_18806);
and U21385 (N_21385,N_18152,N_19087);
nand U21386 (N_21386,N_19330,N_18594);
and U21387 (N_21387,N_19307,N_18454);
nor U21388 (N_21388,N_18191,N_18369);
and U21389 (N_21389,N_19912,N_19509);
nor U21390 (N_21390,N_19145,N_18515);
xor U21391 (N_21391,N_19704,N_19989);
xnor U21392 (N_21392,N_19984,N_19271);
or U21393 (N_21393,N_18837,N_19866);
nand U21394 (N_21394,N_18272,N_19535);
and U21395 (N_21395,N_18292,N_18453);
nor U21396 (N_21396,N_18702,N_18201);
or U21397 (N_21397,N_18100,N_19831);
nor U21398 (N_21398,N_18639,N_19214);
or U21399 (N_21399,N_18661,N_18048);
nor U21400 (N_21400,N_18295,N_18938);
and U21401 (N_21401,N_18462,N_18170);
or U21402 (N_21402,N_19352,N_18720);
xor U21403 (N_21403,N_19331,N_19837);
and U21404 (N_21404,N_19060,N_18920);
nor U21405 (N_21405,N_19348,N_19087);
and U21406 (N_21406,N_19095,N_18537);
and U21407 (N_21407,N_19976,N_18915);
or U21408 (N_21408,N_19974,N_19525);
nand U21409 (N_21409,N_19767,N_18649);
nand U21410 (N_21410,N_18114,N_18870);
and U21411 (N_21411,N_19793,N_18874);
and U21412 (N_21412,N_19477,N_19729);
nand U21413 (N_21413,N_18454,N_19935);
xor U21414 (N_21414,N_19055,N_19326);
or U21415 (N_21415,N_18636,N_19366);
or U21416 (N_21416,N_18459,N_18539);
xor U21417 (N_21417,N_18715,N_18386);
xor U21418 (N_21418,N_19467,N_19001);
xor U21419 (N_21419,N_18284,N_18485);
xor U21420 (N_21420,N_19281,N_18136);
xor U21421 (N_21421,N_18023,N_19609);
or U21422 (N_21422,N_19412,N_19695);
xor U21423 (N_21423,N_19784,N_19544);
and U21424 (N_21424,N_18803,N_19737);
nand U21425 (N_21425,N_18321,N_19135);
and U21426 (N_21426,N_18265,N_19539);
nor U21427 (N_21427,N_18424,N_18990);
nor U21428 (N_21428,N_19161,N_19644);
or U21429 (N_21429,N_18096,N_18082);
nor U21430 (N_21430,N_18819,N_19734);
nor U21431 (N_21431,N_19240,N_18007);
nor U21432 (N_21432,N_18910,N_19211);
xor U21433 (N_21433,N_19318,N_18550);
or U21434 (N_21434,N_18196,N_19141);
or U21435 (N_21435,N_18302,N_18453);
and U21436 (N_21436,N_19605,N_19451);
and U21437 (N_21437,N_19832,N_19000);
or U21438 (N_21438,N_18789,N_19224);
or U21439 (N_21439,N_19097,N_18251);
and U21440 (N_21440,N_18661,N_18283);
nand U21441 (N_21441,N_18823,N_19428);
xnor U21442 (N_21442,N_18339,N_18299);
nand U21443 (N_21443,N_19749,N_18098);
nor U21444 (N_21444,N_19803,N_18026);
and U21445 (N_21445,N_19688,N_19958);
and U21446 (N_21446,N_19349,N_19406);
xor U21447 (N_21447,N_19409,N_19111);
xor U21448 (N_21448,N_18737,N_18603);
xnor U21449 (N_21449,N_18118,N_19834);
nor U21450 (N_21450,N_19728,N_18670);
or U21451 (N_21451,N_18957,N_18822);
nor U21452 (N_21452,N_19009,N_18694);
or U21453 (N_21453,N_18347,N_18890);
xnor U21454 (N_21454,N_18417,N_19026);
nor U21455 (N_21455,N_18463,N_18716);
nand U21456 (N_21456,N_19958,N_19780);
nor U21457 (N_21457,N_18501,N_18236);
nand U21458 (N_21458,N_19358,N_18213);
and U21459 (N_21459,N_18969,N_19194);
and U21460 (N_21460,N_19205,N_19620);
nand U21461 (N_21461,N_18702,N_18659);
or U21462 (N_21462,N_18540,N_18160);
or U21463 (N_21463,N_19316,N_18935);
nand U21464 (N_21464,N_18966,N_19948);
xor U21465 (N_21465,N_18499,N_19974);
nand U21466 (N_21466,N_19709,N_19445);
or U21467 (N_21467,N_18366,N_19917);
nor U21468 (N_21468,N_19097,N_19692);
or U21469 (N_21469,N_18203,N_18146);
xor U21470 (N_21470,N_19788,N_18243);
nor U21471 (N_21471,N_19712,N_18738);
nand U21472 (N_21472,N_18855,N_18856);
nor U21473 (N_21473,N_18015,N_19250);
or U21474 (N_21474,N_19569,N_18143);
and U21475 (N_21475,N_18521,N_18686);
and U21476 (N_21476,N_18817,N_19753);
or U21477 (N_21477,N_19524,N_19662);
nor U21478 (N_21478,N_18875,N_19231);
nor U21479 (N_21479,N_18648,N_18173);
xor U21480 (N_21480,N_19098,N_19611);
or U21481 (N_21481,N_19037,N_19140);
or U21482 (N_21482,N_19706,N_18875);
and U21483 (N_21483,N_19306,N_18588);
nor U21484 (N_21484,N_19773,N_19682);
or U21485 (N_21485,N_18593,N_19272);
xor U21486 (N_21486,N_19255,N_19422);
nand U21487 (N_21487,N_19999,N_18249);
nand U21488 (N_21488,N_18021,N_18554);
xor U21489 (N_21489,N_18959,N_19921);
and U21490 (N_21490,N_18940,N_18130);
nor U21491 (N_21491,N_19565,N_18446);
nand U21492 (N_21492,N_18125,N_18843);
and U21493 (N_21493,N_18747,N_18105);
xnor U21494 (N_21494,N_18283,N_18172);
and U21495 (N_21495,N_19309,N_18405);
nor U21496 (N_21496,N_19285,N_19527);
xnor U21497 (N_21497,N_18608,N_19327);
and U21498 (N_21498,N_18755,N_18416);
and U21499 (N_21499,N_19176,N_19037);
or U21500 (N_21500,N_19769,N_19019);
nor U21501 (N_21501,N_19361,N_19033);
and U21502 (N_21502,N_18002,N_19289);
or U21503 (N_21503,N_18524,N_19544);
nor U21504 (N_21504,N_18159,N_19842);
xor U21505 (N_21505,N_19885,N_19327);
xnor U21506 (N_21506,N_19860,N_19315);
and U21507 (N_21507,N_19583,N_18098);
nor U21508 (N_21508,N_19422,N_18581);
nor U21509 (N_21509,N_18179,N_19820);
and U21510 (N_21510,N_19458,N_18438);
nand U21511 (N_21511,N_19894,N_18354);
and U21512 (N_21512,N_19806,N_18704);
and U21513 (N_21513,N_19701,N_19259);
and U21514 (N_21514,N_19968,N_18052);
and U21515 (N_21515,N_18321,N_18370);
xnor U21516 (N_21516,N_19093,N_18074);
nand U21517 (N_21517,N_19209,N_19057);
xnor U21518 (N_21518,N_18161,N_18273);
or U21519 (N_21519,N_19562,N_18702);
nand U21520 (N_21520,N_18164,N_19054);
nor U21521 (N_21521,N_18964,N_19062);
nor U21522 (N_21522,N_18095,N_19115);
or U21523 (N_21523,N_19307,N_19945);
nand U21524 (N_21524,N_18288,N_19115);
or U21525 (N_21525,N_18162,N_18688);
nor U21526 (N_21526,N_18652,N_19393);
nand U21527 (N_21527,N_18046,N_19465);
xor U21528 (N_21528,N_19096,N_18295);
and U21529 (N_21529,N_18323,N_18748);
nand U21530 (N_21530,N_19988,N_19470);
or U21531 (N_21531,N_18387,N_19032);
nand U21532 (N_21532,N_19747,N_18195);
or U21533 (N_21533,N_19498,N_19341);
and U21534 (N_21534,N_18828,N_18568);
and U21535 (N_21535,N_18455,N_18358);
nand U21536 (N_21536,N_18001,N_19650);
nand U21537 (N_21537,N_18900,N_19867);
nand U21538 (N_21538,N_18621,N_19774);
nand U21539 (N_21539,N_18974,N_18556);
nand U21540 (N_21540,N_18266,N_19669);
or U21541 (N_21541,N_18567,N_19919);
and U21542 (N_21542,N_19446,N_19684);
nor U21543 (N_21543,N_19992,N_18426);
xnor U21544 (N_21544,N_18522,N_18131);
and U21545 (N_21545,N_18401,N_18993);
or U21546 (N_21546,N_19486,N_18584);
and U21547 (N_21547,N_19004,N_18222);
and U21548 (N_21548,N_18028,N_19417);
xor U21549 (N_21549,N_19452,N_19138);
and U21550 (N_21550,N_18581,N_19273);
nor U21551 (N_21551,N_19455,N_19257);
xor U21552 (N_21552,N_18661,N_19231);
and U21553 (N_21553,N_18843,N_19836);
xnor U21554 (N_21554,N_19973,N_19448);
nor U21555 (N_21555,N_18527,N_19598);
and U21556 (N_21556,N_18739,N_18131);
xor U21557 (N_21557,N_19459,N_19008);
nor U21558 (N_21558,N_19781,N_19868);
or U21559 (N_21559,N_18444,N_18617);
and U21560 (N_21560,N_19563,N_18492);
and U21561 (N_21561,N_18038,N_19454);
or U21562 (N_21562,N_18697,N_18254);
or U21563 (N_21563,N_19549,N_19064);
nand U21564 (N_21564,N_19232,N_18359);
or U21565 (N_21565,N_19827,N_18388);
nand U21566 (N_21566,N_18753,N_18955);
xor U21567 (N_21567,N_18315,N_19464);
or U21568 (N_21568,N_19307,N_19419);
nand U21569 (N_21569,N_18623,N_18748);
and U21570 (N_21570,N_18829,N_19546);
and U21571 (N_21571,N_19827,N_18426);
or U21572 (N_21572,N_18289,N_19934);
nor U21573 (N_21573,N_19856,N_19100);
xor U21574 (N_21574,N_19192,N_19277);
xor U21575 (N_21575,N_19737,N_18013);
xnor U21576 (N_21576,N_18668,N_19069);
and U21577 (N_21577,N_18254,N_18257);
nor U21578 (N_21578,N_19347,N_18703);
nand U21579 (N_21579,N_19921,N_19954);
or U21580 (N_21580,N_18754,N_19071);
nor U21581 (N_21581,N_18326,N_18495);
nand U21582 (N_21582,N_19238,N_18584);
xor U21583 (N_21583,N_18709,N_18821);
or U21584 (N_21584,N_19403,N_18402);
or U21585 (N_21585,N_19142,N_19723);
xnor U21586 (N_21586,N_19559,N_19673);
nor U21587 (N_21587,N_18184,N_19677);
nand U21588 (N_21588,N_19035,N_19753);
nor U21589 (N_21589,N_18988,N_18454);
and U21590 (N_21590,N_18636,N_18812);
or U21591 (N_21591,N_18667,N_18808);
or U21592 (N_21592,N_19315,N_19041);
nor U21593 (N_21593,N_19063,N_18726);
nor U21594 (N_21594,N_19352,N_19280);
or U21595 (N_21595,N_19034,N_18315);
xnor U21596 (N_21596,N_19654,N_18201);
nor U21597 (N_21597,N_19697,N_18239);
xor U21598 (N_21598,N_19813,N_19419);
or U21599 (N_21599,N_18838,N_19774);
nor U21600 (N_21600,N_19681,N_18480);
or U21601 (N_21601,N_18298,N_19426);
nor U21602 (N_21602,N_19519,N_19415);
nand U21603 (N_21603,N_19138,N_19847);
or U21604 (N_21604,N_18633,N_19394);
nor U21605 (N_21605,N_19908,N_18278);
nor U21606 (N_21606,N_18999,N_19587);
and U21607 (N_21607,N_19407,N_19173);
or U21608 (N_21608,N_18541,N_18554);
nand U21609 (N_21609,N_18544,N_19037);
nand U21610 (N_21610,N_19430,N_18474);
xor U21611 (N_21611,N_19509,N_19322);
or U21612 (N_21612,N_18624,N_18692);
and U21613 (N_21613,N_19614,N_19411);
or U21614 (N_21614,N_18667,N_19298);
nor U21615 (N_21615,N_18039,N_18409);
or U21616 (N_21616,N_19650,N_19069);
nor U21617 (N_21617,N_19305,N_19087);
or U21618 (N_21618,N_19628,N_18413);
xor U21619 (N_21619,N_18499,N_18808);
or U21620 (N_21620,N_19105,N_18172);
and U21621 (N_21621,N_18475,N_18303);
and U21622 (N_21622,N_18765,N_18198);
nand U21623 (N_21623,N_19382,N_19533);
xnor U21624 (N_21624,N_19312,N_18174);
and U21625 (N_21625,N_19038,N_18218);
or U21626 (N_21626,N_19780,N_19991);
nor U21627 (N_21627,N_19050,N_18669);
or U21628 (N_21628,N_18929,N_18333);
nor U21629 (N_21629,N_19635,N_18876);
xor U21630 (N_21630,N_19611,N_18906);
or U21631 (N_21631,N_19688,N_18884);
nand U21632 (N_21632,N_19311,N_19336);
xnor U21633 (N_21633,N_19419,N_19455);
nor U21634 (N_21634,N_18119,N_19795);
nand U21635 (N_21635,N_19041,N_18254);
nand U21636 (N_21636,N_19056,N_18797);
and U21637 (N_21637,N_18782,N_19998);
or U21638 (N_21638,N_19224,N_19568);
nor U21639 (N_21639,N_19732,N_19146);
nor U21640 (N_21640,N_19678,N_18460);
nand U21641 (N_21641,N_18288,N_19801);
xor U21642 (N_21642,N_19484,N_18997);
nand U21643 (N_21643,N_19739,N_19632);
nor U21644 (N_21644,N_18963,N_19608);
nor U21645 (N_21645,N_18157,N_19776);
nand U21646 (N_21646,N_18957,N_19040);
or U21647 (N_21647,N_19211,N_19370);
nor U21648 (N_21648,N_19520,N_18374);
nand U21649 (N_21649,N_18498,N_18399);
or U21650 (N_21650,N_18343,N_18979);
and U21651 (N_21651,N_18586,N_19004);
nor U21652 (N_21652,N_19209,N_19922);
or U21653 (N_21653,N_19258,N_18390);
nand U21654 (N_21654,N_19832,N_19931);
nor U21655 (N_21655,N_19335,N_19699);
nand U21656 (N_21656,N_19894,N_19732);
and U21657 (N_21657,N_18768,N_19021);
and U21658 (N_21658,N_19029,N_18430);
and U21659 (N_21659,N_19045,N_19983);
nand U21660 (N_21660,N_18182,N_18726);
nand U21661 (N_21661,N_18163,N_18339);
nand U21662 (N_21662,N_19233,N_18478);
and U21663 (N_21663,N_18084,N_19900);
xor U21664 (N_21664,N_18580,N_18484);
nand U21665 (N_21665,N_18564,N_19865);
nor U21666 (N_21666,N_18521,N_19494);
xnor U21667 (N_21667,N_18874,N_19242);
or U21668 (N_21668,N_19111,N_18859);
nor U21669 (N_21669,N_19794,N_19831);
xnor U21670 (N_21670,N_19870,N_18136);
and U21671 (N_21671,N_18102,N_18307);
or U21672 (N_21672,N_19208,N_18857);
xor U21673 (N_21673,N_19686,N_18553);
xnor U21674 (N_21674,N_19621,N_19027);
or U21675 (N_21675,N_19092,N_19552);
xnor U21676 (N_21676,N_19982,N_19331);
nor U21677 (N_21677,N_18452,N_19209);
and U21678 (N_21678,N_19671,N_19983);
nand U21679 (N_21679,N_18494,N_18016);
nand U21680 (N_21680,N_19020,N_19021);
nor U21681 (N_21681,N_18291,N_19631);
and U21682 (N_21682,N_18768,N_18309);
or U21683 (N_21683,N_19366,N_19279);
nand U21684 (N_21684,N_18084,N_19142);
xnor U21685 (N_21685,N_18774,N_18838);
or U21686 (N_21686,N_18273,N_18985);
or U21687 (N_21687,N_18108,N_18368);
nor U21688 (N_21688,N_18832,N_18009);
nand U21689 (N_21689,N_18644,N_19017);
xnor U21690 (N_21690,N_19435,N_19453);
nor U21691 (N_21691,N_19345,N_18012);
and U21692 (N_21692,N_19202,N_18868);
nand U21693 (N_21693,N_18373,N_18810);
and U21694 (N_21694,N_19484,N_18672);
nand U21695 (N_21695,N_18238,N_18852);
nand U21696 (N_21696,N_19061,N_18455);
or U21697 (N_21697,N_18797,N_18873);
and U21698 (N_21698,N_19678,N_19748);
nor U21699 (N_21699,N_18814,N_18057);
or U21700 (N_21700,N_18739,N_18437);
xor U21701 (N_21701,N_18828,N_19849);
and U21702 (N_21702,N_19924,N_18934);
xnor U21703 (N_21703,N_18736,N_18111);
and U21704 (N_21704,N_19350,N_19557);
and U21705 (N_21705,N_19570,N_18005);
or U21706 (N_21706,N_19918,N_19652);
nor U21707 (N_21707,N_19824,N_18123);
and U21708 (N_21708,N_18062,N_18685);
xnor U21709 (N_21709,N_18033,N_19954);
or U21710 (N_21710,N_18176,N_18077);
nand U21711 (N_21711,N_19888,N_19855);
nor U21712 (N_21712,N_18159,N_18827);
and U21713 (N_21713,N_19620,N_19089);
and U21714 (N_21714,N_18518,N_18632);
nand U21715 (N_21715,N_18601,N_19110);
nand U21716 (N_21716,N_18263,N_18109);
and U21717 (N_21717,N_18357,N_19440);
xor U21718 (N_21718,N_18318,N_18498);
nand U21719 (N_21719,N_19587,N_18532);
and U21720 (N_21720,N_18545,N_19485);
nand U21721 (N_21721,N_18835,N_19648);
or U21722 (N_21722,N_18504,N_19522);
nor U21723 (N_21723,N_19439,N_19181);
xor U21724 (N_21724,N_18245,N_19759);
and U21725 (N_21725,N_18022,N_19642);
or U21726 (N_21726,N_18330,N_18054);
nand U21727 (N_21727,N_18928,N_18000);
or U21728 (N_21728,N_18919,N_19956);
or U21729 (N_21729,N_18885,N_18918);
or U21730 (N_21730,N_19257,N_18673);
nand U21731 (N_21731,N_18723,N_18898);
xor U21732 (N_21732,N_19184,N_18384);
nand U21733 (N_21733,N_19437,N_18445);
or U21734 (N_21734,N_19940,N_19574);
xor U21735 (N_21735,N_19384,N_19852);
xor U21736 (N_21736,N_18911,N_18521);
or U21737 (N_21737,N_19445,N_18901);
and U21738 (N_21738,N_18229,N_18047);
xor U21739 (N_21739,N_19290,N_18818);
xor U21740 (N_21740,N_18828,N_19588);
nor U21741 (N_21741,N_19712,N_19449);
nand U21742 (N_21742,N_18540,N_19394);
nand U21743 (N_21743,N_19312,N_18126);
nor U21744 (N_21744,N_19815,N_19197);
nor U21745 (N_21745,N_19703,N_19559);
or U21746 (N_21746,N_19237,N_19332);
nor U21747 (N_21747,N_18094,N_18864);
nor U21748 (N_21748,N_18646,N_18776);
nand U21749 (N_21749,N_18817,N_19486);
nor U21750 (N_21750,N_18831,N_18354);
nor U21751 (N_21751,N_18318,N_18568);
nand U21752 (N_21752,N_19026,N_18590);
or U21753 (N_21753,N_19809,N_19581);
and U21754 (N_21754,N_19753,N_18141);
and U21755 (N_21755,N_19358,N_18294);
and U21756 (N_21756,N_19518,N_19584);
or U21757 (N_21757,N_18827,N_19131);
xnor U21758 (N_21758,N_19125,N_18181);
xor U21759 (N_21759,N_19423,N_18317);
and U21760 (N_21760,N_18845,N_18643);
xnor U21761 (N_21761,N_19078,N_18738);
and U21762 (N_21762,N_19580,N_18766);
and U21763 (N_21763,N_18675,N_18691);
or U21764 (N_21764,N_19370,N_18661);
and U21765 (N_21765,N_19841,N_19810);
or U21766 (N_21766,N_18171,N_18342);
nand U21767 (N_21767,N_18587,N_19152);
nand U21768 (N_21768,N_19844,N_18994);
and U21769 (N_21769,N_19792,N_19014);
xor U21770 (N_21770,N_19807,N_18867);
nor U21771 (N_21771,N_18326,N_18706);
or U21772 (N_21772,N_19075,N_19639);
or U21773 (N_21773,N_18181,N_18604);
or U21774 (N_21774,N_18593,N_19938);
nor U21775 (N_21775,N_19787,N_19083);
nor U21776 (N_21776,N_19016,N_19766);
nor U21777 (N_21777,N_18693,N_18814);
nor U21778 (N_21778,N_19598,N_18067);
xor U21779 (N_21779,N_19653,N_18998);
nand U21780 (N_21780,N_18338,N_19568);
or U21781 (N_21781,N_18323,N_19547);
and U21782 (N_21782,N_19451,N_18460);
or U21783 (N_21783,N_19920,N_18737);
xor U21784 (N_21784,N_18038,N_19746);
and U21785 (N_21785,N_19836,N_18462);
or U21786 (N_21786,N_19389,N_19647);
xor U21787 (N_21787,N_18332,N_19750);
and U21788 (N_21788,N_18129,N_18671);
xnor U21789 (N_21789,N_19816,N_18546);
or U21790 (N_21790,N_19882,N_18320);
and U21791 (N_21791,N_19053,N_19847);
and U21792 (N_21792,N_19248,N_19346);
xor U21793 (N_21793,N_19175,N_18728);
nand U21794 (N_21794,N_19225,N_19401);
xnor U21795 (N_21795,N_19069,N_18727);
xor U21796 (N_21796,N_19183,N_18514);
and U21797 (N_21797,N_19014,N_18998);
nor U21798 (N_21798,N_18163,N_18621);
or U21799 (N_21799,N_19883,N_19918);
nor U21800 (N_21800,N_19911,N_19063);
or U21801 (N_21801,N_19732,N_19018);
and U21802 (N_21802,N_19171,N_18455);
nand U21803 (N_21803,N_19499,N_19398);
nand U21804 (N_21804,N_18887,N_19280);
and U21805 (N_21805,N_19029,N_19859);
and U21806 (N_21806,N_19217,N_18663);
nor U21807 (N_21807,N_18817,N_18856);
and U21808 (N_21808,N_19771,N_18779);
xnor U21809 (N_21809,N_18670,N_18207);
xnor U21810 (N_21810,N_19854,N_19235);
and U21811 (N_21811,N_18076,N_18674);
xnor U21812 (N_21812,N_18627,N_19730);
nor U21813 (N_21813,N_18433,N_19528);
or U21814 (N_21814,N_18952,N_18794);
nand U21815 (N_21815,N_18451,N_19993);
and U21816 (N_21816,N_18323,N_18050);
or U21817 (N_21817,N_19125,N_19729);
xor U21818 (N_21818,N_18861,N_18464);
xor U21819 (N_21819,N_19230,N_19180);
or U21820 (N_21820,N_19161,N_19492);
nor U21821 (N_21821,N_18152,N_19885);
nand U21822 (N_21822,N_18075,N_19791);
xnor U21823 (N_21823,N_18041,N_18621);
nand U21824 (N_21824,N_18055,N_19618);
and U21825 (N_21825,N_18876,N_19299);
or U21826 (N_21826,N_18730,N_19753);
nand U21827 (N_21827,N_19388,N_18153);
or U21828 (N_21828,N_18731,N_18149);
nand U21829 (N_21829,N_18186,N_18676);
and U21830 (N_21830,N_18962,N_18815);
xor U21831 (N_21831,N_18418,N_19592);
nor U21832 (N_21832,N_19419,N_18678);
and U21833 (N_21833,N_19877,N_18884);
and U21834 (N_21834,N_19328,N_19097);
and U21835 (N_21835,N_18407,N_19305);
nor U21836 (N_21836,N_19578,N_19066);
nor U21837 (N_21837,N_19930,N_19653);
nand U21838 (N_21838,N_19525,N_18745);
and U21839 (N_21839,N_18520,N_18408);
and U21840 (N_21840,N_18288,N_19000);
xnor U21841 (N_21841,N_18982,N_18289);
or U21842 (N_21842,N_18696,N_19101);
or U21843 (N_21843,N_19548,N_18442);
or U21844 (N_21844,N_19099,N_19455);
or U21845 (N_21845,N_18955,N_19952);
xor U21846 (N_21846,N_19093,N_19884);
and U21847 (N_21847,N_19966,N_19004);
and U21848 (N_21848,N_19460,N_18428);
and U21849 (N_21849,N_18984,N_18599);
or U21850 (N_21850,N_18443,N_19234);
nand U21851 (N_21851,N_19674,N_18003);
xnor U21852 (N_21852,N_19259,N_19791);
and U21853 (N_21853,N_19655,N_18364);
and U21854 (N_21854,N_18587,N_19727);
xor U21855 (N_21855,N_19265,N_19276);
and U21856 (N_21856,N_19051,N_18255);
and U21857 (N_21857,N_18352,N_19039);
nand U21858 (N_21858,N_19412,N_18610);
nand U21859 (N_21859,N_19650,N_18067);
nor U21860 (N_21860,N_18307,N_19706);
or U21861 (N_21861,N_19730,N_19480);
xor U21862 (N_21862,N_18716,N_19624);
or U21863 (N_21863,N_19602,N_18784);
nand U21864 (N_21864,N_19100,N_19476);
nor U21865 (N_21865,N_19911,N_18046);
nor U21866 (N_21866,N_18919,N_18321);
nor U21867 (N_21867,N_18733,N_18696);
nand U21868 (N_21868,N_18518,N_19170);
nand U21869 (N_21869,N_18934,N_18101);
xor U21870 (N_21870,N_18150,N_19943);
nor U21871 (N_21871,N_19854,N_18130);
nand U21872 (N_21872,N_19890,N_18791);
nor U21873 (N_21873,N_19290,N_18768);
nor U21874 (N_21874,N_18342,N_19315);
nor U21875 (N_21875,N_18528,N_19399);
or U21876 (N_21876,N_19545,N_19350);
and U21877 (N_21877,N_18993,N_18159);
or U21878 (N_21878,N_19939,N_19717);
and U21879 (N_21879,N_18457,N_19397);
and U21880 (N_21880,N_18675,N_19660);
nor U21881 (N_21881,N_19804,N_18785);
nand U21882 (N_21882,N_19083,N_19553);
xnor U21883 (N_21883,N_19826,N_19503);
nor U21884 (N_21884,N_18802,N_19011);
or U21885 (N_21885,N_18632,N_19362);
nor U21886 (N_21886,N_18685,N_18055);
nor U21887 (N_21887,N_18688,N_19323);
nand U21888 (N_21888,N_18581,N_18148);
xnor U21889 (N_21889,N_18405,N_19780);
or U21890 (N_21890,N_19462,N_18124);
nand U21891 (N_21891,N_19630,N_19385);
nand U21892 (N_21892,N_18694,N_19199);
nand U21893 (N_21893,N_19260,N_18256);
and U21894 (N_21894,N_19003,N_19194);
and U21895 (N_21895,N_18359,N_19502);
xor U21896 (N_21896,N_19114,N_19203);
nor U21897 (N_21897,N_18847,N_19297);
xnor U21898 (N_21898,N_19440,N_19465);
nand U21899 (N_21899,N_19188,N_18968);
and U21900 (N_21900,N_18723,N_19286);
and U21901 (N_21901,N_18963,N_19225);
and U21902 (N_21902,N_18662,N_19411);
and U21903 (N_21903,N_18805,N_19011);
nor U21904 (N_21904,N_18578,N_18360);
xor U21905 (N_21905,N_18322,N_19334);
xor U21906 (N_21906,N_19720,N_18796);
nand U21907 (N_21907,N_19975,N_19472);
xor U21908 (N_21908,N_19624,N_18794);
xor U21909 (N_21909,N_18184,N_19746);
nor U21910 (N_21910,N_19251,N_18995);
and U21911 (N_21911,N_18479,N_19121);
nor U21912 (N_21912,N_19829,N_19985);
nor U21913 (N_21913,N_18014,N_18294);
nor U21914 (N_21914,N_19076,N_19711);
or U21915 (N_21915,N_18113,N_18153);
nand U21916 (N_21916,N_19336,N_18493);
nand U21917 (N_21917,N_18253,N_18503);
and U21918 (N_21918,N_18433,N_18109);
nand U21919 (N_21919,N_18584,N_18406);
xor U21920 (N_21920,N_18403,N_19546);
nand U21921 (N_21921,N_19838,N_18392);
xnor U21922 (N_21922,N_19317,N_19468);
or U21923 (N_21923,N_19246,N_19895);
nand U21924 (N_21924,N_19648,N_19733);
or U21925 (N_21925,N_19029,N_19780);
or U21926 (N_21926,N_19085,N_19882);
xor U21927 (N_21927,N_18505,N_18236);
and U21928 (N_21928,N_19150,N_19331);
nand U21929 (N_21929,N_19674,N_19669);
nor U21930 (N_21930,N_18695,N_19605);
nor U21931 (N_21931,N_18750,N_18123);
nand U21932 (N_21932,N_19485,N_18881);
nor U21933 (N_21933,N_19801,N_19797);
nand U21934 (N_21934,N_18350,N_18335);
nor U21935 (N_21935,N_19287,N_18009);
nor U21936 (N_21936,N_18581,N_18425);
nor U21937 (N_21937,N_18310,N_19324);
nor U21938 (N_21938,N_19112,N_18395);
xnor U21939 (N_21939,N_18140,N_19534);
nor U21940 (N_21940,N_19374,N_19541);
xor U21941 (N_21941,N_18876,N_18719);
or U21942 (N_21942,N_19756,N_18617);
xnor U21943 (N_21943,N_18629,N_19194);
and U21944 (N_21944,N_18535,N_18863);
and U21945 (N_21945,N_18487,N_19755);
nor U21946 (N_21946,N_18985,N_19086);
or U21947 (N_21947,N_18918,N_18185);
xnor U21948 (N_21948,N_19007,N_18079);
and U21949 (N_21949,N_18626,N_18882);
nand U21950 (N_21950,N_19928,N_19903);
or U21951 (N_21951,N_18695,N_19795);
or U21952 (N_21952,N_18633,N_18647);
nor U21953 (N_21953,N_18609,N_18261);
nand U21954 (N_21954,N_18889,N_18681);
nor U21955 (N_21955,N_19883,N_18033);
and U21956 (N_21956,N_18795,N_19327);
nand U21957 (N_21957,N_18160,N_19075);
nor U21958 (N_21958,N_18703,N_18275);
and U21959 (N_21959,N_18352,N_19229);
nand U21960 (N_21960,N_18873,N_18388);
and U21961 (N_21961,N_18035,N_19334);
nor U21962 (N_21962,N_19593,N_18527);
xnor U21963 (N_21963,N_18745,N_18445);
or U21964 (N_21964,N_18722,N_18348);
and U21965 (N_21965,N_18068,N_19356);
nor U21966 (N_21966,N_19263,N_19616);
or U21967 (N_21967,N_19756,N_18767);
nand U21968 (N_21968,N_18004,N_19512);
xnor U21969 (N_21969,N_19744,N_18397);
nor U21970 (N_21970,N_19357,N_18331);
and U21971 (N_21971,N_18085,N_18654);
or U21972 (N_21972,N_19670,N_19713);
xnor U21973 (N_21973,N_19006,N_19158);
or U21974 (N_21974,N_19879,N_18982);
and U21975 (N_21975,N_18064,N_19187);
nor U21976 (N_21976,N_18827,N_18028);
or U21977 (N_21977,N_18111,N_19229);
or U21978 (N_21978,N_19185,N_19811);
or U21979 (N_21979,N_19959,N_19869);
or U21980 (N_21980,N_18086,N_18119);
or U21981 (N_21981,N_18542,N_19294);
nand U21982 (N_21982,N_19759,N_18368);
nand U21983 (N_21983,N_18388,N_18889);
and U21984 (N_21984,N_19005,N_18610);
or U21985 (N_21985,N_19900,N_18178);
nand U21986 (N_21986,N_18629,N_19857);
and U21987 (N_21987,N_19132,N_18527);
nand U21988 (N_21988,N_18439,N_18183);
nand U21989 (N_21989,N_19345,N_19679);
or U21990 (N_21990,N_18904,N_19896);
nand U21991 (N_21991,N_18805,N_19891);
xnor U21992 (N_21992,N_19416,N_19549);
and U21993 (N_21993,N_18179,N_19101);
xor U21994 (N_21994,N_18301,N_19503);
nand U21995 (N_21995,N_19876,N_18116);
xor U21996 (N_21996,N_19765,N_18994);
or U21997 (N_21997,N_19114,N_18578);
nand U21998 (N_21998,N_19532,N_19341);
xnor U21999 (N_21999,N_19985,N_19795);
or U22000 (N_22000,N_21365,N_21438);
xnor U22001 (N_22001,N_21425,N_20672);
nor U22002 (N_22002,N_21235,N_20364);
and U22003 (N_22003,N_21732,N_20680);
or U22004 (N_22004,N_21093,N_21561);
nor U22005 (N_22005,N_21480,N_20966);
and U22006 (N_22006,N_20879,N_20895);
xnor U22007 (N_22007,N_21160,N_21088);
or U22008 (N_22008,N_21644,N_20628);
nand U22009 (N_22009,N_21455,N_21866);
nor U22010 (N_22010,N_20337,N_20733);
or U22011 (N_22011,N_21453,N_20410);
nor U22012 (N_22012,N_20185,N_21663);
nand U22013 (N_22013,N_21903,N_20161);
xnor U22014 (N_22014,N_20992,N_20458);
nand U22015 (N_22015,N_20542,N_20502);
or U22016 (N_22016,N_21817,N_21556);
nand U22017 (N_22017,N_20514,N_20774);
and U22018 (N_22018,N_20807,N_21220);
nor U22019 (N_22019,N_20728,N_21163);
nor U22020 (N_22020,N_20102,N_21113);
and U22021 (N_22021,N_21853,N_21970);
or U22022 (N_22022,N_21621,N_20307);
nand U22023 (N_22023,N_21175,N_21413);
nor U22024 (N_22024,N_20990,N_21744);
or U22025 (N_22025,N_20381,N_20689);
or U22026 (N_22026,N_20157,N_20495);
nor U22027 (N_22027,N_20445,N_20105);
nand U22028 (N_22028,N_20974,N_20958);
nand U22029 (N_22029,N_21850,N_21972);
xor U22030 (N_22030,N_20773,N_20581);
xor U22031 (N_22031,N_21386,N_21335);
and U22032 (N_22032,N_20323,N_21071);
nand U22033 (N_22033,N_21822,N_21001);
and U22034 (N_22034,N_21056,N_20694);
nor U22035 (N_22035,N_20266,N_20338);
nor U22036 (N_22036,N_21185,N_20836);
and U22037 (N_22037,N_20249,N_21016);
and U22038 (N_22038,N_20878,N_21796);
and U22039 (N_22039,N_21905,N_21958);
and U22040 (N_22040,N_21594,N_21532);
nor U22041 (N_22041,N_21353,N_20655);
or U22042 (N_22042,N_20621,N_20950);
nand U22043 (N_22043,N_21013,N_21994);
or U22044 (N_22044,N_21389,N_20395);
xor U22045 (N_22045,N_21152,N_21182);
nand U22046 (N_22046,N_21385,N_20016);
nand U22047 (N_22047,N_21026,N_20930);
nor U22048 (N_22048,N_21545,N_21757);
nand U22049 (N_22049,N_21441,N_21526);
and U22050 (N_22050,N_20258,N_21246);
and U22051 (N_22051,N_21833,N_21107);
nor U22052 (N_22052,N_20000,N_20870);
or U22053 (N_22053,N_20500,N_20726);
xnor U22054 (N_22054,N_21697,N_20835);
nand U22055 (N_22055,N_21311,N_20032);
and U22056 (N_22056,N_20729,N_20247);
or U22057 (N_22057,N_20027,N_20420);
and U22058 (N_22058,N_21297,N_20041);
or U22059 (N_22059,N_20312,N_20644);
xnor U22060 (N_22060,N_21483,N_20178);
xnor U22061 (N_22061,N_20480,N_21295);
xor U22062 (N_22062,N_20918,N_20942);
xnor U22063 (N_22063,N_21535,N_21338);
nand U22064 (N_22064,N_21391,N_21890);
and U22065 (N_22065,N_20716,N_21025);
nand U22066 (N_22066,N_20659,N_20685);
nor U22067 (N_22067,N_21178,N_21959);
and U22068 (N_22068,N_21290,N_21166);
and U22069 (N_22069,N_20030,N_21052);
and U22070 (N_22070,N_20798,N_20075);
or U22071 (N_22071,N_20104,N_20664);
xnor U22072 (N_22072,N_21995,N_20885);
or U22073 (N_22073,N_20257,N_20842);
xor U22074 (N_22074,N_21529,N_20417);
nor U22075 (N_22075,N_21352,N_21322);
xor U22076 (N_22076,N_21027,N_21883);
xnor U22077 (N_22077,N_21012,N_21068);
xnor U22078 (N_22078,N_21701,N_21804);
xnor U22079 (N_22079,N_20787,N_20795);
and U22080 (N_22080,N_20704,N_21040);
and U22081 (N_22081,N_20927,N_20781);
nand U22082 (N_22082,N_20822,N_21221);
or U22083 (N_22083,N_21884,N_21775);
nor U22084 (N_22084,N_21601,N_21928);
nand U22085 (N_22085,N_21910,N_20736);
or U22086 (N_22086,N_21437,N_20872);
xnor U22087 (N_22087,N_20993,N_20887);
nor U22088 (N_22088,N_20592,N_21961);
nor U22089 (N_22089,N_20354,N_21269);
nor U22090 (N_22090,N_21622,N_20444);
or U22091 (N_22091,N_21685,N_21493);
and U22092 (N_22092,N_21226,N_20192);
nor U22093 (N_22093,N_21479,N_21579);
xor U22094 (N_22094,N_20864,N_20679);
nor U22095 (N_22095,N_21751,N_20606);
or U22096 (N_22096,N_21294,N_21575);
and U22097 (N_22097,N_20154,N_20675);
or U22098 (N_22098,N_21625,N_20690);
nor U22099 (N_22099,N_20073,N_21608);
or U22100 (N_22100,N_20548,N_21767);
or U22101 (N_22101,N_20439,N_20342);
xnor U22102 (N_22102,N_21860,N_21530);
xor U22103 (N_22103,N_20120,N_21652);
nor U22104 (N_22104,N_20441,N_21123);
and U22105 (N_22105,N_20936,N_21607);
nor U22106 (N_22106,N_21665,N_20335);
xnor U22107 (N_22107,N_20517,N_21129);
nor U22108 (N_22108,N_20768,N_20893);
nand U22109 (N_22109,N_20889,N_20866);
nand U22110 (N_22110,N_20259,N_20479);
nand U22111 (N_22111,N_20788,N_20876);
xor U22112 (N_22112,N_20098,N_21380);
and U22113 (N_22113,N_21296,N_20317);
nand U22114 (N_22114,N_21136,N_20719);
nor U22115 (N_22115,N_20854,N_21733);
nand U22116 (N_22116,N_20806,N_21849);
or U22117 (N_22117,N_21240,N_21315);
nand U22118 (N_22118,N_21042,N_20316);
nand U22119 (N_22119,N_21834,N_21150);
or U22120 (N_22120,N_21891,N_20640);
xnor U22121 (N_22121,N_20633,N_20435);
and U22122 (N_22122,N_21760,N_21555);
nor U22123 (N_22123,N_21251,N_21519);
xor U22124 (N_22124,N_21935,N_20687);
xor U22125 (N_22125,N_20724,N_20196);
xnor U22126 (N_22126,N_21067,N_20860);
nand U22127 (N_22127,N_21004,N_20218);
and U22128 (N_22128,N_21130,N_21907);
nand U22129 (N_22129,N_21643,N_20200);
nand U22130 (N_22130,N_21768,N_20171);
and U22131 (N_22131,N_21727,N_20355);
xnor U22132 (N_22132,N_20845,N_20002);
nor U22133 (N_22133,N_20361,N_21057);
or U22134 (N_22134,N_21139,N_21950);
or U22135 (N_22135,N_21195,N_21162);
nor U22136 (N_22136,N_21761,N_20203);
xor U22137 (N_22137,N_21006,N_20566);
nand U22138 (N_22138,N_20039,N_20666);
nand U22139 (N_22139,N_20841,N_21773);
nand U22140 (N_22140,N_20584,N_20108);
nor U22141 (N_22141,N_20553,N_21576);
nand U22142 (N_22142,N_21401,N_20569);
nand U22143 (N_22143,N_20115,N_20508);
nand U22144 (N_22144,N_21902,N_20824);
and U22145 (N_22145,N_20934,N_21734);
or U22146 (N_22146,N_21547,N_20139);
or U22147 (N_22147,N_20515,N_21362);
and U22148 (N_22148,N_20909,N_20899);
and U22149 (N_22149,N_21770,N_20440);
and U22150 (N_22150,N_20919,N_21921);
nand U22151 (N_22151,N_21037,N_20859);
nand U22152 (N_22152,N_21873,N_21224);
nor U22153 (N_22153,N_20759,N_21716);
nor U22154 (N_22154,N_20292,N_20090);
xor U22155 (N_22155,N_21912,N_20195);
xnor U22156 (N_22156,N_21028,N_20305);
nand U22157 (N_22157,N_21814,N_21914);
nor U22158 (N_22158,N_21254,N_20518);
or U22159 (N_22159,N_20873,N_21359);
nor U22160 (N_22160,N_21939,N_20877);
xor U22161 (N_22161,N_21244,N_21194);
or U22162 (N_22162,N_20910,N_20343);
xnor U22163 (N_22163,N_20250,N_21702);
or U22164 (N_22164,N_21377,N_20949);
nand U22165 (N_22165,N_21097,N_20582);
nand U22166 (N_22166,N_21157,N_21563);
nand U22167 (N_22167,N_20764,N_20176);
nand U22168 (N_22168,N_20756,N_21856);
nand U22169 (N_22169,N_20232,N_21343);
and U22170 (N_22170,N_21542,N_20332);
nand U22171 (N_22171,N_20238,N_21403);
and U22172 (N_22172,N_20983,N_20952);
or U22173 (N_22173,N_21992,N_20632);
and U22174 (N_22174,N_21477,N_21661);
and U22175 (N_22175,N_20868,N_20760);
nand U22176 (N_22176,N_21554,N_20657);
and U22177 (N_22177,N_21500,N_21303);
nor U22178 (N_22178,N_21174,N_21008);
xor U22179 (N_22179,N_21983,N_20604);
nor U22180 (N_22180,N_21475,N_20658);
and U22181 (N_22181,N_20559,N_20600);
or U22182 (N_22182,N_21192,N_21419);
nand U22183 (N_22183,N_20297,N_20168);
xnor U22184 (N_22184,N_21752,N_20838);
nand U22185 (N_22185,N_21741,N_21316);
nand U22186 (N_22186,N_20101,N_21147);
nor U22187 (N_22187,N_21135,N_21895);
and U22188 (N_22188,N_20863,N_20131);
nor U22189 (N_22189,N_20802,N_20057);
xnor U22190 (N_22190,N_20384,N_21806);
and U22191 (N_22191,N_21357,N_20097);
nand U22192 (N_22192,N_21229,N_21824);
nand U22193 (N_22193,N_21981,N_20700);
xnor U22194 (N_22194,N_20701,N_21793);
nand U22195 (N_22195,N_20901,N_20789);
nor U22196 (N_22196,N_20148,N_20284);
nor U22197 (N_22197,N_21830,N_20352);
and U22198 (N_22198,N_20184,N_20085);
xnor U22199 (N_22199,N_21242,N_20091);
xnor U22200 (N_22200,N_21168,N_21937);
xor U22201 (N_22201,N_21639,N_20425);
nand U22202 (N_22202,N_20791,N_21142);
nand U22203 (N_22203,N_21651,N_21670);
or U22204 (N_22204,N_21876,N_20905);
nand U22205 (N_22205,N_21987,N_21376);
nor U22206 (N_22206,N_20394,N_21423);
or U22207 (N_22207,N_20922,N_20496);
nand U22208 (N_22208,N_20483,N_20627);
xnor U22209 (N_22209,N_20086,N_21034);
nor U22210 (N_22210,N_20886,N_20603);
nand U22211 (N_22211,N_21906,N_20221);
or U22212 (N_22212,N_20572,N_20010);
or U22213 (N_22213,N_21282,N_20540);
nand U22214 (N_22214,N_21250,N_21739);
xor U22215 (N_22215,N_20782,N_21451);
and U22216 (N_22216,N_20466,N_20817);
and U22217 (N_22217,N_20706,N_21094);
xnor U22218 (N_22218,N_21213,N_21120);
or U22219 (N_22219,N_21589,N_20298);
xor U22220 (N_22220,N_20277,N_21759);
nor U22221 (N_22221,N_20235,N_21838);
xnor U22222 (N_22222,N_21997,N_20947);
and U22223 (N_22223,N_21946,N_21118);
xor U22224 (N_22224,N_20434,N_20299);
nor U22225 (N_22225,N_20437,N_21691);
xnor U22226 (N_22226,N_20286,N_21859);
nor U22227 (N_22227,N_20830,N_20071);
nand U22228 (N_22228,N_20984,N_21449);
and U22229 (N_22229,N_20662,N_20538);
xnor U22230 (N_22230,N_20275,N_20350);
nor U22231 (N_22231,N_20937,N_20892);
nor U22232 (N_22232,N_20376,N_20641);
and U22233 (N_22233,N_20507,N_20982);
nand U22234 (N_22234,N_20869,N_20147);
nor U22235 (N_22235,N_21688,N_21099);
or U22236 (N_22236,N_20180,N_20403);
nand U22237 (N_22237,N_21600,N_20767);
or U22238 (N_22238,N_20433,N_20094);
nor U22239 (N_22239,N_21565,N_20516);
nand U22240 (N_22240,N_20593,N_20233);
or U22241 (N_22241,N_21126,N_20194);
and U22242 (N_22242,N_21682,N_21267);
xor U22243 (N_22243,N_21301,N_21617);
and U22244 (N_22244,N_21999,N_20610);
nor U22245 (N_22245,N_20179,N_20401);
and U22246 (N_22246,N_20953,N_20251);
and U22247 (N_22247,N_20551,N_21948);
xnor U22248 (N_22248,N_21717,N_21172);
nand U22249 (N_22249,N_20771,N_21924);
nor U22250 (N_22250,N_21991,N_20109);
and U22251 (N_22251,N_21405,N_20575);
or U22252 (N_22252,N_21698,N_21144);
nor U22253 (N_22253,N_20279,N_21394);
nand U22254 (N_22254,N_21388,N_21979);
xnor U22255 (N_22255,N_20205,N_20311);
nand U22256 (N_22256,N_20143,N_20599);
and U22257 (N_22257,N_21803,N_21851);
nor U22258 (N_22258,N_20329,N_20678);
xnor U22259 (N_22259,N_21434,N_20028);
nor U22260 (N_22260,N_20545,N_20945);
and U22261 (N_22261,N_21146,N_21331);
xor U22262 (N_22262,N_20489,N_21882);
nor U22263 (N_22263,N_20754,N_20177);
nand U22264 (N_22264,N_21019,N_20254);
xor U22265 (N_22265,N_20182,N_21422);
or U22266 (N_22266,N_20749,N_20210);
nor U22267 (N_22267,N_21553,N_20363);
and U22268 (N_22268,N_21134,N_21543);
and U22269 (N_22269,N_20585,N_21075);
or U22270 (N_22270,N_20744,N_21925);
nor U22271 (N_22271,N_20819,N_20049);
nor U22272 (N_22272,N_20714,N_21597);
nand U22273 (N_22273,N_20734,N_21638);
xnor U22274 (N_22274,N_20081,N_21944);
or U22275 (N_22275,N_21472,N_20160);
nor U22276 (N_22276,N_20587,N_21725);
and U22277 (N_22277,N_21179,N_21742);
nor U22278 (N_22278,N_21230,N_21580);
nand U22279 (N_22279,N_21109,N_21257);
or U22280 (N_22280,N_21930,N_21679);
nor U22281 (N_22281,N_21392,N_21030);
and U22282 (N_22282,N_20225,N_20612);
or U22283 (N_22283,N_20067,N_21464);
or U22284 (N_22284,N_21762,N_21326);
nand U22285 (N_22285,N_21786,N_21193);
or U22286 (N_22286,N_21933,N_21497);
or U22287 (N_22287,N_20477,N_20698);
and U22288 (N_22288,N_20637,N_21033);
or U22289 (N_22289,N_21839,N_20301);
and U22290 (N_22290,N_21264,N_21096);
xnor U22291 (N_22291,N_20442,N_21103);
or U22292 (N_22292,N_20228,N_20047);
nand U22293 (N_22293,N_21707,N_21354);
nand U22294 (N_22294,N_20427,N_20943);
nor U22295 (N_22295,N_20867,N_20981);
xor U22296 (N_22296,N_21674,N_20274);
or U22297 (N_22297,N_20828,N_21511);
nand U22298 (N_22298,N_21374,N_21533);
nor U22299 (N_22299,N_20718,N_20539);
and U22300 (N_22300,N_20215,N_21916);
nand U22301 (N_22301,N_21754,N_20935);
and U22302 (N_22302,N_21031,N_21206);
nand U22303 (N_22303,N_21342,N_21684);
xor U22304 (N_22304,N_21239,N_20325);
and U22305 (N_22305,N_21957,N_21054);
or U22306 (N_22306,N_20890,N_20271);
nand U22307 (N_22307,N_20705,N_21410);
or U22308 (N_22308,N_20955,N_20809);
or U22309 (N_22309,N_20797,N_21785);
xnor U22310 (N_22310,N_21119,N_21585);
xor U22311 (N_22311,N_21274,N_21708);
nand U22312 (N_22312,N_20188,N_21582);
xor U22313 (N_22313,N_21678,N_20630);
and U22314 (N_22314,N_21366,N_20407);
or U22315 (N_22315,N_21515,N_20529);
nor U22316 (N_22316,N_21044,N_20330);
nand U22317 (N_22317,N_21211,N_21400);
and U22318 (N_22318,N_20327,N_21417);
nor U22319 (N_22319,N_20884,N_20751);
nor U22320 (N_22320,N_20524,N_20907);
nand U22321 (N_22321,N_20080,N_20206);
nor U22322 (N_22322,N_21677,N_21635);
or U22323 (N_22323,N_21932,N_21631);
nand U22324 (N_22324,N_21781,N_21911);
nand U22325 (N_22325,N_21996,N_20422);
nand U22326 (N_22326,N_20055,N_21842);
and U22327 (N_22327,N_21623,N_20971);
xnor U22328 (N_22328,N_21323,N_21484);
xor U22329 (N_22329,N_20117,N_20370);
and U22330 (N_22330,N_20834,N_20999);
nor U22331 (N_22331,N_21909,N_20263);
nor U22332 (N_22332,N_20643,N_20416);
or U22333 (N_22333,N_20378,N_20940);
or U22334 (N_22334,N_20673,N_21976);
nor U22335 (N_22335,N_20283,N_21966);
or U22336 (N_22336,N_21985,N_20563);
and U22337 (N_22337,N_21436,N_20615);
xnor U22338 (N_22338,N_20898,N_20505);
xnor U22339 (N_22339,N_20391,N_21955);
nand U22340 (N_22340,N_20366,N_21117);
and U22341 (N_22341,N_20207,N_20805);
or U22342 (N_22342,N_20324,N_20969);
or U22343 (N_22343,N_20405,N_20462);
or U22344 (N_22344,N_21686,N_21514);
nor U22345 (N_22345,N_20519,N_20007);
xor U22346 (N_22346,N_21372,N_21021);
nor U22347 (N_22347,N_20239,N_21774);
and U22348 (N_22348,N_20722,N_21210);
and U22349 (N_22349,N_20320,N_20036);
or U22350 (N_22350,N_21358,N_20290);
or U22351 (N_22351,N_21270,N_21720);
and U22352 (N_22352,N_20045,N_20231);
nor U22353 (N_22353,N_21812,N_20111);
nand U22354 (N_22354,N_21149,N_20093);
xor U22355 (N_22355,N_21495,N_21779);
xnor U22356 (N_22356,N_20699,N_21942);
or U22357 (N_22357,N_21836,N_20491);
and U22358 (N_22358,N_21855,N_21947);
xor U22359 (N_22359,N_20793,N_20124);
and U22360 (N_22360,N_20762,N_21956);
xnor U22361 (N_22361,N_20758,N_20784);
or U22362 (N_22362,N_20060,N_21110);
nor U22363 (N_22363,N_20443,N_21186);
or U22364 (N_22364,N_21281,N_20591);
nor U22365 (N_22365,N_20107,N_21080);
nor U22366 (N_22366,N_21344,N_21023);
nand U22367 (N_22367,N_20608,N_21102);
xnor U22368 (N_22368,N_21593,N_21191);
or U22369 (N_22369,N_21381,N_21258);
nand U22370 (N_22370,N_20022,N_21225);
xnor U22371 (N_22371,N_21587,N_21507);
and U22372 (N_22372,N_21571,N_20133);
xnor U22373 (N_22373,N_21485,N_20216);
nand U22374 (N_22374,N_20880,N_20645);
xor U22375 (N_22375,N_21705,N_20114);
nor U22376 (N_22376,N_21628,N_21990);
nor U22377 (N_22377,N_20386,N_21675);
or U22378 (N_22378,N_20362,N_21747);
and U22379 (N_22379,N_20588,N_20163);
nor U22380 (N_22380,N_20721,N_21444);
or U22381 (N_22381,N_20488,N_20684);
and U22382 (N_22382,N_20775,N_20810);
nand U22383 (N_22383,N_21592,N_20796);
and U22384 (N_22384,N_21847,N_21443);
nor U22385 (N_22385,N_21393,N_21518);
nand U22386 (N_22386,N_21818,N_20913);
and U22387 (N_22387,N_20451,N_21821);
and U22388 (N_22388,N_21208,N_21633);
and U22389 (N_22389,N_21840,N_21098);
nand U22390 (N_22390,N_20837,N_20492);
nand U22391 (N_22391,N_20471,N_20304);
nand U22392 (N_22392,N_20786,N_20211);
and U22393 (N_22393,N_20356,N_20478);
or U22394 (N_22394,N_20513,N_20219);
xnor U22395 (N_22395,N_20638,N_20341);
nand U22396 (N_22396,N_20865,N_20322);
nor U22397 (N_22397,N_20268,N_20103);
and U22398 (N_22398,N_20564,N_20008);
nand U22399 (N_22399,N_20253,N_20654);
or U22400 (N_22400,N_20815,N_21649);
or U22401 (N_22401,N_20393,N_20503);
or U22402 (N_22402,N_20962,N_21746);
nor U22403 (N_22403,N_21433,N_21159);
and U22404 (N_22404,N_20397,N_20723);
and U22405 (N_22405,N_21487,N_21308);
nor U22406 (N_22406,N_21435,N_20289);
and U22407 (N_22407,N_21161,N_20647);
nand U22408 (N_22408,N_21993,N_21370);
nand U22409 (N_22409,N_20006,N_20601);
or U22410 (N_22410,N_21878,N_21396);
xnor U22411 (N_22411,N_20270,N_21085);
xor U22412 (N_22412,N_20533,N_20162);
and U22413 (N_22413,N_20135,N_20994);
nor U22414 (N_22414,N_21414,N_21945);
nand U22415 (N_22415,N_21462,N_20560);
or U22416 (N_22416,N_20512,N_21823);
xnor U22417 (N_22417,N_20453,N_20926);
xor U22418 (N_22418,N_20522,N_21466);
or U22419 (N_22419,N_20025,N_21799);
nor U22420 (N_22420,N_20476,N_21629);
or U22421 (N_22421,N_20129,N_21153);
nor U22422 (N_22422,N_20346,N_21750);
and U22423 (N_22423,N_21671,N_20506);
or U22424 (N_22424,N_20713,N_20765);
nand U22425 (N_22425,N_21700,N_20291);
and U22426 (N_22426,N_20063,N_21090);
nand U22427 (N_22427,N_21897,N_20596);
and U22428 (N_22428,N_20302,N_21079);
xnor U22429 (N_22429,N_21486,N_20340);
and U22430 (N_22430,N_20318,N_21035);
and U22431 (N_22431,N_20382,N_20475);
nand U22432 (N_22432,N_20928,N_21969);
and U22433 (N_22433,N_21805,N_20455);
nor U22434 (N_22434,N_20446,N_21205);
xor U22435 (N_22435,N_21041,N_21900);
nor U22436 (N_22436,N_21478,N_21527);
nand U22437 (N_22437,N_20747,N_20121);
nand U22438 (N_22438,N_21364,N_20020);
nand U22439 (N_22439,N_21673,N_20636);
xnor U22440 (N_22440,N_20237,N_21003);
nand U22441 (N_22441,N_20255,N_20487);
nor U22442 (N_22442,N_21634,N_20799);
and U22443 (N_22443,N_20681,N_21846);
xor U22444 (N_22444,N_20853,N_20167);
or U22445 (N_22445,N_20465,N_20697);
nand U22446 (N_22446,N_20653,N_21397);
nand U22447 (N_22447,N_20042,N_21577);
and U22448 (N_22448,N_21207,N_20883);
nand U22449 (N_22449,N_20313,N_21782);
xor U22450 (N_22450,N_20198,N_20183);
xor U22451 (N_22451,N_21726,N_21284);
nand U22452 (N_22452,N_20383,N_21885);
or U22453 (N_22453,N_21304,N_20164);
nor U22454 (N_22454,N_21442,N_21963);
xnor U22455 (N_22455,N_21356,N_21769);
nor U22456 (N_22456,N_20688,N_21062);
and U22457 (N_22457,N_20494,N_21913);
or U22458 (N_22458,N_20474,N_20616);
nor U22459 (N_22459,N_20558,N_21169);
nor U22460 (N_22460,N_20421,N_21681);
xor U22461 (N_22461,N_20939,N_20482);
nor U22462 (N_22462,N_20264,N_21567);
nor U22463 (N_22463,N_20294,N_20613);
or U22464 (N_22464,N_20776,N_20504);
nor U22465 (N_22465,N_20938,N_20151);
or U22466 (N_22466,N_20709,N_20046);
nand U22467 (N_22467,N_20191,N_21181);
or U22468 (N_22468,N_21875,N_21668);
xnor U22469 (N_22469,N_21710,N_21133);
nor U22470 (N_22470,N_20881,N_20261);
nor U22471 (N_22471,N_21073,N_21415);
nand U22472 (N_22472,N_21534,N_20061);
or U22473 (N_22473,N_20521,N_21457);
nand U22474 (N_22474,N_21263,N_21501);
or U22475 (N_22475,N_21887,N_21378);
nor U22476 (N_22476,N_20336,N_20523);
and U22477 (N_22477,N_21862,N_21584);
nor U22478 (N_22478,N_21285,N_21190);
xnor U22479 (N_22479,N_20078,N_20084);
and U22480 (N_22480,N_21893,N_21491);
xnor U22481 (N_22481,N_20448,N_21908);
xnor U22482 (N_22482,N_21375,N_21641);
nand U22483 (N_22483,N_21266,N_21857);
xnor U22484 (N_22484,N_21586,N_20932);
xor U22485 (N_22485,N_21615,N_21596);
nor U22486 (N_22486,N_21346,N_21662);
or U22487 (N_22487,N_20400,N_20464);
or U22488 (N_22488,N_20024,N_21813);
xnor U22489 (N_22489,N_20976,N_20753);
and U22490 (N_22490,N_20497,N_21940);
xor U22491 (N_22491,N_21771,N_20068);
xnor U22492 (N_22492,N_20725,N_20743);
nand U22493 (N_22493,N_20511,N_20349);
nor U22494 (N_22494,N_21919,N_21347);
xor U22495 (N_22495,N_21299,N_21171);
and U22496 (N_22496,N_21384,N_20650);
nand U22497 (N_22497,N_20611,N_20348);
and U22498 (N_22498,N_21305,N_21986);
or U22499 (N_22499,N_20029,N_20429);
nand U22500 (N_22500,N_21063,N_20833);
nand U22501 (N_22501,N_20037,N_21872);
xnor U22502 (N_22502,N_21792,N_20306);
and U22503 (N_22503,N_20894,N_21780);
and U22504 (N_22504,N_21982,N_21998);
and U22505 (N_22505,N_20856,N_21703);
nor U22506 (N_22506,N_20169,N_21217);
xor U22507 (N_22507,N_21917,N_20328);
or U22508 (N_22508,N_20671,N_20963);
nor U22509 (N_22509,N_21516,N_21201);
nand U22510 (N_22510,N_21049,N_21772);
nand U22511 (N_22511,N_20402,N_21595);
and U22512 (N_22512,N_21055,N_21604);
nor U22513 (N_22513,N_21260,N_21470);
and U22514 (N_22514,N_20739,N_21245);
nand U22515 (N_22515,N_20965,N_20457);
xnor U22516 (N_22516,N_20674,N_20931);
xor U22517 (N_22517,N_20871,N_21047);
xnor U22518 (N_22518,N_20321,N_21233);
xor U22519 (N_22519,N_21431,N_21758);
nor U22520 (N_22520,N_21825,N_20447);
and U22521 (N_22521,N_21496,N_21606);
or U22522 (N_22522,N_20142,N_21029);
nor U22523 (N_22523,N_21588,N_21454);
nor U22524 (N_22524,N_21611,N_21014);
or U22525 (N_22525,N_21361,N_20351);
or U22526 (N_22526,N_20537,N_20096);
nand U22527 (N_22527,N_20490,N_20532);
and U22528 (N_22528,N_20738,N_21829);
nor U22529 (N_22529,N_20732,N_20314);
xnor U22530 (N_22530,N_20379,N_21790);
or U22531 (N_22531,N_20574,N_21317);
xor U22532 (N_22532,N_21398,N_21077);
or U22533 (N_22533,N_21699,N_21418);
xnor U22534 (N_22534,N_20549,N_21329);
and U22535 (N_22535,N_21791,N_21420);
nand U22536 (N_22536,N_20594,N_21915);
xor U22537 (N_22537,N_20347,N_21340);
nor U22538 (N_22538,N_20223,N_20048);
or U22539 (N_22539,N_20175,N_21520);
nor U22540 (N_22540,N_21574,N_20849);
xor U22541 (N_22541,N_20552,N_20531);
or U22542 (N_22542,N_21952,N_21632);
and U22543 (N_22543,N_21901,N_20141);
nand U22544 (N_22544,N_20399,N_21801);
or U22545 (N_22545,N_21390,N_20083);
nor U22546 (N_22546,N_20074,N_20667);
nor U22547 (N_22547,N_21072,N_21043);
and U22548 (N_22548,N_21570,N_21974);
or U22549 (N_22549,N_20988,N_21938);
and U22550 (N_22550,N_20668,N_21541);
nor U22551 (N_22551,N_21177,N_21881);
and U22552 (N_22552,N_21411,N_21517);
xnor U22553 (N_22553,N_21749,N_20916);
or U22554 (N_22554,N_21984,N_21714);
or U22555 (N_22555,N_20929,N_20509);
nand U22556 (N_22556,N_20648,N_20902);
and U22557 (N_22557,N_20064,N_20573);
and U22558 (N_22558,N_21241,N_20419);
or U22559 (N_22559,N_20742,N_20345);
xor U22560 (N_22560,N_21800,N_21557);
and U22561 (N_22561,N_20546,N_21572);
nor U22562 (N_22562,N_20213,N_21788);
or U22563 (N_22563,N_21558,N_20229);
and U22564 (N_22564,N_21655,N_21598);
nand U22565 (N_22565,N_21624,N_20125);
nand U22566 (N_22566,N_21463,N_21763);
nand U22567 (N_22567,N_21721,N_21100);
nor U22568 (N_22568,N_21278,N_21988);
or U22569 (N_22569,N_20498,N_20252);
or U22570 (N_22570,N_21735,N_21332);
nor U22571 (N_22571,N_20486,N_20780);
nor U22572 (N_22572,N_21091,N_20209);
xnor U22573 (N_22573,N_20197,N_20035);
xor U22574 (N_22574,N_20385,N_21568);
and U22575 (N_22575,N_20220,N_21636);
nor U22576 (N_22576,N_21197,N_20374);
and U22577 (N_22577,N_20053,N_20159);
nor U22578 (N_22578,N_21599,N_20050);
and U22579 (N_22579,N_20745,N_21868);
nor U22580 (N_22580,N_20906,N_21215);
and U22581 (N_22581,N_21283,N_21170);
and U22582 (N_22582,N_20665,N_20821);
nand U22583 (N_22583,N_21870,N_21505);
nor U22584 (N_22584,N_21499,N_20772);
xor U22585 (N_22585,N_20077,N_20763);
or U22586 (N_22586,N_21645,N_20707);
xnor U22587 (N_22587,N_20390,N_21711);
xor U22588 (N_22588,N_21059,N_20319);
or U22589 (N_22589,N_21022,N_20550);
nand U22590 (N_22590,N_20598,N_21508);
or U22591 (N_22591,N_21719,N_20100);
xor U22592 (N_22592,N_21184,N_20280);
and U22593 (N_22593,N_21083,N_20960);
xnor U22594 (N_22594,N_21148,N_21368);
xnor U22595 (N_22595,N_21832,N_20583);
and U22596 (N_22596,N_20079,N_21355);
nand U22597 (N_22597,N_21494,N_21863);
xor U22598 (N_22598,N_20779,N_20415);
or U22599 (N_22599,N_20165,N_21407);
and U22600 (N_22600,N_21865,N_21256);
nand U22601 (N_22601,N_21776,N_21605);
xor U22602 (N_22602,N_21523,N_21539);
and U22603 (N_22603,N_20561,N_20189);
and U22604 (N_22604,N_20034,N_21053);
or U22605 (N_22605,N_20663,N_21271);
nor U22606 (N_22606,N_21069,N_21469);
nor U22607 (N_22607,N_20534,N_20851);
xnor U22608 (N_22608,N_21765,N_20387);
nor U22609 (N_22609,N_21045,N_20832);
and U22610 (N_22610,N_20891,N_20012);
and U22611 (N_22611,N_21248,N_20282);
or U22612 (N_22612,N_21559,N_21816);
nor U22613 (N_22613,N_20411,N_21756);
and U22614 (N_22614,N_20003,N_21656);
xnor U22615 (N_22615,N_20438,N_21307);
or U22616 (N_22616,N_21124,N_20735);
nand U22617 (N_22617,N_21715,N_20624);
and U22618 (N_22618,N_20740,N_21659);
nand U22619 (N_22619,N_21082,N_20526);
nand U22620 (N_22620,N_20556,N_20839);
xor U22621 (N_22621,N_20278,N_21802);
or U22622 (N_22622,N_21723,N_21748);
nand U22623 (N_22623,N_20472,N_20956);
nor U22624 (N_22624,N_20652,N_20857);
or U22625 (N_22625,N_20847,N_20954);
xnor U22626 (N_22626,N_21445,N_21328);
and U22627 (N_22627,N_21432,N_20018);
xnor U22628 (N_22628,N_21005,N_20412);
or U22629 (N_22629,N_20011,N_21989);
or U22630 (N_22630,N_21618,N_21777);
or U22631 (N_22631,N_20882,N_20288);
nor U22632 (N_22632,N_20112,N_20146);
xnor U22633 (N_22633,N_20145,N_21828);
or U22634 (N_22634,N_20398,N_20651);
and U22635 (N_22635,N_21809,N_21287);
nor U22636 (N_22636,N_20501,N_20661);
xor U22637 (N_22637,N_21941,N_21864);
and U22638 (N_22638,N_21373,N_21578);
xor U22639 (N_22639,N_20536,N_21273);
nor U22640 (N_22640,N_20911,N_20995);
nor U22641 (N_22641,N_21877,N_21488);
nand U22642 (N_22642,N_20243,N_20755);
nor U22643 (N_22643,N_21789,N_20944);
and U22644 (N_22644,N_20731,N_21018);
and U22645 (N_22645,N_20256,N_20752);
nor U22646 (N_22646,N_21132,N_20975);
nand U22647 (N_22647,N_20941,N_21448);
or U22648 (N_22648,N_20373,N_21440);
xor U22649 (N_22649,N_20908,N_20964);
nor U22650 (N_22650,N_20682,N_21010);
nand U22651 (N_22651,N_20800,N_21081);
nor U22652 (N_22652,N_20333,N_20691);
xor U22653 (N_22653,N_21669,N_21784);
nand U22654 (N_22654,N_21614,N_20541);
or U22655 (N_22655,N_21319,N_20009);
nand U22656 (N_22656,N_21404,N_20043);
or U22657 (N_22657,N_20785,N_20470);
or U22658 (N_22658,N_21764,N_21613);
nor U22659 (N_22659,N_20089,N_21158);
nand U22660 (N_22660,N_21167,N_20156);
and U22661 (N_22661,N_20242,N_21819);
nand U22662 (N_22662,N_21122,N_21498);
and U22663 (N_22663,N_20158,N_20001);
or U22664 (N_22664,N_21871,N_20520);
and U22665 (N_22665,N_21231,N_20269);
and U22666 (N_22666,N_20309,N_20748);
and U22667 (N_22667,N_21712,N_21713);
nand U22668 (N_22668,N_21426,N_21074);
nand U22669 (N_22669,N_21513,N_20737);
xnor U22670 (N_22670,N_20190,N_20172);
xnor U22671 (N_22671,N_21648,N_20017);
nand U22672 (N_22672,N_21473,N_21218);
and U22673 (N_22673,N_21198,N_20578);
or U22674 (N_22674,N_21324,N_21280);
or U22675 (N_22675,N_20991,N_20459);
and U22676 (N_22676,N_20750,N_21039);
nand U22677 (N_22677,N_21934,N_20912);
or U22678 (N_22678,N_20485,N_21402);
or U22679 (N_22679,N_21371,N_21731);
nor U22680 (N_22680,N_20375,N_20149);
nand U22681 (N_22681,N_20484,N_20979);
nor U22682 (N_22682,N_21894,N_20669);
xor U22683 (N_22683,N_21874,N_20717);
nand U22684 (N_22684,N_21642,N_20367);
nor U22685 (N_22685,N_20528,N_21951);
nor U22686 (N_22686,N_21536,N_21549);
nor U22687 (N_22687,N_21918,N_21637);
nand U22688 (N_22688,N_20136,N_20814);
nor U22689 (N_22689,N_21692,N_20977);
and U22690 (N_22690,N_20631,N_21196);
xor U22691 (N_22691,N_20917,N_21430);
and U22692 (N_22692,N_21808,N_21143);
nor U22693 (N_22693,N_21564,N_21521);
or U22694 (N_22694,N_21603,N_20082);
nor U22695 (N_22695,N_20850,N_20804);
and U22696 (N_22696,N_21630,N_20070);
and U22697 (N_22697,N_20344,N_20510);
nand U22698 (N_22698,N_20676,N_21095);
and U22699 (N_22699,N_20059,N_21105);
or U22700 (N_22700,N_21212,N_21412);
and U22701 (N_22701,N_21204,N_20609);
xor U22702 (N_22702,N_21330,N_21923);
nand U22703 (N_22703,N_20460,N_20122);
xnor U22704 (N_22704,N_20054,N_21227);
nand U22705 (N_22705,N_21108,N_20371);
or U22706 (N_22706,N_20224,N_21078);
nand U22707 (N_22707,N_20595,N_20741);
nand U22708 (N_22708,N_20076,N_20248);
nand U22709 (N_22709,N_21620,N_21309);
nor U22710 (N_22710,N_21658,N_21156);
nand U22711 (N_22711,N_20293,N_21476);
or U22712 (N_22712,N_21509,N_20826);
xnor U22713 (N_22713,N_21237,N_20757);
or U22714 (N_22714,N_21187,N_20015);
and U22715 (N_22715,N_20123,N_20986);
nand U22716 (N_22716,N_21695,N_21844);
xor U22717 (N_22717,N_20715,N_20946);
or U22718 (N_22718,N_20670,N_20924);
and U22719 (N_22719,N_20044,N_21693);
nand U22720 (N_22720,N_20920,N_21209);
and U22721 (N_22721,N_21943,N_20088);
xnor U22722 (N_22722,N_21960,N_21164);
xor U22723 (N_22723,N_21173,N_21456);
and U22724 (N_22724,N_21089,N_20778);
xnor U22725 (N_22725,N_21428,N_21116);
nand U22726 (N_22726,N_20128,N_20110);
or U22727 (N_22727,N_20406,N_21743);
or U22728 (N_22728,N_21383,N_21798);
or U22729 (N_22729,N_20727,N_21544);
or U22730 (N_22730,N_20281,N_21540);
nand U22731 (N_22731,N_21616,N_21408);
or U22732 (N_22732,N_20711,N_20296);
and U22733 (N_22733,N_20454,N_20888);
or U22734 (N_22734,N_21766,N_20260);
nand U22735 (N_22735,N_21612,N_20428);
nand U22736 (N_22736,N_20418,N_21778);
or U22737 (N_22737,N_20987,N_20703);
and U22738 (N_22738,N_20996,N_20062);
and U22739 (N_22739,N_21060,N_21140);
nand U22740 (N_22740,N_21718,N_20170);
nand U22741 (N_22741,N_20377,N_20087);
nor U22742 (N_22742,N_20557,N_20858);
nand U22743 (N_22743,N_21811,N_20245);
nor U22744 (N_22744,N_21036,N_20618);
or U22745 (N_22745,N_21203,N_20202);
and U22746 (N_22746,N_20808,N_21017);
nand U22747 (N_22747,N_21234,N_20597);
xor U22748 (N_22748,N_20204,N_20855);
nor U22749 (N_22749,N_20530,N_21826);
xnor U22750 (N_22750,N_20423,N_21573);
or U22751 (N_22751,N_21660,N_21740);
and U22752 (N_22752,N_21138,N_21064);
nor U22753 (N_22753,N_21537,N_21787);
nand U22754 (N_22754,N_21076,N_21722);
nand U22755 (N_22755,N_21471,N_21728);
or U22756 (N_22756,N_21896,N_20985);
and U22757 (N_22757,N_20449,N_21000);
and U22758 (N_22758,N_20310,N_21155);
nor U22759 (N_22759,N_20246,N_21382);
nand U22760 (N_22760,N_20031,N_20212);
or U22761 (N_22761,N_21551,N_20033);
and U22762 (N_22762,N_20761,N_20456);
nand U22763 (N_22763,N_20262,N_20696);
and U22764 (N_22764,N_20130,N_20276);
nand U22765 (N_22765,N_20392,N_21672);
or U22766 (N_22766,N_20013,N_21293);
and U22767 (N_22767,N_20467,N_21199);
and U22768 (N_22768,N_21232,N_21046);
or U22769 (N_22769,N_20380,N_20998);
xnor U22770 (N_22770,N_20660,N_20607);
and U22771 (N_22771,N_21333,N_21510);
and U22772 (N_22772,N_21854,N_20535);
xor U22773 (N_22773,N_21222,N_20978);
nor U22774 (N_22774,N_20181,N_21867);
nor U22775 (N_22775,N_20113,N_21341);
nand U22776 (N_22776,N_21680,N_20914);
or U22777 (N_22777,N_21446,N_20577);
and U22778 (N_22778,N_21964,N_21627);
xor U22779 (N_22779,N_21350,N_20625);
and U22780 (N_22780,N_21709,N_20617);
nor U22781 (N_22781,N_21704,N_20589);
nand U22782 (N_22782,N_20925,N_20369);
xnor U22783 (N_22783,N_20683,N_21845);
and U22784 (N_22784,N_20052,N_20357);
and U22785 (N_22785,N_21255,N_21978);
xnor U22786 (N_22786,N_21538,N_20968);
nand U22787 (N_22787,N_21503,N_20730);
and U22788 (N_22788,N_21111,N_21467);
nand U22789 (N_22789,N_21929,N_21038);
nand U22790 (N_22790,N_21861,N_21706);
nor U22791 (N_22791,N_20746,N_20623);
xnor U22792 (N_22792,N_21954,N_20915);
nor U22793 (N_22793,N_20127,N_21736);
and U22794 (N_22794,N_20138,N_20783);
and U22795 (N_22795,N_21276,N_21827);
nand U22796 (N_22796,N_21602,N_21837);
nor U22797 (N_22797,N_21265,N_21020);
or U22798 (N_22798,N_20639,N_21310);
and U22799 (N_22799,N_20436,N_20525);
nor U22800 (N_22800,N_21395,N_20770);
xor U22801 (N_22801,N_20635,N_20896);
or U22802 (N_22802,N_20622,N_21252);
and U22803 (N_22803,N_21188,N_21898);
nor U22804 (N_22804,N_21524,N_20173);
nand U22805 (N_22805,N_21880,N_20816);
and U22806 (N_22806,N_20201,N_21279);
and U22807 (N_22807,N_21367,N_21216);
nor U22808 (N_22808,N_20900,N_21345);
nor U22809 (N_22809,N_21975,N_21115);
xnor U22810 (N_22810,N_20222,N_21755);
nand U22811 (N_22811,N_20285,N_21581);
or U22812 (N_22812,N_21848,N_21061);
and U22813 (N_22813,N_21141,N_20021);
xnor U22814 (N_22814,N_20140,N_20199);
nor U22815 (N_22815,N_20642,N_20693);
xor U22816 (N_22816,N_20921,N_21512);
and U22817 (N_22817,N_21458,N_20527);
nand U22818 (N_22818,N_21977,N_20961);
and U22819 (N_22819,N_21737,N_21249);
or U22820 (N_22820,N_21452,N_21653);
and U22821 (N_22821,N_21300,N_20493);
and U22822 (N_22822,N_21272,N_20214);
xnor U22823 (N_22823,N_21683,N_21106);
and U22824 (N_22824,N_21236,N_20287);
nand U22825 (N_22825,N_21334,N_21321);
xnor U22826 (N_22826,N_21127,N_20404);
nand U22827 (N_22827,N_20646,N_20801);
or U22828 (N_22828,N_20846,N_21447);
or U22829 (N_22829,N_21238,N_21502);
nand U22830 (N_22830,N_21506,N_21640);
or U22831 (N_22831,N_21569,N_21690);
nand U22832 (N_22832,N_21406,N_21666);
or U22833 (N_22833,N_21609,N_21327);
or U22834 (N_22834,N_21590,N_21525);
xor U22835 (N_22835,N_20095,N_21489);
and U22836 (N_22836,N_21831,N_21011);
or U22837 (N_22837,N_20241,N_20134);
and U22838 (N_22838,N_20554,N_21729);
and U22839 (N_22839,N_20951,N_21399);
xnor U22840 (N_22840,N_21051,N_20058);
and U22841 (N_22841,N_20408,N_21980);
nand U22842 (N_22842,N_20562,N_21753);
nor U22843 (N_22843,N_20295,N_20997);
nand U22844 (N_22844,N_21730,N_21288);
xor U22845 (N_22845,N_21253,N_21626);
nand U22846 (N_22846,N_21654,N_21325);
or U22847 (N_22847,N_21949,N_21465);
nand U22848 (N_22848,N_21869,N_21292);
nand U22849 (N_22849,N_21490,N_21899);
and U22850 (N_22850,N_21810,N_20818);
and U22851 (N_22851,N_20353,N_20244);
and U22852 (N_22852,N_21657,N_20092);
nand U22853 (N_22853,N_20368,N_21504);
nand U22854 (N_22854,N_20234,N_20118);
nand U22855 (N_22855,N_20580,N_20686);
nand U22856 (N_22856,N_20973,N_20019);
xor U22857 (N_22857,N_20473,N_21262);
nand U22858 (N_22858,N_21125,N_21421);
nand U22859 (N_22859,N_20315,N_21360);
nor U22860 (N_22860,N_20056,N_21528);
nor U22861 (N_22861,N_21531,N_20132);
xor U22862 (N_22862,N_20848,N_21687);
or U22863 (N_22863,N_21409,N_20372);
nand U22864 (N_22864,N_21114,N_21450);
nand U22865 (N_22865,N_21566,N_20852);
xor U22866 (N_22866,N_21667,N_20619);
nor U22867 (N_22867,N_21048,N_20360);
and U22868 (N_22868,N_21289,N_21313);
xnor U22869 (N_22869,N_20861,N_21835);
or U22870 (N_22870,N_21696,N_21087);
and U22871 (N_22871,N_20777,N_21920);
nand U22872 (N_22872,N_21348,N_21349);
nand U22873 (N_22873,N_21092,N_21298);
and U22874 (N_22874,N_21228,N_21336);
nand U22875 (N_22875,N_20634,N_20144);
or U22876 (N_22876,N_20576,N_21351);
nor U22877 (N_22877,N_20414,N_20794);
nand U22878 (N_22878,N_21427,N_21387);
or U22879 (N_22879,N_20365,N_21416);
nor U22880 (N_22880,N_21965,N_20308);
and U22881 (N_22881,N_20236,N_21050);
and U22882 (N_22882,N_21971,N_21128);
xnor U22883 (N_22883,N_21369,N_21318);
xnor U22884 (N_22884,N_21219,N_21967);
xor U22885 (N_22885,N_21889,N_21807);
nand U22886 (N_22886,N_21104,N_21492);
xor U22887 (N_22887,N_21904,N_20174);
nand U22888 (N_22888,N_20933,N_20567);
or U22889 (N_22889,N_21002,N_21202);
nor U22890 (N_22890,N_20605,N_20904);
or U22891 (N_22891,N_20614,N_21154);
and U22892 (N_22892,N_20813,N_20602);
xnor U22893 (N_22893,N_21086,N_21032);
and U22894 (N_22894,N_21689,N_21646);
or U22895 (N_22895,N_20326,N_20409);
nand U22896 (N_22896,N_21815,N_21552);
and U22897 (N_22897,N_20677,N_21223);
nor U22898 (N_22898,N_20166,N_20481);
and U22899 (N_22899,N_20544,N_21015);
xor U22900 (N_22900,N_20267,N_21189);
xor U22901 (N_22901,N_21676,N_21066);
nor U22902 (N_22902,N_21121,N_20568);
and U22903 (N_22903,N_21200,N_20186);
nor U22904 (N_22904,N_21548,N_20463);
and U22905 (N_22905,N_20331,N_21936);
nand U22906 (N_22906,N_21275,N_21058);
or U22907 (N_22907,N_21145,N_20844);
nor U22908 (N_22908,N_20843,N_20358);
nor U22909 (N_22909,N_20766,N_20862);
nor U22910 (N_22910,N_20066,N_21583);
or U22911 (N_22911,N_21009,N_20026);
xnor U22912 (N_22912,N_21724,N_21259);
and U22913 (N_22913,N_20072,N_21591);
or U22914 (N_22914,N_20710,N_21461);
xnor U22915 (N_22915,N_21843,N_20137);
or U22916 (N_22916,N_21363,N_21858);
nor U22917 (N_22917,N_20980,N_21795);
xnor U22918 (N_22918,N_20208,N_20579);
nor U22919 (N_22919,N_21481,N_20970);
nand U22920 (N_22920,N_20413,N_20187);
nand U22921 (N_22921,N_20300,N_21312);
and U22922 (N_22922,N_20069,N_20629);
and U22923 (N_22923,N_21968,N_21460);
or U22924 (N_22924,N_20875,N_20272);
xnor U22925 (N_22925,N_20959,N_21176);
or U22926 (N_22926,N_20702,N_20099);
nand U22927 (N_22927,N_21302,N_20334);
or U22928 (N_22928,N_21007,N_20547);
or U22929 (N_22929,N_20265,N_20570);
nand U22930 (N_22930,N_20790,N_20153);
xor U22931 (N_22931,N_20792,N_20119);
xor U22932 (N_22932,N_21738,N_21745);
nor U22933 (N_22933,N_21277,N_20155);
xor U22934 (N_22934,N_20586,N_20720);
nand U22935 (N_22935,N_20468,N_20005);
nand U22936 (N_22936,N_20106,N_21664);
xnor U22937 (N_22937,N_21522,N_20590);
and U22938 (N_22938,N_20065,N_20923);
nor U22939 (N_22939,N_20499,N_20620);
or U22940 (N_22940,N_21468,N_21783);
and U22941 (N_22941,N_21953,N_20126);
xnor U22942 (N_22942,N_20389,N_20972);
and U22943 (N_22943,N_21841,N_20825);
and U22944 (N_22944,N_20967,N_21562);
and U22945 (N_22945,N_21291,N_21180);
nand U22946 (N_22946,N_21962,N_20469);
xor U22947 (N_22947,N_21647,N_21926);
or U22948 (N_22948,N_21439,N_20831);
and U22949 (N_22949,N_20116,N_21922);
nand U22950 (N_22950,N_20829,N_21151);
nor U22951 (N_22951,N_20708,N_20626);
or U22952 (N_22952,N_20424,N_21794);
or U22953 (N_22953,N_20014,N_21474);
xor U22954 (N_22954,N_21892,N_21137);
nor U22955 (N_22955,N_20957,N_20903);
or U22956 (N_22956,N_20461,N_21247);
nand U22957 (N_22957,N_21183,N_21339);
nor U22958 (N_22958,N_20023,N_21165);
or U22959 (N_22959,N_20240,N_21852);
and U22960 (N_22960,N_21070,N_20695);
nand U22961 (N_22961,N_21243,N_21973);
or U22962 (N_22962,N_20692,N_21931);
and U22963 (N_22963,N_20426,N_20897);
nor U22964 (N_22964,N_20543,N_20226);
nor U22965 (N_22965,N_20388,N_21694);
xnor U22966 (N_22966,N_20450,N_20359);
xnor U22967 (N_22967,N_21879,N_20004);
and U22968 (N_22968,N_20051,N_21024);
nor U22969 (N_22969,N_21429,N_20571);
xnor U22970 (N_22970,N_20565,N_20038);
nor U22971 (N_22971,N_20989,N_21886);
nand U22972 (N_22972,N_20217,N_21131);
xor U22973 (N_22973,N_20193,N_21268);
nand U22974 (N_22974,N_20431,N_20040);
and U22975 (N_22975,N_21888,N_21546);
xnor U22976 (N_22976,N_20430,N_21650);
nor U22977 (N_22977,N_21610,N_20823);
nand U22978 (N_22978,N_21820,N_20555);
or U22979 (N_22979,N_20712,N_21101);
nor U22980 (N_22980,N_21084,N_21459);
or U22981 (N_22981,N_21550,N_20273);
and U22982 (N_22982,N_21320,N_20150);
and U22983 (N_22983,N_20874,N_21261);
and U22984 (N_22984,N_21065,N_20230);
and U22985 (N_22985,N_20432,N_21927);
nand U22986 (N_22986,N_21337,N_21314);
or U22987 (N_22987,N_20812,N_20840);
nor U22988 (N_22988,N_21424,N_20769);
nor U22989 (N_22989,N_20303,N_21797);
nor U22990 (N_22990,N_20827,N_21560);
or U22991 (N_22991,N_21306,N_20152);
nor U22992 (N_22992,N_20649,N_20339);
nand U22993 (N_22993,N_20452,N_21286);
or U22994 (N_22994,N_21619,N_21482);
xnor U22995 (N_22995,N_20811,N_21112);
or U22996 (N_22996,N_20227,N_20396);
nor U22997 (N_22997,N_20803,N_20656);
and U22998 (N_22998,N_21379,N_20820);
or U22999 (N_22999,N_21214,N_20948);
and U23000 (N_23000,N_21571,N_21700);
nor U23001 (N_23001,N_20132,N_21799);
xnor U23002 (N_23002,N_20683,N_21618);
or U23003 (N_23003,N_20100,N_20137);
xnor U23004 (N_23004,N_20216,N_21548);
and U23005 (N_23005,N_20982,N_20369);
nand U23006 (N_23006,N_20777,N_21462);
nand U23007 (N_23007,N_21936,N_21179);
nor U23008 (N_23008,N_21554,N_21678);
or U23009 (N_23009,N_21493,N_21390);
nor U23010 (N_23010,N_21294,N_20381);
nand U23011 (N_23011,N_21329,N_20169);
or U23012 (N_23012,N_20455,N_21251);
nand U23013 (N_23013,N_21433,N_20738);
and U23014 (N_23014,N_20289,N_20777);
nand U23015 (N_23015,N_21560,N_21213);
xnor U23016 (N_23016,N_20051,N_20468);
nor U23017 (N_23017,N_21773,N_20213);
nor U23018 (N_23018,N_20482,N_21625);
nand U23019 (N_23019,N_20476,N_21809);
or U23020 (N_23020,N_21913,N_21781);
nor U23021 (N_23021,N_20068,N_20628);
xnor U23022 (N_23022,N_21743,N_21156);
nor U23023 (N_23023,N_21981,N_21232);
or U23024 (N_23024,N_20519,N_20241);
nor U23025 (N_23025,N_20571,N_20670);
xnor U23026 (N_23026,N_21377,N_20677);
nor U23027 (N_23027,N_20219,N_21542);
xor U23028 (N_23028,N_21996,N_20757);
xor U23029 (N_23029,N_20682,N_21080);
xnor U23030 (N_23030,N_20978,N_21208);
xor U23031 (N_23031,N_21063,N_21900);
xnor U23032 (N_23032,N_21265,N_20357);
xor U23033 (N_23033,N_20696,N_21927);
xnor U23034 (N_23034,N_20573,N_20952);
or U23035 (N_23035,N_21227,N_20891);
or U23036 (N_23036,N_21332,N_21448);
or U23037 (N_23037,N_21694,N_20881);
or U23038 (N_23038,N_21448,N_21123);
nand U23039 (N_23039,N_20571,N_20119);
nor U23040 (N_23040,N_20386,N_20825);
nor U23041 (N_23041,N_20845,N_21849);
and U23042 (N_23042,N_20805,N_20417);
nand U23043 (N_23043,N_21421,N_20778);
or U23044 (N_23044,N_20926,N_20104);
xnor U23045 (N_23045,N_20560,N_20648);
xnor U23046 (N_23046,N_21570,N_21855);
xor U23047 (N_23047,N_21163,N_21064);
and U23048 (N_23048,N_21059,N_20435);
nor U23049 (N_23049,N_20759,N_21620);
or U23050 (N_23050,N_20003,N_20822);
nand U23051 (N_23051,N_21515,N_20649);
nand U23052 (N_23052,N_21767,N_21549);
nand U23053 (N_23053,N_21095,N_20058);
nand U23054 (N_23054,N_20303,N_21946);
or U23055 (N_23055,N_20459,N_21722);
or U23056 (N_23056,N_20784,N_20048);
nand U23057 (N_23057,N_20430,N_21059);
nand U23058 (N_23058,N_20721,N_21872);
nand U23059 (N_23059,N_21829,N_21842);
nor U23060 (N_23060,N_21822,N_20989);
nand U23061 (N_23061,N_21271,N_21700);
nand U23062 (N_23062,N_20141,N_20420);
nor U23063 (N_23063,N_21778,N_20512);
and U23064 (N_23064,N_20553,N_20985);
nor U23065 (N_23065,N_21370,N_21764);
xnor U23066 (N_23066,N_21055,N_21632);
nand U23067 (N_23067,N_21464,N_20055);
or U23068 (N_23068,N_20841,N_21613);
or U23069 (N_23069,N_21042,N_20459);
and U23070 (N_23070,N_20711,N_20932);
nand U23071 (N_23071,N_21330,N_20955);
and U23072 (N_23072,N_20208,N_21012);
xnor U23073 (N_23073,N_20027,N_21670);
nor U23074 (N_23074,N_20552,N_21138);
nand U23075 (N_23075,N_21113,N_20635);
nand U23076 (N_23076,N_20864,N_20094);
nor U23077 (N_23077,N_21954,N_21014);
or U23078 (N_23078,N_21123,N_21200);
nand U23079 (N_23079,N_21261,N_20098);
and U23080 (N_23080,N_20068,N_21423);
and U23081 (N_23081,N_21878,N_21097);
nor U23082 (N_23082,N_21824,N_20098);
or U23083 (N_23083,N_21504,N_21520);
or U23084 (N_23084,N_20437,N_21910);
nor U23085 (N_23085,N_20279,N_21218);
nand U23086 (N_23086,N_21464,N_20512);
nand U23087 (N_23087,N_21409,N_20527);
and U23088 (N_23088,N_20676,N_21203);
xnor U23089 (N_23089,N_21912,N_20137);
nor U23090 (N_23090,N_20740,N_21306);
nor U23091 (N_23091,N_21756,N_20206);
nand U23092 (N_23092,N_20872,N_21726);
xnor U23093 (N_23093,N_21719,N_20722);
or U23094 (N_23094,N_21248,N_21105);
xor U23095 (N_23095,N_21705,N_21059);
nor U23096 (N_23096,N_21491,N_21910);
and U23097 (N_23097,N_20998,N_21488);
xor U23098 (N_23098,N_21222,N_20640);
nand U23099 (N_23099,N_20556,N_20238);
xor U23100 (N_23100,N_20620,N_21043);
nor U23101 (N_23101,N_21622,N_21052);
and U23102 (N_23102,N_20002,N_20079);
nor U23103 (N_23103,N_20407,N_21472);
nand U23104 (N_23104,N_21344,N_21021);
nor U23105 (N_23105,N_20331,N_21265);
xnor U23106 (N_23106,N_21744,N_20803);
nor U23107 (N_23107,N_21153,N_20952);
and U23108 (N_23108,N_20476,N_21091);
and U23109 (N_23109,N_20727,N_21155);
nand U23110 (N_23110,N_21974,N_21689);
nand U23111 (N_23111,N_20392,N_20632);
or U23112 (N_23112,N_21389,N_20922);
and U23113 (N_23113,N_21400,N_20246);
nor U23114 (N_23114,N_21886,N_21071);
nor U23115 (N_23115,N_21436,N_20464);
or U23116 (N_23116,N_21611,N_20863);
nand U23117 (N_23117,N_20999,N_20144);
xnor U23118 (N_23118,N_21393,N_21678);
nand U23119 (N_23119,N_20914,N_21155);
or U23120 (N_23120,N_21663,N_20959);
xor U23121 (N_23121,N_21652,N_21757);
xor U23122 (N_23122,N_20672,N_20937);
and U23123 (N_23123,N_20654,N_20729);
and U23124 (N_23124,N_20380,N_20400);
nor U23125 (N_23125,N_20192,N_21711);
nand U23126 (N_23126,N_20996,N_20920);
nand U23127 (N_23127,N_20831,N_21850);
or U23128 (N_23128,N_20190,N_21641);
nand U23129 (N_23129,N_21353,N_21589);
xor U23130 (N_23130,N_20582,N_20094);
or U23131 (N_23131,N_20942,N_21114);
xor U23132 (N_23132,N_20962,N_21365);
or U23133 (N_23133,N_21967,N_21049);
xor U23134 (N_23134,N_21681,N_20114);
xnor U23135 (N_23135,N_21931,N_20908);
or U23136 (N_23136,N_20678,N_20180);
and U23137 (N_23137,N_21276,N_21716);
nand U23138 (N_23138,N_20879,N_20878);
or U23139 (N_23139,N_21142,N_21393);
and U23140 (N_23140,N_20588,N_20922);
nor U23141 (N_23141,N_20962,N_20810);
xor U23142 (N_23142,N_21671,N_20381);
and U23143 (N_23143,N_20598,N_20762);
nor U23144 (N_23144,N_21336,N_21053);
xnor U23145 (N_23145,N_21577,N_20557);
xnor U23146 (N_23146,N_20280,N_20217);
nor U23147 (N_23147,N_21763,N_20686);
nor U23148 (N_23148,N_21358,N_21024);
xor U23149 (N_23149,N_20519,N_21441);
and U23150 (N_23150,N_21210,N_20420);
or U23151 (N_23151,N_20072,N_21708);
or U23152 (N_23152,N_21995,N_21744);
nor U23153 (N_23153,N_21962,N_20792);
nor U23154 (N_23154,N_21386,N_20533);
and U23155 (N_23155,N_20523,N_20670);
nand U23156 (N_23156,N_20682,N_20075);
nor U23157 (N_23157,N_21158,N_20027);
or U23158 (N_23158,N_20646,N_20763);
nor U23159 (N_23159,N_21261,N_20657);
or U23160 (N_23160,N_21284,N_20030);
nor U23161 (N_23161,N_21195,N_21047);
xor U23162 (N_23162,N_21779,N_21996);
or U23163 (N_23163,N_20460,N_21311);
or U23164 (N_23164,N_21363,N_21231);
nor U23165 (N_23165,N_20290,N_20631);
nand U23166 (N_23166,N_21784,N_21956);
nand U23167 (N_23167,N_20179,N_20303);
nor U23168 (N_23168,N_21095,N_21220);
nand U23169 (N_23169,N_20622,N_20102);
and U23170 (N_23170,N_20820,N_21244);
or U23171 (N_23171,N_21483,N_21235);
or U23172 (N_23172,N_21712,N_21998);
nor U23173 (N_23173,N_20232,N_21872);
or U23174 (N_23174,N_21924,N_21245);
or U23175 (N_23175,N_21450,N_20193);
xnor U23176 (N_23176,N_21069,N_20802);
and U23177 (N_23177,N_20930,N_20993);
or U23178 (N_23178,N_20216,N_21096);
and U23179 (N_23179,N_21149,N_21289);
or U23180 (N_23180,N_21011,N_21752);
and U23181 (N_23181,N_20906,N_20874);
nand U23182 (N_23182,N_20367,N_21655);
nand U23183 (N_23183,N_21274,N_20311);
nor U23184 (N_23184,N_21584,N_20264);
nor U23185 (N_23185,N_20076,N_21440);
xnor U23186 (N_23186,N_21186,N_20167);
nor U23187 (N_23187,N_21532,N_21699);
nor U23188 (N_23188,N_20949,N_20423);
xnor U23189 (N_23189,N_20940,N_20066);
and U23190 (N_23190,N_20203,N_21556);
or U23191 (N_23191,N_21468,N_20475);
or U23192 (N_23192,N_20721,N_20855);
or U23193 (N_23193,N_20811,N_21198);
nor U23194 (N_23194,N_20766,N_20871);
and U23195 (N_23195,N_20121,N_21878);
and U23196 (N_23196,N_20248,N_20247);
xnor U23197 (N_23197,N_21717,N_20639);
nand U23198 (N_23198,N_20001,N_20938);
nand U23199 (N_23199,N_21242,N_21548);
and U23200 (N_23200,N_21468,N_21316);
and U23201 (N_23201,N_20475,N_21134);
nand U23202 (N_23202,N_21262,N_21890);
nor U23203 (N_23203,N_21786,N_20177);
nand U23204 (N_23204,N_21280,N_20804);
nor U23205 (N_23205,N_21666,N_21099);
or U23206 (N_23206,N_21028,N_20529);
and U23207 (N_23207,N_21821,N_20231);
or U23208 (N_23208,N_21978,N_20520);
or U23209 (N_23209,N_21689,N_21692);
or U23210 (N_23210,N_21807,N_21938);
nand U23211 (N_23211,N_20083,N_21991);
or U23212 (N_23212,N_21832,N_21511);
nand U23213 (N_23213,N_20399,N_20368);
or U23214 (N_23214,N_21073,N_20184);
or U23215 (N_23215,N_20923,N_21285);
nor U23216 (N_23216,N_21684,N_20366);
or U23217 (N_23217,N_21664,N_20644);
nor U23218 (N_23218,N_20184,N_20377);
nand U23219 (N_23219,N_21908,N_20849);
nand U23220 (N_23220,N_20030,N_21623);
or U23221 (N_23221,N_21397,N_20617);
nor U23222 (N_23222,N_20489,N_21316);
nor U23223 (N_23223,N_20632,N_20770);
xnor U23224 (N_23224,N_20422,N_21693);
and U23225 (N_23225,N_20921,N_20799);
nor U23226 (N_23226,N_20088,N_21516);
nand U23227 (N_23227,N_20513,N_21236);
nand U23228 (N_23228,N_21535,N_20089);
nor U23229 (N_23229,N_21132,N_21722);
xnor U23230 (N_23230,N_20519,N_21065);
nor U23231 (N_23231,N_21708,N_20460);
nor U23232 (N_23232,N_20637,N_21521);
or U23233 (N_23233,N_21232,N_20162);
or U23234 (N_23234,N_20450,N_21468);
xor U23235 (N_23235,N_21582,N_20364);
or U23236 (N_23236,N_20771,N_20419);
nor U23237 (N_23237,N_20780,N_20933);
nor U23238 (N_23238,N_21334,N_20126);
nand U23239 (N_23239,N_21453,N_20749);
or U23240 (N_23240,N_21798,N_20392);
nor U23241 (N_23241,N_21491,N_21935);
xnor U23242 (N_23242,N_20770,N_20766);
and U23243 (N_23243,N_21576,N_21920);
and U23244 (N_23244,N_20689,N_20189);
nand U23245 (N_23245,N_20753,N_20735);
and U23246 (N_23246,N_21061,N_21085);
nand U23247 (N_23247,N_20692,N_21897);
nor U23248 (N_23248,N_21970,N_20987);
xor U23249 (N_23249,N_21648,N_20068);
nand U23250 (N_23250,N_21414,N_21083);
xnor U23251 (N_23251,N_21099,N_21682);
or U23252 (N_23252,N_20524,N_20291);
and U23253 (N_23253,N_20388,N_20851);
and U23254 (N_23254,N_21689,N_20581);
nor U23255 (N_23255,N_21083,N_20589);
nor U23256 (N_23256,N_21423,N_20975);
and U23257 (N_23257,N_20336,N_20451);
or U23258 (N_23258,N_21108,N_20466);
nor U23259 (N_23259,N_20742,N_21848);
and U23260 (N_23260,N_21281,N_21799);
and U23261 (N_23261,N_21266,N_21720);
nor U23262 (N_23262,N_20404,N_21961);
or U23263 (N_23263,N_20081,N_20749);
or U23264 (N_23264,N_20291,N_21799);
nand U23265 (N_23265,N_20391,N_21103);
xor U23266 (N_23266,N_20497,N_20041);
xnor U23267 (N_23267,N_21824,N_21156);
and U23268 (N_23268,N_21281,N_21546);
and U23269 (N_23269,N_21319,N_20854);
xor U23270 (N_23270,N_20356,N_21719);
or U23271 (N_23271,N_21811,N_21924);
and U23272 (N_23272,N_20624,N_20250);
nor U23273 (N_23273,N_20623,N_21943);
nand U23274 (N_23274,N_21128,N_20538);
or U23275 (N_23275,N_21412,N_20269);
and U23276 (N_23276,N_21347,N_20448);
xnor U23277 (N_23277,N_21142,N_20932);
nand U23278 (N_23278,N_21701,N_20742);
nor U23279 (N_23279,N_20163,N_20678);
nor U23280 (N_23280,N_20999,N_20802);
or U23281 (N_23281,N_20952,N_21529);
nor U23282 (N_23282,N_21345,N_21448);
or U23283 (N_23283,N_20072,N_21790);
xor U23284 (N_23284,N_21827,N_21013);
or U23285 (N_23285,N_20658,N_21442);
nand U23286 (N_23286,N_21947,N_21338);
nor U23287 (N_23287,N_21872,N_20154);
nand U23288 (N_23288,N_20310,N_21843);
nor U23289 (N_23289,N_20789,N_20923);
xor U23290 (N_23290,N_20651,N_21374);
nor U23291 (N_23291,N_21266,N_20685);
nand U23292 (N_23292,N_21843,N_20574);
nor U23293 (N_23293,N_20772,N_20580);
nor U23294 (N_23294,N_21541,N_21872);
or U23295 (N_23295,N_21872,N_20164);
xnor U23296 (N_23296,N_21122,N_20918);
nand U23297 (N_23297,N_20799,N_21843);
nand U23298 (N_23298,N_21155,N_21822);
or U23299 (N_23299,N_21462,N_20145);
xnor U23300 (N_23300,N_21469,N_20718);
xnor U23301 (N_23301,N_21358,N_20673);
and U23302 (N_23302,N_21123,N_21836);
nor U23303 (N_23303,N_20672,N_21591);
nand U23304 (N_23304,N_20589,N_20746);
xnor U23305 (N_23305,N_21821,N_21153);
xnor U23306 (N_23306,N_20957,N_20134);
nor U23307 (N_23307,N_20917,N_20207);
or U23308 (N_23308,N_21529,N_20313);
and U23309 (N_23309,N_20283,N_21123);
nand U23310 (N_23310,N_21537,N_20237);
nor U23311 (N_23311,N_21347,N_20231);
xnor U23312 (N_23312,N_20263,N_21275);
or U23313 (N_23313,N_20467,N_20098);
nor U23314 (N_23314,N_21292,N_21092);
or U23315 (N_23315,N_21367,N_20906);
and U23316 (N_23316,N_20948,N_20091);
nand U23317 (N_23317,N_20789,N_20559);
xnor U23318 (N_23318,N_20869,N_20007);
or U23319 (N_23319,N_20763,N_20533);
or U23320 (N_23320,N_21848,N_20549);
nor U23321 (N_23321,N_21010,N_21736);
and U23322 (N_23322,N_20804,N_20040);
nand U23323 (N_23323,N_20069,N_21200);
and U23324 (N_23324,N_20897,N_20072);
and U23325 (N_23325,N_21219,N_21080);
or U23326 (N_23326,N_20088,N_20923);
nor U23327 (N_23327,N_20232,N_20233);
nor U23328 (N_23328,N_21484,N_21932);
xor U23329 (N_23329,N_21818,N_21051);
or U23330 (N_23330,N_21716,N_21641);
nor U23331 (N_23331,N_21491,N_21567);
nand U23332 (N_23332,N_21221,N_21601);
nand U23333 (N_23333,N_21340,N_21984);
and U23334 (N_23334,N_21659,N_20728);
or U23335 (N_23335,N_20217,N_20771);
or U23336 (N_23336,N_20624,N_20112);
or U23337 (N_23337,N_21027,N_20415);
and U23338 (N_23338,N_20567,N_20675);
nand U23339 (N_23339,N_20414,N_20024);
nand U23340 (N_23340,N_20895,N_21185);
nor U23341 (N_23341,N_21392,N_20839);
xnor U23342 (N_23342,N_21857,N_20692);
nor U23343 (N_23343,N_20051,N_21288);
nand U23344 (N_23344,N_20214,N_20581);
xnor U23345 (N_23345,N_21181,N_21119);
xor U23346 (N_23346,N_21195,N_20743);
nor U23347 (N_23347,N_20626,N_21399);
xnor U23348 (N_23348,N_21110,N_21888);
and U23349 (N_23349,N_20973,N_21927);
and U23350 (N_23350,N_20184,N_21634);
or U23351 (N_23351,N_21168,N_20727);
xor U23352 (N_23352,N_21602,N_21524);
and U23353 (N_23353,N_21131,N_20939);
xnor U23354 (N_23354,N_21985,N_20495);
xor U23355 (N_23355,N_20850,N_20028);
nand U23356 (N_23356,N_20048,N_21114);
and U23357 (N_23357,N_21653,N_21632);
or U23358 (N_23358,N_21741,N_20949);
nand U23359 (N_23359,N_20130,N_20021);
or U23360 (N_23360,N_20474,N_21691);
nor U23361 (N_23361,N_21346,N_21044);
nor U23362 (N_23362,N_21478,N_20709);
nand U23363 (N_23363,N_20531,N_20321);
or U23364 (N_23364,N_21668,N_20550);
nand U23365 (N_23365,N_21564,N_21351);
and U23366 (N_23366,N_20584,N_21944);
nand U23367 (N_23367,N_21455,N_20523);
nand U23368 (N_23368,N_21731,N_20585);
and U23369 (N_23369,N_21356,N_20808);
nor U23370 (N_23370,N_21573,N_20190);
nor U23371 (N_23371,N_20021,N_20613);
nor U23372 (N_23372,N_21482,N_20945);
xor U23373 (N_23373,N_20874,N_21612);
xnor U23374 (N_23374,N_20778,N_21843);
and U23375 (N_23375,N_20119,N_20447);
nand U23376 (N_23376,N_21543,N_20483);
or U23377 (N_23377,N_20551,N_20053);
and U23378 (N_23378,N_21287,N_21901);
nand U23379 (N_23379,N_21072,N_20653);
nand U23380 (N_23380,N_21506,N_21656);
nor U23381 (N_23381,N_21242,N_21579);
xor U23382 (N_23382,N_20448,N_21618);
and U23383 (N_23383,N_20130,N_20011);
nor U23384 (N_23384,N_21374,N_21607);
and U23385 (N_23385,N_21718,N_21023);
or U23386 (N_23386,N_21933,N_20915);
xor U23387 (N_23387,N_21729,N_21358);
xnor U23388 (N_23388,N_20718,N_21869);
and U23389 (N_23389,N_20308,N_20899);
nor U23390 (N_23390,N_21831,N_20581);
xor U23391 (N_23391,N_20477,N_20691);
nand U23392 (N_23392,N_21307,N_21629);
or U23393 (N_23393,N_21847,N_21671);
nand U23394 (N_23394,N_21887,N_21999);
or U23395 (N_23395,N_21952,N_20932);
nor U23396 (N_23396,N_20141,N_20350);
xor U23397 (N_23397,N_20159,N_20174);
or U23398 (N_23398,N_20338,N_20365);
nor U23399 (N_23399,N_20889,N_20459);
and U23400 (N_23400,N_21934,N_20361);
and U23401 (N_23401,N_21332,N_21258);
xnor U23402 (N_23402,N_20990,N_21271);
and U23403 (N_23403,N_20827,N_21299);
xnor U23404 (N_23404,N_20315,N_20179);
and U23405 (N_23405,N_20265,N_21614);
xor U23406 (N_23406,N_20160,N_21993);
nor U23407 (N_23407,N_21918,N_21526);
nor U23408 (N_23408,N_21427,N_20703);
or U23409 (N_23409,N_20687,N_20549);
and U23410 (N_23410,N_21141,N_20363);
nand U23411 (N_23411,N_20643,N_21092);
nand U23412 (N_23412,N_21531,N_21189);
xor U23413 (N_23413,N_20861,N_21695);
nand U23414 (N_23414,N_21639,N_21392);
nand U23415 (N_23415,N_20964,N_21385);
nand U23416 (N_23416,N_21184,N_20429);
and U23417 (N_23417,N_21680,N_20899);
xnor U23418 (N_23418,N_20659,N_20217);
xor U23419 (N_23419,N_21404,N_20606);
or U23420 (N_23420,N_20625,N_20133);
and U23421 (N_23421,N_21611,N_21879);
and U23422 (N_23422,N_21155,N_21387);
and U23423 (N_23423,N_20180,N_21372);
xnor U23424 (N_23424,N_21631,N_21686);
nand U23425 (N_23425,N_21339,N_20038);
and U23426 (N_23426,N_20848,N_20601);
nand U23427 (N_23427,N_21755,N_21397);
nand U23428 (N_23428,N_21339,N_20799);
xor U23429 (N_23429,N_21887,N_21126);
nand U23430 (N_23430,N_20036,N_20374);
and U23431 (N_23431,N_20088,N_21599);
and U23432 (N_23432,N_21446,N_21982);
and U23433 (N_23433,N_21294,N_21375);
xor U23434 (N_23434,N_20140,N_20935);
nand U23435 (N_23435,N_21844,N_21170);
or U23436 (N_23436,N_21839,N_21547);
xnor U23437 (N_23437,N_21839,N_20818);
or U23438 (N_23438,N_20872,N_20429);
and U23439 (N_23439,N_21861,N_20947);
nor U23440 (N_23440,N_21206,N_21590);
nand U23441 (N_23441,N_20097,N_21897);
or U23442 (N_23442,N_20814,N_20072);
nor U23443 (N_23443,N_20271,N_21647);
and U23444 (N_23444,N_21649,N_21676);
xor U23445 (N_23445,N_21679,N_21289);
xor U23446 (N_23446,N_21965,N_20371);
nand U23447 (N_23447,N_20439,N_21947);
nor U23448 (N_23448,N_21307,N_21135);
and U23449 (N_23449,N_21765,N_20580);
nand U23450 (N_23450,N_21997,N_20849);
or U23451 (N_23451,N_20800,N_20736);
nor U23452 (N_23452,N_21042,N_20666);
nor U23453 (N_23453,N_20902,N_20016);
nand U23454 (N_23454,N_21401,N_21903);
or U23455 (N_23455,N_21590,N_21827);
nand U23456 (N_23456,N_20156,N_20370);
or U23457 (N_23457,N_21490,N_21999);
and U23458 (N_23458,N_20269,N_20562);
xor U23459 (N_23459,N_21115,N_21058);
nand U23460 (N_23460,N_20444,N_20443);
nor U23461 (N_23461,N_21426,N_20936);
nand U23462 (N_23462,N_20967,N_20169);
xnor U23463 (N_23463,N_20243,N_20948);
and U23464 (N_23464,N_20786,N_20756);
nand U23465 (N_23465,N_21873,N_20593);
xnor U23466 (N_23466,N_20433,N_21276);
nor U23467 (N_23467,N_21800,N_21008);
and U23468 (N_23468,N_20839,N_20923);
or U23469 (N_23469,N_20970,N_21260);
or U23470 (N_23470,N_21068,N_21149);
nor U23471 (N_23471,N_20950,N_20905);
or U23472 (N_23472,N_20113,N_20565);
xnor U23473 (N_23473,N_20509,N_20727);
nand U23474 (N_23474,N_20178,N_21534);
and U23475 (N_23475,N_20539,N_20704);
and U23476 (N_23476,N_21991,N_20858);
nand U23477 (N_23477,N_20207,N_21664);
or U23478 (N_23478,N_20492,N_20336);
nor U23479 (N_23479,N_21480,N_20243);
or U23480 (N_23480,N_21239,N_20840);
nand U23481 (N_23481,N_20314,N_20200);
and U23482 (N_23482,N_20974,N_20789);
or U23483 (N_23483,N_20312,N_20603);
and U23484 (N_23484,N_20903,N_20817);
and U23485 (N_23485,N_21186,N_21855);
xnor U23486 (N_23486,N_21819,N_21979);
nor U23487 (N_23487,N_20459,N_20773);
nand U23488 (N_23488,N_20116,N_21816);
and U23489 (N_23489,N_21531,N_21228);
and U23490 (N_23490,N_20351,N_21382);
and U23491 (N_23491,N_21607,N_21606);
or U23492 (N_23492,N_20252,N_20451);
nand U23493 (N_23493,N_21674,N_21671);
xnor U23494 (N_23494,N_21086,N_20871);
nor U23495 (N_23495,N_20952,N_21326);
or U23496 (N_23496,N_21821,N_21020);
and U23497 (N_23497,N_21525,N_21233);
xnor U23498 (N_23498,N_21566,N_20273);
or U23499 (N_23499,N_21721,N_20288);
or U23500 (N_23500,N_21322,N_21125);
nor U23501 (N_23501,N_21206,N_20461);
nand U23502 (N_23502,N_21146,N_20035);
xor U23503 (N_23503,N_20205,N_21456);
and U23504 (N_23504,N_21152,N_20389);
or U23505 (N_23505,N_20508,N_21680);
nor U23506 (N_23506,N_21010,N_20172);
nand U23507 (N_23507,N_21021,N_21667);
nand U23508 (N_23508,N_21520,N_20728);
xor U23509 (N_23509,N_20772,N_20001);
nor U23510 (N_23510,N_20300,N_21552);
nand U23511 (N_23511,N_20249,N_20857);
nand U23512 (N_23512,N_21168,N_20460);
xor U23513 (N_23513,N_21523,N_21590);
or U23514 (N_23514,N_20940,N_20517);
nor U23515 (N_23515,N_20594,N_21988);
nor U23516 (N_23516,N_21506,N_21965);
and U23517 (N_23517,N_20716,N_21114);
nor U23518 (N_23518,N_21626,N_21195);
nor U23519 (N_23519,N_21772,N_20226);
and U23520 (N_23520,N_20404,N_21040);
and U23521 (N_23521,N_20158,N_21437);
nand U23522 (N_23522,N_21561,N_21403);
xnor U23523 (N_23523,N_20127,N_20866);
and U23524 (N_23524,N_21005,N_20209);
and U23525 (N_23525,N_20586,N_21377);
nor U23526 (N_23526,N_21919,N_20134);
and U23527 (N_23527,N_20297,N_20284);
nor U23528 (N_23528,N_21517,N_20049);
or U23529 (N_23529,N_21032,N_21217);
nor U23530 (N_23530,N_21995,N_20511);
nor U23531 (N_23531,N_21288,N_21018);
nand U23532 (N_23532,N_21572,N_21926);
xnor U23533 (N_23533,N_21831,N_20702);
xor U23534 (N_23534,N_21769,N_20681);
xor U23535 (N_23535,N_20625,N_20687);
nor U23536 (N_23536,N_21514,N_21122);
nand U23537 (N_23537,N_21406,N_20761);
xnor U23538 (N_23538,N_21470,N_20240);
nor U23539 (N_23539,N_20251,N_21253);
and U23540 (N_23540,N_20017,N_21219);
nand U23541 (N_23541,N_20625,N_20618);
xnor U23542 (N_23542,N_20254,N_20899);
or U23543 (N_23543,N_20836,N_20746);
nand U23544 (N_23544,N_21867,N_21701);
or U23545 (N_23545,N_20215,N_21071);
nand U23546 (N_23546,N_20592,N_21183);
nor U23547 (N_23547,N_20790,N_21833);
nor U23548 (N_23548,N_20630,N_21776);
nor U23549 (N_23549,N_21947,N_20691);
or U23550 (N_23550,N_20918,N_21968);
nand U23551 (N_23551,N_21868,N_20467);
xor U23552 (N_23552,N_21609,N_20015);
or U23553 (N_23553,N_20005,N_20853);
and U23554 (N_23554,N_21391,N_20442);
and U23555 (N_23555,N_21127,N_20813);
or U23556 (N_23556,N_21912,N_21190);
xnor U23557 (N_23557,N_20279,N_20116);
and U23558 (N_23558,N_21633,N_21982);
or U23559 (N_23559,N_21906,N_21555);
xor U23560 (N_23560,N_20796,N_21862);
or U23561 (N_23561,N_21920,N_20353);
nand U23562 (N_23562,N_21852,N_21742);
nor U23563 (N_23563,N_20862,N_21330);
or U23564 (N_23564,N_20744,N_21582);
or U23565 (N_23565,N_20668,N_21904);
nor U23566 (N_23566,N_20806,N_21429);
nand U23567 (N_23567,N_21491,N_21020);
or U23568 (N_23568,N_20096,N_20705);
or U23569 (N_23569,N_20865,N_20232);
xnor U23570 (N_23570,N_20164,N_20183);
nand U23571 (N_23571,N_20816,N_20703);
and U23572 (N_23572,N_20944,N_20738);
nand U23573 (N_23573,N_20815,N_20604);
or U23574 (N_23574,N_21412,N_21858);
xnor U23575 (N_23575,N_21618,N_21311);
xnor U23576 (N_23576,N_20881,N_21930);
or U23577 (N_23577,N_20820,N_21403);
nor U23578 (N_23578,N_21180,N_20601);
xnor U23579 (N_23579,N_20557,N_20639);
or U23580 (N_23580,N_20259,N_20499);
nor U23581 (N_23581,N_20006,N_21634);
and U23582 (N_23582,N_21444,N_21697);
or U23583 (N_23583,N_21579,N_20755);
xor U23584 (N_23584,N_21022,N_21006);
or U23585 (N_23585,N_21491,N_20862);
nand U23586 (N_23586,N_21099,N_21422);
or U23587 (N_23587,N_21357,N_21913);
xor U23588 (N_23588,N_20170,N_21023);
and U23589 (N_23589,N_20658,N_20787);
or U23590 (N_23590,N_21191,N_21222);
or U23591 (N_23591,N_20712,N_21090);
and U23592 (N_23592,N_21187,N_21293);
nand U23593 (N_23593,N_20796,N_20985);
nand U23594 (N_23594,N_20304,N_21525);
nand U23595 (N_23595,N_20078,N_21153);
and U23596 (N_23596,N_20065,N_21157);
nor U23597 (N_23597,N_21603,N_20448);
xnor U23598 (N_23598,N_21862,N_20928);
and U23599 (N_23599,N_20651,N_21145);
or U23600 (N_23600,N_20193,N_21601);
or U23601 (N_23601,N_20890,N_21928);
and U23602 (N_23602,N_21447,N_21684);
xor U23603 (N_23603,N_20011,N_20383);
nand U23604 (N_23604,N_21320,N_20325);
nor U23605 (N_23605,N_20798,N_21610);
xnor U23606 (N_23606,N_20358,N_20708);
and U23607 (N_23607,N_20739,N_20851);
nor U23608 (N_23608,N_21831,N_20279);
nand U23609 (N_23609,N_20307,N_21862);
nor U23610 (N_23610,N_21667,N_20024);
xor U23611 (N_23611,N_21476,N_21401);
xnor U23612 (N_23612,N_21008,N_21205);
nor U23613 (N_23613,N_21183,N_21685);
nor U23614 (N_23614,N_20479,N_20237);
nor U23615 (N_23615,N_21882,N_20397);
nor U23616 (N_23616,N_20914,N_21070);
xor U23617 (N_23617,N_21539,N_21669);
nand U23618 (N_23618,N_20750,N_21687);
nor U23619 (N_23619,N_20131,N_21327);
and U23620 (N_23620,N_21407,N_20586);
nand U23621 (N_23621,N_20301,N_21181);
xor U23622 (N_23622,N_21451,N_20861);
xnor U23623 (N_23623,N_21228,N_21022);
and U23624 (N_23624,N_20642,N_21755);
xnor U23625 (N_23625,N_20424,N_20310);
and U23626 (N_23626,N_20942,N_21393);
or U23627 (N_23627,N_21035,N_21940);
or U23628 (N_23628,N_20036,N_21849);
nand U23629 (N_23629,N_20490,N_20153);
and U23630 (N_23630,N_20032,N_20079);
xnor U23631 (N_23631,N_20897,N_20891);
nor U23632 (N_23632,N_20323,N_21627);
or U23633 (N_23633,N_20595,N_21571);
xor U23634 (N_23634,N_21315,N_21852);
nand U23635 (N_23635,N_21951,N_20376);
or U23636 (N_23636,N_21053,N_21081);
nor U23637 (N_23637,N_20898,N_20429);
xor U23638 (N_23638,N_21902,N_20870);
and U23639 (N_23639,N_20505,N_20301);
xnor U23640 (N_23640,N_21649,N_20608);
xor U23641 (N_23641,N_20263,N_21243);
nor U23642 (N_23642,N_21463,N_20981);
or U23643 (N_23643,N_20780,N_20460);
xnor U23644 (N_23644,N_21179,N_20612);
or U23645 (N_23645,N_20210,N_21413);
and U23646 (N_23646,N_21606,N_21363);
and U23647 (N_23647,N_20335,N_20905);
xor U23648 (N_23648,N_20750,N_21196);
xnor U23649 (N_23649,N_21438,N_21295);
nand U23650 (N_23650,N_20366,N_20885);
xnor U23651 (N_23651,N_21631,N_21259);
or U23652 (N_23652,N_21177,N_21178);
and U23653 (N_23653,N_21016,N_21588);
and U23654 (N_23654,N_20900,N_20030);
nand U23655 (N_23655,N_21550,N_20741);
or U23656 (N_23656,N_21842,N_20493);
xnor U23657 (N_23657,N_21840,N_21761);
nor U23658 (N_23658,N_21261,N_21854);
and U23659 (N_23659,N_20708,N_20296);
nand U23660 (N_23660,N_20112,N_21668);
xnor U23661 (N_23661,N_21353,N_20041);
and U23662 (N_23662,N_20262,N_21690);
or U23663 (N_23663,N_21434,N_20498);
or U23664 (N_23664,N_21116,N_21846);
xor U23665 (N_23665,N_21116,N_20259);
nand U23666 (N_23666,N_20198,N_21213);
or U23667 (N_23667,N_20671,N_20166);
or U23668 (N_23668,N_20306,N_21834);
and U23669 (N_23669,N_21279,N_21908);
and U23670 (N_23670,N_20081,N_20437);
nor U23671 (N_23671,N_21934,N_21373);
and U23672 (N_23672,N_20790,N_20495);
and U23673 (N_23673,N_20269,N_20565);
nand U23674 (N_23674,N_20249,N_21031);
or U23675 (N_23675,N_20903,N_21821);
xnor U23676 (N_23676,N_21136,N_20794);
nor U23677 (N_23677,N_20139,N_21915);
nor U23678 (N_23678,N_20220,N_20061);
or U23679 (N_23679,N_21003,N_20947);
nor U23680 (N_23680,N_21556,N_20658);
or U23681 (N_23681,N_21409,N_20688);
nor U23682 (N_23682,N_20475,N_20524);
nor U23683 (N_23683,N_21518,N_20562);
and U23684 (N_23684,N_21916,N_21070);
or U23685 (N_23685,N_21820,N_20615);
nand U23686 (N_23686,N_21458,N_20648);
xor U23687 (N_23687,N_21582,N_20420);
nor U23688 (N_23688,N_21897,N_20803);
and U23689 (N_23689,N_21675,N_21508);
xor U23690 (N_23690,N_21963,N_21056);
and U23691 (N_23691,N_20990,N_21132);
and U23692 (N_23692,N_20279,N_21903);
or U23693 (N_23693,N_20067,N_20590);
nand U23694 (N_23694,N_20928,N_20705);
nand U23695 (N_23695,N_21910,N_20398);
xor U23696 (N_23696,N_20158,N_20091);
or U23697 (N_23697,N_20878,N_21419);
or U23698 (N_23698,N_21974,N_20335);
xor U23699 (N_23699,N_21356,N_21407);
and U23700 (N_23700,N_20241,N_21596);
xor U23701 (N_23701,N_21691,N_21233);
nand U23702 (N_23702,N_21951,N_21994);
or U23703 (N_23703,N_21387,N_21533);
or U23704 (N_23704,N_21614,N_20211);
nor U23705 (N_23705,N_21882,N_20996);
nand U23706 (N_23706,N_21123,N_20329);
or U23707 (N_23707,N_21098,N_20884);
and U23708 (N_23708,N_21314,N_21566);
nand U23709 (N_23709,N_21705,N_21680);
or U23710 (N_23710,N_21540,N_21220);
nor U23711 (N_23711,N_21025,N_20935);
nor U23712 (N_23712,N_20444,N_20213);
or U23713 (N_23713,N_20320,N_21360);
nor U23714 (N_23714,N_20005,N_21609);
nand U23715 (N_23715,N_20921,N_21683);
or U23716 (N_23716,N_20840,N_20991);
nor U23717 (N_23717,N_21371,N_21874);
and U23718 (N_23718,N_21148,N_21406);
xor U23719 (N_23719,N_20677,N_20484);
nand U23720 (N_23720,N_21476,N_20153);
nor U23721 (N_23721,N_20224,N_21139);
nor U23722 (N_23722,N_21698,N_20404);
xor U23723 (N_23723,N_20283,N_20870);
nor U23724 (N_23724,N_20557,N_21500);
nand U23725 (N_23725,N_20378,N_21403);
or U23726 (N_23726,N_20682,N_21720);
and U23727 (N_23727,N_20149,N_21188);
nand U23728 (N_23728,N_21695,N_20554);
and U23729 (N_23729,N_21388,N_20351);
and U23730 (N_23730,N_20763,N_20796);
nand U23731 (N_23731,N_21897,N_20552);
and U23732 (N_23732,N_20516,N_21885);
and U23733 (N_23733,N_20663,N_21019);
nand U23734 (N_23734,N_21671,N_20033);
or U23735 (N_23735,N_20543,N_21193);
or U23736 (N_23736,N_21022,N_21193);
nand U23737 (N_23737,N_20532,N_20211);
and U23738 (N_23738,N_21229,N_21199);
and U23739 (N_23739,N_21413,N_20890);
nand U23740 (N_23740,N_20959,N_20086);
or U23741 (N_23741,N_21477,N_20441);
or U23742 (N_23742,N_21157,N_21178);
nor U23743 (N_23743,N_21258,N_20351);
nand U23744 (N_23744,N_21740,N_21356);
nand U23745 (N_23745,N_21762,N_20076);
nor U23746 (N_23746,N_21822,N_21302);
nand U23747 (N_23747,N_20451,N_20438);
nor U23748 (N_23748,N_21075,N_21765);
nor U23749 (N_23749,N_20254,N_20060);
nand U23750 (N_23750,N_20343,N_20189);
xor U23751 (N_23751,N_21571,N_21022);
nor U23752 (N_23752,N_21682,N_20508);
or U23753 (N_23753,N_20798,N_21793);
nand U23754 (N_23754,N_21642,N_20147);
xor U23755 (N_23755,N_20009,N_20879);
and U23756 (N_23756,N_21076,N_20232);
or U23757 (N_23757,N_21273,N_20944);
xor U23758 (N_23758,N_21704,N_21293);
nor U23759 (N_23759,N_21083,N_21974);
and U23760 (N_23760,N_20188,N_20759);
or U23761 (N_23761,N_20438,N_20571);
nor U23762 (N_23762,N_20379,N_20097);
or U23763 (N_23763,N_21026,N_21423);
nor U23764 (N_23764,N_20411,N_21666);
or U23765 (N_23765,N_20608,N_20986);
and U23766 (N_23766,N_21441,N_20307);
nor U23767 (N_23767,N_20234,N_20609);
xnor U23768 (N_23768,N_20247,N_20710);
xor U23769 (N_23769,N_21814,N_21855);
nor U23770 (N_23770,N_21058,N_20460);
or U23771 (N_23771,N_20911,N_21642);
nor U23772 (N_23772,N_20455,N_21317);
nor U23773 (N_23773,N_20666,N_21544);
nand U23774 (N_23774,N_21353,N_21658);
and U23775 (N_23775,N_20566,N_20758);
and U23776 (N_23776,N_20174,N_20674);
xnor U23777 (N_23777,N_21583,N_20399);
and U23778 (N_23778,N_20553,N_21831);
xnor U23779 (N_23779,N_20861,N_21382);
nor U23780 (N_23780,N_21224,N_20629);
or U23781 (N_23781,N_20116,N_20131);
nand U23782 (N_23782,N_21634,N_21258);
nor U23783 (N_23783,N_21532,N_20879);
nand U23784 (N_23784,N_21792,N_21079);
or U23785 (N_23785,N_20420,N_20477);
nor U23786 (N_23786,N_21255,N_21958);
nor U23787 (N_23787,N_21358,N_20325);
nor U23788 (N_23788,N_21182,N_21978);
and U23789 (N_23789,N_20152,N_20126);
xnor U23790 (N_23790,N_20425,N_20611);
xor U23791 (N_23791,N_21931,N_21506);
nand U23792 (N_23792,N_20595,N_21641);
or U23793 (N_23793,N_21914,N_21687);
or U23794 (N_23794,N_20178,N_20282);
or U23795 (N_23795,N_20016,N_21611);
nor U23796 (N_23796,N_20723,N_20423);
xnor U23797 (N_23797,N_20854,N_21395);
and U23798 (N_23798,N_21954,N_21143);
xor U23799 (N_23799,N_21900,N_21420);
and U23800 (N_23800,N_21386,N_21425);
and U23801 (N_23801,N_21464,N_21756);
or U23802 (N_23802,N_20845,N_20730);
nor U23803 (N_23803,N_20183,N_21652);
nor U23804 (N_23804,N_20168,N_21184);
nand U23805 (N_23805,N_20918,N_20039);
or U23806 (N_23806,N_21159,N_20972);
nand U23807 (N_23807,N_21643,N_21598);
xor U23808 (N_23808,N_20843,N_20576);
xnor U23809 (N_23809,N_21584,N_21454);
xor U23810 (N_23810,N_21720,N_20747);
xor U23811 (N_23811,N_21541,N_20165);
xor U23812 (N_23812,N_20677,N_20676);
and U23813 (N_23813,N_21512,N_20526);
or U23814 (N_23814,N_20240,N_20335);
nor U23815 (N_23815,N_20016,N_21070);
nor U23816 (N_23816,N_21936,N_20603);
xor U23817 (N_23817,N_21418,N_20354);
nand U23818 (N_23818,N_20604,N_20347);
nor U23819 (N_23819,N_21553,N_21231);
and U23820 (N_23820,N_20628,N_21666);
or U23821 (N_23821,N_21616,N_20995);
nand U23822 (N_23822,N_21568,N_21338);
and U23823 (N_23823,N_21089,N_21568);
nand U23824 (N_23824,N_21891,N_21333);
nor U23825 (N_23825,N_21884,N_20091);
or U23826 (N_23826,N_20972,N_21485);
xor U23827 (N_23827,N_20808,N_21615);
nand U23828 (N_23828,N_20373,N_20059);
nor U23829 (N_23829,N_20380,N_21509);
nand U23830 (N_23830,N_20287,N_20011);
and U23831 (N_23831,N_20111,N_21313);
and U23832 (N_23832,N_21977,N_21190);
nor U23833 (N_23833,N_20290,N_20747);
nor U23834 (N_23834,N_20952,N_21120);
nor U23835 (N_23835,N_21559,N_21696);
nand U23836 (N_23836,N_21087,N_20716);
nand U23837 (N_23837,N_20124,N_21274);
nor U23838 (N_23838,N_21058,N_20064);
and U23839 (N_23839,N_20097,N_21592);
nand U23840 (N_23840,N_20843,N_20028);
nand U23841 (N_23841,N_20976,N_21064);
xor U23842 (N_23842,N_20895,N_21868);
or U23843 (N_23843,N_20392,N_21475);
and U23844 (N_23844,N_20460,N_21041);
or U23845 (N_23845,N_21631,N_20205);
xor U23846 (N_23846,N_20244,N_20634);
or U23847 (N_23847,N_21054,N_21852);
or U23848 (N_23848,N_21210,N_20387);
nand U23849 (N_23849,N_21305,N_20611);
or U23850 (N_23850,N_20456,N_20968);
and U23851 (N_23851,N_21384,N_21009);
and U23852 (N_23852,N_21507,N_20306);
and U23853 (N_23853,N_20668,N_20694);
nand U23854 (N_23854,N_20109,N_20839);
nand U23855 (N_23855,N_21549,N_20357);
and U23856 (N_23856,N_20135,N_20348);
xnor U23857 (N_23857,N_21535,N_20181);
nor U23858 (N_23858,N_20926,N_20965);
or U23859 (N_23859,N_21096,N_20932);
or U23860 (N_23860,N_20831,N_21444);
nand U23861 (N_23861,N_21106,N_21997);
and U23862 (N_23862,N_20782,N_21959);
nor U23863 (N_23863,N_20076,N_20514);
xnor U23864 (N_23864,N_20511,N_21242);
or U23865 (N_23865,N_20068,N_20531);
nand U23866 (N_23866,N_21909,N_21275);
and U23867 (N_23867,N_21002,N_20513);
nand U23868 (N_23868,N_20331,N_21791);
nand U23869 (N_23869,N_20475,N_20621);
and U23870 (N_23870,N_21790,N_21310);
nand U23871 (N_23871,N_21950,N_20191);
xor U23872 (N_23872,N_20558,N_20430);
nand U23873 (N_23873,N_20160,N_21454);
xor U23874 (N_23874,N_20523,N_20302);
xnor U23875 (N_23875,N_21545,N_20663);
nor U23876 (N_23876,N_21043,N_20254);
nand U23877 (N_23877,N_21224,N_20111);
and U23878 (N_23878,N_21056,N_21290);
nor U23879 (N_23879,N_21907,N_20001);
nor U23880 (N_23880,N_20814,N_20052);
nand U23881 (N_23881,N_20090,N_20162);
and U23882 (N_23882,N_20242,N_20621);
nand U23883 (N_23883,N_21762,N_21408);
or U23884 (N_23884,N_21753,N_20002);
nor U23885 (N_23885,N_20513,N_20992);
nand U23886 (N_23886,N_20599,N_20762);
nor U23887 (N_23887,N_20048,N_20112);
or U23888 (N_23888,N_21394,N_20869);
and U23889 (N_23889,N_21991,N_21735);
and U23890 (N_23890,N_20740,N_20323);
xnor U23891 (N_23891,N_20974,N_20587);
nor U23892 (N_23892,N_21573,N_20175);
xor U23893 (N_23893,N_21290,N_21387);
xor U23894 (N_23894,N_21653,N_21355);
xnor U23895 (N_23895,N_21100,N_20336);
nand U23896 (N_23896,N_21583,N_21206);
nand U23897 (N_23897,N_21575,N_20507);
xor U23898 (N_23898,N_20331,N_20655);
and U23899 (N_23899,N_20066,N_20653);
or U23900 (N_23900,N_21137,N_21329);
nand U23901 (N_23901,N_20420,N_21909);
nor U23902 (N_23902,N_21408,N_21005);
nor U23903 (N_23903,N_20047,N_20856);
xor U23904 (N_23904,N_21615,N_20299);
and U23905 (N_23905,N_20185,N_20536);
or U23906 (N_23906,N_21515,N_20092);
and U23907 (N_23907,N_20421,N_20332);
nor U23908 (N_23908,N_21811,N_20107);
nand U23909 (N_23909,N_21830,N_20558);
nor U23910 (N_23910,N_21256,N_20742);
nor U23911 (N_23911,N_21732,N_20176);
xor U23912 (N_23912,N_20198,N_21479);
nor U23913 (N_23913,N_21354,N_21464);
nor U23914 (N_23914,N_20743,N_21828);
or U23915 (N_23915,N_20356,N_21898);
or U23916 (N_23916,N_21614,N_20469);
xnor U23917 (N_23917,N_20743,N_21805);
xor U23918 (N_23918,N_21820,N_20496);
nor U23919 (N_23919,N_21088,N_21843);
nand U23920 (N_23920,N_21455,N_21617);
nor U23921 (N_23921,N_21795,N_21610);
xnor U23922 (N_23922,N_21623,N_20578);
and U23923 (N_23923,N_21830,N_21195);
xor U23924 (N_23924,N_21974,N_20116);
nand U23925 (N_23925,N_21153,N_21164);
nand U23926 (N_23926,N_21332,N_20391);
or U23927 (N_23927,N_20065,N_20646);
nor U23928 (N_23928,N_21348,N_21970);
nor U23929 (N_23929,N_21403,N_20070);
or U23930 (N_23930,N_20497,N_20459);
and U23931 (N_23931,N_20924,N_20085);
nand U23932 (N_23932,N_21263,N_20662);
or U23933 (N_23933,N_20264,N_20796);
or U23934 (N_23934,N_21052,N_21597);
and U23935 (N_23935,N_20904,N_20758);
nor U23936 (N_23936,N_20494,N_21575);
nor U23937 (N_23937,N_21065,N_21929);
and U23938 (N_23938,N_21661,N_21149);
or U23939 (N_23939,N_20934,N_20968);
or U23940 (N_23940,N_21112,N_21650);
or U23941 (N_23941,N_20154,N_20299);
xnor U23942 (N_23942,N_20553,N_21478);
or U23943 (N_23943,N_20173,N_20889);
nand U23944 (N_23944,N_20182,N_20528);
nor U23945 (N_23945,N_20622,N_20993);
xor U23946 (N_23946,N_21341,N_20678);
xnor U23947 (N_23947,N_21157,N_21169);
or U23948 (N_23948,N_21221,N_21248);
nand U23949 (N_23949,N_21511,N_20226);
nor U23950 (N_23950,N_20947,N_20922);
nand U23951 (N_23951,N_20155,N_20717);
and U23952 (N_23952,N_21913,N_20011);
and U23953 (N_23953,N_21469,N_21837);
and U23954 (N_23954,N_21278,N_21178);
or U23955 (N_23955,N_20958,N_21644);
xor U23956 (N_23956,N_21130,N_21334);
and U23957 (N_23957,N_20525,N_20511);
or U23958 (N_23958,N_21786,N_20051);
or U23959 (N_23959,N_21424,N_21759);
nor U23960 (N_23960,N_20335,N_21155);
nor U23961 (N_23961,N_20590,N_20579);
nor U23962 (N_23962,N_20120,N_20144);
or U23963 (N_23963,N_21780,N_21867);
xor U23964 (N_23964,N_20335,N_20973);
nand U23965 (N_23965,N_21998,N_21720);
and U23966 (N_23966,N_21181,N_21430);
or U23967 (N_23967,N_21719,N_20608);
nand U23968 (N_23968,N_21751,N_20390);
nand U23969 (N_23969,N_21340,N_20805);
or U23970 (N_23970,N_20015,N_20313);
nand U23971 (N_23971,N_20693,N_20398);
nand U23972 (N_23972,N_20813,N_21629);
and U23973 (N_23973,N_21078,N_20036);
and U23974 (N_23974,N_21781,N_20412);
nand U23975 (N_23975,N_21165,N_20512);
xnor U23976 (N_23976,N_20123,N_20995);
xnor U23977 (N_23977,N_20663,N_21638);
nand U23978 (N_23978,N_21636,N_21514);
xor U23979 (N_23979,N_21955,N_21918);
or U23980 (N_23980,N_20407,N_21382);
nand U23981 (N_23981,N_21328,N_21257);
or U23982 (N_23982,N_20835,N_21631);
nand U23983 (N_23983,N_20501,N_20031);
nand U23984 (N_23984,N_21960,N_20149);
xor U23985 (N_23985,N_20445,N_20654);
nor U23986 (N_23986,N_20854,N_20927);
and U23987 (N_23987,N_20593,N_21757);
nor U23988 (N_23988,N_20693,N_20004);
nor U23989 (N_23989,N_20802,N_21170);
xor U23990 (N_23990,N_21466,N_20147);
or U23991 (N_23991,N_20114,N_20214);
xnor U23992 (N_23992,N_20767,N_21802);
or U23993 (N_23993,N_20046,N_21311);
and U23994 (N_23994,N_20305,N_21151);
nor U23995 (N_23995,N_21686,N_21443);
or U23996 (N_23996,N_20628,N_20704);
nor U23997 (N_23997,N_21650,N_21938);
or U23998 (N_23998,N_20105,N_20121);
xor U23999 (N_23999,N_21456,N_20258);
or U24000 (N_24000,N_23239,N_23390);
nand U24001 (N_24001,N_22165,N_23443);
or U24002 (N_24002,N_22612,N_23056);
xnor U24003 (N_24003,N_23541,N_23894);
nor U24004 (N_24004,N_23023,N_22474);
xnor U24005 (N_24005,N_22753,N_23185);
or U24006 (N_24006,N_22330,N_23581);
xnor U24007 (N_24007,N_23005,N_23888);
nand U24008 (N_24008,N_22705,N_23471);
nor U24009 (N_24009,N_23168,N_22056);
or U24010 (N_24010,N_23523,N_22600);
or U24011 (N_24011,N_23515,N_22573);
nand U24012 (N_24012,N_23638,N_23205);
nor U24013 (N_24013,N_22763,N_22201);
nand U24014 (N_24014,N_23403,N_22316);
nand U24015 (N_24015,N_22537,N_23223);
nor U24016 (N_24016,N_22438,N_22200);
xnor U24017 (N_24017,N_23867,N_23870);
xor U24018 (N_24018,N_23626,N_23357);
or U24019 (N_24019,N_22656,N_23221);
or U24020 (N_24020,N_23649,N_22334);
nor U24021 (N_24021,N_22677,N_22363);
and U24022 (N_24022,N_23635,N_22583);
xor U24023 (N_24023,N_22733,N_22308);
and U24024 (N_24024,N_22014,N_23359);
or U24025 (N_24025,N_23257,N_22571);
or U24026 (N_24026,N_23863,N_23200);
nor U24027 (N_24027,N_23866,N_22079);
nor U24028 (N_24028,N_23982,N_22728);
nand U24029 (N_24029,N_23254,N_22473);
nand U24030 (N_24030,N_23587,N_23828);
nor U24031 (N_24031,N_22364,N_23445);
nand U24032 (N_24032,N_22163,N_23646);
or U24033 (N_24033,N_23464,N_23779);
nor U24034 (N_24034,N_23801,N_22935);
or U24035 (N_24035,N_22749,N_22027);
xor U24036 (N_24036,N_22682,N_23608);
and U24037 (N_24037,N_22619,N_23874);
xor U24038 (N_24038,N_22383,N_23266);
and U24039 (N_24039,N_23376,N_22517);
nor U24040 (N_24040,N_23776,N_23291);
and U24041 (N_24041,N_23662,N_23524);
and U24042 (N_24042,N_23188,N_22215);
nor U24043 (N_24043,N_23909,N_22767);
or U24044 (N_24044,N_22693,N_23313);
nand U24045 (N_24045,N_22930,N_23891);
xnor U24046 (N_24046,N_23955,N_22429);
nor U24047 (N_24047,N_23980,N_22178);
nand U24048 (N_24048,N_23630,N_23184);
nor U24049 (N_24049,N_23788,N_23969);
or U24050 (N_24050,N_22957,N_23526);
nor U24051 (N_24051,N_22807,N_22620);
nor U24052 (N_24052,N_23512,N_23500);
nor U24053 (N_24053,N_23468,N_23873);
xor U24054 (N_24054,N_22333,N_22147);
nor U24055 (N_24055,N_22124,N_23309);
nand U24056 (N_24056,N_23908,N_22060);
nor U24057 (N_24057,N_22506,N_22412);
and U24058 (N_24058,N_22596,N_22526);
xnor U24059 (N_24059,N_23098,N_23077);
xnor U24060 (N_24060,N_22755,N_22367);
and U24061 (N_24061,N_23858,N_22536);
and U24062 (N_24062,N_23379,N_22845);
nand U24063 (N_24063,N_22959,N_23099);
and U24064 (N_24064,N_22575,N_23162);
or U24065 (N_24065,N_22657,N_23108);
nor U24066 (N_24066,N_23210,N_22666);
nor U24067 (N_24067,N_23582,N_23632);
or U24068 (N_24068,N_23502,N_22616);
xor U24069 (N_24069,N_22437,N_23112);
or U24070 (N_24070,N_23277,N_22221);
xnor U24071 (N_24071,N_23220,N_23835);
nand U24072 (N_24072,N_22050,N_23265);
or U24073 (N_24073,N_22582,N_22439);
xor U24074 (N_24074,N_22874,N_22727);
xor U24075 (N_24075,N_22916,N_23804);
and U24076 (N_24076,N_23556,N_23737);
nand U24077 (N_24077,N_22695,N_22402);
xor U24078 (N_24078,N_23449,N_23620);
nand U24079 (N_24079,N_22503,N_22488);
and U24080 (N_24080,N_23007,N_22237);
xnor U24081 (N_24081,N_22016,N_22501);
or U24082 (N_24082,N_22835,N_23451);
nand U24083 (N_24083,N_22740,N_22726);
or U24084 (N_24084,N_23900,N_23038);
and U24085 (N_24085,N_22100,N_22812);
xnor U24086 (N_24086,N_22272,N_23611);
nor U24087 (N_24087,N_22183,N_23740);
or U24088 (N_24088,N_23422,N_22343);
and U24089 (N_24089,N_23217,N_23871);
or U24090 (N_24090,N_22990,N_23362);
nand U24091 (N_24091,N_22299,N_23938);
xnor U24092 (N_24092,N_23329,N_23404);
nor U24093 (N_24093,N_22779,N_22551);
or U24094 (N_24094,N_22114,N_22149);
nor U24095 (N_24095,N_23631,N_22660);
or U24096 (N_24096,N_22256,N_23009);
and U24097 (N_24097,N_22271,N_22670);
and U24098 (N_24098,N_23042,N_22837);
xnor U24099 (N_24099,N_22855,N_23957);
and U24100 (N_24100,N_22524,N_22735);
or U24101 (N_24101,N_22039,N_22170);
nand U24102 (N_24102,N_23881,N_23805);
or U24103 (N_24103,N_22138,N_22385);
or U24104 (N_24104,N_22640,N_22672);
nor U24105 (N_24105,N_23692,N_23853);
or U24106 (N_24106,N_22794,N_22372);
xor U24107 (N_24107,N_22344,N_23561);
or U24108 (N_24108,N_23657,N_22382);
nor U24109 (N_24109,N_23732,N_23886);
and U24110 (N_24110,N_22643,N_23063);
and U24111 (N_24111,N_23034,N_23979);
and U24112 (N_24112,N_23130,N_23251);
nor U24113 (N_24113,N_23171,N_23141);
or U24114 (N_24114,N_22264,N_22665);
nand U24115 (N_24115,N_22997,N_22152);
nand U24116 (N_24116,N_22309,N_23558);
or U24117 (N_24117,N_23480,N_23694);
or U24118 (N_24118,N_23714,N_23961);
and U24119 (N_24119,N_22618,N_22157);
nor U24120 (N_24120,N_22956,N_22588);
xor U24121 (N_24121,N_22131,N_22718);
or U24122 (N_24122,N_23644,N_23547);
or U24123 (N_24123,N_23044,N_22066);
and U24124 (N_24124,N_23510,N_23902);
or U24125 (N_24125,N_23229,N_23519);
xor U24126 (N_24126,N_23267,N_22781);
nand U24127 (N_24127,N_22465,N_23363);
or U24128 (N_24128,N_22830,N_22750);
and U24129 (N_24129,N_22456,N_23400);
and U24130 (N_24130,N_23456,N_23378);
or U24131 (N_24131,N_22389,N_22988);
or U24132 (N_24132,N_22717,N_23018);
and U24133 (N_24133,N_23474,N_22846);
nor U24134 (N_24134,N_22336,N_22758);
or U24135 (N_24135,N_22743,N_23916);
nand U24136 (N_24136,N_22253,N_23452);
xor U24137 (N_24137,N_23967,N_23546);
and U24138 (N_24138,N_22730,N_22240);
nor U24139 (N_24139,N_23335,N_23648);
and U24140 (N_24140,N_22199,N_22135);
or U24141 (N_24141,N_22798,N_23094);
xor U24142 (N_24142,N_23534,N_23743);
xor U24143 (N_24143,N_23415,N_22939);
nand U24144 (N_24144,N_22391,N_23962);
or U24145 (N_24145,N_23917,N_22606);
or U24146 (N_24146,N_22556,N_22917);
nand U24147 (N_24147,N_22088,N_22623);
nand U24148 (N_24148,N_23535,N_22914);
or U24149 (N_24149,N_22980,N_23933);
and U24150 (N_24150,N_23585,N_22707);
xor U24151 (N_24151,N_22599,N_23211);
nand U24152 (N_24152,N_23292,N_22058);
xnor U24153 (N_24153,N_22565,N_23769);
nand U24154 (N_24154,N_22622,N_23450);
nor U24155 (N_24155,N_23919,N_22942);
nand U24156 (N_24156,N_23436,N_23570);
nor U24157 (N_24157,N_22994,N_23301);
nand U24158 (N_24158,N_23704,N_23166);
xor U24159 (N_24159,N_23518,N_23525);
nor U24160 (N_24160,N_22828,N_23149);
or U24161 (N_24161,N_23808,N_22952);
nor U24162 (N_24162,N_22244,N_23670);
xnor U24163 (N_24163,N_23781,N_23627);
and U24164 (N_24164,N_22928,N_22674);
nand U24165 (N_24165,N_23384,N_23813);
or U24166 (N_24166,N_23549,N_22972);
or U24167 (N_24167,N_22061,N_22948);
nand U24168 (N_24168,N_22865,N_22844);
and U24169 (N_24169,N_22184,N_23127);
xnor U24170 (N_24170,N_22720,N_23574);
xor U24171 (N_24171,N_22105,N_22987);
nor U24172 (N_24172,N_22232,N_22592);
xor U24173 (N_24173,N_23106,N_22975);
or U24174 (N_24174,N_22715,N_22734);
xor U24175 (N_24175,N_22587,N_22196);
or U24176 (N_24176,N_22132,N_23231);
nor U24177 (N_24177,N_23173,N_22546);
or U24178 (N_24178,N_22283,N_23531);
nand U24179 (N_24179,N_22801,N_23407);
and U24180 (N_24180,N_23847,N_22408);
nor U24181 (N_24181,N_23444,N_22087);
nand U24182 (N_24182,N_22971,N_23744);
and U24183 (N_24183,N_22228,N_22034);
or U24184 (N_24184,N_23457,N_23928);
xnor U24185 (N_24185,N_23071,N_22772);
nand U24186 (N_24186,N_22598,N_23307);
nand U24187 (N_24187,N_23589,N_22858);
xor U24188 (N_24188,N_22929,N_23840);
nand U24189 (N_24189,N_22561,N_23181);
and U24190 (N_24190,N_23975,N_23613);
and U24191 (N_24191,N_23113,N_22166);
nand U24192 (N_24192,N_23599,N_22529);
xnor U24193 (N_24193,N_22477,N_23537);
nor U24194 (N_24194,N_23489,N_23432);
nor U24195 (N_24195,N_22151,N_23678);
and U24196 (N_24196,N_23138,N_22589);
and U24197 (N_24197,N_23976,N_23745);
xor U24198 (N_24198,N_23616,N_23533);
nor U24199 (N_24199,N_23253,N_22193);
nor U24200 (N_24200,N_22329,N_22968);
nor U24201 (N_24201,N_22202,N_23330);
nor U24202 (N_24202,N_23072,N_22632);
or U24203 (N_24203,N_22886,N_23666);
and U24204 (N_24204,N_22922,N_23084);
nand U24205 (N_24205,N_23892,N_23517);
xor U24206 (N_24206,N_22044,N_22864);
nor U24207 (N_24207,N_22508,N_23696);
nor U24208 (N_24208,N_22624,N_23712);
or U24209 (N_24209,N_23597,N_22799);
and U24210 (N_24210,N_22721,N_22073);
xor U24211 (N_24211,N_22441,N_23062);
nor U24212 (N_24212,N_23380,N_22577);
and U24213 (N_24213,N_23219,N_23821);
nand U24214 (N_24214,N_23566,N_23983);
nor U24215 (N_24215,N_22000,N_23538);
xnor U24216 (N_24216,N_23945,N_22945);
nor U24217 (N_24217,N_23553,N_23275);
or U24218 (N_24218,N_23987,N_23758);
xor U24219 (N_24219,N_23684,N_22366);
xnor U24220 (N_24220,N_23985,N_23941);
nor U24221 (N_24221,N_22615,N_22913);
and U24222 (N_24222,N_22511,N_23771);
xnor U24223 (N_24223,N_22171,N_23722);
nand U24224 (N_24224,N_22017,N_23573);
and U24225 (N_24225,N_22494,N_22908);
nand U24226 (N_24226,N_22198,N_23773);
xor U24227 (N_24227,N_22159,N_22530);
nand U24228 (N_24228,N_22744,N_22607);
xor U24229 (N_24229,N_23332,N_23504);
nor U24230 (N_24230,N_23943,N_23529);
xor U24231 (N_24231,N_22230,N_23775);
nor U24232 (N_24232,N_22901,N_23910);
nor U24233 (N_24233,N_22609,N_23922);
nor U24234 (N_24234,N_23875,N_23802);
nor U24235 (N_24235,N_22368,N_23183);
xor U24236 (N_24236,N_23925,N_22761);
nor U24237 (N_24237,N_23798,N_22045);
nor U24238 (N_24238,N_22466,N_23651);
nor U24239 (N_24239,N_22673,N_23483);
or U24240 (N_24240,N_23230,N_23395);
and U24241 (N_24241,N_22081,N_22424);
and U24242 (N_24242,N_23114,N_22030);
or U24243 (N_24243,N_22703,N_23389);
nand U24244 (N_24244,N_22031,N_22013);
xor U24245 (N_24245,N_23706,N_23559);
nor U24246 (N_24246,N_22295,N_22160);
nand U24247 (N_24247,N_23145,N_22651);
nor U24248 (N_24248,N_22578,N_23350);
nand U24249 (N_24249,N_22586,N_22921);
or U24250 (N_24250,N_22963,N_22273);
and U24251 (N_24251,N_22722,N_23841);
nand U24252 (N_24252,N_23927,N_22502);
xnor U24253 (N_24253,N_22820,N_22162);
xor U24254 (N_24254,N_23476,N_22348);
xnor U24255 (N_24255,N_22791,N_23695);
nor U24256 (N_24256,N_23199,N_22784);
and U24257 (N_24257,N_23026,N_23469);
nand U24258 (N_24258,N_23844,N_23564);
nor U24259 (N_24259,N_22307,N_22291);
or U24260 (N_24260,N_23133,N_22380);
nor U24261 (N_24261,N_23795,N_22225);
xnor U24262 (N_24262,N_23673,N_23037);
xor U24263 (N_24263,N_23912,N_23787);
xnor U24264 (N_24264,N_23467,N_22970);
and U24265 (N_24265,N_22690,N_22895);
xor U24266 (N_24266,N_23033,N_22821);
xnor U24267 (N_24267,N_23315,N_22590);
xor U24268 (N_24268,N_23655,N_22214);
nor U24269 (N_24269,N_22787,N_22259);
nand U24270 (N_24270,N_22966,N_22154);
xor U24271 (N_24271,N_22018,N_22675);
nand U24272 (N_24272,N_23375,N_22853);
nand U24273 (N_24273,N_22411,N_23940);
nor U24274 (N_24274,N_23270,N_22552);
nand U24275 (N_24275,N_22685,N_23012);
or U24276 (N_24276,N_23930,N_22435);
or U24277 (N_24277,N_23609,N_22332);
or U24278 (N_24278,N_22752,N_22759);
or U24279 (N_24279,N_22926,N_22448);
xnor U24280 (N_24280,N_23715,N_23341);
xnor U24281 (N_24281,N_22669,N_23258);
or U24282 (N_24282,N_23920,N_23972);
or U24283 (N_24283,N_22033,N_23242);
and U24284 (N_24284,N_23061,N_23391);
nor U24285 (N_24285,N_23069,N_23700);
or U24286 (N_24286,N_23232,N_23859);
and U24287 (N_24287,N_23355,N_22248);
or U24288 (N_24288,N_23179,N_23667);
nor U24289 (N_24289,N_22738,N_23100);
and U24290 (N_24290,N_22584,N_22732);
and U24291 (N_24291,N_23111,N_23165);
or U24292 (N_24292,N_22832,N_23539);
nand U24293 (N_24293,N_22369,N_23294);
xor U24294 (N_24294,N_23414,N_22139);
and U24295 (N_24295,N_22683,N_23707);
and U24296 (N_24296,N_22993,N_22370);
or U24297 (N_24297,N_23261,N_22986);
nand U24298 (N_24298,N_23435,N_22514);
nor U24299 (N_24299,N_22814,N_22115);
xor U24300 (N_24300,N_23194,N_23346);
xnor U24301 (N_24301,N_23348,N_23675);
nand U24302 (N_24302,N_22011,N_23750);
xnor U24303 (N_24303,N_23506,N_22444);
nand U24304 (N_24304,N_22324,N_22498);
xor U24305 (N_24305,N_23080,N_23093);
and U24306 (N_24306,N_22455,N_22318);
nand U24307 (N_24307,N_23883,N_22554);
xnor U24308 (N_24308,N_22491,N_22143);
nand U24309 (N_24309,N_23503,N_22112);
nand U24310 (N_24310,N_23461,N_23586);
xnor U24311 (N_24311,N_23697,N_23437);
nor U24312 (N_24312,N_23498,N_23322);
nand U24313 (N_24313,N_23090,N_22724);
nand U24314 (N_24314,N_22219,N_22133);
nor U24315 (N_24315,N_23830,N_23421);
or U24316 (N_24316,N_23103,N_23834);
and U24317 (N_24317,N_23175,N_22300);
nand U24318 (N_24318,N_22863,N_22881);
and U24319 (N_24319,N_22247,N_22827);
nand U24320 (N_24320,N_23893,N_22177);
and U24321 (N_24321,N_23899,N_23334);
xnor U24322 (N_24322,N_22775,N_22155);
or U24323 (N_24323,N_23371,N_22856);
xnor U24324 (N_24324,N_23392,N_22636);
xor U24325 (N_24325,N_23575,N_22242);
and U24326 (N_24326,N_23833,N_22797);
or U24327 (N_24327,N_23323,N_23720);
or U24328 (N_24328,N_22175,N_23699);
or U24329 (N_24329,N_23584,N_22442);
nor U24330 (N_24330,N_22420,N_22218);
nor U24331 (N_24331,N_23992,N_23050);
and U24332 (N_24332,N_22946,N_22611);
and U24333 (N_24333,N_23430,N_23478);
nor U24334 (N_24334,N_23351,N_23014);
or U24335 (N_24335,N_23727,N_23022);
and U24336 (N_24336,N_22976,N_23460);
nand U24337 (N_24337,N_23458,N_22037);
nor U24338 (N_24338,N_22723,N_23497);
and U24339 (N_24339,N_23295,N_23466);
xnor U24340 (N_24340,N_22495,N_23550);
and U24341 (N_24341,N_23206,N_23356);
xnor U24342 (N_24342,N_23028,N_23260);
and U24343 (N_24343,N_23079,N_23352);
xor U24344 (N_24344,N_22415,N_22663);
and U24345 (N_24345,N_22436,N_22181);
xor U24346 (N_24346,N_22413,N_22449);
or U24347 (N_24347,N_23793,N_23511);
and U24348 (N_24348,N_23247,N_22704);
and U24349 (N_24349,N_23595,N_23994);
and U24350 (N_24350,N_22729,N_22453);
and U24351 (N_24351,N_23197,N_23016);
or U24352 (N_24352,N_22516,N_22462);
and U24353 (N_24353,N_23192,N_22168);
nor U24354 (N_24354,N_23396,N_22484);
xnor U24355 (N_24355,N_22388,N_23153);
nor U24356 (N_24356,N_23622,N_22089);
nor U24357 (N_24357,N_22207,N_22634);
xnor U24358 (N_24358,N_23532,N_22072);
nor U24359 (N_24359,N_23241,N_23520);
and U24360 (N_24360,N_23685,N_23721);
nor U24361 (N_24361,N_22051,N_23470);
nor U24362 (N_24362,N_23496,N_23193);
xnor U24363 (N_24363,N_23705,N_22542);
nor U24364 (N_24364,N_23059,N_23701);
or U24365 (N_24365,N_23827,N_22505);
nand U24366 (N_24366,N_23011,N_22331);
and U24367 (N_24367,N_22940,N_22579);
xor U24368 (N_24368,N_23687,N_22766);
or U24369 (N_24369,N_23932,N_23191);
nor U24370 (N_24370,N_22595,N_23856);
nor U24371 (N_24371,N_23693,N_23039);
or U24372 (N_24372,N_23484,N_23372);
nor U24373 (N_24373,N_23008,N_22706);
and U24374 (N_24374,N_23385,N_22741);
nand U24375 (N_24375,N_23164,N_22648);
nor U24376 (N_24376,N_23639,N_22375);
xor U24377 (N_24377,N_22338,N_22818);
nor U24378 (N_24378,N_23148,N_23868);
xor U24379 (N_24379,N_23325,N_23121);
nand U24380 (N_24380,N_23854,N_22387);
nor U24381 (N_24381,N_22077,N_22048);
and U24382 (N_24382,N_23250,N_22128);
nand U24383 (N_24383,N_22541,N_23144);
or U24384 (N_24384,N_22545,N_23652);
nor U24385 (N_24385,N_23102,N_23297);
xnor U24386 (N_24386,N_22628,N_22631);
xor U24387 (N_24387,N_22947,N_22645);
xor U24388 (N_24388,N_23681,N_23462);
nand U24389 (N_24389,N_22129,N_22626);
xnor U24390 (N_24390,N_22189,N_22093);
nand U24391 (N_24391,N_23086,N_22550);
xor U24392 (N_24392,N_22062,N_22398);
xnor U24393 (N_24393,N_22274,N_23293);
and U24394 (N_24394,N_22978,N_22239);
or U24395 (N_24395,N_22304,N_22261);
xnor U24396 (N_24396,N_23645,N_22843);
nand U24397 (N_24397,N_23860,N_22602);
nand U24398 (N_24398,N_23851,N_22662);
nand U24399 (N_24399,N_23736,N_23799);
nand U24400 (N_24400,N_23562,N_22136);
xor U24401 (N_24401,N_23934,N_23846);
nand U24402 (N_24402,N_23176,N_22604);
nor U24403 (N_24403,N_22995,N_23249);
xor U24404 (N_24404,N_22739,N_23683);
nand U24405 (N_24405,N_22418,N_23410);
or U24406 (N_24406,N_23600,N_22776);
and U24407 (N_24407,N_22684,N_23746);
nand U24408 (N_24408,N_22659,N_23654);
nor U24409 (N_24409,N_22255,N_22401);
xnor U24410 (N_24410,N_23327,N_22702);
nor U24411 (N_24411,N_23901,N_23953);
or U24412 (N_24412,N_22267,N_22475);
nand U24413 (N_24413,N_22123,N_22637);
xor U24414 (N_24414,N_22172,N_23988);
xnor U24415 (N_24415,N_22053,N_22294);
nand U24416 (N_24416,N_22376,N_23317);
nor U24417 (N_24417,N_23719,N_22173);
xnor U24418 (N_24418,N_22190,N_22325);
nor U24419 (N_24419,N_22771,N_22633);
xor U24420 (N_24420,N_23441,N_22601);
and U24421 (N_24421,N_23215,N_22394);
or U24422 (N_24422,N_23619,N_22802);
or U24423 (N_24423,N_22906,N_23996);
and U24424 (N_24424,N_23676,N_22454);
nor U24425 (N_24425,N_23151,N_23660);
or U24426 (N_24426,N_23861,N_23155);
nand U24427 (N_24427,N_23066,N_23713);
nor U24428 (N_24428,N_22927,N_22410);
nor U24429 (N_24429,N_22967,N_23156);
and U24430 (N_24430,N_22650,N_22937);
and U24431 (N_24431,N_23020,N_22909);
nand U24432 (N_24432,N_23058,N_23288);
and U24433 (N_24433,N_22712,N_23664);
or U24434 (N_24434,N_22688,N_22831);
nor U24435 (N_24435,N_23826,N_22915);
and U24436 (N_24436,N_22156,N_23105);
xor U24437 (N_24437,N_22236,N_22841);
and U24438 (N_24438,N_22098,N_22266);
or U24439 (N_24439,N_22400,N_23358);
xor U24440 (N_24440,N_22384,N_22737);
or U24441 (N_24441,N_22041,N_23110);
or U24442 (N_24442,N_23245,N_23528);
xnor U24443 (N_24443,N_22500,N_22358);
or U24444 (N_24444,N_23650,N_22276);
nor U24445 (N_24445,N_23051,N_23843);
xor U24446 (N_24446,N_22130,N_22187);
nand U24447 (N_24447,N_23321,N_22686);
and U24448 (N_24448,N_23601,N_23944);
and U24449 (N_24449,N_23680,N_22641);
or U24450 (N_24450,N_23576,N_22497);
and U24451 (N_24451,N_23954,N_22019);
nor U24452 (N_24452,N_23641,N_23420);
nand U24453 (N_24453,N_23999,N_23424);
and U24454 (N_24454,N_22340,N_22315);
nor U24455 (N_24455,N_23568,N_23839);
nand U24456 (N_24456,N_22951,N_23225);
or U24457 (N_24457,N_23485,N_22119);
nand U24458 (N_24458,N_23274,N_22337);
xor U24459 (N_24459,N_22907,N_23139);
or U24460 (N_24460,N_23882,N_22713);
nand U24461 (N_24461,N_22806,N_22839);
nor U24462 (N_24462,N_23088,N_22751);
nor U24463 (N_24463,N_22852,N_23820);
or U24464 (N_24464,N_22714,N_23971);
or U24465 (N_24465,N_23494,N_23198);
or U24466 (N_24466,N_23089,N_23491);
and U24467 (N_24467,N_22842,N_22095);
nand U24468 (N_24468,N_23083,N_23926);
nand U24469 (N_24469,N_23981,N_22532);
or U24470 (N_24470,N_22121,N_22293);
nor U24471 (N_24471,N_22654,N_23006);
and U24472 (N_24472,N_22811,N_22208);
and U24473 (N_24473,N_22479,N_22169);
xnor U24474 (N_24474,N_22876,N_23019);
or U24475 (N_24475,N_22848,N_23091);
and U24476 (N_24476,N_23505,N_23495);
and U24477 (N_24477,N_23739,N_23136);
and U24478 (N_24478,N_22538,N_22883);
xnor U24479 (N_24479,N_22804,N_23381);
xor U24480 (N_24480,N_22793,N_22492);
nor U24481 (N_24481,N_23998,N_23025);
and U24482 (N_24482,N_22911,N_23878);
nor U24483 (N_24483,N_23310,N_23448);
nand U24484 (N_24484,N_22485,N_22134);
xnor U24485 (N_24485,N_23316,N_22323);
nor U24486 (N_24486,N_22305,N_23542);
or U24487 (N_24487,N_22360,N_23688);
nand U24488 (N_24488,N_22211,N_23942);
xnor U24489 (N_24489,N_23774,N_22817);
nor U24490 (N_24490,N_23222,N_23203);
xnor U24491 (N_24491,N_22658,N_22185);
nor U24492 (N_24492,N_23213,N_22862);
nor U24493 (N_24493,N_23836,N_23767);
and U24494 (N_24494,N_22238,N_23447);
and U24495 (N_24495,N_23101,N_22047);
or U24496 (N_24496,N_23658,N_23730);
nand U24497 (N_24497,N_23053,N_22824);
nand U24498 (N_24498,N_22188,N_23463);
and U24499 (N_24499,N_23973,N_23780);
nor U24500 (N_24500,N_22765,N_22700);
xor U24501 (N_24501,N_22671,N_22074);
nand U24502 (N_24502,N_22719,N_23904);
xor U24503 (N_24503,N_22629,N_22871);
or U24504 (N_24504,N_23140,N_23852);
nand U24505 (N_24505,N_23428,N_23751);
or U24506 (N_24506,N_22287,N_23308);
nor U24507 (N_24507,N_22430,N_22581);
xnor U24508 (N_24508,N_22227,N_23929);
nor U24509 (N_24509,N_23208,N_22191);
xor U24510 (N_24510,N_23965,N_22192);
and U24511 (N_24511,N_22306,N_23741);
or U24512 (N_24512,N_22515,N_22083);
xnor U24513 (N_24513,N_22954,N_22481);
xnor U24514 (N_24514,N_22046,N_22025);
xor U24515 (N_24515,N_23508,N_22569);
nand U24516 (N_24516,N_22009,N_23426);
xor U24517 (N_24517,N_22711,N_23606);
nor U24518 (N_24518,N_22894,N_22667);
or U24519 (N_24519,N_22161,N_22148);
or U24520 (N_24520,N_23117,N_23021);
xor U24521 (N_24521,N_23097,N_23552);
nand U24522 (N_24522,N_23540,N_23482);
nand U24523 (N_24523,N_23823,N_22458);
and U24524 (N_24524,N_23119,N_22285);
and U24525 (N_24525,N_23320,N_23015);
xnor U24526 (N_24526,N_22647,N_22851);
nor U24527 (N_24527,N_22745,N_23060);
nand U24528 (N_24528,N_23734,N_23374);
nor U24529 (N_24529,N_23952,N_22164);
nand U24530 (N_24530,N_23995,N_22534);
and U24531 (N_24531,N_22603,N_22955);
nor U24532 (N_24532,N_22923,N_23545);
or U24533 (N_24533,N_23324,N_23885);
xor U24534 (N_24534,N_22483,N_23731);
and U24535 (N_24535,N_22860,N_23132);
nand U24536 (N_24536,N_23416,N_23280);
or U24537 (N_24537,N_22269,N_23551);
or U24538 (N_24538,N_23339,N_23340);
or U24539 (N_24539,N_23342,N_23347);
xor U24540 (N_24540,N_23488,N_22872);
nand U24541 (N_24541,N_23784,N_23825);
nand U24542 (N_24542,N_23439,N_23472);
or U24543 (N_24543,N_23783,N_23236);
or U24544 (N_24544,N_22086,N_22101);
nor U24545 (N_24545,N_23465,N_22346);
and U24546 (N_24546,N_23178,N_23530);
or U24547 (N_24547,N_23349,N_22560);
and U24548 (N_24548,N_23186,N_23234);
xor U24549 (N_24549,N_22471,N_22985);
nand U24550 (N_24550,N_23583,N_22301);
or U24551 (N_24551,N_23147,N_23202);
or U24552 (N_24552,N_23169,N_23163);
and U24553 (N_24553,N_22891,N_23262);
nor U24554 (N_24554,N_23306,N_22661);
xor U24555 (N_24555,N_23305,N_23742);
or U24556 (N_24556,N_22496,N_23876);
or U24557 (N_24557,N_22613,N_23240);
xor U24558 (N_24558,N_22823,N_22887);
nand U24559 (N_24559,N_23377,N_22889);
xnor U24560 (N_24560,N_22610,N_23233);
xor U24561 (N_24561,N_22280,N_22407);
and U24562 (N_24562,N_22697,N_22625);
nand U24563 (N_24563,N_23991,N_23216);
or U24564 (N_24564,N_23300,N_22878);
nand U24565 (N_24565,N_23244,N_23064);
nand U24566 (N_24566,N_22094,N_23024);
xor U24567 (N_24567,N_23710,N_22819);
and U24568 (N_24568,N_22938,N_22392);
or U24569 (N_24569,N_23344,N_22694);
nand U24570 (N_24570,N_23728,N_23182);
nor U24571 (N_24571,N_23046,N_22962);
and U24572 (N_24572,N_23278,N_23509);
and U24573 (N_24573,N_23521,N_23590);
and U24574 (N_24574,N_22800,N_22371);
or U24575 (N_24575,N_22126,N_23725);
nand U24576 (N_24576,N_23554,N_23076);
nand U24577 (N_24577,N_23669,N_23049);
nor U24578 (N_24578,N_23490,N_23142);
xor U24579 (N_24579,N_23180,N_23459);
nand U24580 (N_24580,N_22194,N_22576);
or U24581 (N_24581,N_23778,N_22850);
xor U24582 (N_24582,N_23029,N_23411);
nand U24583 (N_24583,N_23000,N_23890);
or U24584 (N_24584,N_23653,N_22680);
nand U24585 (N_24585,N_23207,N_22140);
or U24586 (N_24586,N_22489,N_22097);
and U24587 (N_24587,N_23898,N_23759);
or U24588 (N_24588,N_23337,N_22222);
nand U24589 (N_24589,N_23791,N_23235);
xnor U24590 (N_24590,N_23711,N_22055);
or U24591 (N_24591,N_22012,N_22639);
xnor U24592 (N_24592,N_22224,N_22983);
nand U24593 (N_24593,N_22996,N_22374);
or U24594 (N_24594,N_22974,N_23237);
and U24595 (N_24595,N_23897,N_22250);
nand U24596 (N_24596,N_23418,N_23811);
nor U24597 (N_24597,N_22288,N_22757);
and U24598 (N_24598,N_23656,N_23296);
nand U24599 (N_24599,N_23977,N_23455);
nor U24600 (N_24600,N_22432,N_22965);
nor U24601 (N_24601,N_23032,N_22270);
and U24602 (N_24602,N_22118,N_22897);
or U24603 (N_24603,N_23748,N_23984);
xor U24604 (N_24604,N_22810,N_22167);
nand U24605 (N_24605,N_23272,N_22960);
or U24606 (N_24606,N_22989,N_22574);
and U24607 (N_24607,N_23122,N_22953);
nor U24608 (N_24608,N_23757,N_23939);
and U24609 (N_24609,N_22099,N_22092);
or U24610 (N_24610,N_23361,N_22040);
xor U24611 (N_24611,N_22258,N_23906);
nor U24612 (N_24612,N_23336,N_22768);
and U24613 (N_24613,N_22805,N_22969);
nor U24614 (N_24614,N_23368,N_22347);
nor U24615 (N_24615,N_22290,N_22007);
xor U24616 (N_24616,N_23312,N_22888);
nor U24617 (N_24617,N_23544,N_22941);
xor U24618 (N_24618,N_23747,N_22365);
nor U24619 (N_24619,N_22877,N_23045);
xnor U24620 (N_24620,N_23040,N_22652);
xnor U24621 (N_24621,N_23259,N_22345);
nand U24622 (N_24622,N_22570,N_22022);
xnor U24623 (N_24623,N_22203,N_22900);
nand U24624 (N_24624,N_22137,N_22427);
and U24625 (N_24625,N_23286,N_23703);
nor U24626 (N_24626,N_23143,N_23951);
or U24627 (N_24627,N_22958,N_22052);
or U24628 (N_24628,N_23078,N_22857);
nor U24629 (N_24629,N_22527,N_22080);
nand U24630 (N_24630,N_23486,N_23580);
xnor U24631 (N_24631,N_22557,N_22523);
or U24632 (N_24632,N_23958,N_23252);
nand U24633 (N_24633,N_22698,N_22866);
xnor U24634 (N_24634,N_22838,N_23075);
or U24635 (N_24635,N_22472,N_23864);
nor U24636 (N_24636,N_23157,N_23054);
or U24637 (N_24637,N_22795,N_23360);
xor U24638 (N_24638,N_22210,N_22068);
or U24639 (N_24639,N_23903,N_22326);
nand U24640 (N_24640,N_22404,N_22186);
and U24641 (N_24641,N_23159,N_22764);
nor U24642 (N_24642,N_23665,N_23765);
nand U24643 (N_24643,N_22423,N_23161);
xnor U24644 (N_24644,N_22687,N_23615);
or U24645 (N_24645,N_22245,N_22499);
nand U24646 (N_24646,N_22327,N_23679);
and U24647 (N_24647,N_22519,N_23760);
nor U24648 (N_24648,N_23043,N_23263);
xnor U24649 (N_24649,N_23067,N_22770);
xor U24650 (N_24650,N_22182,N_23850);
and U24651 (N_24651,N_23514,N_23382);
xnor U24652 (N_24652,N_22825,N_22355);
nor U24653 (N_24653,N_22174,N_22390);
nand U24654 (N_24654,N_22936,N_22145);
xnor U24655 (N_24655,N_23818,N_22004);
nor U24656 (N_24656,N_23803,N_22254);
or U24657 (N_24657,N_22563,N_23723);
nand U24658 (N_24658,N_22459,N_22447);
nand U24659 (N_24659,N_22065,N_23499);
or U24660 (N_24660,N_22090,N_23735);
nand U24661 (N_24661,N_22328,N_22070);
nor U24662 (N_24662,N_23682,N_23082);
or U24663 (N_24663,N_22998,N_22277);
nand U24664 (N_24664,N_23433,N_23588);
and U24665 (N_24665,N_23201,N_22950);
nand U24666 (N_24666,N_22836,N_23107);
xnor U24667 (N_24667,N_23831,N_22028);
or U24668 (N_24668,N_23227,N_22059);
nand U24669 (N_24669,N_22206,N_23877);
nor U24670 (N_24670,N_23624,N_23884);
nor U24671 (N_24671,N_23817,N_23052);
nor U24672 (N_24672,N_22696,N_22681);
or U24673 (N_24673,N_23264,N_23663);
and U24674 (N_24674,N_22414,N_22486);
xnor U24675 (N_24675,N_22023,N_23284);
nor U24676 (N_24676,N_23170,N_22567);
and U24677 (N_24677,N_23848,N_23733);
and U24678 (N_24678,N_22109,N_23593);
nand U24679 (N_24679,N_23081,N_23949);
nor U24680 (N_24680,N_22566,N_23289);
xor U24681 (N_24681,N_22540,N_22445);
or U24682 (N_24682,N_22405,N_22813);
nor U24683 (N_24683,N_23671,N_22885);
and U24684 (N_24684,N_23152,N_23555);
nor U24685 (N_24685,N_23096,N_23989);
xor U24686 (N_24686,N_23172,N_23255);
and U24687 (N_24687,N_22020,N_23842);
nor U24688 (N_24688,N_22614,N_23970);
and U24689 (N_24689,N_23131,N_23109);
xnor U24690 (N_24690,N_22892,N_23364);
nor U24691 (N_24691,N_23406,N_23214);
or U24692 (N_24692,N_22533,N_22470);
and U24693 (N_24693,N_22867,N_23978);
and U24694 (N_24694,N_23388,N_23283);
xnor U24695 (N_24695,N_23633,N_22428);
or U24696 (N_24696,N_22890,N_22932);
nor U24697 (N_24697,N_22226,N_22731);
or U24698 (N_24698,N_22463,N_22434);
or U24699 (N_24699,N_23116,N_22547);
nor U24700 (N_24700,N_22834,N_22103);
nand U24701 (N_24701,N_23209,N_23268);
or U24702 (N_24702,N_22010,N_23605);
and U24703 (N_24703,N_23493,N_23475);
and U24704 (N_24704,N_23677,N_23095);
nand U24705 (N_24705,N_23668,N_23409);
xor U24706 (N_24706,N_22854,N_22469);
or U24707 (N_24707,N_22487,N_22555);
nor U24708 (N_24708,N_23782,N_22476);
and U24709 (N_24709,N_23212,N_22531);
nand U24710 (N_24710,N_23634,N_22773);
nor U24711 (N_24711,N_22521,N_22252);
and U24712 (N_24712,N_23298,N_23446);
xor U24713 (N_24713,N_22233,N_22443);
nor U24714 (N_24714,N_23387,N_22880);
and U24715 (N_24715,N_22919,N_23786);
and U24716 (N_24716,N_22510,N_23762);
or U24717 (N_24717,N_22049,N_22106);
xnor U24718 (N_24718,N_23569,N_22635);
and U24719 (N_24719,N_22847,N_23726);
xor U24720 (N_24720,N_22668,N_22679);
nor U24721 (N_24721,N_22507,N_23686);
nor U24722 (N_24722,N_22359,N_23516);
nor U24723 (N_24723,N_23572,N_23918);
nand U24724 (N_24724,N_23709,N_23592);
nand U24725 (N_24725,N_22335,N_23124);
xnor U24726 (N_24726,N_22961,N_22630);
nand U24727 (N_24727,N_22924,N_23328);
or U24728 (N_24728,N_22216,N_23314);
or U24729 (N_24729,N_23806,N_23338);
nor U24730 (N_24730,N_23548,N_22422);
or U24731 (N_24731,N_22111,N_23578);
or U24732 (N_24732,N_23010,N_23238);
and U24733 (N_24733,N_22243,N_22783);
xor U24734 (N_24734,N_22869,N_23947);
and U24735 (N_24735,N_23889,N_22262);
nand U24736 (N_24736,N_23567,N_23343);
xor U24737 (N_24737,N_22001,N_23560);
or U24738 (N_24738,N_23647,N_23013);
and U24739 (N_24739,N_23068,N_23819);
or U24740 (N_24740,N_23689,N_22528);
nand U24741 (N_24741,N_22063,N_22522);
nand U24742 (N_24742,N_23158,N_23913);
xor U24743 (N_24743,N_22071,N_22403);
xnor U24744 (N_24744,N_23303,N_23271);
or U24745 (N_24745,N_23822,N_22350);
or U24746 (N_24746,N_23438,N_23123);
or U24747 (N_24747,N_22117,N_22317);
or U24748 (N_24748,N_23370,N_23246);
and U24749 (N_24749,N_22341,N_22725);
and U24750 (N_24750,N_23331,N_23276);
and U24751 (N_24751,N_22653,N_23003);
xnor U24752 (N_24752,N_23764,N_23753);
or U24753 (N_24753,N_23964,N_22769);
or U24754 (N_24754,N_22816,N_23935);
and U24755 (N_24755,N_23408,N_22912);
or U24756 (N_24756,N_23150,N_22220);
nand U24757 (N_24757,N_23146,N_23812);
nand U24758 (N_24758,N_23907,N_23800);
and U24759 (N_24759,N_23429,N_23189);
nor U24760 (N_24760,N_22217,N_22054);
xor U24761 (N_24761,N_22084,N_22379);
nand U24762 (N_24762,N_23434,N_22461);
or U24763 (N_24763,N_23637,N_22279);
nand U24764 (N_24764,N_23880,N_22029);
and U24765 (N_24765,N_22689,N_23118);
nor U24766 (N_24766,N_22746,N_22833);
or U24767 (N_24767,N_22568,N_23224);
nand U24768 (N_24768,N_22231,N_22518);
nor U24769 (N_24769,N_23326,N_22464);
or U24770 (N_24770,N_22008,N_23612);
and U24771 (N_24771,N_23055,N_23423);
nand U24772 (N_24772,N_23968,N_22896);
nor U24773 (N_24773,N_22490,N_23129);
and U24774 (N_24774,N_23001,N_23617);
nand U24775 (N_24775,N_23290,N_23281);
or U24776 (N_24776,N_23065,N_23950);
and U24777 (N_24777,N_23104,N_23865);
nor U24778 (N_24778,N_22257,N_23785);
nor U24779 (N_24779,N_23974,N_23862);
or U24780 (N_24780,N_23397,N_22796);
or U24781 (N_24781,N_23501,N_22113);
nor U24782 (N_24782,N_22747,N_22627);
xnor U24783 (N_24783,N_22153,N_23594);
nor U24784 (N_24784,N_23807,N_22905);
and U24785 (N_24785,N_23837,N_22482);
xnor U24786 (N_24786,N_22544,N_23756);
xnor U24787 (N_24787,N_22241,N_23674);
nand U24788 (N_24788,N_23770,N_23824);
nor U24789 (N_24789,N_23070,N_23273);
or U24790 (N_24790,N_23218,N_22642);
xor U24791 (N_24791,N_22281,N_23373);
nor U24792 (N_24792,N_22580,N_22638);
and U24793 (N_24793,N_22110,N_23196);
nor U24794 (N_24794,N_23993,N_23128);
nor U24795 (N_24795,N_23857,N_23887);
and U24796 (N_24796,N_22525,N_22933);
or U24797 (N_24797,N_22042,N_22756);
xnor U24798 (N_24798,N_22535,N_22320);
nor U24799 (N_24799,N_22512,N_22078);
xnor U24800 (N_24800,N_23571,N_23393);
nor U24801 (N_24801,N_23966,N_23419);
nor U24802 (N_24802,N_22785,N_22934);
or U24803 (N_24803,N_23248,N_22005);
nor U24804 (N_24804,N_23937,N_23986);
or U24805 (N_24805,N_23797,N_22205);
nor U24806 (N_24806,N_22664,N_22585);
nand U24807 (N_24807,N_23794,N_22342);
nand U24808 (N_24808,N_23724,N_22548);
nand U24809 (N_24809,N_23174,N_22513);
or U24810 (N_24810,N_23923,N_22091);
nand U24811 (N_24811,N_23557,N_22925);
or U24812 (N_24812,N_22792,N_22425);
nand U24813 (N_24813,N_23367,N_22451);
xnor U24814 (N_24814,N_22296,N_22964);
xnor U24815 (N_24815,N_22754,N_22158);
nand U24816 (N_24816,N_22125,N_23963);
and U24817 (N_24817,N_22902,N_22899);
nand U24818 (N_24818,N_22275,N_22562);
xor U24819 (N_24819,N_22235,N_23598);
or U24820 (N_24820,N_23177,N_23440);
or U24821 (N_24821,N_22144,N_22035);
xnor U24822 (N_24822,N_22597,N_23618);
nand U24823 (N_24823,N_23716,N_22879);
and U24824 (N_24824,N_23302,N_23256);
and U24825 (N_24825,N_22107,N_22409);
xor U24826 (N_24826,N_23855,N_23369);
or U24827 (N_24827,N_23454,N_22303);
nor U24828 (N_24828,N_22419,N_23492);
nor U24829 (N_24829,N_22782,N_23738);
and U24830 (N_24830,N_23629,N_23563);
or U24831 (N_24831,N_22085,N_23698);
or U24832 (N_24832,N_22903,N_23614);
or U24833 (N_24833,N_22572,N_22716);
nand U24834 (N_24834,N_22361,N_22354);
and U24835 (N_24835,N_22559,N_22116);
nand U24836 (N_24836,N_23956,N_23838);
nor U24837 (N_24837,N_22195,N_23035);
or U24838 (N_24838,N_23412,N_22314);
and U24839 (N_24839,N_22180,N_23004);
nor U24840 (N_24840,N_22692,N_22617);
nand U24841 (N_24841,N_22780,N_22748);
nor U24842 (N_24842,N_22339,N_23405);
and U24843 (N_24843,N_23394,N_22381);
nor U24844 (N_24844,N_22868,N_22608);
nand U24845 (N_24845,N_22043,N_23135);
and U24846 (N_24846,N_22399,N_22265);
xor U24847 (N_24847,N_22102,N_23386);
nor U24848 (N_24848,N_23997,N_22778);
and U24849 (N_24849,N_22142,N_22920);
nor U24850 (N_24850,N_22910,N_22815);
nand U24851 (N_24851,N_23120,N_22357);
nand U24852 (N_24852,N_23643,N_23507);
and U24853 (N_24853,N_22351,N_22127);
xnor U24854 (N_24854,N_22803,N_23002);
and U24855 (N_24855,N_22742,N_23718);
or U24856 (N_24856,N_22708,N_23816);
nor U24857 (N_24857,N_22840,N_23311);
xor U24858 (N_24858,N_22786,N_23345);
nand U24859 (N_24859,N_23477,N_23154);
xor U24860 (N_24860,N_23383,N_23879);
or U24861 (N_24861,N_22179,N_22981);
or U24862 (N_24862,N_23279,N_22312);
or U24863 (N_24863,N_22564,N_22893);
xor U24864 (N_24864,N_22736,N_23402);
nand U24865 (N_24865,N_22710,N_23914);
nor U24866 (N_24866,N_22691,N_22002);
and U24867 (N_24867,N_22038,N_22701);
nand U24868 (N_24868,N_22356,N_23754);
or U24869 (N_24869,N_22973,N_22069);
xnor U24870 (N_24870,N_23134,N_22605);
nor U24871 (N_24871,N_23137,N_23073);
nor U24872 (N_24872,N_22467,N_23425);
nand U24873 (N_24873,N_22064,N_23936);
nand U24874 (N_24874,N_22246,N_23768);
nand U24875 (N_24875,N_22678,N_22212);
and U24876 (N_24876,N_22146,N_23661);
nand U24877 (N_24877,N_22875,N_23299);
nor U24878 (N_24878,N_22026,N_22762);
and U24879 (N_24879,N_22504,N_23659);
nand U24880 (N_24880,N_22991,N_22015);
xor U24881 (N_24881,N_22433,N_23481);
xor U24882 (N_24882,N_22861,N_23522);
xnor U24883 (N_24883,N_23911,N_22298);
nor U24884 (N_24884,N_22021,N_23872);
xor U24885 (N_24885,N_22251,N_22644);
nand U24886 (N_24886,N_22918,N_23603);
nand U24887 (N_24887,N_22353,N_23792);
nand U24888 (N_24888,N_22292,N_22543);
and U24889 (N_24889,N_23125,N_23417);
and U24890 (N_24890,N_23623,N_23047);
nand U24891 (N_24891,N_23401,N_22594);
xor U24892 (N_24892,N_23030,N_22709);
nor U24893 (N_24893,N_23473,N_23579);
nand U24894 (N_24894,N_22621,N_23365);
nand U24895 (N_24895,N_23636,N_23895);
and U24896 (N_24896,N_23832,N_22310);
xnor U24897 (N_24897,N_22075,N_22789);
nand U24898 (N_24898,N_22377,N_22992);
and U24899 (N_24899,N_23915,N_23228);
and U24900 (N_24900,N_22943,N_22006);
or U24901 (N_24901,N_22176,N_23690);
or U24902 (N_24902,N_23702,N_22944);
or U24903 (N_24903,N_23814,N_23431);
nand U24904 (N_24904,N_23442,N_23243);
nor U24905 (N_24905,N_23755,N_22760);
nand U24906 (N_24906,N_22204,N_22539);
nor U24907 (N_24907,N_23960,N_23729);
nor U24908 (N_24908,N_22898,N_22826);
and U24909 (N_24909,N_22104,N_23640);
nor U24910 (N_24910,N_22297,N_23772);
or U24911 (N_24911,N_23789,N_23604);
nand U24912 (N_24912,N_23031,N_23628);
nor U24913 (N_24913,N_23708,N_22378);
and U24914 (N_24914,N_22349,N_22829);
nand U24915 (N_24915,N_23621,N_23036);
xnor U24916 (N_24916,N_22268,N_23607);
or U24917 (N_24917,N_22286,N_23761);
xnor U24918 (N_24918,N_23160,N_23333);
nand U24919 (N_24919,N_22395,N_23319);
or U24920 (N_24920,N_23087,N_23849);
or U24921 (N_24921,N_23366,N_22067);
or U24922 (N_24922,N_23074,N_22082);
or U24923 (N_24923,N_23115,N_22076);
nand U24924 (N_24924,N_22032,N_22809);
nor U24925 (N_24925,N_22416,N_23591);
xor U24926 (N_24926,N_23869,N_23602);
or U24927 (N_24927,N_23905,N_23085);
xnor U24928 (N_24928,N_22260,N_22057);
nor U24929 (N_24929,N_23190,N_23427);
nand U24930 (N_24930,N_23527,N_22108);
nor U24931 (N_24931,N_23829,N_22646);
xor U24932 (N_24932,N_22984,N_22036);
xor U24933 (N_24933,N_22478,N_22452);
nand U24934 (N_24934,N_22777,N_22873);
and U24935 (N_24935,N_22421,N_23282);
or U24936 (N_24936,N_23717,N_23398);
nand U24937 (N_24937,N_23777,N_22278);
xnor U24938 (N_24938,N_22468,N_22311);
xor U24939 (N_24939,N_22822,N_23536);
and U24940 (N_24940,N_22321,N_23596);
nor U24941 (N_24941,N_22520,N_22319);
or U24942 (N_24942,N_22284,N_23790);
xor U24943 (N_24943,N_23796,N_22446);
or U24944 (N_24944,N_23353,N_23763);
xor U24945 (N_24945,N_22904,N_22120);
and U24946 (N_24946,N_22223,N_23204);
and U24947 (N_24947,N_22676,N_23921);
xor U24948 (N_24948,N_23896,N_23226);
or U24949 (N_24949,N_22493,N_23931);
or U24950 (N_24950,N_22593,N_22558);
nor U24951 (N_24951,N_23815,N_22790);
xnor U24952 (N_24952,N_23948,N_22406);
nand U24953 (N_24953,N_23399,N_22480);
nor U24954 (N_24954,N_22417,N_23513);
and U24955 (N_24955,N_22352,N_22882);
nor U24956 (N_24956,N_23990,N_23543);
or U24957 (N_24957,N_22808,N_22999);
xnor U24958 (N_24958,N_23565,N_22213);
or U24959 (N_24959,N_22373,N_22982);
and U24960 (N_24960,N_23287,N_23810);
and U24961 (N_24961,N_22450,N_22397);
nand U24962 (N_24962,N_22460,N_23187);
nor U24963 (N_24963,N_22979,N_22229);
nor U24964 (N_24964,N_22431,N_22655);
nor U24965 (N_24965,N_22949,N_23479);
nand U24966 (N_24966,N_22553,N_22141);
and U24967 (N_24967,N_23809,N_22150);
and U24968 (N_24968,N_22249,N_22096);
nor U24969 (N_24969,N_22263,N_22362);
and U24970 (N_24970,N_22393,N_23413);
xor U24971 (N_24971,N_23625,N_23318);
xor U24972 (N_24972,N_22426,N_23269);
nand U24973 (N_24973,N_23749,N_23487);
nand U24974 (N_24974,N_22386,N_23057);
and U24975 (N_24975,N_23195,N_22457);
xnor U24976 (N_24976,N_22302,N_22699);
and U24977 (N_24977,N_23924,N_23126);
xnor U24978 (N_24978,N_22931,N_23672);
xnor U24979 (N_24979,N_22870,N_22313);
and U24980 (N_24980,N_22884,N_22859);
or U24981 (N_24981,N_22122,N_23453);
or U24982 (N_24982,N_23959,N_23304);
and U24983 (N_24983,N_22282,N_23017);
or U24984 (N_24984,N_23285,N_22849);
and U24985 (N_24985,N_22003,N_23610);
xor U24986 (N_24986,N_22440,N_23167);
and U24987 (N_24987,N_22209,N_22977);
or U24988 (N_24988,N_22509,N_23845);
and U24989 (N_24989,N_23577,N_22197);
xor U24990 (N_24990,N_23048,N_22234);
and U24991 (N_24991,N_22788,N_22024);
xnor U24992 (N_24992,N_22591,N_22774);
nand U24993 (N_24993,N_23354,N_23752);
nor U24994 (N_24994,N_22322,N_22289);
xor U24995 (N_24995,N_23946,N_23092);
nand U24996 (N_24996,N_22549,N_23041);
or U24997 (N_24997,N_23766,N_23691);
and U24998 (N_24998,N_22649,N_23642);
nor U24999 (N_24999,N_23027,N_22396);
nor U25000 (N_25000,N_22600,N_22920);
xnor U25001 (N_25001,N_23307,N_22451);
or U25002 (N_25002,N_23279,N_23347);
or U25003 (N_25003,N_22699,N_23580);
nand U25004 (N_25004,N_22937,N_22218);
nand U25005 (N_25005,N_22030,N_23699);
or U25006 (N_25006,N_23166,N_23356);
xnor U25007 (N_25007,N_23186,N_23753);
nor U25008 (N_25008,N_22761,N_23935);
xor U25009 (N_25009,N_23709,N_22937);
nor U25010 (N_25010,N_23676,N_23004);
nand U25011 (N_25011,N_22139,N_22696);
or U25012 (N_25012,N_22490,N_22296);
xor U25013 (N_25013,N_23509,N_23167);
and U25014 (N_25014,N_22402,N_23029);
or U25015 (N_25015,N_22864,N_22255);
or U25016 (N_25016,N_23602,N_23796);
xnor U25017 (N_25017,N_23431,N_22954);
nor U25018 (N_25018,N_22953,N_22427);
and U25019 (N_25019,N_22751,N_22863);
nand U25020 (N_25020,N_22586,N_22619);
nand U25021 (N_25021,N_23619,N_23493);
and U25022 (N_25022,N_23425,N_22274);
nor U25023 (N_25023,N_22864,N_23488);
nor U25024 (N_25024,N_22581,N_23223);
and U25025 (N_25025,N_22419,N_22941);
nand U25026 (N_25026,N_23398,N_22123);
or U25027 (N_25027,N_23518,N_23606);
nand U25028 (N_25028,N_23568,N_22276);
or U25029 (N_25029,N_22997,N_22789);
nor U25030 (N_25030,N_22616,N_22964);
xnor U25031 (N_25031,N_22840,N_22671);
xnor U25032 (N_25032,N_22329,N_22888);
nor U25033 (N_25033,N_22512,N_23774);
xor U25034 (N_25034,N_23464,N_22692);
nand U25035 (N_25035,N_23614,N_22915);
xnor U25036 (N_25036,N_23713,N_23352);
or U25037 (N_25037,N_22821,N_22455);
and U25038 (N_25038,N_23707,N_22770);
xor U25039 (N_25039,N_22079,N_23187);
or U25040 (N_25040,N_22105,N_22031);
or U25041 (N_25041,N_22723,N_22084);
and U25042 (N_25042,N_22624,N_23295);
nand U25043 (N_25043,N_23653,N_23081);
nand U25044 (N_25044,N_23842,N_22893);
and U25045 (N_25045,N_22241,N_23968);
and U25046 (N_25046,N_23539,N_23788);
nand U25047 (N_25047,N_22537,N_23604);
nand U25048 (N_25048,N_22390,N_22347);
nor U25049 (N_25049,N_23566,N_23921);
and U25050 (N_25050,N_22565,N_22872);
or U25051 (N_25051,N_23201,N_23901);
nand U25052 (N_25052,N_22105,N_22448);
and U25053 (N_25053,N_22596,N_23376);
and U25054 (N_25054,N_23414,N_23511);
nor U25055 (N_25055,N_23571,N_23567);
nor U25056 (N_25056,N_22273,N_22592);
nand U25057 (N_25057,N_23528,N_23274);
and U25058 (N_25058,N_23771,N_22466);
or U25059 (N_25059,N_22818,N_23008);
xnor U25060 (N_25060,N_23749,N_22362);
or U25061 (N_25061,N_22341,N_23219);
nor U25062 (N_25062,N_23955,N_22879);
nor U25063 (N_25063,N_22091,N_23079);
or U25064 (N_25064,N_22353,N_23658);
nand U25065 (N_25065,N_22895,N_23947);
nand U25066 (N_25066,N_23584,N_22331);
nand U25067 (N_25067,N_23089,N_23444);
xor U25068 (N_25068,N_22230,N_23127);
and U25069 (N_25069,N_22235,N_22920);
nor U25070 (N_25070,N_23539,N_22753);
or U25071 (N_25071,N_22629,N_23929);
xor U25072 (N_25072,N_22200,N_22385);
and U25073 (N_25073,N_23064,N_23476);
xnor U25074 (N_25074,N_23750,N_23702);
nand U25075 (N_25075,N_22177,N_22496);
nor U25076 (N_25076,N_22122,N_22390);
nand U25077 (N_25077,N_22910,N_22631);
xor U25078 (N_25078,N_23503,N_22177);
or U25079 (N_25079,N_23325,N_23197);
or U25080 (N_25080,N_23780,N_22852);
xnor U25081 (N_25081,N_23886,N_22529);
xnor U25082 (N_25082,N_23446,N_22555);
nand U25083 (N_25083,N_22369,N_23704);
nand U25084 (N_25084,N_23198,N_22635);
nor U25085 (N_25085,N_23757,N_23024);
or U25086 (N_25086,N_23280,N_22033);
nor U25087 (N_25087,N_23766,N_22300);
xor U25088 (N_25088,N_22410,N_22974);
and U25089 (N_25089,N_22855,N_23353);
xor U25090 (N_25090,N_23785,N_22025);
and U25091 (N_25091,N_23176,N_22446);
xnor U25092 (N_25092,N_22006,N_22708);
nor U25093 (N_25093,N_23308,N_23361);
xnor U25094 (N_25094,N_23167,N_22857);
xor U25095 (N_25095,N_22721,N_22445);
nand U25096 (N_25096,N_22407,N_22826);
and U25097 (N_25097,N_23362,N_23357);
nor U25098 (N_25098,N_22764,N_22353);
and U25099 (N_25099,N_23460,N_23845);
nor U25100 (N_25100,N_23330,N_22510);
nand U25101 (N_25101,N_23856,N_22999);
nand U25102 (N_25102,N_22708,N_23038);
and U25103 (N_25103,N_23381,N_22815);
xnor U25104 (N_25104,N_23062,N_22185);
nand U25105 (N_25105,N_22886,N_22874);
nor U25106 (N_25106,N_23047,N_23727);
or U25107 (N_25107,N_22056,N_22221);
or U25108 (N_25108,N_22463,N_22578);
and U25109 (N_25109,N_23279,N_22933);
nor U25110 (N_25110,N_22902,N_22228);
and U25111 (N_25111,N_22135,N_22353);
xnor U25112 (N_25112,N_23720,N_22923);
or U25113 (N_25113,N_22603,N_23905);
nand U25114 (N_25114,N_22920,N_22514);
nor U25115 (N_25115,N_23304,N_22457);
nand U25116 (N_25116,N_23403,N_22158);
nor U25117 (N_25117,N_23274,N_23430);
nand U25118 (N_25118,N_22679,N_22433);
nand U25119 (N_25119,N_22335,N_22917);
nor U25120 (N_25120,N_22783,N_23315);
and U25121 (N_25121,N_23281,N_22612);
or U25122 (N_25122,N_22289,N_22781);
xor U25123 (N_25123,N_22770,N_22135);
and U25124 (N_25124,N_22897,N_22849);
and U25125 (N_25125,N_22708,N_23579);
xor U25126 (N_25126,N_23941,N_22014);
xor U25127 (N_25127,N_22684,N_23161);
or U25128 (N_25128,N_23382,N_23955);
nor U25129 (N_25129,N_22784,N_23613);
nor U25130 (N_25130,N_22206,N_22074);
and U25131 (N_25131,N_22153,N_23378);
nor U25132 (N_25132,N_23620,N_23758);
nand U25133 (N_25133,N_22529,N_22568);
nand U25134 (N_25134,N_22962,N_23340);
and U25135 (N_25135,N_23478,N_22243);
or U25136 (N_25136,N_22858,N_22963);
nand U25137 (N_25137,N_22846,N_23641);
xor U25138 (N_25138,N_22628,N_22322);
nor U25139 (N_25139,N_22239,N_22261);
nand U25140 (N_25140,N_22582,N_23822);
and U25141 (N_25141,N_23376,N_22881);
nor U25142 (N_25142,N_22044,N_23762);
or U25143 (N_25143,N_22989,N_22058);
xnor U25144 (N_25144,N_23057,N_22373);
nand U25145 (N_25145,N_22715,N_23484);
or U25146 (N_25146,N_22289,N_23731);
xnor U25147 (N_25147,N_22262,N_22229);
or U25148 (N_25148,N_23255,N_22768);
or U25149 (N_25149,N_22544,N_22866);
nor U25150 (N_25150,N_23123,N_22223);
or U25151 (N_25151,N_22269,N_23628);
xnor U25152 (N_25152,N_23755,N_23334);
nand U25153 (N_25153,N_22266,N_22929);
nand U25154 (N_25154,N_22968,N_22518);
nor U25155 (N_25155,N_22213,N_23230);
nor U25156 (N_25156,N_22843,N_23200);
or U25157 (N_25157,N_22248,N_22603);
xor U25158 (N_25158,N_22508,N_23426);
and U25159 (N_25159,N_22524,N_23339);
nor U25160 (N_25160,N_23205,N_23727);
or U25161 (N_25161,N_22582,N_23893);
or U25162 (N_25162,N_23671,N_22232);
xor U25163 (N_25163,N_23035,N_23546);
or U25164 (N_25164,N_22856,N_23278);
xnor U25165 (N_25165,N_22727,N_23058);
xnor U25166 (N_25166,N_22365,N_22716);
xor U25167 (N_25167,N_22491,N_22241);
nor U25168 (N_25168,N_23294,N_23754);
xnor U25169 (N_25169,N_23072,N_22385);
xnor U25170 (N_25170,N_23860,N_23880);
nor U25171 (N_25171,N_22825,N_23153);
nand U25172 (N_25172,N_23264,N_23470);
nand U25173 (N_25173,N_22887,N_23567);
xor U25174 (N_25174,N_22151,N_23584);
nor U25175 (N_25175,N_23495,N_23894);
xor U25176 (N_25176,N_22852,N_22729);
and U25177 (N_25177,N_22127,N_22162);
and U25178 (N_25178,N_23245,N_23124);
nor U25179 (N_25179,N_23621,N_22872);
xnor U25180 (N_25180,N_23081,N_22612);
xor U25181 (N_25181,N_22387,N_22812);
or U25182 (N_25182,N_23686,N_22479);
nor U25183 (N_25183,N_22536,N_23292);
and U25184 (N_25184,N_22887,N_23576);
nor U25185 (N_25185,N_23771,N_22486);
or U25186 (N_25186,N_23730,N_22035);
xnor U25187 (N_25187,N_23871,N_22879);
nand U25188 (N_25188,N_23917,N_23958);
nor U25189 (N_25189,N_22889,N_23624);
nand U25190 (N_25190,N_23191,N_22842);
xor U25191 (N_25191,N_22044,N_23605);
xor U25192 (N_25192,N_23684,N_23582);
and U25193 (N_25193,N_23624,N_23921);
xnor U25194 (N_25194,N_23292,N_23459);
and U25195 (N_25195,N_22555,N_22710);
xor U25196 (N_25196,N_23033,N_22221);
nand U25197 (N_25197,N_22473,N_23341);
and U25198 (N_25198,N_22230,N_23810);
nor U25199 (N_25199,N_23831,N_22477);
and U25200 (N_25200,N_22935,N_22244);
nand U25201 (N_25201,N_23885,N_23177);
nor U25202 (N_25202,N_23834,N_23918);
or U25203 (N_25203,N_23905,N_22537);
and U25204 (N_25204,N_22172,N_22655);
nand U25205 (N_25205,N_22748,N_23413);
nand U25206 (N_25206,N_22242,N_22484);
or U25207 (N_25207,N_22333,N_23904);
and U25208 (N_25208,N_22755,N_22649);
or U25209 (N_25209,N_23258,N_23753);
nand U25210 (N_25210,N_23607,N_22637);
xor U25211 (N_25211,N_23422,N_22508);
and U25212 (N_25212,N_23459,N_22572);
and U25213 (N_25213,N_22850,N_22625);
nor U25214 (N_25214,N_22248,N_23678);
nor U25215 (N_25215,N_22394,N_23809);
xor U25216 (N_25216,N_22845,N_22507);
xnor U25217 (N_25217,N_23505,N_22529);
xor U25218 (N_25218,N_22619,N_22205);
nor U25219 (N_25219,N_23064,N_22102);
or U25220 (N_25220,N_22744,N_23625);
and U25221 (N_25221,N_22417,N_23495);
and U25222 (N_25222,N_23580,N_22720);
xnor U25223 (N_25223,N_23094,N_23989);
and U25224 (N_25224,N_23029,N_23911);
and U25225 (N_25225,N_23273,N_22877);
nor U25226 (N_25226,N_22547,N_23843);
and U25227 (N_25227,N_22273,N_22439);
or U25228 (N_25228,N_22992,N_23504);
nand U25229 (N_25229,N_23186,N_23330);
nor U25230 (N_25230,N_22286,N_23440);
nand U25231 (N_25231,N_23473,N_22167);
nor U25232 (N_25232,N_22735,N_23258);
and U25233 (N_25233,N_22705,N_23148);
and U25234 (N_25234,N_23253,N_23496);
or U25235 (N_25235,N_23822,N_23170);
nor U25236 (N_25236,N_23527,N_23170);
nand U25237 (N_25237,N_22329,N_23886);
nor U25238 (N_25238,N_22677,N_22047);
xor U25239 (N_25239,N_23520,N_23312);
xnor U25240 (N_25240,N_23296,N_22597);
xor U25241 (N_25241,N_23156,N_23436);
nor U25242 (N_25242,N_23087,N_22866);
xnor U25243 (N_25243,N_22810,N_22782);
nand U25244 (N_25244,N_22171,N_22331);
nand U25245 (N_25245,N_23708,N_23793);
nor U25246 (N_25246,N_23462,N_22944);
and U25247 (N_25247,N_23409,N_23382);
xor U25248 (N_25248,N_23249,N_23315);
nand U25249 (N_25249,N_23225,N_22829);
xor U25250 (N_25250,N_23165,N_23193);
xor U25251 (N_25251,N_22777,N_23769);
xor U25252 (N_25252,N_23674,N_23813);
and U25253 (N_25253,N_22719,N_22836);
xnor U25254 (N_25254,N_22159,N_23620);
and U25255 (N_25255,N_23462,N_22855);
nor U25256 (N_25256,N_23242,N_23192);
or U25257 (N_25257,N_23903,N_23234);
or U25258 (N_25258,N_22389,N_22929);
nand U25259 (N_25259,N_22995,N_22923);
nor U25260 (N_25260,N_22399,N_22169);
and U25261 (N_25261,N_22951,N_23145);
nor U25262 (N_25262,N_23738,N_22025);
xnor U25263 (N_25263,N_23522,N_23626);
or U25264 (N_25264,N_23222,N_23959);
or U25265 (N_25265,N_23739,N_23168);
and U25266 (N_25266,N_22829,N_23297);
xnor U25267 (N_25267,N_23789,N_22163);
nor U25268 (N_25268,N_23556,N_22720);
or U25269 (N_25269,N_23702,N_22821);
nand U25270 (N_25270,N_22642,N_22490);
nor U25271 (N_25271,N_23376,N_23504);
nor U25272 (N_25272,N_23262,N_22072);
nor U25273 (N_25273,N_22931,N_23717);
and U25274 (N_25274,N_22541,N_23513);
nand U25275 (N_25275,N_22939,N_22683);
xnor U25276 (N_25276,N_23848,N_23103);
nor U25277 (N_25277,N_23399,N_23330);
nand U25278 (N_25278,N_23869,N_22847);
and U25279 (N_25279,N_23597,N_22944);
or U25280 (N_25280,N_23702,N_23864);
and U25281 (N_25281,N_22549,N_22389);
nor U25282 (N_25282,N_23012,N_23243);
and U25283 (N_25283,N_22741,N_22311);
nor U25284 (N_25284,N_22652,N_23152);
nor U25285 (N_25285,N_22308,N_23026);
nand U25286 (N_25286,N_23658,N_22851);
nor U25287 (N_25287,N_22904,N_22619);
xor U25288 (N_25288,N_22585,N_23394);
nand U25289 (N_25289,N_23878,N_23256);
nand U25290 (N_25290,N_22990,N_22552);
and U25291 (N_25291,N_22451,N_22967);
nand U25292 (N_25292,N_23316,N_23394);
nor U25293 (N_25293,N_22146,N_22864);
xnor U25294 (N_25294,N_22890,N_23819);
nand U25295 (N_25295,N_23564,N_22280);
nor U25296 (N_25296,N_23815,N_22588);
nor U25297 (N_25297,N_23021,N_22738);
or U25298 (N_25298,N_23322,N_22349);
nand U25299 (N_25299,N_22880,N_22518);
nand U25300 (N_25300,N_23289,N_22768);
or U25301 (N_25301,N_23638,N_22968);
and U25302 (N_25302,N_23534,N_23574);
and U25303 (N_25303,N_22309,N_22094);
nor U25304 (N_25304,N_23881,N_23590);
nand U25305 (N_25305,N_22074,N_22993);
or U25306 (N_25306,N_22868,N_23335);
nor U25307 (N_25307,N_22940,N_23008);
or U25308 (N_25308,N_23962,N_22715);
xnor U25309 (N_25309,N_23477,N_22712);
nor U25310 (N_25310,N_23743,N_23423);
nand U25311 (N_25311,N_23512,N_22370);
or U25312 (N_25312,N_22295,N_23463);
and U25313 (N_25313,N_23849,N_23158);
or U25314 (N_25314,N_22802,N_23722);
xnor U25315 (N_25315,N_22982,N_23317);
and U25316 (N_25316,N_22323,N_23265);
nor U25317 (N_25317,N_22288,N_22747);
nor U25318 (N_25318,N_23221,N_22073);
nand U25319 (N_25319,N_23977,N_22511);
and U25320 (N_25320,N_23474,N_23632);
or U25321 (N_25321,N_23112,N_22826);
or U25322 (N_25322,N_22988,N_23054);
nor U25323 (N_25323,N_22760,N_22171);
nor U25324 (N_25324,N_23509,N_23704);
or U25325 (N_25325,N_22388,N_23645);
and U25326 (N_25326,N_22683,N_22858);
or U25327 (N_25327,N_22365,N_22836);
or U25328 (N_25328,N_22696,N_23058);
nand U25329 (N_25329,N_23789,N_22390);
nor U25330 (N_25330,N_23500,N_22795);
xnor U25331 (N_25331,N_23555,N_23610);
nor U25332 (N_25332,N_23045,N_23899);
xnor U25333 (N_25333,N_23489,N_23472);
xnor U25334 (N_25334,N_23314,N_23535);
or U25335 (N_25335,N_22632,N_22112);
xnor U25336 (N_25336,N_22514,N_23830);
nor U25337 (N_25337,N_23637,N_22293);
or U25338 (N_25338,N_22264,N_22029);
and U25339 (N_25339,N_23149,N_22346);
and U25340 (N_25340,N_22537,N_22343);
nor U25341 (N_25341,N_22940,N_22125);
xor U25342 (N_25342,N_22025,N_22925);
or U25343 (N_25343,N_23536,N_22047);
and U25344 (N_25344,N_23125,N_22380);
nor U25345 (N_25345,N_23282,N_22288);
nand U25346 (N_25346,N_22825,N_23744);
nor U25347 (N_25347,N_22735,N_23319);
nor U25348 (N_25348,N_22236,N_23996);
and U25349 (N_25349,N_22721,N_23292);
xnor U25350 (N_25350,N_23560,N_22765);
nor U25351 (N_25351,N_23069,N_23079);
and U25352 (N_25352,N_22703,N_23314);
nand U25353 (N_25353,N_22520,N_22587);
or U25354 (N_25354,N_23707,N_22572);
nor U25355 (N_25355,N_23491,N_23730);
nor U25356 (N_25356,N_22884,N_23916);
nand U25357 (N_25357,N_23320,N_22505);
or U25358 (N_25358,N_23571,N_22444);
xor U25359 (N_25359,N_22612,N_22746);
nand U25360 (N_25360,N_23745,N_23366);
xnor U25361 (N_25361,N_22942,N_23329);
nand U25362 (N_25362,N_23953,N_22853);
xnor U25363 (N_25363,N_22157,N_23196);
xor U25364 (N_25364,N_22183,N_23637);
nor U25365 (N_25365,N_22100,N_22290);
nand U25366 (N_25366,N_23629,N_23672);
nor U25367 (N_25367,N_23618,N_22395);
nor U25368 (N_25368,N_23978,N_23868);
and U25369 (N_25369,N_22235,N_23736);
xnor U25370 (N_25370,N_23719,N_22894);
nor U25371 (N_25371,N_23410,N_23662);
xor U25372 (N_25372,N_23248,N_23900);
and U25373 (N_25373,N_22565,N_23573);
or U25374 (N_25374,N_22323,N_23818);
nand U25375 (N_25375,N_23098,N_23150);
xor U25376 (N_25376,N_22268,N_22590);
nor U25377 (N_25377,N_22990,N_23228);
and U25378 (N_25378,N_23695,N_23309);
xnor U25379 (N_25379,N_22733,N_23282);
or U25380 (N_25380,N_22229,N_23145);
or U25381 (N_25381,N_22333,N_22301);
xor U25382 (N_25382,N_22677,N_23820);
nor U25383 (N_25383,N_22051,N_22877);
or U25384 (N_25384,N_23902,N_22874);
nor U25385 (N_25385,N_22829,N_22353);
and U25386 (N_25386,N_22858,N_23840);
xor U25387 (N_25387,N_22537,N_22908);
nand U25388 (N_25388,N_22145,N_22921);
nand U25389 (N_25389,N_22419,N_23910);
or U25390 (N_25390,N_22261,N_23261);
nor U25391 (N_25391,N_23474,N_22276);
xnor U25392 (N_25392,N_23645,N_22897);
or U25393 (N_25393,N_23125,N_22111);
and U25394 (N_25394,N_23717,N_22819);
and U25395 (N_25395,N_22407,N_22056);
nor U25396 (N_25396,N_23982,N_22426);
nor U25397 (N_25397,N_23675,N_23887);
nand U25398 (N_25398,N_22856,N_23313);
and U25399 (N_25399,N_22727,N_22931);
nand U25400 (N_25400,N_23534,N_22018);
or U25401 (N_25401,N_22448,N_23258);
nor U25402 (N_25402,N_23081,N_22661);
nor U25403 (N_25403,N_23496,N_23685);
nand U25404 (N_25404,N_22783,N_23723);
or U25405 (N_25405,N_22588,N_22173);
xor U25406 (N_25406,N_22455,N_22488);
xor U25407 (N_25407,N_23800,N_23152);
xor U25408 (N_25408,N_22080,N_22733);
xor U25409 (N_25409,N_23033,N_22385);
and U25410 (N_25410,N_23206,N_23529);
nand U25411 (N_25411,N_22033,N_23633);
or U25412 (N_25412,N_22660,N_22670);
or U25413 (N_25413,N_22504,N_23314);
nand U25414 (N_25414,N_23887,N_23297);
nand U25415 (N_25415,N_22925,N_23429);
xnor U25416 (N_25416,N_23293,N_22466);
nand U25417 (N_25417,N_22782,N_23643);
xnor U25418 (N_25418,N_23605,N_23857);
and U25419 (N_25419,N_22677,N_23644);
xnor U25420 (N_25420,N_22791,N_23543);
or U25421 (N_25421,N_22887,N_22319);
or U25422 (N_25422,N_23050,N_23145);
nor U25423 (N_25423,N_22179,N_22386);
or U25424 (N_25424,N_22391,N_23157);
nor U25425 (N_25425,N_22503,N_23688);
nor U25426 (N_25426,N_22148,N_23770);
nand U25427 (N_25427,N_22511,N_23883);
nand U25428 (N_25428,N_22935,N_22451);
and U25429 (N_25429,N_23196,N_23941);
or U25430 (N_25430,N_23841,N_23476);
nand U25431 (N_25431,N_22314,N_22237);
xor U25432 (N_25432,N_23304,N_23143);
xor U25433 (N_25433,N_23870,N_23688);
nor U25434 (N_25434,N_22320,N_23537);
nor U25435 (N_25435,N_23778,N_22650);
nand U25436 (N_25436,N_22088,N_23175);
and U25437 (N_25437,N_23437,N_22881);
xor U25438 (N_25438,N_22460,N_23244);
nor U25439 (N_25439,N_23929,N_23202);
and U25440 (N_25440,N_22076,N_22074);
or U25441 (N_25441,N_23060,N_22405);
nand U25442 (N_25442,N_23468,N_23921);
xor U25443 (N_25443,N_22202,N_23887);
nand U25444 (N_25444,N_23676,N_22894);
nand U25445 (N_25445,N_23395,N_22295);
nor U25446 (N_25446,N_22902,N_23531);
nor U25447 (N_25447,N_22280,N_22030);
nor U25448 (N_25448,N_22685,N_22430);
nor U25449 (N_25449,N_23760,N_23810);
nand U25450 (N_25450,N_23196,N_23587);
nand U25451 (N_25451,N_23657,N_23314);
and U25452 (N_25452,N_22048,N_23932);
xor U25453 (N_25453,N_23322,N_22449);
or U25454 (N_25454,N_22860,N_23926);
and U25455 (N_25455,N_23971,N_23363);
or U25456 (N_25456,N_23332,N_22471);
and U25457 (N_25457,N_23486,N_23260);
xor U25458 (N_25458,N_23522,N_22986);
or U25459 (N_25459,N_22103,N_22275);
and U25460 (N_25460,N_23070,N_22664);
xnor U25461 (N_25461,N_23246,N_22136);
nand U25462 (N_25462,N_22828,N_23357);
nand U25463 (N_25463,N_22823,N_22267);
xnor U25464 (N_25464,N_23960,N_22170);
and U25465 (N_25465,N_23832,N_23050);
xnor U25466 (N_25466,N_23997,N_22289);
or U25467 (N_25467,N_22431,N_22216);
nand U25468 (N_25468,N_22988,N_22895);
xnor U25469 (N_25469,N_23191,N_23576);
xnor U25470 (N_25470,N_23627,N_22427);
xor U25471 (N_25471,N_22524,N_22831);
nor U25472 (N_25472,N_22099,N_22869);
xnor U25473 (N_25473,N_22084,N_22163);
nor U25474 (N_25474,N_23823,N_22731);
nor U25475 (N_25475,N_23628,N_23225);
xnor U25476 (N_25476,N_23076,N_23577);
xnor U25477 (N_25477,N_23794,N_22313);
and U25478 (N_25478,N_22534,N_22570);
nor U25479 (N_25479,N_23945,N_22629);
nand U25480 (N_25480,N_22603,N_22818);
nor U25481 (N_25481,N_23836,N_23097);
xor U25482 (N_25482,N_22357,N_23309);
or U25483 (N_25483,N_23933,N_22462);
xnor U25484 (N_25484,N_22756,N_23146);
and U25485 (N_25485,N_23609,N_23668);
and U25486 (N_25486,N_23778,N_23936);
xor U25487 (N_25487,N_23344,N_22170);
and U25488 (N_25488,N_22142,N_23107);
or U25489 (N_25489,N_23137,N_23093);
nand U25490 (N_25490,N_22691,N_23825);
xor U25491 (N_25491,N_23295,N_23132);
and U25492 (N_25492,N_23229,N_22348);
or U25493 (N_25493,N_22436,N_23972);
and U25494 (N_25494,N_23452,N_22032);
or U25495 (N_25495,N_23347,N_23443);
and U25496 (N_25496,N_22850,N_22130);
xnor U25497 (N_25497,N_22314,N_23464);
nor U25498 (N_25498,N_23863,N_22634);
and U25499 (N_25499,N_23188,N_22194);
nand U25500 (N_25500,N_23120,N_23475);
and U25501 (N_25501,N_23342,N_23899);
nor U25502 (N_25502,N_23678,N_22009);
nor U25503 (N_25503,N_23440,N_22890);
and U25504 (N_25504,N_22620,N_23821);
and U25505 (N_25505,N_22592,N_23932);
xor U25506 (N_25506,N_22850,N_23788);
nand U25507 (N_25507,N_23394,N_22905);
nand U25508 (N_25508,N_23012,N_23291);
and U25509 (N_25509,N_23780,N_22666);
nor U25510 (N_25510,N_23687,N_22767);
nand U25511 (N_25511,N_22703,N_22764);
xnor U25512 (N_25512,N_23358,N_22406);
nor U25513 (N_25513,N_23611,N_23450);
nand U25514 (N_25514,N_23686,N_23440);
or U25515 (N_25515,N_22426,N_23801);
xnor U25516 (N_25516,N_22939,N_22022);
xnor U25517 (N_25517,N_22746,N_23186);
nor U25518 (N_25518,N_22176,N_22665);
nand U25519 (N_25519,N_23463,N_23024);
xor U25520 (N_25520,N_23961,N_23167);
nand U25521 (N_25521,N_23232,N_22308);
and U25522 (N_25522,N_23018,N_22159);
xor U25523 (N_25523,N_22628,N_22838);
nand U25524 (N_25524,N_23952,N_23641);
nand U25525 (N_25525,N_23214,N_22902);
or U25526 (N_25526,N_22706,N_22988);
nor U25527 (N_25527,N_23038,N_23242);
xnor U25528 (N_25528,N_22048,N_22128);
nor U25529 (N_25529,N_23513,N_23490);
nand U25530 (N_25530,N_22671,N_22995);
nand U25531 (N_25531,N_23924,N_23215);
or U25532 (N_25532,N_22744,N_23453);
nand U25533 (N_25533,N_23889,N_23150);
nand U25534 (N_25534,N_23963,N_22325);
and U25535 (N_25535,N_23423,N_23677);
nand U25536 (N_25536,N_23305,N_23414);
xor U25537 (N_25537,N_23431,N_22284);
and U25538 (N_25538,N_23973,N_22377);
nand U25539 (N_25539,N_23680,N_23693);
nand U25540 (N_25540,N_22264,N_22015);
or U25541 (N_25541,N_22247,N_23839);
xor U25542 (N_25542,N_22639,N_23653);
or U25543 (N_25543,N_23909,N_22031);
nor U25544 (N_25544,N_22388,N_22054);
and U25545 (N_25545,N_23065,N_22500);
nor U25546 (N_25546,N_22604,N_23581);
nand U25547 (N_25547,N_22475,N_23587);
and U25548 (N_25548,N_22469,N_23555);
nand U25549 (N_25549,N_22120,N_23711);
nand U25550 (N_25550,N_22499,N_22985);
and U25551 (N_25551,N_23396,N_23646);
and U25552 (N_25552,N_22883,N_23439);
nand U25553 (N_25553,N_23926,N_22897);
nor U25554 (N_25554,N_23538,N_23191);
and U25555 (N_25555,N_22480,N_23523);
and U25556 (N_25556,N_22702,N_23175);
nand U25557 (N_25557,N_23691,N_23379);
xor U25558 (N_25558,N_22248,N_22363);
or U25559 (N_25559,N_22046,N_23726);
xnor U25560 (N_25560,N_22575,N_22867);
nand U25561 (N_25561,N_22631,N_23462);
nor U25562 (N_25562,N_22757,N_22936);
or U25563 (N_25563,N_22325,N_23174);
xor U25564 (N_25564,N_23751,N_23463);
and U25565 (N_25565,N_22759,N_23339);
nor U25566 (N_25566,N_22371,N_22470);
and U25567 (N_25567,N_23971,N_23821);
or U25568 (N_25568,N_22827,N_22818);
or U25569 (N_25569,N_23455,N_22274);
and U25570 (N_25570,N_22896,N_23097);
xor U25571 (N_25571,N_23454,N_23715);
nor U25572 (N_25572,N_22778,N_22055);
and U25573 (N_25573,N_23955,N_23628);
nand U25574 (N_25574,N_23826,N_23920);
nor U25575 (N_25575,N_22589,N_22990);
nand U25576 (N_25576,N_22674,N_22648);
nor U25577 (N_25577,N_22982,N_22480);
xor U25578 (N_25578,N_22429,N_23900);
or U25579 (N_25579,N_23927,N_22643);
and U25580 (N_25580,N_22682,N_22328);
and U25581 (N_25581,N_22118,N_23679);
or U25582 (N_25582,N_22579,N_23484);
xnor U25583 (N_25583,N_22466,N_23615);
nor U25584 (N_25584,N_23049,N_23485);
xor U25585 (N_25585,N_23680,N_23514);
or U25586 (N_25586,N_23095,N_22313);
or U25587 (N_25587,N_22736,N_22379);
xnor U25588 (N_25588,N_22266,N_23464);
nor U25589 (N_25589,N_22562,N_22769);
nand U25590 (N_25590,N_23652,N_22114);
or U25591 (N_25591,N_22379,N_22540);
nor U25592 (N_25592,N_23116,N_22618);
nand U25593 (N_25593,N_22919,N_23412);
nand U25594 (N_25594,N_23028,N_23375);
or U25595 (N_25595,N_22565,N_22086);
and U25596 (N_25596,N_22776,N_22175);
xnor U25597 (N_25597,N_23875,N_23427);
or U25598 (N_25598,N_22771,N_22146);
nand U25599 (N_25599,N_22617,N_22991);
nor U25600 (N_25600,N_22009,N_23886);
nand U25601 (N_25601,N_22328,N_23397);
or U25602 (N_25602,N_22388,N_23016);
and U25603 (N_25603,N_23537,N_22262);
nand U25604 (N_25604,N_22335,N_22937);
and U25605 (N_25605,N_23182,N_22378);
or U25606 (N_25606,N_22703,N_23194);
and U25607 (N_25607,N_22902,N_22701);
and U25608 (N_25608,N_22031,N_22430);
or U25609 (N_25609,N_23643,N_22973);
nand U25610 (N_25610,N_23566,N_23684);
or U25611 (N_25611,N_22695,N_23823);
or U25612 (N_25612,N_22728,N_22477);
or U25613 (N_25613,N_23302,N_23744);
nand U25614 (N_25614,N_22387,N_22273);
or U25615 (N_25615,N_22591,N_22432);
xor U25616 (N_25616,N_22211,N_23319);
or U25617 (N_25617,N_23655,N_23381);
nand U25618 (N_25618,N_23156,N_23306);
or U25619 (N_25619,N_22418,N_23804);
xor U25620 (N_25620,N_23549,N_22818);
xnor U25621 (N_25621,N_22660,N_22803);
nor U25622 (N_25622,N_22496,N_22094);
or U25623 (N_25623,N_22948,N_22237);
nor U25624 (N_25624,N_23898,N_23403);
nand U25625 (N_25625,N_22832,N_22512);
and U25626 (N_25626,N_23731,N_23609);
and U25627 (N_25627,N_22434,N_22155);
and U25628 (N_25628,N_22261,N_22195);
nor U25629 (N_25629,N_22339,N_22037);
and U25630 (N_25630,N_23125,N_23985);
nand U25631 (N_25631,N_22352,N_22698);
or U25632 (N_25632,N_22609,N_23080);
xnor U25633 (N_25633,N_23348,N_23632);
or U25634 (N_25634,N_23197,N_22699);
nor U25635 (N_25635,N_22735,N_23994);
and U25636 (N_25636,N_22711,N_22550);
nand U25637 (N_25637,N_22580,N_22359);
xor U25638 (N_25638,N_22050,N_22901);
xor U25639 (N_25639,N_22757,N_23741);
and U25640 (N_25640,N_22777,N_23307);
nor U25641 (N_25641,N_22655,N_22630);
and U25642 (N_25642,N_23105,N_23721);
nor U25643 (N_25643,N_23466,N_23801);
xor U25644 (N_25644,N_22112,N_23108);
nand U25645 (N_25645,N_22807,N_22765);
nand U25646 (N_25646,N_23490,N_22681);
xnor U25647 (N_25647,N_23881,N_22890);
nor U25648 (N_25648,N_22514,N_23691);
and U25649 (N_25649,N_23331,N_22737);
or U25650 (N_25650,N_23686,N_23857);
nor U25651 (N_25651,N_23885,N_22770);
nand U25652 (N_25652,N_23681,N_23216);
and U25653 (N_25653,N_23076,N_22600);
and U25654 (N_25654,N_22291,N_22934);
xnor U25655 (N_25655,N_22211,N_22995);
and U25656 (N_25656,N_22179,N_23310);
or U25657 (N_25657,N_23606,N_23342);
and U25658 (N_25658,N_22770,N_23149);
nand U25659 (N_25659,N_23285,N_23981);
nand U25660 (N_25660,N_23349,N_22388);
nand U25661 (N_25661,N_22811,N_23856);
nand U25662 (N_25662,N_22648,N_22884);
or U25663 (N_25663,N_23692,N_22887);
and U25664 (N_25664,N_23143,N_22442);
nand U25665 (N_25665,N_23517,N_23430);
or U25666 (N_25666,N_23676,N_23282);
xnor U25667 (N_25667,N_22513,N_23647);
nand U25668 (N_25668,N_23103,N_23883);
nor U25669 (N_25669,N_22787,N_23907);
nor U25670 (N_25670,N_22391,N_23091);
or U25671 (N_25671,N_22924,N_23061);
nor U25672 (N_25672,N_22990,N_22363);
and U25673 (N_25673,N_23048,N_22779);
nand U25674 (N_25674,N_23434,N_23582);
nor U25675 (N_25675,N_23572,N_23713);
xor U25676 (N_25676,N_22177,N_23552);
and U25677 (N_25677,N_23143,N_22540);
nor U25678 (N_25678,N_22103,N_22937);
nand U25679 (N_25679,N_23992,N_23209);
xor U25680 (N_25680,N_22588,N_23902);
nand U25681 (N_25681,N_23048,N_23213);
nand U25682 (N_25682,N_23052,N_23629);
nor U25683 (N_25683,N_22567,N_22275);
nor U25684 (N_25684,N_23610,N_23237);
nor U25685 (N_25685,N_22485,N_23911);
nand U25686 (N_25686,N_23466,N_23783);
or U25687 (N_25687,N_23318,N_23244);
nor U25688 (N_25688,N_22116,N_23915);
and U25689 (N_25689,N_22014,N_23213);
and U25690 (N_25690,N_23257,N_22087);
xor U25691 (N_25691,N_22149,N_22355);
nand U25692 (N_25692,N_22623,N_22920);
nand U25693 (N_25693,N_23824,N_22153);
and U25694 (N_25694,N_23996,N_23015);
or U25695 (N_25695,N_22929,N_22540);
xor U25696 (N_25696,N_23681,N_23187);
nor U25697 (N_25697,N_22871,N_22884);
and U25698 (N_25698,N_23424,N_23993);
nor U25699 (N_25699,N_22260,N_23074);
or U25700 (N_25700,N_23532,N_22375);
nand U25701 (N_25701,N_23932,N_22026);
xnor U25702 (N_25702,N_22211,N_22249);
nand U25703 (N_25703,N_23709,N_22312);
or U25704 (N_25704,N_23811,N_22368);
nor U25705 (N_25705,N_22191,N_22024);
nand U25706 (N_25706,N_22647,N_22725);
xnor U25707 (N_25707,N_22158,N_23851);
or U25708 (N_25708,N_23917,N_22830);
and U25709 (N_25709,N_22348,N_23352);
xor U25710 (N_25710,N_22338,N_23683);
and U25711 (N_25711,N_23366,N_23227);
nand U25712 (N_25712,N_22140,N_22357);
nor U25713 (N_25713,N_23172,N_22516);
and U25714 (N_25714,N_22728,N_22005);
nand U25715 (N_25715,N_23224,N_23145);
or U25716 (N_25716,N_22093,N_23587);
nor U25717 (N_25717,N_23338,N_23312);
or U25718 (N_25718,N_23574,N_23468);
or U25719 (N_25719,N_22401,N_22682);
or U25720 (N_25720,N_22962,N_23686);
nand U25721 (N_25721,N_23130,N_23006);
or U25722 (N_25722,N_22730,N_22157);
nor U25723 (N_25723,N_22466,N_22577);
or U25724 (N_25724,N_23295,N_22660);
or U25725 (N_25725,N_22684,N_22501);
xor U25726 (N_25726,N_22863,N_23109);
xnor U25727 (N_25727,N_23627,N_23355);
and U25728 (N_25728,N_23779,N_22393);
or U25729 (N_25729,N_23667,N_23464);
nor U25730 (N_25730,N_22085,N_22769);
xnor U25731 (N_25731,N_22811,N_22964);
xnor U25732 (N_25732,N_23187,N_23429);
or U25733 (N_25733,N_23493,N_23156);
nor U25734 (N_25734,N_23627,N_22714);
and U25735 (N_25735,N_22108,N_23590);
xnor U25736 (N_25736,N_23471,N_23131);
nand U25737 (N_25737,N_23353,N_23977);
xnor U25738 (N_25738,N_22423,N_22813);
and U25739 (N_25739,N_23396,N_22151);
or U25740 (N_25740,N_22004,N_22660);
nand U25741 (N_25741,N_23032,N_23842);
and U25742 (N_25742,N_22409,N_22635);
or U25743 (N_25743,N_23288,N_22465);
and U25744 (N_25744,N_22072,N_23801);
nand U25745 (N_25745,N_22357,N_23197);
or U25746 (N_25746,N_23193,N_22817);
nand U25747 (N_25747,N_23697,N_23917);
nor U25748 (N_25748,N_23037,N_22945);
and U25749 (N_25749,N_22264,N_23524);
and U25750 (N_25750,N_23666,N_22252);
and U25751 (N_25751,N_22092,N_23523);
and U25752 (N_25752,N_23997,N_22776);
xor U25753 (N_25753,N_23160,N_23714);
xor U25754 (N_25754,N_22428,N_23380);
nor U25755 (N_25755,N_22792,N_23897);
nor U25756 (N_25756,N_23373,N_23582);
nand U25757 (N_25757,N_23093,N_22411);
or U25758 (N_25758,N_22541,N_23361);
xnor U25759 (N_25759,N_22190,N_23061);
and U25760 (N_25760,N_22315,N_22107);
and U25761 (N_25761,N_22886,N_22096);
nand U25762 (N_25762,N_22942,N_22944);
xor U25763 (N_25763,N_23875,N_23578);
and U25764 (N_25764,N_22801,N_23516);
and U25765 (N_25765,N_22064,N_22171);
nand U25766 (N_25766,N_22909,N_22277);
or U25767 (N_25767,N_22977,N_23956);
xor U25768 (N_25768,N_22572,N_23455);
and U25769 (N_25769,N_22843,N_23497);
xor U25770 (N_25770,N_23154,N_23300);
or U25771 (N_25771,N_22345,N_22842);
and U25772 (N_25772,N_23104,N_23430);
xor U25773 (N_25773,N_22938,N_22540);
or U25774 (N_25774,N_23792,N_22431);
or U25775 (N_25775,N_23008,N_22582);
xnor U25776 (N_25776,N_22770,N_23341);
xnor U25777 (N_25777,N_22754,N_22634);
nor U25778 (N_25778,N_23802,N_23457);
xnor U25779 (N_25779,N_23513,N_23574);
xnor U25780 (N_25780,N_23560,N_23542);
nor U25781 (N_25781,N_22724,N_23929);
nor U25782 (N_25782,N_23750,N_22420);
nor U25783 (N_25783,N_22876,N_23225);
and U25784 (N_25784,N_23941,N_22578);
nor U25785 (N_25785,N_22381,N_23011);
and U25786 (N_25786,N_22026,N_23519);
or U25787 (N_25787,N_23800,N_22369);
xnor U25788 (N_25788,N_23853,N_22430);
or U25789 (N_25789,N_22483,N_22004);
and U25790 (N_25790,N_22629,N_22730);
nand U25791 (N_25791,N_23623,N_23187);
xor U25792 (N_25792,N_23894,N_22502);
or U25793 (N_25793,N_23783,N_23089);
nand U25794 (N_25794,N_22458,N_22601);
xor U25795 (N_25795,N_23531,N_23365);
nand U25796 (N_25796,N_23677,N_23608);
nand U25797 (N_25797,N_23536,N_23734);
xor U25798 (N_25798,N_23499,N_22839);
nor U25799 (N_25799,N_23283,N_22602);
and U25800 (N_25800,N_23374,N_23506);
and U25801 (N_25801,N_23651,N_22000);
nor U25802 (N_25802,N_22501,N_23492);
and U25803 (N_25803,N_23058,N_22100);
or U25804 (N_25804,N_23724,N_23680);
nor U25805 (N_25805,N_22417,N_22603);
xor U25806 (N_25806,N_22121,N_22867);
and U25807 (N_25807,N_22387,N_22185);
and U25808 (N_25808,N_22557,N_23534);
and U25809 (N_25809,N_22275,N_23702);
xor U25810 (N_25810,N_22839,N_22849);
xnor U25811 (N_25811,N_23717,N_22949);
nand U25812 (N_25812,N_22690,N_23840);
xor U25813 (N_25813,N_22839,N_23948);
and U25814 (N_25814,N_22934,N_22066);
or U25815 (N_25815,N_22422,N_23039);
nor U25816 (N_25816,N_22387,N_22718);
and U25817 (N_25817,N_23323,N_23610);
and U25818 (N_25818,N_22179,N_23166);
xor U25819 (N_25819,N_22059,N_22257);
nand U25820 (N_25820,N_23196,N_22247);
xor U25821 (N_25821,N_22955,N_22429);
and U25822 (N_25822,N_23444,N_23476);
or U25823 (N_25823,N_23616,N_23410);
or U25824 (N_25824,N_23999,N_23889);
xor U25825 (N_25825,N_23644,N_22442);
and U25826 (N_25826,N_22361,N_23902);
or U25827 (N_25827,N_23780,N_23394);
xnor U25828 (N_25828,N_23545,N_22557);
or U25829 (N_25829,N_22961,N_22312);
nand U25830 (N_25830,N_23866,N_22461);
nand U25831 (N_25831,N_23715,N_22870);
nor U25832 (N_25832,N_23643,N_23348);
xnor U25833 (N_25833,N_22992,N_23700);
and U25834 (N_25834,N_23156,N_22634);
xor U25835 (N_25835,N_23216,N_23952);
and U25836 (N_25836,N_22712,N_23011);
nor U25837 (N_25837,N_22505,N_22518);
xor U25838 (N_25838,N_22864,N_23059);
xnor U25839 (N_25839,N_23789,N_22434);
nand U25840 (N_25840,N_23314,N_22923);
or U25841 (N_25841,N_22821,N_23045);
nand U25842 (N_25842,N_23361,N_22662);
or U25843 (N_25843,N_22383,N_23207);
nand U25844 (N_25844,N_22260,N_23948);
nor U25845 (N_25845,N_23589,N_22161);
nand U25846 (N_25846,N_23818,N_22034);
xor U25847 (N_25847,N_23703,N_22037);
or U25848 (N_25848,N_23338,N_23595);
or U25849 (N_25849,N_23630,N_22045);
and U25850 (N_25850,N_23172,N_22287);
nand U25851 (N_25851,N_22100,N_23957);
or U25852 (N_25852,N_23141,N_22564);
nor U25853 (N_25853,N_22132,N_22435);
nor U25854 (N_25854,N_23787,N_23049);
and U25855 (N_25855,N_22170,N_22122);
and U25856 (N_25856,N_22657,N_22036);
nor U25857 (N_25857,N_22280,N_23460);
nor U25858 (N_25858,N_23421,N_22685);
xnor U25859 (N_25859,N_23464,N_22596);
or U25860 (N_25860,N_22039,N_22458);
and U25861 (N_25861,N_23324,N_22658);
nor U25862 (N_25862,N_22733,N_22669);
xnor U25863 (N_25863,N_23296,N_22824);
xnor U25864 (N_25864,N_23386,N_22750);
xnor U25865 (N_25865,N_22780,N_23692);
or U25866 (N_25866,N_22714,N_22967);
or U25867 (N_25867,N_22126,N_22264);
or U25868 (N_25868,N_22030,N_22008);
and U25869 (N_25869,N_22997,N_23850);
xnor U25870 (N_25870,N_22105,N_23072);
nand U25871 (N_25871,N_23818,N_22211);
nor U25872 (N_25872,N_22361,N_23231);
and U25873 (N_25873,N_22951,N_22443);
and U25874 (N_25874,N_22211,N_22100);
and U25875 (N_25875,N_23689,N_23051);
xor U25876 (N_25876,N_22138,N_23330);
or U25877 (N_25877,N_23883,N_22498);
nor U25878 (N_25878,N_23616,N_23540);
xnor U25879 (N_25879,N_23313,N_22304);
nand U25880 (N_25880,N_23665,N_22698);
nand U25881 (N_25881,N_22921,N_23714);
nor U25882 (N_25882,N_23073,N_22755);
nand U25883 (N_25883,N_22149,N_22973);
and U25884 (N_25884,N_23511,N_22413);
and U25885 (N_25885,N_23423,N_22500);
nand U25886 (N_25886,N_22695,N_23209);
nor U25887 (N_25887,N_22435,N_23234);
nand U25888 (N_25888,N_23288,N_23216);
nand U25889 (N_25889,N_23507,N_22571);
nand U25890 (N_25890,N_22106,N_23326);
and U25891 (N_25891,N_22495,N_22929);
nor U25892 (N_25892,N_22703,N_22273);
xnor U25893 (N_25893,N_22760,N_23651);
nor U25894 (N_25894,N_22260,N_22882);
and U25895 (N_25895,N_22804,N_22024);
or U25896 (N_25896,N_22711,N_23674);
or U25897 (N_25897,N_23380,N_23317);
nand U25898 (N_25898,N_22300,N_23075);
and U25899 (N_25899,N_22278,N_22819);
nand U25900 (N_25900,N_22508,N_23634);
nand U25901 (N_25901,N_22177,N_23695);
nand U25902 (N_25902,N_22746,N_23090);
or U25903 (N_25903,N_22343,N_22740);
or U25904 (N_25904,N_22553,N_23542);
or U25905 (N_25905,N_22177,N_23012);
or U25906 (N_25906,N_22991,N_23298);
xnor U25907 (N_25907,N_23878,N_23271);
nor U25908 (N_25908,N_22004,N_22189);
or U25909 (N_25909,N_22727,N_22091);
or U25910 (N_25910,N_22990,N_23836);
and U25911 (N_25911,N_23845,N_22572);
and U25912 (N_25912,N_22010,N_23831);
nand U25913 (N_25913,N_22359,N_22563);
xnor U25914 (N_25914,N_22412,N_23569);
nor U25915 (N_25915,N_22760,N_23388);
or U25916 (N_25916,N_22838,N_22815);
xnor U25917 (N_25917,N_23330,N_23484);
nor U25918 (N_25918,N_23281,N_22627);
or U25919 (N_25919,N_23008,N_22487);
and U25920 (N_25920,N_22121,N_23336);
and U25921 (N_25921,N_23422,N_22923);
nor U25922 (N_25922,N_23783,N_23445);
or U25923 (N_25923,N_22426,N_22869);
and U25924 (N_25924,N_23094,N_23434);
xnor U25925 (N_25925,N_22700,N_23314);
or U25926 (N_25926,N_23652,N_22561);
and U25927 (N_25927,N_23145,N_23176);
xnor U25928 (N_25928,N_22796,N_22125);
nor U25929 (N_25929,N_23415,N_23556);
nor U25930 (N_25930,N_23248,N_23088);
xor U25931 (N_25931,N_22154,N_22572);
nand U25932 (N_25932,N_22520,N_22999);
and U25933 (N_25933,N_22306,N_22379);
xor U25934 (N_25934,N_23724,N_23187);
or U25935 (N_25935,N_23111,N_22146);
and U25936 (N_25936,N_22206,N_23370);
or U25937 (N_25937,N_23087,N_23494);
and U25938 (N_25938,N_23582,N_22869);
and U25939 (N_25939,N_22793,N_22676);
nor U25940 (N_25940,N_22035,N_22838);
and U25941 (N_25941,N_22120,N_23570);
xnor U25942 (N_25942,N_23070,N_22793);
xor U25943 (N_25943,N_23146,N_22085);
nor U25944 (N_25944,N_22286,N_22246);
nor U25945 (N_25945,N_23121,N_23646);
xor U25946 (N_25946,N_22383,N_22844);
nand U25947 (N_25947,N_23362,N_23317);
xnor U25948 (N_25948,N_22269,N_22513);
nor U25949 (N_25949,N_22229,N_23635);
or U25950 (N_25950,N_22593,N_22035);
or U25951 (N_25951,N_22186,N_22392);
xnor U25952 (N_25952,N_23926,N_23006);
or U25953 (N_25953,N_22792,N_22094);
xor U25954 (N_25954,N_23301,N_23276);
and U25955 (N_25955,N_22198,N_22382);
nor U25956 (N_25956,N_22869,N_22387);
and U25957 (N_25957,N_22049,N_22572);
or U25958 (N_25958,N_22752,N_22410);
and U25959 (N_25959,N_23148,N_23107);
nand U25960 (N_25960,N_22878,N_23783);
nand U25961 (N_25961,N_23336,N_22492);
nor U25962 (N_25962,N_22584,N_23110);
nor U25963 (N_25963,N_22140,N_22517);
nor U25964 (N_25964,N_23808,N_22275);
or U25965 (N_25965,N_23978,N_22156);
nand U25966 (N_25966,N_23678,N_23793);
or U25967 (N_25967,N_23752,N_22011);
nor U25968 (N_25968,N_22854,N_22290);
or U25969 (N_25969,N_23494,N_22773);
xnor U25970 (N_25970,N_22273,N_22335);
nand U25971 (N_25971,N_22151,N_23490);
xnor U25972 (N_25972,N_22574,N_22770);
xor U25973 (N_25973,N_22663,N_22630);
nand U25974 (N_25974,N_23368,N_23461);
and U25975 (N_25975,N_22342,N_23329);
and U25976 (N_25976,N_23571,N_23276);
or U25977 (N_25977,N_23850,N_22054);
or U25978 (N_25978,N_23747,N_23253);
xor U25979 (N_25979,N_22261,N_23734);
or U25980 (N_25980,N_22884,N_23814);
and U25981 (N_25981,N_23508,N_22535);
or U25982 (N_25982,N_23661,N_23428);
xor U25983 (N_25983,N_22908,N_23070);
nand U25984 (N_25984,N_23586,N_23036);
or U25985 (N_25985,N_22990,N_23789);
and U25986 (N_25986,N_23563,N_23926);
or U25987 (N_25987,N_22418,N_23533);
xnor U25988 (N_25988,N_22525,N_23811);
xnor U25989 (N_25989,N_22914,N_23229);
and U25990 (N_25990,N_22145,N_23528);
nand U25991 (N_25991,N_23430,N_22953);
xor U25992 (N_25992,N_23409,N_22369);
nand U25993 (N_25993,N_23946,N_22961);
xnor U25994 (N_25994,N_22580,N_23262);
nor U25995 (N_25995,N_23159,N_22938);
and U25996 (N_25996,N_23208,N_23126);
nor U25997 (N_25997,N_22909,N_23464);
nand U25998 (N_25998,N_22389,N_23964);
nand U25999 (N_25999,N_22387,N_22517);
nand U26000 (N_26000,N_25673,N_25129);
nor U26001 (N_26001,N_25636,N_24499);
xnor U26002 (N_26002,N_24535,N_25366);
and U26003 (N_26003,N_25604,N_24220);
nand U26004 (N_26004,N_24918,N_24808);
xnor U26005 (N_26005,N_25995,N_24880);
xnor U26006 (N_26006,N_24762,N_25944);
nand U26007 (N_26007,N_25009,N_25736);
xnor U26008 (N_26008,N_24182,N_25706);
nor U26009 (N_26009,N_25000,N_25428);
nor U26010 (N_26010,N_25715,N_25796);
and U26011 (N_26011,N_25478,N_24299);
and U26012 (N_26012,N_25739,N_24171);
nand U26013 (N_26013,N_24640,N_25466);
or U26014 (N_26014,N_25066,N_25927);
and U26015 (N_26015,N_25998,N_24391);
or U26016 (N_26016,N_24687,N_24533);
xnor U26017 (N_26017,N_24928,N_25514);
nor U26018 (N_26018,N_24083,N_24604);
nand U26019 (N_26019,N_24317,N_24045);
or U26020 (N_26020,N_24834,N_25856);
nand U26021 (N_26021,N_24094,N_25443);
nor U26022 (N_26022,N_24704,N_25726);
or U26023 (N_26023,N_24081,N_25777);
and U26024 (N_26024,N_25089,N_25106);
nor U26025 (N_26025,N_25907,N_24207);
or U26026 (N_26026,N_25900,N_24683);
xor U26027 (N_26027,N_25071,N_24658);
nand U26028 (N_26028,N_24224,N_24034);
and U26029 (N_26029,N_25245,N_25839);
xnor U26030 (N_26030,N_24944,N_24297);
nor U26031 (N_26031,N_25210,N_24088);
and U26032 (N_26032,N_25462,N_25672);
and U26033 (N_26033,N_24457,N_25234);
or U26034 (N_26034,N_24619,N_25842);
and U26035 (N_26035,N_25580,N_24885);
and U26036 (N_26036,N_24819,N_25127);
or U26037 (N_26037,N_24164,N_24799);
and U26038 (N_26038,N_24823,N_24179);
xor U26039 (N_26039,N_24400,N_24483);
and U26040 (N_26040,N_24650,N_24096);
and U26041 (N_26041,N_25869,N_25097);
xor U26042 (N_26042,N_25033,N_24411);
or U26043 (N_26043,N_25812,N_24945);
or U26044 (N_26044,N_24929,N_24690);
xnor U26045 (N_26045,N_24187,N_24957);
nand U26046 (N_26046,N_24739,N_24904);
nand U26047 (N_26047,N_25390,N_25427);
nor U26048 (N_26048,N_24024,N_24442);
nand U26049 (N_26049,N_24730,N_25408);
xnor U26050 (N_26050,N_25924,N_24318);
nor U26051 (N_26051,N_25566,N_24169);
nor U26052 (N_26052,N_24788,N_25710);
or U26053 (N_26053,N_25136,N_24884);
and U26054 (N_26054,N_24544,N_25511);
nand U26055 (N_26055,N_24802,N_25759);
nor U26056 (N_26056,N_24502,N_25996);
nor U26057 (N_26057,N_25772,N_25393);
nor U26058 (N_26058,N_25161,N_24315);
xnor U26059 (N_26059,N_24981,N_24900);
nor U26060 (N_26060,N_24584,N_24899);
or U26061 (N_26061,N_25296,N_25980);
nand U26062 (N_26062,N_25001,N_24719);
and U26063 (N_26063,N_24370,N_25958);
or U26064 (N_26064,N_25148,N_24891);
nand U26065 (N_26065,N_24051,N_24350);
nor U26066 (N_26066,N_24377,N_25452);
or U26067 (N_26067,N_24939,N_24506);
nand U26068 (N_26068,N_25740,N_25769);
nand U26069 (N_26069,N_25553,N_25118);
xor U26070 (N_26070,N_24489,N_25676);
or U26071 (N_26071,N_25645,N_25548);
or U26072 (N_26072,N_25974,N_25467);
nor U26073 (N_26073,N_25936,N_25444);
or U26074 (N_26074,N_24610,N_25120);
nor U26075 (N_26075,N_24763,N_24272);
or U26076 (N_26076,N_25690,N_25101);
and U26077 (N_26077,N_25252,N_24048);
nand U26078 (N_26078,N_24638,N_24564);
nor U26079 (N_26079,N_24826,N_24410);
nor U26080 (N_26080,N_25577,N_24890);
xnor U26081 (N_26081,N_24425,N_25701);
and U26082 (N_26082,N_25145,N_25850);
and U26083 (N_26083,N_24919,N_24732);
or U26084 (N_26084,N_25258,N_24901);
nand U26085 (N_26085,N_25809,N_24571);
nand U26086 (N_26086,N_24398,N_24897);
or U26087 (N_26087,N_25200,N_25217);
or U26088 (N_26088,N_24557,N_25949);
nand U26089 (N_26089,N_25158,N_25853);
nor U26090 (N_26090,N_25620,N_25574);
xnor U26091 (N_26091,N_24809,N_24173);
nor U26092 (N_26092,N_24432,N_25080);
nor U26093 (N_26093,N_25347,N_25599);
and U26094 (N_26094,N_25205,N_24602);
and U26095 (N_26095,N_24351,N_24682);
xnor U26096 (N_26096,N_24313,N_24942);
or U26097 (N_26097,N_25332,N_25659);
or U26098 (N_26098,N_25587,N_24750);
nor U26099 (N_26099,N_25179,N_24634);
or U26100 (N_26100,N_24274,N_25218);
and U26101 (N_26101,N_25261,N_24217);
xnor U26102 (N_26102,N_25045,N_24283);
xnor U26103 (N_26103,N_24741,N_24563);
and U26104 (N_26104,N_24192,N_24586);
nor U26105 (N_26105,N_24941,N_25373);
and U26106 (N_26106,N_24241,N_24184);
or U26107 (N_26107,N_25058,N_24303);
xnor U26108 (N_26108,N_24117,N_24159);
and U26109 (N_26109,N_24293,N_24233);
and U26110 (N_26110,N_25350,N_25729);
nor U26111 (N_26111,N_25978,N_25895);
xor U26112 (N_26112,N_24488,N_24416);
or U26113 (N_26113,N_25251,N_24744);
nor U26114 (N_26114,N_25563,N_25680);
nor U26115 (N_26115,N_24764,N_25922);
nor U26116 (N_26116,N_25932,N_24577);
xnor U26117 (N_26117,N_25592,N_24703);
and U26118 (N_26118,N_25381,N_24145);
and U26119 (N_26119,N_24617,N_25727);
and U26120 (N_26120,N_24212,N_24349);
and U26121 (N_26121,N_25888,N_24701);
or U26122 (N_26122,N_24327,N_24140);
or U26123 (N_26123,N_25133,N_24195);
nor U26124 (N_26124,N_24820,N_25440);
nand U26125 (N_26125,N_24996,N_24210);
xnor U26126 (N_26126,N_24025,N_25551);
nor U26127 (N_26127,N_24080,N_24468);
or U26128 (N_26128,N_25400,N_24242);
nand U26129 (N_26129,N_25988,N_25913);
nand U26130 (N_26130,N_25696,N_24917);
and U26131 (N_26131,N_25215,N_24320);
or U26132 (N_26132,N_25230,N_25171);
xor U26133 (N_26133,N_24490,N_25685);
or U26134 (N_26134,N_24209,N_25151);
and U26135 (N_26135,N_24659,N_25448);
nor U26136 (N_26136,N_25273,N_25439);
nand U26137 (N_26137,N_25947,N_25199);
or U26138 (N_26138,N_25090,N_24837);
xnor U26139 (N_26139,N_24681,N_24494);
and U26140 (N_26140,N_24958,N_25723);
nand U26141 (N_26141,N_25733,N_24403);
xor U26142 (N_26142,N_25425,N_25530);
or U26143 (N_26143,N_25705,N_25681);
and U26144 (N_26144,N_24628,N_24839);
xor U26145 (N_26145,N_25337,N_25675);
nor U26146 (N_26146,N_24545,N_24838);
nand U26147 (N_26147,N_24177,N_25309);
xnor U26148 (N_26148,N_25072,N_24911);
or U26149 (N_26149,N_24438,N_25067);
nand U26150 (N_26150,N_24865,N_25233);
nand U26151 (N_26151,N_25892,N_25250);
xor U26152 (N_26152,N_25979,N_25880);
nand U26153 (N_26153,N_24050,N_25486);
or U26154 (N_26154,N_24765,N_24962);
nand U26155 (N_26155,N_25510,N_25256);
and U26156 (N_26156,N_25203,N_25552);
nor U26157 (N_26157,N_24673,N_25983);
xor U26158 (N_26158,N_25292,N_25507);
xnor U26159 (N_26159,N_25087,N_25785);
nor U26160 (N_26160,N_24576,N_25483);
xor U26161 (N_26161,N_24841,N_25718);
and U26162 (N_26162,N_24481,N_24835);
and U26163 (N_26163,N_25355,N_24593);
nand U26164 (N_26164,N_24742,N_24269);
xnor U26165 (N_26165,N_24692,N_24952);
or U26166 (N_26166,N_24896,N_24150);
xor U26167 (N_26167,N_25214,N_24062);
xor U26168 (N_26168,N_24013,N_24832);
nor U26169 (N_26169,N_24568,N_24976);
xor U26170 (N_26170,N_24655,N_24086);
nand U26171 (N_26171,N_24705,N_24870);
xnor U26172 (N_26172,N_25891,N_24389);
or U26173 (N_26173,N_25805,N_24231);
and U26174 (N_26174,N_25588,N_25018);
nand U26175 (N_26175,N_24553,N_25352);
xor U26176 (N_26176,N_25190,N_25135);
and U26177 (N_26177,N_24590,N_24455);
nand U26178 (N_26178,N_24424,N_25854);
and U26179 (N_26179,N_24772,N_25914);
and U26180 (N_26180,N_24740,N_25073);
nor U26181 (N_26181,N_25055,N_24654);
xnor U26182 (N_26182,N_24125,N_24232);
nand U26183 (N_26183,N_25160,N_24412);
and U26184 (N_26184,N_24613,N_25325);
nand U26185 (N_26185,N_25545,N_24148);
xnor U26186 (N_26186,N_25982,N_25557);
or U26187 (N_26187,N_25833,N_24469);
xnor U26188 (N_26188,N_24873,N_25847);
nand U26189 (N_26189,N_24038,N_24206);
nor U26190 (N_26190,N_24259,N_25871);
xnor U26191 (N_26191,N_25874,N_25040);
nor U26192 (N_26192,N_24382,N_25322);
nor U26193 (N_26193,N_25225,N_25797);
nor U26194 (N_26194,N_24436,N_25801);
nand U26195 (N_26195,N_25930,N_24229);
or U26196 (N_26196,N_25802,N_24374);
xnor U26197 (N_26197,N_24189,N_24591);
xnor U26198 (N_26198,N_25986,N_25059);
or U26199 (N_26199,N_24782,N_25265);
or U26200 (N_26200,N_24912,N_24116);
xor U26201 (N_26201,N_25820,N_24922);
or U26202 (N_26202,N_25761,N_24265);
xnor U26203 (N_26203,N_25344,N_24768);
nand U26204 (N_26204,N_24243,N_24844);
and U26205 (N_26205,N_24336,N_25298);
nor U26206 (N_26206,N_24697,N_25572);
nor U26207 (N_26207,N_25311,N_24193);
xor U26208 (N_26208,N_24185,N_24367);
nor U26209 (N_26209,N_25743,N_25893);
nor U26210 (N_26210,N_24898,N_25321);
and U26211 (N_26211,N_25267,N_25867);
nand U26212 (N_26212,N_24017,N_25091);
or U26213 (N_26213,N_25519,N_25206);
or U26214 (N_26214,N_24459,N_25315);
and U26215 (N_26215,N_24827,N_24810);
nor U26216 (N_26216,N_24234,N_24724);
and U26217 (N_26217,N_25969,N_25236);
or U26218 (N_26218,N_24097,N_25491);
and U26219 (N_26219,N_24186,N_24005);
or U26220 (N_26220,N_25078,N_24126);
xor U26221 (N_26221,N_25951,N_25872);
xor U26222 (N_26222,N_24933,N_24905);
nor U26223 (N_26223,N_24258,N_24363);
or U26224 (N_26224,N_24871,N_25260);
and U26225 (N_26225,N_25392,N_24644);
nor U26226 (N_26226,N_24920,N_24277);
nor U26227 (N_26227,N_25735,N_24848);
and U26228 (N_26228,N_25846,N_25167);
nand U26229 (N_26229,N_24579,N_25968);
and U26230 (N_26230,N_25342,N_24369);
or U26231 (N_26231,N_25372,N_25612);
and U26232 (N_26232,N_24138,N_24757);
nor U26233 (N_26233,N_25196,N_25808);
and U26234 (N_26234,N_24202,N_25442);
nand U26235 (N_26235,N_25037,N_25704);
nor U26236 (N_26236,N_25354,N_25682);
nand U26237 (N_26237,N_25541,N_25535);
and U26238 (N_26238,N_24894,N_24018);
or U26239 (N_26239,N_25115,N_25760);
nor U26240 (N_26240,N_24307,N_24226);
or U26241 (N_26241,N_25235,N_24358);
or U26242 (N_26242,N_24789,N_24444);
xnor U26243 (N_26243,N_24803,N_24228);
nand U26244 (N_26244,N_25665,N_24044);
nor U26245 (N_26245,N_25902,N_25790);
and U26246 (N_26246,N_24329,N_24609);
nand U26247 (N_26247,N_25629,N_25211);
nand U26248 (N_26248,N_25901,N_25697);
or U26249 (N_26249,N_24262,N_25131);
nand U26250 (N_26250,N_24354,N_25413);
nand U26251 (N_26251,N_25543,N_24910);
or U26252 (N_26252,N_25301,N_25633);
or U26253 (N_26253,N_24294,N_25320);
xor U26254 (N_26254,N_24636,N_25691);
or U26255 (N_26255,N_25560,N_25879);
nor U26256 (N_26256,N_25578,N_24937);
nand U26257 (N_26257,N_24089,N_24032);
xor U26258 (N_26258,N_24046,N_25505);
xor U26259 (N_26259,N_25667,N_25013);
xor U26260 (N_26260,N_24688,N_25684);
nor U26261 (N_26261,N_24647,N_25475);
nor U26262 (N_26262,N_24585,N_25928);
and U26263 (N_26263,N_24282,N_25108);
nand U26264 (N_26264,N_24850,N_24989);
nand U26265 (N_26265,N_24693,N_25119);
xor U26266 (N_26266,N_24561,N_25765);
and U26267 (N_26267,N_25806,N_25942);
nand U26268 (N_26268,N_24422,N_24271);
or U26269 (N_26269,N_24497,N_24596);
or U26270 (N_26270,N_24264,N_25096);
xnor U26271 (N_26271,N_25766,N_25186);
and U26272 (N_26272,N_25613,N_25644);
xnor U26273 (N_26273,N_24940,N_25004);
or U26274 (N_26274,N_25600,N_24605);
nor U26275 (N_26275,N_25461,N_25589);
nor U26276 (N_26276,N_24227,N_24621);
and U26277 (N_26277,N_24304,N_25399);
and U26278 (N_26278,N_24774,N_24566);
nand U26279 (N_26279,N_25410,N_24181);
or U26280 (N_26280,N_24333,N_25420);
nor U26281 (N_26281,N_25012,N_25547);
and U26282 (N_26282,N_25212,N_25652);
nand U26283 (N_26283,N_25534,N_24601);
xor U26284 (N_26284,N_25126,N_24405);
nor U26285 (N_26285,N_24646,N_24131);
nor U26286 (N_26286,N_24430,N_24113);
or U26287 (N_26287,N_25188,N_24895);
and U26288 (N_26288,N_24501,N_24831);
xnor U26289 (N_26289,N_25493,N_25387);
nand U26290 (N_26290,N_24378,N_25559);
nor U26291 (N_26291,N_25085,N_24443);
or U26292 (N_26292,N_24979,N_24295);
and U26293 (N_26293,N_25747,N_25904);
nand U26294 (N_26294,N_25228,N_24332);
nor U26295 (N_26295,N_24015,N_24678);
nand U26296 (N_26296,N_25502,N_25484);
xor U26297 (N_26297,N_25182,N_25906);
nor U26298 (N_26298,N_24063,N_25005);
or U26299 (N_26299,N_25776,N_24624);
nand U26300 (N_26300,N_24699,N_24984);
nand U26301 (N_26301,N_24101,N_25639);
and U26302 (N_26302,N_25109,N_24538);
nand U26303 (N_26303,N_25885,N_24176);
nand U26304 (N_26304,N_24846,N_24129);
nand U26305 (N_26305,N_25051,N_24861);
or U26306 (N_26306,N_25795,N_24066);
xnor U26307 (N_26307,N_24067,N_25147);
and U26308 (N_26308,N_24092,N_24666);
xor U26309 (N_26309,N_24010,N_25751);
xnor U26310 (N_26310,N_25702,N_25700);
or U26311 (N_26311,N_24540,N_25630);
or U26312 (N_26312,N_25987,N_25015);
nor U26313 (N_26313,N_24251,N_25935);
or U26314 (N_26314,N_24775,N_25434);
xnor U26315 (N_26315,N_25364,N_24770);
xor U26316 (N_26316,N_25829,N_24934);
nand U26317 (N_26317,N_24334,N_24555);
nand U26318 (N_26318,N_25162,N_25827);
and U26319 (N_26319,N_25458,N_25993);
nand U26320 (N_26320,N_24057,N_24649);
or U26321 (N_26321,N_25172,N_24375);
or U26322 (N_26322,N_25635,N_24419);
nand U26323 (N_26323,N_25384,N_24951);
or U26324 (N_26324,N_24214,N_24569);
or U26325 (N_26325,N_24023,N_25029);
nor U26326 (N_26326,N_24451,N_25583);
and U26327 (N_26327,N_25417,N_24060);
and U26328 (N_26328,N_25426,N_24281);
and U26329 (N_26329,N_24751,N_24932);
xnor U26330 (N_26330,N_25446,N_25666);
or U26331 (N_26331,N_24152,N_24132);
or U26332 (N_26332,N_24467,N_25554);
nor U26333 (N_26333,N_24883,N_25770);
and U26334 (N_26334,N_24999,N_24280);
nor U26335 (N_26335,N_24990,N_25940);
or U26336 (N_26336,N_24298,N_25287);
nand U26337 (N_26337,N_24053,N_25423);
nand U26338 (N_26338,N_24392,N_24921);
nor U26339 (N_26339,N_24760,N_25441);
or U26340 (N_26340,N_24084,N_24480);
or U26341 (N_26341,N_24859,N_25204);
xor U26342 (N_26342,N_24589,N_24039);
or U26343 (N_26343,N_24780,N_25201);
xnor U26344 (N_26344,N_25377,N_25116);
nor U26345 (N_26345,N_25388,N_24863);
or U26346 (N_26346,N_25289,N_25991);
or U26347 (N_26347,N_24465,N_25688);
nor U26348 (N_26348,N_25338,N_25544);
or U26349 (N_26349,N_24626,N_25607);
or U26350 (N_26350,N_25890,N_25349);
nand U26351 (N_26351,N_24508,N_24828);
nor U26352 (N_26352,N_24671,N_25368);
nand U26353 (N_26353,N_25093,N_25631);
xnor U26354 (N_26354,N_24698,N_24851);
nand U26355 (N_26355,N_24474,N_25095);
xnor U26356 (N_26356,N_24409,N_24098);
xor U26357 (N_26357,N_25937,N_24364);
or U26358 (N_26358,N_24515,N_24845);
or U26359 (N_26359,N_24548,N_25584);
nand U26360 (N_26360,N_24752,N_24893);
and U26361 (N_26361,N_24273,N_24118);
and U26362 (N_26362,N_24103,N_24792);
xnor U26363 (N_26363,N_25834,N_24759);
xnor U26364 (N_26364,N_25878,N_25436);
nand U26365 (N_26365,N_24971,N_24689);
nor U26366 (N_26366,N_25130,N_25734);
and U26367 (N_26367,N_25006,N_25915);
nor U26368 (N_26368,N_25389,N_24208);
nor U26369 (N_26369,N_24380,N_25961);
or U26370 (N_26370,N_24580,N_24439);
nand U26371 (N_26371,N_24559,N_24001);
and U26372 (N_26372,N_24523,N_25835);
nand U26373 (N_26373,N_24082,N_24479);
nor U26374 (N_26374,N_24927,N_24592);
nand U26375 (N_26375,N_24435,N_24583);
or U26376 (N_26376,N_24221,N_25243);
nor U26377 (N_26377,N_24987,N_24423);
and U26378 (N_26378,N_25189,N_25207);
xor U26379 (N_26379,N_24814,N_25720);
and U26380 (N_26380,N_25169,N_24413);
nand U26381 (N_26381,N_25282,N_25602);
nor U26382 (N_26382,N_25568,N_24384);
xor U26383 (N_26383,N_25717,N_24805);
nor U26384 (N_26384,N_25110,N_25278);
nor U26385 (N_26385,N_25506,N_24200);
and U26386 (N_26386,N_24135,N_24886);
and U26387 (N_26387,N_24721,N_24471);
nand U26388 (N_26388,N_24041,N_25242);
nor U26389 (N_26389,N_25336,N_25333);
or U26390 (N_26390,N_24031,N_25821);
and U26391 (N_26391,N_25002,N_24278);
or U26392 (N_26392,N_24461,N_24387);
or U26393 (N_26393,N_24249,N_25339);
or U26394 (N_26394,N_25429,N_24661);
and U26395 (N_26395,N_24055,N_24174);
xor U26396 (N_26396,N_25971,N_25905);
xor U26397 (N_26397,N_24505,N_24973);
nand U26398 (N_26398,N_24395,N_25451);
and U26399 (N_26399,N_24924,N_24767);
nor U26400 (N_26400,N_24528,N_24729);
nor U26401 (N_26401,N_24344,N_25625);
or U26402 (N_26402,N_24997,N_25582);
xnor U26403 (N_26403,N_24255,N_24720);
xor U26404 (N_26404,N_25076,N_25889);
nor U26405 (N_26405,N_25084,N_24575);
and U26406 (N_26406,N_24341,N_25517);
or U26407 (N_26407,N_24529,N_24037);
nor U26408 (N_26408,N_24753,N_25330);
and U26409 (N_26409,N_24194,N_25619);
nor U26410 (N_26410,N_25855,N_24473);
nor U26411 (N_26411,N_25774,N_25124);
nor U26412 (N_26412,N_24611,N_25657);
nor U26413 (N_26413,N_24340,N_24250);
nand U26414 (N_26414,N_25816,N_24361);
and U26415 (N_26415,N_25341,N_24141);
nand U26416 (N_26416,N_25678,N_24755);
xor U26417 (N_26417,N_25860,N_25537);
and U26418 (N_26418,N_24256,N_24087);
or U26419 (N_26419,N_24028,N_24285);
and U26420 (N_26420,N_24582,N_25596);
or U26421 (N_26421,N_24966,N_25496);
and U26422 (N_26422,N_25570,N_25353);
xor U26423 (N_26423,N_25787,N_24965);
nand U26424 (N_26424,N_24402,N_25374);
nor U26425 (N_26425,N_24160,N_24606);
and U26426 (N_26426,N_24049,N_24977);
nor U26427 (N_26427,N_25480,N_25938);
and U26428 (N_26428,N_24030,N_25039);
or U26429 (N_26429,N_25818,N_24709);
nand U26430 (N_26430,N_25522,N_25088);
xor U26431 (N_26431,N_25683,N_24953);
nand U26432 (N_26432,N_24620,N_25314);
nor U26433 (N_26433,N_24290,N_24817);
xnor U26434 (N_26434,N_24029,N_25571);
nand U26435 (N_26435,N_25221,N_24829);
nand U26436 (N_26436,N_24735,N_25793);
nand U26437 (N_26437,N_24597,N_25224);
and U26438 (N_26438,N_25663,N_25745);
and U26439 (N_26439,N_25102,N_25043);
nor U26440 (N_26440,N_24458,N_24065);
and U26441 (N_26441,N_25773,N_25634);
nand U26442 (N_26442,N_25371,N_25753);
and U26443 (N_26443,N_24429,N_25918);
and U26444 (N_26444,N_24335,N_24175);
or U26445 (N_26445,N_25007,N_25495);
or U26446 (N_26446,N_25020,N_25208);
and U26447 (N_26447,N_25213,N_24314);
nor U26448 (N_26448,N_25868,N_24236);
or U26449 (N_26449,N_24622,N_25963);
nor U26450 (N_26450,N_24993,N_25497);
nand U26451 (N_26451,N_24068,N_24246);
or U26452 (N_26452,N_25788,N_25057);
xor U26453 (N_26453,N_25750,N_24860);
nor U26454 (N_26454,N_24261,N_24248);
nor U26455 (N_26455,N_25246,N_25293);
and U26456 (N_26456,N_24383,N_24935);
nor U26457 (N_26457,N_25970,N_25356);
and U26458 (N_26458,N_25654,N_25358);
or U26459 (N_26459,N_25359,N_24162);
and U26460 (N_26460,N_25792,N_25724);
xnor U26461 (N_26461,N_24309,N_24858);
and U26462 (N_26462,N_25783,N_24223);
or U26463 (N_26463,N_25456,N_24059);
nand U26464 (N_26464,N_25409,N_24887);
or U26465 (N_26465,N_25194,N_24245);
xor U26466 (N_26466,N_24632,N_24254);
nor U26467 (N_26467,N_24806,N_25113);
nand U26468 (N_26468,N_24180,N_24914);
or U26469 (N_26469,N_24727,N_25437);
and U26470 (N_26470,N_24915,N_25756);
nor U26471 (N_26471,N_24748,N_24676);
or U26472 (N_26472,N_25259,N_25404);
and U26473 (N_26473,N_25990,N_24836);
nor U26474 (N_26474,N_25603,N_25117);
nand U26475 (N_26475,N_25653,N_25295);
or U26476 (N_26476,N_25624,N_25762);
xnor U26477 (N_26477,N_25608,N_25290);
nor U26478 (N_26478,N_25421,N_25693);
and U26479 (N_26479,N_25082,N_25403);
or U26480 (N_26480,N_25558,N_24988);
nand U26481 (N_26481,N_25238,N_25165);
xor U26482 (N_26482,N_25053,N_25192);
or U26483 (N_26483,N_24456,N_24058);
nor U26484 (N_26484,N_24756,N_25722);
xnor U26485 (N_26485,N_25379,N_25955);
and U26486 (N_26486,N_24270,N_24095);
nor U26487 (N_26487,N_24326,N_24627);
or U26488 (N_26488,N_24426,N_25643);
or U26489 (N_26489,N_24840,N_24478);
xor U26490 (N_26490,N_24075,N_25143);
and U26491 (N_26491,N_25616,N_25447);
or U26492 (N_26492,N_24417,N_24711);
nor U26493 (N_26493,N_25929,N_25432);
and U26494 (N_26494,N_24311,N_25593);
and U26495 (N_26495,N_24907,N_25692);
or U26496 (N_26496,N_25516,N_24726);
xnor U26497 (N_26497,N_24795,N_24629);
xnor U26498 (N_26498,N_25957,N_24600);
nand U26499 (N_26499,N_24930,N_25324);
or U26500 (N_26500,N_24486,N_25527);
and U26501 (N_26501,N_24824,N_25763);
nand U26502 (N_26502,N_25876,N_24908);
or U26503 (N_26503,N_24874,N_25026);
and U26504 (N_26504,N_24122,N_25032);
and U26505 (N_26505,N_25948,N_25367);
and U26506 (N_26506,N_25490,N_24670);
and U26507 (N_26507,N_24696,N_25424);
xor U26508 (N_26508,N_24519,N_25836);
xnor U26509 (N_26509,N_24510,N_24042);
nor U26510 (N_26510,N_25146,N_25193);
and U26511 (N_26511,N_24948,N_24434);
nor U26512 (N_26512,N_25515,N_25457);
or U26513 (N_26513,N_24791,N_24734);
or U26514 (N_26514,N_25916,N_25781);
and U26515 (N_26515,N_25863,N_24260);
or U26516 (N_26516,N_25656,N_24496);
and U26517 (N_26517,N_25877,N_25976);
and U26518 (N_26518,N_24825,N_25615);
and U26519 (N_26519,N_24842,N_25524);
and U26520 (N_26520,N_25370,N_25755);
and U26521 (N_26521,N_24855,N_25828);
nor U26522 (N_26522,N_25782,N_24121);
xor U26523 (N_26523,N_25946,N_25931);
xor U26524 (N_26524,N_25272,N_24972);
and U26525 (N_26525,N_24807,N_24147);
or U26526 (N_26526,N_25317,N_24440);
xnor U26527 (N_26527,N_24257,N_24725);
nand U26528 (N_26528,N_25865,N_24244);
or U26529 (N_26529,N_25798,N_25291);
nor U26530 (N_26530,N_25385,N_24156);
and U26531 (N_26531,N_25549,N_25041);
nor U26532 (N_26532,N_24485,N_25065);
nand U26533 (N_26533,N_24110,N_24960);
and U26534 (N_26534,N_24339,N_25859);
nand U26535 (N_26535,N_24252,N_24736);
or U26536 (N_26536,N_24776,N_25492);
nand U26537 (N_26537,N_25741,N_24394);
or U26538 (N_26538,N_25128,N_25539);
nor U26539 (N_26539,N_24085,N_24833);
and U26540 (N_26540,N_24572,N_25870);
or U26541 (N_26541,N_25757,N_24631);
nor U26542 (N_26542,N_24128,N_24872);
and U26543 (N_26543,N_25595,N_24338);
or U26544 (N_26544,N_25326,N_25270);
xnor U26545 (N_26545,N_24012,N_24503);
and U26546 (N_26546,N_24718,N_25953);
or U26547 (N_26547,N_24950,N_25383);
xnor U26548 (N_26548,N_25241,N_25925);
nor U26549 (N_26549,N_24302,N_24595);
nor U26550 (N_26550,N_24864,N_25894);
nand U26551 (N_26551,N_25542,N_24399);
and U26552 (N_26552,N_24286,N_25921);
nand U26553 (N_26553,N_25651,N_25881);
or U26554 (N_26554,N_25132,N_25838);
and U26555 (N_26555,N_25375,N_25679);
nor U26556 (N_26556,N_25716,N_25822);
or U26557 (N_26557,N_24964,N_25811);
and U26558 (N_26558,N_24672,N_25327);
and U26559 (N_26559,N_24731,N_25079);
nor U26560 (N_26560,N_24888,N_24869);
xor U26561 (N_26561,N_24961,N_25837);
nor U26562 (N_26562,N_25485,N_24454);
and U26563 (N_26563,N_24504,N_24665);
nor U26564 (N_26564,N_24276,N_25284);
nand U26565 (N_26565,N_24360,N_25197);
or U26566 (N_26566,N_25474,N_25416);
nand U26567 (N_26567,N_24500,N_24794);
and U26568 (N_26568,N_25335,N_25391);
and U26569 (N_26569,N_25768,N_24211);
xnor U26570 (N_26570,N_24567,N_24040);
xor U26571 (N_26571,N_25830,N_24552);
or U26572 (N_26572,N_25939,N_25732);
or U26573 (N_26573,N_24205,N_25134);
nand U26574 (N_26574,N_24204,N_24573);
or U26575 (N_26575,N_24714,N_24139);
xnor U26576 (N_26576,N_25841,N_25275);
nand U26577 (N_26577,N_24786,N_25477);
or U26578 (N_26578,N_25899,N_25689);
nand U26579 (N_26579,N_24168,N_24056);
nor U26580 (N_26580,N_24766,N_25329);
or U26581 (N_26581,N_24982,N_24279);
nand U26582 (N_26582,N_24133,N_24587);
nand U26583 (N_26583,N_24702,N_25494);
and U26584 (N_26584,N_24574,N_24284);
xor U26585 (N_26585,N_24633,N_25686);
or U26586 (N_26586,N_24643,N_25310);
or U26587 (N_26587,N_24522,N_25468);
or U26588 (N_26588,N_25011,N_24674);
and U26589 (N_26589,N_25470,N_24542);
and U26590 (N_26590,N_24639,N_25857);
xor U26591 (N_26591,N_24877,N_24959);
and U26592 (N_26592,N_25300,N_25274);
nor U26593 (N_26593,N_24530,N_25460);
nor U26594 (N_26594,N_25911,N_25528);
nor U26595 (N_26595,N_24172,N_25307);
xor U26596 (N_26596,N_25671,N_25884);
nor U26597 (N_26597,N_25112,N_25565);
nand U26598 (N_26598,N_25984,N_24099);
and U26599 (N_26599,N_25521,N_25471);
nand U26600 (N_26600,N_25401,N_25981);
and U26601 (N_26601,N_25786,N_25887);
or U26602 (N_26602,N_24306,N_24009);
nor U26603 (N_26603,N_24091,N_25178);
nor U26604 (N_26604,N_25489,N_24968);
xor U26605 (N_26605,N_24143,N_24054);
nor U26606 (N_26606,N_25323,N_24007);
and U26607 (N_26607,N_24615,N_25008);
or U26608 (N_26608,N_25861,N_24524);
nor U26609 (N_26609,N_24728,N_25122);
and U26610 (N_26610,N_25973,N_25183);
nand U26611 (N_26611,N_24777,N_24319);
and U26612 (N_26612,N_25056,N_25025);
or U26613 (N_26613,N_25155,N_25281);
xor U26614 (N_26614,N_25019,N_25357);
nor U26615 (N_26615,N_24453,N_24026);
or U26616 (N_26616,N_24651,N_25606);
nand U26617 (N_26617,N_25909,N_25209);
xor U26618 (N_26618,N_24635,N_24511);
nand U26619 (N_26619,N_24783,N_24291);
nand U26620 (N_26620,N_25504,N_25331);
xor U26621 (N_26621,N_25849,N_24630);
xnor U26622 (N_26622,N_25637,N_25223);
xnor U26623 (N_26623,N_24366,N_24800);
and U26624 (N_26624,N_24079,N_25775);
nand U26625 (N_26625,N_24513,N_25523);
and U26626 (N_26626,N_25237,N_24178);
and U26627 (N_26627,N_24267,N_25297);
and U26628 (N_26628,N_25573,N_25140);
and U26629 (N_26629,N_24867,N_24594);
nor U26630 (N_26630,N_24372,N_24356);
nor U26631 (N_26631,N_24487,N_25114);
xnor U26632 (N_26632,N_24695,N_25737);
nor U26633 (N_26633,N_24324,N_25744);
nand U26634 (N_26634,N_24365,N_25453);
and U26635 (N_26635,N_25754,N_25070);
nor U26636 (N_26636,N_25569,N_24123);
and U26637 (N_26637,N_24645,N_25555);
nand U26638 (N_26638,N_24104,N_25075);
nand U26639 (N_26639,N_25999,N_25382);
nor U26640 (N_26640,N_25176,N_24447);
nand U26641 (N_26641,N_24796,N_24052);
nand U26642 (N_26642,N_25016,N_24337);
xor U26643 (N_26643,N_24761,N_25276);
nand U26644 (N_26644,N_25014,N_24663);
or U26645 (N_26645,N_24985,N_25994);
xnor U26646 (N_26646,N_25170,N_24931);
and U26647 (N_26647,N_25866,N_24157);
nor U26648 (N_26648,N_25778,N_24925);
nor U26649 (N_26649,N_25185,N_24263);
nand U26650 (N_26650,N_24797,N_24607);
and U26651 (N_26651,N_25017,N_25585);
nor U26652 (N_26652,N_25934,N_25858);
and U26653 (N_26653,N_25173,N_24581);
nand U26654 (N_26654,N_25526,N_24947);
xnor U26655 (N_26655,N_24653,N_25253);
nor U26656 (N_26656,N_24866,N_24452);
xnor U26657 (N_26657,N_25419,N_25061);
xnor U26658 (N_26658,N_24849,N_25174);
nor U26659 (N_26659,N_25714,N_24983);
or U26660 (N_26660,N_25529,N_25229);
nor U26661 (N_26661,N_25826,N_24011);
nand U26662 (N_26662,N_24700,N_24675);
xor U26663 (N_26663,N_24969,N_24685);
or U26664 (N_26664,N_24343,N_25711);
and U26665 (N_26665,N_24556,N_24493);
nor U26666 (N_26666,N_24801,N_25658);
nor U26667 (N_26667,N_24196,N_24450);
and U26668 (N_26668,N_25840,N_24061);
xor U26669 (N_26669,N_24136,N_25023);
nor U26670 (N_26670,N_25920,N_24428);
or U26671 (N_26671,N_25640,N_25513);
xnor U26672 (N_26672,N_24562,N_25823);
or U26673 (N_26673,N_25749,N_24153);
or U26674 (N_26674,N_25181,N_25546);
nand U26675 (N_26675,N_24385,N_24612);
nor U26676 (N_26676,N_24637,N_25137);
nand U26677 (N_26677,N_25343,N_25954);
nand U26678 (N_26678,N_25348,N_24745);
nor U26679 (N_26679,N_24124,N_25459);
nand U26680 (N_26680,N_24514,N_25641);
and U26681 (N_26681,N_25268,N_25719);
nor U26682 (N_26682,N_24712,N_25219);
or U26683 (N_26683,N_25731,N_24812);
nor U26684 (N_26684,N_25157,N_24570);
nor U26685 (N_26685,N_24393,N_25154);
nand U26686 (N_26686,N_25077,N_25030);
and U26687 (N_26687,N_25063,N_24625);
or U26688 (N_26688,N_25227,N_25518);
nor U26689 (N_26689,N_24287,N_24362);
or U26690 (N_26690,N_25163,N_25713);
xor U26691 (N_26691,N_25959,N_25479);
and U26692 (N_26692,N_24433,N_24388);
or U26693 (N_26693,N_25650,N_25156);
or U26694 (N_26694,N_25648,N_25628);
or U26695 (N_26695,N_25472,N_24946);
or U26696 (N_26696,N_24390,N_24238);
nor U26697 (N_26697,N_24954,N_25216);
xor U26698 (N_26698,N_24821,N_24408);
and U26699 (N_26699,N_24158,N_24427);
nand U26700 (N_26700,N_25415,N_24371);
nand U26701 (N_26701,N_25844,N_24652);
xnor U26702 (N_26702,N_24549,N_25361);
nand U26703 (N_26703,N_24289,N_25908);
nor U26704 (N_26704,N_25255,N_24137);
or U26705 (N_26705,N_24151,N_24347);
or U26706 (N_26706,N_25638,N_25698);
or U26707 (N_26707,N_24142,N_25263);
nor U26708 (N_26708,N_25964,N_25674);
and U26709 (N_26709,N_25034,N_24847);
xor U26710 (N_26710,N_25285,N_25299);
nor U26711 (N_26711,N_25804,N_25220);
nand U26712 (N_26712,N_25550,N_25661);
xor U26713 (N_26713,N_24240,N_25397);
xnor U26714 (N_26714,N_24437,N_24926);
xnor U26715 (N_26715,N_25824,N_25042);
and U26716 (N_26716,N_24420,N_24149);
xor U26717 (N_26717,N_25254,N_24546);
xnor U26718 (N_26718,N_25875,N_24680);
or U26719 (N_26719,N_24991,N_24520);
nor U26720 (N_26720,N_24648,N_24328);
nor U26721 (N_26721,N_24308,N_24554);
or U26722 (N_26722,N_24418,N_25621);
nand U26723 (N_26723,N_24955,N_24198);
and U26724 (N_26724,N_25138,N_25469);
and U26725 (N_26725,N_24183,N_24716);
nor U26726 (N_26726,N_24477,N_24713);
or U26727 (N_26727,N_24491,N_24167);
nand U26728 (N_26728,N_24275,N_24401);
and U26729 (N_26729,N_25360,N_25780);
or U26730 (N_26730,N_25815,N_25027);
and U26731 (N_26731,N_25561,N_25590);
or U26732 (N_26732,N_24108,N_25531);
nand U26733 (N_26733,N_25501,N_24441);
nand U26734 (N_26734,N_25831,N_24036);
xnor U26735 (N_26735,N_25139,N_24219);
and U26736 (N_26736,N_25028,N_24660);
nor U26737 (N_26737,N_24074,N_25746);
or U26738 (N_26738,N_24623,N_25992);
xnor U26739 (N_26739,N_25152,N_25742);
nor U26740 (N_26740,N_25111,N_25465);
or U26741 (N_26741,N_25153,N_24197);
or U26742 (N_26742,N_25271,N_24998);
or U26743 (N_26743,N_24686,N_25060);
xor U26744 (N_26744,N_24902,N_25283);
nor U26745 (N_26745,N_25977,N_24330);
xor U26746 (N_26746,N_24445,N_25807);
or U26747 (N_26747,N_25226,N_25222);
xnor U26748 (N_26748,N_24710,N_25610);
or U26749 (N_26749,N_24813,N_25677);
or U26750 (N_26750,N_24881,N_24203);
nand U26751 (N_26751,N_25476,N_25707);
nor U26752 (N_26752,N_24352,N_24239);
nand U26753 (N_26753,N_24266,N_24043);
and U26754 (N_26754,N_25049,N_25664);
nand U26755 (N_26755,N_24154,N_25398);
xor U26756 (N_26756,N_24856,N_25532);
and U26757 (N_26757,N_25655,N_25883);
nor U26758 (N_26758,N_25454,N_24790);
or U26759 (N_26759,N_24875,N_25302);
nand U26760 (N_26760,N_25365,N_24463);
xor U26761 (N_26761,N_24879,N_24414);
and U26762 (N_26762,N_24614,N_25074);
xor U26763 (N_26763,N_24550,N_24102);
and U26764 (N_26764,N_24359,N_25943);
and U26765 (N_26765,N_25721,N_24588);
or U26766 (N_26766,N_24464,N_24170);
and U26767 (N_26767,N_24551,N_25810);
nor U26768 (N_26768,N_25695,N_24397);
nand U26769 (N_26769,N_25803,N_25306);
and U26770 (N_26770,N_24292,N_25304);
nand U26771 (N_26771,N_24516,N_24033);
xnor U26772 (N_26772,N_24975,N_25509);
nand U26773 (N_26773,N_24532,N_25280);
nor U26774 (N_26774,N_24852,N_24738);
xnor U26775 (N_26775,N_24003,N_24404);
and U26776 (N_26776,N_25626,N_25198);
or U26777 (N_26777,N_24995,N_25738);
or U26778 (N_26778,N_24733,N_25989);
nand U26779 (N_26779,N_25601,N_24379);
or U26780 (N_26780,N_24743,N_25886);
nand U26781 (N_26781,N_24321,N_24035);
or U26782 (N_26782,N_25898,N_25498);
nand U26783 (N_26783,N_25896,N_25422);
xnor U26784 (N_26784,N_25031,N_24793);
or U26785 (N_26785,N_25177,N_25611);
or U26786 (N_26786,N_25662,N_24342);
or U26787 (N_26787,N_24472,N_24247);
and U26788 (N_26788,N_25614,N_25345);
xor U26789 (N_26789,N_24090,N_25279);
or U26790 (N_26790,N_25328,N_24857);
or U26791 (N_26791,N_24541,N_24027);
or U26792 (N_26792,N_25266,N_25168);
xnor U26793 (N_26793,N_24111,N_24213);
or U26794 (N_26794,N_24373,N_24008);
or U26795 (N_26795,N_25594,N_25418);
xnor U26796 (N_26796,N_25972,N_24708);
xnor U26797 (N_26797,N_25240,N_25623);
nand U26798 (N_26798,N_24002,N_25402);
and U26799 (N_26799,N_25617,N_24679);
or U26800 (N_26800,N_25239,N_24754);
nor U26801 (N_26801,N_24903,N_25487);
xnor U26802 (N_26802,N_24268,N_24449);
xnor U26803 (N_26803,N_24218,N_24021);
xor U26804 (N_26804,N_24355,N_25694);
nand U26805 (N_26805,N_25597,N_24737);
and U26806 (N_26806,N_24521,N_24599);
and U26807 (N_26807,N_24779,N_24527);
and U26808 (N_26808,N_24707,N_25412);
xnor U26809 (N_26809,N_25618,N_25411);
nor U26810 (N_26810,N_24876,N_24717);
nand U26811 (N_26811,N_24004,N_25103);
or U26812 (N_26812,N_24161,N_24146);
and U26813 (N_26813,N_24476,N_25503);
or U26814 (N_26814,N_25340,N_24300);
nor U26815 (N_26815,N_25380,N_25430);
nand U26816 (N_26816,N_25202,N_25264);
xnor U26817 (N_26817,N_24916,N_25149);
xor U26818 (N_26818,N_24667,N_24492);
xnor U26819 (N_26819,N_24069,N_25997);
nand U26820 (N_26820,N_25832,N_25294);
nand U26821 (N_26821,N_25010,N_24657);
and U26822 (N_26822,N_25910,N_25598);
nand U26823 (N_26823,N_25752,N_24305);
nand U26824 (N_26824,N_24526,N_24518);
nand U26825 (N_26825,N_25789,N_24862);
nand U26826 (N_26826,N_25873,N_24155);
xor U26827 (N_26827,N_24119,N_25141);
and U26828 (N_26828,N_25660,N_24822);
or U26829 (N_26829,N_25395,N_25632);
nor U26830 (N_26830,N_25845,N_24346);
and U26831 (N_26831,N_25748,N_24070);
xnor U26832 (N_26832,N_25142,N_24543);
and U26833 (N_26833,N_25730,N_24956);
and U26834 (N_26834,N_25455,N_25463);
nor U26835 (N_26835,N_25396,N_24909);
nand U26836 (N_26836,N_24237,N_25047);
or U26837 (N_26837,N_25813,N_25647);
xnor U26838 (N_26838,N_24201,N_25508);
xor U26839 (N_26839,N_25068,N_25575);
nor U26840 (N_26840,N_24992,N_24804);
nor U26841 (N_26841,N_24642,N_24323);
and U26842 (N_26842,N_25044,N_24565);
nand U26843 (N_26843,N_25912,N_24507);
nor U26844 (N_26844,N_25819,N_25862);
nand U26845 (N_26845,N_25346,N_24190);
nand U26846 (N_26846,N_24235,N_25414);
nand U26847 (N_26847,N_24466,N_25450);
xnor U26848 (N_26848,N_25779,N_25581);
nand U26849 (N_26849,N_24115,N_24191);
xor U26850 (N_26850,N_25187,N_25435);
or U26851 (N_26851,N_24000,N_25945);
xor U26852 (N_26852,N_25562,N_25316);
nor U26853 (N_26853,N_25567,N_25054);
or U26854 (N_26854,N_24798,N_25649);
or U26855 (N_26855,N_25482,N_25670);
nor U26856 (N_26856,N_24560,N_24509);
and U26857 (N_26857,N_25622,N_24722);
nor U26858 (N_26858,N_25851,N_25191);
nor U26859 (N_26859,N_24407,N_25556);
nor U26860 (N_26860,N_25334,N_24706);
nand U26861 (N_26861,N_24778,N_24165);
nor U26862 (N_26862,N_24114,N_24406);
xor U26863 (N_26863,N_24073,N_24495);
and U26864 (N_26864,N_25758,N_25708);
xnor U26865 (N_26865,N_24773,N_24784);
nor U26866 (N_26866,N_25540,N_24022);
nand U26867 (N_26867,N_25107,N_24906);
or U26868 (N_26868,N_25277,N_25092);
nor U26869 (N_26869,N_24446,N_24892);
nor U26870 (N_26870,N_25965,N_25791);
nand U26871 (N_26871,N_24376,N_24868);
or U26872 (N_26872,N_24771,N_24694);
and U26873 (N_26873,N_25852,N_25099);
or U26874 (N_26874,N_25771,N_25903);
nor U26875 (N_26875,N_24093,N_24723);
and U26876 (N_26876,N_24078,N_25257);
or U26877 (N_26877,N_25104,N_24938);
nand U26878 (N_26878,N_24889,N_24230);
nor U26879 (N_26879,N_24854,N_24288);
nor U26880 (N_26880,N_25449,N_25728);
and U26881 (N_26881,N_25923,N_25488);
and U26882 (N_26882,N_25050,N_25288);
nor U26883 (N_26883,N_24127,N_25605);
xnor U26884 (N_26884,N_25035,N_24769);
nand U26885 (N_26885,N_25520,N_25897);
nand U26886 (N_26886,N_25985,N_25308);
xnor U26887 (N_26887,N_24936,N_24967);
nand U26888 (N_26888,N_24475,N_24105);
and U26889 (N_26889,N_24448,N_24994);
nand U26890 (N_26890,N_25882,N_24830);
nor U26891 (N_26891,N_24130,N_24970);
xnor U26892 (N_26892,N_25579,N_24641);
or U26893 (N_26893,N_25564,N_24758);
or U26894 (N_26894,N_25919,N_24014);
xnor U26895 (N_26895,N_25712,N_24357);
nand U26896 (N_26896,N_24064,N_24016);
xor U26897 (N_26897,N_25499,N_24785);
and U26898 (N_26898,N_24310,N_24747);
and U26899 (N_26899,N_25312,N_25036);
and U26900 (N_26900,N_25843,N_25046);
nor U26901 (N_26901,N_24882,N_24100);
and U26902 (N_26902,N_24325,N_24301);
and U26903 (N_26903,N_24980,N_25286);
or U26904 (N_26904,N_25407,N_24166);
xor U26905 (N_26905,N_24525,N_24537);
or U26906 (N_26906,N_25933,N_24019);
or U26907 (N_26907,N_24348,N_24386);
nand U26908 (N_26908,N_24949,N_24216);
and U26909 (N_26909,N_25105,N_25022);
or U26910 (N_26910,N_24781,N_25319);
nand U26911 (N_26911,N_25642,N_24396);
and U26912 (N_26912,N_25445,N_25917);
xnor U26913 (N_26913,N_25512,N_24225);
and U26914 (N_26914,N_24986,N_25003);
or U26915 (N_26915,N_25627,N_25699);
nor U26916 (N_26916,N_25394,N_25473);
nor U26917 (N_26917,N_25249,N_25538);
nand U26918 (N_26918,N_24322,N_25175);
or U26919 (N_26919,N_25262,N_24749);
nor U26920 (N_26920,N_25363,N_25048);
and U26921 (N_26921,N_24878,N_24020);
or U26922 (N_26922,N_24199,N_24072);
nand U26923 (N_26923,N_24047,N_24818);
nand U26924 (N_26924,N_24188,N_24656);
xnor U26925 (N_26925,N_25244,N_25405);
or U26926 (N_26926,N_24974,N_25166);
and U26927 (N_26927,N_24421,N_25814);
nor U26928 (N_26928,N_24222,N_25962);
nor U26929 (N_26929,N_24598,N_25083);
nand U26930 (N_26930,N_25431,N_25533);
and U26931 (N_26931,N_24616,N_24531);
xor U26932 (N_26932,N_24669,N_25351);
and U26933 (N_26933,N_24815,N_25668);
and U26934 (N_26934,N_24462,N_24006);
and U26935 (N_26935,N_24482,N_24215);
nand U26936 (N_26936,N_25150,N_25232);
nor U26937 (N_26937,N_25646,N_25064);
xor U26938 (N_26938,N_25764,N_25121);
xnor U26939 (N_26939,N_24578,N_24558);
or U26940 (N_26940,N_24107,N_24353);
nor U26941 (N_26941,N_25038,N_24664);
xor U26942 (N_26942,N_25481,N_24470);
xor U26943 (N_26943,N_24662,N_24076);
nand U26944 (N_26944,N_24677,N_25024);
nand U26945 (N_26945,N_25536,N_25975);
xor U26946 (N_26946,N_25794,N_24816);
or U26947 (N_26947,N_24253,N_24144);
and U26948 (N_26948,N_25159,N_24312);
nor U26949 (N_26949,N_25586,N_24715);
nand U26950 (N_26950,N_25248,N_25052);
or U26951 (N_26951,N_24381,N_24963);
nor U26952 (N_26952,N_25438,N_25952);
xor U26953 (N_26953,N_25303,N_25966);
nand U26954 (N_26954,N_24668,N_25767);
nand U26955 (N_26955,N_25848,N_25164);
nor U26956 (N_26956,N_25062,N_24853);
or U26957 (N_26957,N_24943,N_24431);
or U26958 (N_26958,N_24603,N_25086);
and U26959 (N_26959,N_24120,N_25609);
xor U26960 (N_26960,N_24843,N_24978);
or U26961 (N_26961,N_25525,N_25369);
or U26962 (N_26962,N_25926,N_25144);
or U26963 (N_26963,N_24746,N_25669);
nand U26964 (N_26964,N_25305,N_25406);
and U26965 (N_26965,N_25195,N_25825);
xor U26966 (N_26966,N_24539,N_24536);
nor U26967 (N_26967,N_24691,N_25386);
nor U26968 (N_26968,N_24923,N_25784);
or U26969 (N_26969,N_24811,N_25180);
and U26970 (N_26970,N_25021,N_24368);
nor U26971 (N_26971,N_25950,N_25464);
nand U26972 (N_26972,N_25864,N_24484);
nand U26973 (N_26973,N_24316,N_25500);
xor U26974 (N_26974,N_24109,N_25184);
xor U26975 (N_26975,N_25318,N_24077);
xnor U26976 (N_26976,N_25591,N_25817);
and U26977 (N_26977,N_25799,N_25576);
or U26978 (N_26978,N_25376,N_25094);
or U26979 (N_26979,N_25967,N_25081);
or U26980 (N_26980,N_25378,N_24787);
xnor U26981 (N_26981,N_25703,N_25247);
and U26982 (N_26982,N_24163,N_24106);
nand U26983 (N_26983,N_24517,N_25709);
xor U26984 (N_26984,N_25098,N_25100);
or U26985 (N_26985,N_25941,N_25125);
nand U26986 (N_26986,N_24331,N_25069);
or U26987 (N_26987,N_24460,N_25362);
nor U26988 (N_26988,N_25313,N_25231);
xnor U26989 (N_26989,N_25800,N_24071);
nand U26990 (N_26990,N_25433,N_25687);
and U26991 (N_26991,N_25960,N_24134);
xnor U26992 (N_26992,N_24415,N_25123);
nand U26993 (N_26993,N_24913,N_24547);
nand U26994 (N_26994,N_25725,N_24684);
nand U26995 (N_26995,N_24618,N_25956);
and U26996 (N_26996,N_24112,N_24534);
and U26997 (N_26997,N_25269,N_24498);
nand U26998 (N_26998,N_24512,N_24296);
nor U26999 (N_26999,N_24608,N_24345);
or U27000 (N_27000,N_24718,N_25639);
and U27001 (N_27001,N_24802,N_25680);
nor U27002 (N_27002,N_24056,N_25450);
or U27003 (N_27003,N_24034,N_24508);
nand U27004 (N_27004,N_24771,N_25930);
xnor U27005 (N_27005,N_24241,N_24939);
nand U27006 (N_27006,N_25766,N_24667);
nor U27007 (N_27007,N_24178,N_25954);
nand U27008 (N_27008,N_24868,N_24090);
and U27009 (N_27009,N_24213,N_24460);
nand U27010 (N_27010,N_25807,N_25502);
and U27011 (N_27011,N_24372,N_24486);
xnor U27012 (N_27012,N_24697,N_24506);
xnor U27013 (N_27013,N_24687,N_25499);
or U27014 (N_27014,N_24427,N_25085);
nand U27015 (N_27015,N_24721,N_25261);
or U27016 (N_27016,N_24908,N_25536);
or U27017 (N_27017,N_25737,N_25449);
xor U27018 (N_27018,N_25565,N_24359);
nor U27019 (N_27019,N_24546,N_24543);
and U27020 (N_27020,N_24464,N_24585);
or U27021 (N_27021,N_24426,N_25591);
and U27022 (N_27022,N_24505,N_25429);
xnor U27023 (N_27023,N_25884,N_24530);
or U27024 (N_27024,N_25158,N_25537);
nor U27025 (N_27025,N_25077,N_25860);
xor U27026 (N_27026,N_25113,N_25287);
and U27027 (N_27027,N_24672,N_25670);
or U27028 (N_27028,N_25594,N_25192);
nand U27029 (N_27029,N_25470,N_25734);
nand U27030 (N_27030,N_25179,N_24438);
and U27031 (N_27031,N_25583,N_25692);
xor U27032 (N_27032,N_24871,N_24586);
xor U27033 (N_27033,N_24938,N_24160);
xor U27034 (N_27034,N_25884,N_24667);
or U27035 (N_27035,N_24992,N_24562);
or U27036 (N_27036,N_25583,N_25839);
and U27037 (N_27037,N_25232,N_24959);
xnor U27038 (N_27038,N_24188,N_25028);
and U27039 (N_27039,N_25772,N_25227);
xnor U27040 (N_27040,N_24743,N_24084);
or U27041 (N_27041,N_24176,N_24795);
or U27042 (N_27042,N_25651,N_25049);
xor U27043 (N_27043,N_25288,N_25721);
nor U27044 (N_27044,N_25117,N_25387);
and U27045 (N_27045,N_25230,N_25972);
nand U27046 (N_27046,N_25551,N_24744);
or U27047 (N_27047,N_25603,N_24698);
nor U27048 (N_27048,N_25027,N_24808);
and U27049 (N_27049,N_24116,N_25950);
or U27050 (N_27050,N_24026,N_24688);
nand U27051 (N_27051,N_25865,N_24787);
nor U27052 (N_27052,N_24800,N_25970);
nor U27053 (N_27053,N_25938,N_24226);
and U27054 (N_27054,N_24387,N_24788);
and U27055 (N_27055,N_25204,N_24912);
nor U27056 (N_27056,N_24991,N_24594);
nor U27057 (N_27057,N_25181,N_24566);
or U27058 (N_27058,N_24543,N_25076);
nand U27059 (N_27059,N_24154,N_25775);
xor U27060 (N_27060,N_25718,N_25876);
or U27061 (N_27061,N_25061,N_24336);
and U27062 (N_27062,N_25406,N_25736);
xnor U27063 (N_27063,N_25717,N_24089);
nor U27064 (N_27064,N_25848,N_24061);
xor U27065 (N_27065,N_24879,N_24689);
xnor U27066 (N_27066,N_24217,N_24451);
xnor U27067 (N_27067,N_24506,N_24451);
or U27068 (N_27068,N_25850,N_25702);
and U27069 (N_27069,N_24960,N_25287);
nor U27070 (N_27070,N_25407,N_24567);
nor U27071 (N_27071,N_25914,N_25561);
or U27072 (N_27072,N_25966,N_25869);
and U27073 (N_27073,N_25325,N_24064);
nor U27074 (N_27074,N_24673,N_25743);
or U27075 (N_27075,N_25954,N_24868);
nand U27076 (N_27076,N_25572,N_24058);
xor U27077 (N_27077,N_25874,N_24477);
or U27078 (N_27078,N_24526,N_24500);
nor U27079 (N_27079,N_24924,N_24482);
and U27080 (N_27080,N_24067,N_25627);
nand U27081 (N_27081,N_25414,N_24754);
xor U27082 (N_27082,N_24514,N_24821);
and U27083 (N_27083,N_25795,N_25415);
xnor U27084 (N_27084,N_24061,N_24197);
xnor U27085 (N_27085,N_24259,N_24703);
xor U27086 (N_27086,N_25894,N_25431);
nand U27087 (N_27087,N_25639,N_24711);
nand U27088 (N_27088,N_24509,N_24976);
xnor U27089 (N_27089,N_25777,N_24043);
xor U27090 (N_27090,N_24687,N_25937);
xnor U27091 (N_27091,N_24393,N_25344);
nand U27092 (N_27092,N_25444,N_25291);
and U27093 (N_27093,N_24553,N_24252);
or U27094 (N_27094,N_24652,N_24273);
or U27095 (N_27095,N_24260,N_25111);
xnor U27096 (N_27096,N_25561,N_25688);
nor U27097 (N_27097,N_24197,N_24311);
nand U27098 (N_27098,N_25922,N_24419);
xnor U27099 (N_27099,N_24458,N_25453);
nor U27100 (N_27100,N_25258,N_25399);
or U27101 (N_27101,N_25465,N_25594);
xor U27102 (N_27102,N_25258,N_25286);
or U27103 (N_27103,N_25481,N_24190);
nand U27104 (N_27104,N_24037,N_25922);
or U27105 (N_27105,N_25833,N_25690);
nor U27106 (N_27106,N_25515,N_24011);
or U27107 (N_27107,N_24717,N_24218);
nand U27108 (N_27108,N_24978,N_24517);
nand U27109 (N_27109,N_25245,N_24832);
or U27110 (N_27110,N_25293,N_25661);
or U27111 (N_27111,N_24965,N_24064);
or U27112 (N_27112,N_24891,N_24577);
and U27113 (N_27113,N_25192,N_24324);
xnor U27114 (N_27114,N_25705,N_24456);
xnor U27115 (N_27115,N_24303,N_24737);
xor U27116 (N_27116,N_25355,N_24050);
nand U27117 (N_27117,N_24645,N_25986);
and U27118 (N_27118,N_25974,N_24294);
xnor U27119 (N_27119,N_25638,N_24867);
and U27120 (N_27120,N_24497,N_24580);
nand U27121 (N_27121,N_25698,N_25489);
and U27122 (N_27122,N_24356,N_25838);
xor U27123 (N_27123,N_24087,N_25655);
nand U27124 (N_27124,N_24148,N_25412);
or U27125 (N_27125,N_25075,N_25679);
nor U27126 (N_27126,N_24278,N_24572);
nor U27127 (N_27127,N_24848,N_24775);
and U27128 (N_27128,N_25220,N_25207);
xor U27129 (N_27129,N_25099,N_25483);
xnor U27130 (N_27130,N_24891,N_25439);
xor U27131 (N_27131,N_24241,N_25232);
xnor U27132 (N_27132,N_24120,N_25064);
xnor U27133 (N_27133,N_24364,N_25741);
and U27134 (N_27134,N_25419,N_24708);
nand U27135 (N_27135,N_25621,N_24330);
nand U27136 (N_27136,N_25884,N_24903);
and U27137 (N_27137,N_24262,N_25688);
nand U27138 (N_27138,N_24981,N_25619);
nor U27139 (N_27139,N_24027,N_25440);
and U27140 (N_27140,N_24500,N_25001);
and U27141 (N_27141,N_24571,N_24431);
nand U27142 (N_27142,N_25891,N_24620);
nand U27143 (N_27143,N_25347,N_24400);
and U27144 (N_27144,N_24125,N_25237);
and U27145 (N_27145,N_24751,N_24744);
nand U27146 (N_27146,N_24878,N_24211);
or U27147 (N_27147,N_24423,N_24024);
nand U27148 (N_27148,N_24429,N_24885);
or U27149 (N_27149,N_25849,N_25112);
and U27150 (N_27150,N_25066,N_25141);
nand U27151 (N_27151,N_24845,N_25668);
nor U27152 (N_27152,N_25498,N_25909);
or U27153 (N_27153,N_24600,N_25248);
nand U27154 (N_27154,N_25384,N_25093);
nand U27155 (N_27155,N_24319,N_24156);
and U27156 (N_27156,N_24236,N_25744);
or U27157 (N_27157,N_24120,N_24724);
nand U27158 (N_27158,N_25148,N_25277);
nor U27159 (N_27159,N_25711,N_24133);
nand U27160 (N_27160,N_24602,N_25104);
and U27161 (N_27161,N_25826,N_24232);
or U27162 (N_27162,N_24174,N_24673);
xor U27163 (N_27163,N_25301,N_24990);
or U27164 (N_27164,N_25598,N_25879);
xnor U27165 (N_27165,N_25331,N_24949);
and U27166 (N_27166,N_25821,N_25042);
nand U27167 (N_27167,N_24325,N_24415);
xnor U27168 (N_27168,N_25582,N_24483);
xor U27169 (N_27169,N_24001,N_24894);
and U27170 (N_27170,N_25227,N_25805);
xnor U27171 (N_27171,N_25287,N_25997);
or U27172 (N_27172,N_24048,N_25809);
or U27173 (N_27173,N_24142,N_24333);
nand U27174 (N_27174,N_25905,N_25347);
xor U27175 (N_27175,N_25830,N_24400);
nand U27176 (N_27176,N_25387,N_24121);
or U27177 (N_27177,N_25258,N_24492);
and U27178 (N_27178,N_25630,N_25547);
nand U27179 (N_27179,N_24436,N_25642);
nor U27180 (N_27180,N_24267,N_24546);
or U27181 (N_27181,N_25942,N_24213);
and U27182 (N_27182,N_25900,N_25584);
or U27183 (N_27183,N_25434,N_24145);
or U27184 (N_27184,N_25462,N_24577);
nand U27185 (N_27185,N_25241,N_24043);
or U27186 (N_27186,N_24770,N_24205);
and U27187 (N_27187,N_25914,N_25759);
nand U27188 (N_27188,N_24060,N_24588);
nand U27189 (N_27189,N_25323,N_24606);
xor U27190 (N_27190,N_24235,N_24165);
xnor U27191 (N_27191,N_25331,N_24619);
nand U27192 (N_27192,N_25834,N_24516);
or U27193 (N_27193,N_25284,N_25663);
xnor U27194 (N_27194,N_24313,N_24102);
and U27195 (N_27195,N_24476,N_25267);
nor U27196 (N_27196,N_25731,N_24724);
nand U27197 (N_27197,N_24536,N_24914);
or U27198 (N_27198,N_25825,N_25573);
nand U27199 (N_27199,N_25812,N_24046);
nor U27200 (N_27200,N_24099,N_25202);
nor U27201 (N_27201,N_25626,N_24033);
nand U27202 (N_27202,N_25318,N_25826);
and U27203 (N_27203,N_24519,N_25162);
nand U27204 (N_27204,N_24816,N_24333);
nor U27205 (N_27205,N_25484,N_25626);
xor U27206 (N_27206,N_25681,N_24528);
nor U27207 (N_27207,N_25350,N_24300);
and U27208 (N_27208,N_24440,N_25196);
xor U27209 (N_27209,N_25076,N_25721);
nor U27210 (N_27210,N_25047,N_25066);
nand U27211 (N_27211,N_24230,N_25769);
or U27212 (N_27212,N_24724,N_25658);
or U27213 (N_27213,N_25790,N_25072);
xnor U27214 (N_27214,N_25060,N_25564);
and U27215 (N_27215,N_24471,N_24778);
nand U27216 (N_27216,N_24956,N_25081);
xnor U27217 (N_27217,N_25638,N_24858);
nand U27218 (N_27218,N_25494,N_25599);
xnor U27219 (N_27219,N_24517,N_24710);
or U27220 (N_27220,N_24918,N_25499);
nand U27221 (N_27221,N_25300,N_24686);
nor U27222 (N_27222,N_24393,N_24427);
xnor U27223 (N_27223,N_24150,N_25383);
nand U27224 (N_27224,N_24714,N_24398);
or U27225 (N_27225,N_25956,N_25392);
nand U27226 (N_27226,N_25254,N_24333);
xor U27227 (N_27227,N_24753,N_25713);
xnor U27228 (N_27228,N_25765,N_25736);
xnor U27229 (N_27229,N_25656,N_24326);
and U27230 (N_27230,N_24203,N_25114);
xnor U27231 (N_27231,N_25065,N_24170);
nand U27232 (N_27232,N_25428,N_25993);
nand U27233 (N_27233,N_25796,N_25134);
nor U27234 (N_27234,N_24497,N_25113);
or U27235 (N_27235,N_25855,N_25538);
xnor U27236 (N_27236,N_25842,N_24711);
nand U27237 (N_27237,N_24401,N_25160);
nand U27238 (N_27238,N_24046,N_25440);
xnor U27239 (N_27239,N_24916,N_25033);
and U27240 (N_27240,N_24217,N_24982);
nor U27241 (N_27241,N_24679,N_24127);
or U27242 (N_27242,N_25162,N_24483);
nor U27243 (N_27243,N_25058,N_24360);
nor U27244 (N_27244,N_25204,N_24551);
nor U27245 (N_27245,N_24258,N_25032);
or U27246 (N_27246,N_25532,N_25033);
or U27247 (N_27247,N_25729,N_25575);
nand U27248 (N_27248,N_24231,N_24703);
xnor U27249 (N_27249,N_25432,N_24100);
or U27250 (N_27250,N_25193,N_25015);
nand U27251 (N_27251,N_24731,N_25921);
and U27252 (N_27252,N_24015,N_25019);
xnor U27253 (N_27253,N_25919,N_24895);
and U27254 (N_27254,N_24942,N_24718);
and U27255 (N_27255,N_25645,N_25098);
nand U27256 (N_27256,N_25393,N_24077);
and U27257 (N_27257,N_25188,N_24373);
nor U27258 (N_27258,N_25867,N_25278);
nor U27259 (N_27259,N_24603,N_24833);
xnor U27260 (N_27260,N_24861,N_25208);
nor U27261 (N_27261,N_24340,N_25274);
xnor U27262 (N_27262,N_24602,N_25057);
or U27263 (N_27263,N_25135,N_25140);
or U27264 (N_27264,N_24862,N_24115);
xnor U27265 (N_27265,N_25133,N_24822);
nand U27266 (N_27266,N_24921,N_24540);
and U27267 (N_27267,N_24915,N_25642);
and U27268 (N_27268,N_25584,N_24524);
and U27269 (N_27269,N_24595,N_24046);
xor U27270 (N_27270,N_25933,N_24072);
xnor U27271 (N_27271,N_24819,N_24192);
and U27272 (N_27272,N_24476,N_24523);
or U27273 (N_27273,N_24672,N_25815);
nor U27274 (N_27274,N_24381,N_25280);
nand U27275 (N_27275,N_24361,N_25257);
and U27276 (N_27276,N_24301,N_25403);
and U27277 (N_27277,N_25747,N_25887);
nor U27278 (N_27278,N_25591,N_24693);
nand U27279 (N_27279,N_25165,N_25493);
and U27280 (N_27280,N_25180,N_25741);
nand U27281 (N_27281,N_25451,N_25773);
or U27282 (N_27282,N_25028,N_24979);
nor U27283 (N_27283,N_25511,N_25368);
nand U27284 (N_27284,N_24989,N_24694);
nand U27285 (N_27285,N_24734,N_24139);
nor U27286 (N_27286,N_25527,N_24819);
nand U27287 (N_27287,N_24846,N_24148);
nor U27288 (N_27288,N_25012,N_24554);
or U27289 (N_27289,N_24453,N_25986);
and U27290 (N_27290,N_25037,N_25623);
or U27291 (N_27291,N_24880,N_24115);
or U27292 (N_27292,N_24410,N_24024);
xnor U27293 (N_27293,N_25142,N_24972);
nor U27294 (N_27294,N_24770,N_25940);
nand U27295 (N_27295,N_25618,N_25013);
nand U27296 (N_27296,N_24372,N_25369);
nand U27297 (N_27297,N_25242,N_24368);
nor U27298 (N_27298,N_24154,N_25157);
nor U27299 (N_27299,N_24505,N_25997);
nor U27300 (N_27300,N_25141,N_24510);
and U27301 (N_27301,N_25171,N_24790);
nand U27302 (N_27302,N_25585,N_25646);
and U27303 (N_27303,N_25503,N_25386);
nor U27304 (N_27304,N_25062,N_25053);
or U27305 (N_27305,N_24171,N_25341);
nor U27306 (N_27306,N_24026,N_25891);
and U27307 (N_27307,N_24018,N_24768);
nor U27308 (N_27308,N_25261,N_24343);
nand U27309 (N_27309,N_25153,N_25977);
and U27310 (N_27310,N_25766,N_24460);
or U27311 (N_27311,N_24824,N_25654);
and U27312 (N_27312,N_25249,N_25156);
xor U27313 (N_27313,N_25016,N_24402);
nor U27314 (N_27314,N_25512,N_24644);
nor U27315 (N_27315,N_24562,N_25001);
and U27316 (N_27316,N_25894,N_24047);
nor U27317 (N_27317,N_25593,N_24667);
and U27318 (N_27318,N_25683,N_24763);
or U27319 (N_27319,N_24560,N_24553);
nor U27320 (N_27320,N_25902,N_24687);
nor U27321 (N_27321,N_25135,N_24420);
or U27322 (N_27322,N_25039,N_24004);
nor U27323 (N_27323,N_25624,N_24724);
nand U27324 (N_27324,N_25821,N_24741);
xor U27325 (N_27325,N_24947,N_24323);
or U27326 (N_27326,N_25623,N_25473);
or U27327 (N_27327,N_24699,N_25929);
nand U27328 (N_27328,N_25850,N_25986);
and U27329 (N_27329,N_24836,N_25480);
nand U27330 (N_27330,N_25852,N_25355);
or U27331 (N_27331,N_25210,N_24670);
nor U27332 (N_27332,N_25639,N_24136);
nand U27333 (N_27333,N_25319,N_24091);
xor U27334 (N_27334,N_25743,N_25749);
or U27335 (N_27335,N_24973,N_25355);
nor U27336 (N_27336,N_24010,N_25585);
xor U27337 (N_27337,N_25879,N_24854);
nand U27338 (N_27338,N_24731,N_24251);
xor U27339 (N_27339,N_24874,N_24340);
or U27340 (N_27340,N_25594,N_24482);
nor U27341 (N_27341,N_25875,N_24240);
nand U27342 (N_27342,N_24100,N_25062);
or U27343 (N_27343,N_25100,N_24619);
or U27344 (N_27344,N_25741,N_24672);
and U27345 (N_27345,N_24656,N_25318);
nor U27346 (N_27346,N_24810,N_25716);
nor U27347 (N_27347,N_25220,N_24578);
nand U27348 (N_27348,N_24236,N_24368);
nand U27349 (N_27349,N_25921,N_24511);
nor U27350 (N_27350,N_25964,N_24067);
and U27351 (N_27351,N_24242,N_24950);
xnor U27352 (N_27352,N_25207,N_24975);
nor U27353 (N_27353,N_25644,N_25076);
and U27354 (N_27354,N_24773,N_25488);
or U27355 (N_27355,N_25612,N_25264);
xnor U27356 (N_27356,N_25904,N_25944);
or U27357 (N_27357,N_24123,N_25852);
xor U27358 (N_27358,N_25523,N_25355);
nand U27359 (N_27359,N_25809,N_24834);
nand U27360 (N_27360,N_24658,N_24294);
nor U27361 (N_27361,N_24914,N_25951);
nand U27362 (N_27362,N_24857,N_25635);
and U27363 (N_27363,N_25288,N_24205);
and U27364 (N_27364,N_24898,N_25347);
and U27365 (N_27365,N_25027,N_24852);
and U27366 (N_27366,N_24225,N_24554);
xnor U27367 (N_27367,N_24276,N_24636);
or U27368 (N_27368,N_24519,N_25770);
xnor U27369 (N_27369,N_24477,N_24178);
nor U27370 (N_27370,N_24158,N_24350);
nor U27371 (N_27371,N_25138,N_24664);
and U27372 (N_27372,N_25315,N_25183);
and U27373 (N_27373,N_24320,N_25959);
xor U27374 (N_27374,N_25056,N_24431);
or U27375 (N_27375,N_25551,N_25189);
nor U27376 (N_27376,N_25061,N_24564);
xor U27377 (N_27377,N_25552,N_25057);
xnor U27378 (N_27378,N_25677,N_24848);
or U27379 (N_27379,N_24590,N_24753);
nand U27380 (N_27380,N_25034,N_24190);
or U27381 (N_27381,N_25595,N_25076);
nand U27382 (N_27382,N_24074,N_24340);
nor U27383 (N_27383,N_24253,N_24465);
or U27384 (N_27384,N_25171,N_24796);
and U27385 (N_27385,N_25860,N_25603);
nand U27386 (N_27386,N_24688,N_24352);
or U27387 (N_27387,N_25351,N_24719);
xnor U27388 (N_27388,N_24807,N_24475);
and U27389 (N_27389,N_25899,N_25129);
nor U27390 (N_27390,N_24623,N_25709);
or U27391 (N_27391,N_24748,N_24654);
xnor U27392 (N_27392,N_24421,N_24945);
or U27393 (N_27393,N_25094,N_25167);
and U27394 (N_27394,N_25767,N_24944);
nand U27395 (N_27395,N_24283,N_25036);
and U27396 (N_27396,N_24298,N_24655);
or U27397 (N_27397,N_25129,N_24798);
nor U27398 (N_27398,N_24662,N_24378);
and U27399 (N_27399,N_24842,N_24460);
xnor U27400 (N_27400,N_24284,N_24176);
nand U27401 (N_27401,N_25543,N_25118);
nor U27402 (N_27402,N_24589,N_24602);
and U27403 (N_27403,N_25618,N_24086);
nand U27404 (N_27404,N_24720,N_25337);
xor U27405 (N_27405,N_24133,N_25413);
nor U27406 (N_27406,N_24832,N_24716);
nor U27407 (N_27407,N_24821,N_25380);
nand U27408 (N_27408,N_25744,N_24016);
xnor U27409 (N_27409,N_25887,N_25721);
nor U27410 (N_27410,N_25345,N_24980);
nand U27411 (N_27411,N_24156,N_24691);
or U27412 (N_27412,N_24938,N_24053);
nand U27413 (N_27413,N_24242,N_24553);
nand U27414 (N_27414,N_24407,N_24339);
nor U27415 (N_27415,N_24182,N_24366);
xor U27416 (N_27416,N_24721,N_24808);
and U27417 (N_27417,N_25058,N_24287);
and U27418 (N_27418,N_24731,N_25134);
xnor U27419 (N_27419,N_25216,N_24782);
or U27420 (N_27420,N_24695,N_24008);
or U27421 (N_27421,N_25154,N_25804);
xnor U27422 (N_27422,N_24806,N_25216);
nor U27423 (N_27423,N_25498,N_25780);
or U27424 (N_27424,N_25046,N_24036);
xor U27425 (N_27425,N_24998,N_24437);
nand U27426 (N_27426,N_25609,N_24261);
and U27427 (N_27427,N_25744,N_25472);
xor U27428 (N_27428,N_25291,N_25273);
nor U27429 (N_27429,N_25922,N_25009);
nor U27430 (N_27430,N_25787,N_24851);
or U27431 (N_27431,N_25177,N_25309);
or U27432 (N_27432,N_24184,N_24674);
nor U27433 (N_27433,N_24663,N_24743);
nand U27434 (N_27434,N_25321,N_25405);
nor U27435 (N_27435,N_24551,N_25273);
or U27436 (N_27436,N_24869,N_24691);
and U27437 (N_27437,N_24141,N_25538);
nor U27438 (N_27438,N_24002,N_25468);
nand U27439 (N_27439,N_25135,N_24616);
nand U27440 (N_27440,N_25106,N_24778);
nor U27441 (N_27441,N_25905,N_24334);
nor U27442 (N_27442,N_24595,N_24597);
nand U27443 (N_27443,N_24819,N_25718);
or U27444 (N_27444,N_25689,N_25840);
or U27445 (N_27445,N_24654,N_25040);
xnor U27446 (N_27446,N_25166,N_24753);
nor U27447 (N_27447,N_25212,N_25274);
and U27448 (N_27448,N_24427,N_24968);
or U27449 (N_27449,N_24843,N_25211);
xor U27450 (N_27450,N_25451,N_24515);
nand U27451 (N_27451,N_25510,N_25746);
nor U27452 (N_27452,N_24165,N_25278);
nand U27453 (N_27453,N_25032,N_24206);
or U27454 (N_27454,N_24596,N_24436);
and U27455 (N_27455,N_25217,N_24843);
nor U27456 (N_27456,N_25406,N_24400);
xnor U27457 (N_27457,N_25250,N_24797);
xor U27458 (N_27458,N_24422,N_24284);
and U27459 (N_27459,N_24356,N_25731);
nor U27460 (N_27460,N_24623,N_24124);
nor U27461 (N_27461,N_24528,N_25313);
xor U27462 (N_27462,N_25671,N_25560);
xnor U27463 (N_27463,N_25875,N_25028);
nand U27464 (N_27464,N_25566,N_25729);
and U27465 (N_27465,N_24050,N_25272);
or U27466 (N_27466,N_24970,N_25718);
or U27467 (N_27467,N_25113,N_24996);
and U27468 (N_27468,N_24925,N_24713);
or U27469 (N_27469,N_24171,N_24030);
and U27470 (N_27470,N_25785,N_25968);
and U27471 (N_27471,N_24484,N_24218);
and U27472 (N_27472,N_25175,N_25762);
nor U27473 (N_27473,N_24341,N_24434);
and U27474 (N_27474,N_24644,N_24296);
xnor U27475 (N_27475,N_25795,N_24185);
xor U27476 (N_27476,N_25337,N_25836);
and U27477 (N_27477,N_24165,N_24998);
nand U27478 (N_27478,N_24254,N_24129);
nor U27479 (N_27479,N_24223,N_24314);
xor U27480 (N_27480,N_25595,N_25214);
nor U27481 (N_27481,N_25126,N_24533);
nand U27482 (N_27482,N_25989,N_25408);
nor U27483 (N_27483,N_25064,N_24423);
nand U27484 (N_27484,N_25976,N_24026);
or U27485 (N_27485,N_25335,N_25240);
or U27486 (N_27486,N_24203,N_25624);
nor U27487 (N_27487,N_24582,N_24319);
and U27488 (N_27488,N_25441,N_24044);
xor U27489 (N_27489,N_25048,N_24786);
xor U27490 (N_27490,N_25464,N_25102);
nor U27491 (N_27491,N_24474,N_25680);
nor U27492 (N_27492,N_24972,N_24149);
and U27493 (N_27493,N_24061,N_24718);
nor U27494 (N_27494,N_24430,N_24744);
nand U27495 (N_27495,N_24700,N_24009);
and U27496 (N_27496,N_24459,N_25781);
xor U27497 (N_27497,N_24978,N_25762);
nand U27498 (N_27498,N_24902,N_25737);
or U27499 (N_27499,N_24118,N_25267);
or U27500 (N_27500,N_24756,N_24766);
and U27501 (N_27501,N_24695,N_25673);
or U27502 (N_27502,N_24577,N_25691);
nand U27503 (N_27503,N_24759,N_24569);
or U27504 (N_27504,N_24533,N_24620);
and U27505 (N_27505,N_25901,N_24470);
nor U27506 (N_27506,N_24205,N_25546);
or U27507 (N_27507,N_24151,N_24699);
and U27508 (N_27508,N_24266,N_24074);
or U27509 (N_27509,N_25547,N_25658);
or U27510 (N_27510,N_25224,N_24203);
or U27511 (N_27511,N_24317,N_24982);
and U27512 (N_27512,N_24351,N_24353);
nor U27513 (N_27513,N_24767,N_24989);
nor U27514 (N_27514,N_24031,N_24928);
and U27515 (N_27515,N_24365,N_24742);
or U27516 (N_27516,N_24490,N_25130);
and U27517 (N_27517,N_25163,N_25435);
nor U27518 (N_27518,N_25035,N_25038);
nand U27519 (N_27519,N_25155,N_25552);
or U27520 (N_27520,N_25284,N_25424);
or U27521 (N_27521,N_25043,N_24178);
nor U27522 (N_27522,N_25048,N_24389);
nor U27523 (N_27523,N_24521,N_25572);
xnor U27524 (N_27524,N_25402,N_25545);
or U27525 (N_27525,N_25068,N_24535);
and U27526 (N_27526,N_24518,N_25752);
and U27527 (N_27527,N_25254,N_25893);
nor U27528 (N_27528,N_24052,N_25240);
nor U27529 (N_27529,N_25081,N_24921);
nor U27530 (N_27530,N_24557,N_25059);
nor U27531 (N_27531,N_25490,N_24438);
or U27532 (N_27532,N_25932,N_24796);
nor U27533 (N_27533,N_25105,N_25348);
nand U27534 (N_27534,N_24080,N_25531);
xnor U27535 (N_27535,N_25011,N_24203);
nor U27536 (N_27536,N_24100,N_24343);
xor U27537 (N_27537,N_24846,N_25915);
nor U27538 (N_27538,N_24050,N_25929);
nor U27539 (N_27539,N_24720,N_24323);
nand U27540 (N_27540,N_25342,N_25163);
nand U27541 (N_27541,N_24863,N_24077);
nand U27542 (N_27542,N_24836,N_25890);
nand U27543 (N_27543,N_24711,N_25116);
nor U27544 (N_27544,N_24393,N_24455);
nor U27545 (N_27545,N_25353,N_24801);
xnor U27546 (N_27546,N_24532,N_25438);
and U27547 (N_27547,N_25645,N_24864);
xor U27548 (N_27548,N_25551,N_24844);
nor U27549 (N_27549,N_24087,N_24943);
nor U27550 (N_27550,N_24920,N_25890);
and U27551 (N_27551,N_24197,N_24147);
or U27552 (N_27552,N_25082,N_25382);
nor U27553 (N_27553,N_25154,N_24147);
xor U27554 (N_27554,N_25576,N_24762);
nand U27555 (N_27555,N_24512,N_25627);
and U27556 (N_27556,N_24637,N_24977);
nor U27557 (N_27557,N_25406,N_25409);
and U27558 (N_27558,N_25395,N_25209);
or U27559 (N_27559,N_24930,N_24949);
or U27560 (N_27560,N_24462,N_25619);
nor U27561 (N_27561,N_24427,N_24261);
or U27562 (N_27562,N_24640,N_24350);
or U27563 (N_27563,N_24432,N_24535);
nor U27564 (N_27564,N_24957,N_24955);
nand U27565 (N_27565,N_25078,N_24972);
or U27566 (N_27566,N_25022,N_25093);
or U27567 (N_27567,N_25679,N_25911);
nand U27568 (N_27568,N_25967,N_24845);
xnor U27569 (N_27569,N_25005,N_24604);
nor U27570 (N_27570,N_24951,N_25507);
nand U27571 (N_27571,N_24709,N_25198);
and U27572 (N_27572,N_24126,N_25440);
nor U27573 (N_27573,N_25531,N_24319);
nand U27574 (N_27574,N_25051,N_24292);
xor U27575 (N_27575,N_24182,N_25220);
xnor U27576 (N_27576,N_25947,N_24701);
xnor U27577 (N_27577,N_25179,N_24727);
nor U27578 (N_27578,N_25240,N_24337);
or U27579 (N_27579,N_24202,N_25468);
nor U27580 (N_27580,N_24740,N_25930);
xnor U27581 (N_27581,N_24396,N_25126);
and U27582 (N_27582,N_24706,N_24545);
and U27583 (N_27583,N_24556,N_25301);
and U27584 (N_27584,N_25448,N_24799);
and U27585 (N_27585,N_25746,N_25193);
nor U27586 (N_27586,N_25577,N_25988);
xor U27587 (N_27587,N_24309,N_24017);
and U27588 (N_27588,N_25627,N_24751);
and U27589 (N_27589,N_24313,N_25549);
nand U27590 (N_27590,N_24660,N_25390);
xor U27591 (N_27591,N_24813,N_24831);
or U27592 (N_27592,N_24522,N_24105);
xnor U27593 (N_27593,N_25863,N_24686);
and U27594 (N_27594,N_24456,N_24908);
nor U27595 (N_27595,N_24807,N_24371);
or U27596 (N_27596,N_25077,N_25151);
nor U27597 (N_27597,N_25969,N_24931);
xnor U27598 (N_27598,N_25172,N_24655);
or U27599 (N_27599,N_24923,N_25625);
or U27600 (N_27600,N_25789,N_25128);
nand U27601 (N_27601,N_24737,N_24339);
or U27602 (N_27602,N_25360,N_24698);
xor U27603 (N_27603,N_24367,N_25492);
xnor U27604 (N_27604,N_24796,N_24087);
or U27605 (N_27605,N_25374,N_24746);
or U27606 (N_27606,N_25537,N_24034);
and U27607 (N_27607,N_25495,N_25061);
or U27608 (N_27608,N_25813,N_25050);
xnor U27609 (N_27609,N_24533,N_24084);
nor U27610 (N_27610,N_24507,N_25147);
nor U27611 (N_27611,N_25737,N_24966);
or U27612 (N_27612,N_24118,N_25720);
xor U27613 (N_27613,N_24810,N_25141);
nand U27614 (N_27614,N_25513,N_25190);
and U27615 (N_27615,N_24035,N_25856);
and U27616 (N_27616,N_25046,N_24408);
nor U27617 (N_27617,N_25620,N_25194);
nor U27618 (N_27618,N_24855,N_25899);
and U27619 (N_27619,N_24860,N_24280);
nand U27620 (N_27620,N_24155,N_25150);
or U27621 (N_27621,N_24365,N_25115);
xnor U27622 (N_27622,N_25446,N_24065);
xor U27623 (N_27623,N_24895,N_25834);
nor U27624 (N_27624,N_24592,N_24760);
or U27625 (N_27625,N_25932,N_24372);
and U27626 (N_27626,N_25071,N_24143);
or U27627 (N_27627,N_25616,N_24877);
nor U27628 (N_27628,N_24381,N_24447);
or U27629 (N_27629,N_25174,N_24941);
and U27630 (N_27630,N_25211,N_24937);
xor U27631 (N_27631,N_25070,N_25338);
or U27632 (N_27632,N_25895,N_25379);
or U27633 (N_27633,N_25254,N_24797);
and U27634 (N_27634,N_24812,N_25534);
nand U27635 (N_27635,N_24518,N_24590);
xnor U27636 (N_27636,N_25484,N_24029);
nand U27637 (N_27637,N_24421,N_24800);
or U27638 (N_27638,N_24610,N_24245);
xnor U27639 (N_27639,N_24201,N_24024);
or U27640 (N_27640,N_24016,N_24789);
xnor U27641 (N_27641,N_24048,N_24623);
or U27642 (N_27642,N_25050,N_25780);
nand U27643 (N_27643,N_24965,N_24399);
or U27644 (N_27644,N_25325,N_25893);
nand U27645 (N_27645,N_25130,N_25600);
xnor U27646 (N_27646,N_24244,N_24261);
and U27647 (N_27647,N_25867,N_24062);
xnor U27648 (N_27648,N_25237,N_24776);
xor U27649 (N_27649,N_25171,N_24244);
nand U27650 (N_27650,N_25087,N_25889);
nor U27651 (N_27651,N_25995,N_25581);
nor U27652 (N_27652,N_25120,N_24151);
nor U27653 (N_27653,N_24350,N_24592);
nor U27654 (N_27654,N_25818,N_24893);
or U27655 (N_27655,N_25811,N_25590);
xnor U27656 (N_27656,N_25502,N_25131);
or U27657 (N_27657,N_25221,N_24851);
xnor U27658 (N_27658,N_24194,N_25031);
nor U27659 (N_27659,N_25253,N_24491);
and U27660 (N_27660,N_25984,N_24507);
nor U27661 (N_27661,N_25610,N_25819);
nor U27662 (N_27662,N_25414,N_25681);
or U27663 (N_27663,N_25844,N_25003);
nand U27664 (N_27664,N_24212,N_25215);
nand U27665 (N_27665,N_25027,N_24656);
xnor U27666 (N_27666,N_24734,N_24428);
nor U27667 (N_27667,N_24130,N_25268);
xnor U27668 (N_27668,N_25572,N_25196);
xor U27669 (N_27669,N_25613,N_25602);
and U27670 (N_27670,N_24143,N_24201);
nand U27671 (N_27671,N_25088,N_25206);
nor U27672 (N_27672,N_24500,N_25779);
xnor U27673 (N_27673,N_25840,N_25096);
and U27674 (N_27674,N_25052,N_25763);
or U27675 (N_27675,N_24038,N_24894);
nor U27676 (N_27676,N_24558,N_25373);
xnor U27677 (N_27677,N_25702,N_24940);
nand U27678 (N_27678,N_24173,N_24501);
xnor U27679 (N_27679,N_25099,N_24414);
or U27680 (N_27680,N_25727,N_25644);
and U27681 (N_27681,N_25559,N_25731);
nand U27682 (N_27682,N_25633,N_25975);
and U27683 (N_27683,N_25980,N_25139);
nand U27684 (N_27684,N_25808,N_25490);
nor U27685 (N_27685,N_25571,N_25086);
nand U27686 (N_27686,N_24304,N_24375);
or U27687 (N_27687,N_25818,N_24734);
nand U27688 (N_27688,N_25587,N_25603);
nand U27689 (N_27689,N_25251,N_25195);
xor U27690 (N_27690,N_25463,N_24373);
xor U27691 (N_27691,N_25359,N_24227);
or U27692 (N_27692,N_24679,N_24188);
or U27693 (N_27693,N_25179,N_24805);
or U27694 (N_27694,N_25732,N_24583);
nand U27695 (N_27695,N_25797,N_25400);
and U27696 (N_27696,N_25889,N_25448);
xnor U27697 (N_27697,N_25681,N_25589);
and U27698 (N_27698,N_25990,N_25837);
nor U27699 (N_27699,N_24252,N_24601);
nor U27700 (N_27700,N_25033,N_25573);
and U27701 (N_27701,N_25081,N_25725);
nand U27702 (N_27702,N_24013,N_24396);
nor U27703 (N_27703,N_24982,N_25006);
nand U27704 (N_27704,N_24021,N_24730);
nand U27705 (N_27705,N_25010,N_25583);
and U27706 (N_27706,N_25812,N_25832);
nor U27707 (N_27707,N_24995,N_24045);
nand U27708 (N_27708,N_25108,N_25919);
nor U27709 (N_27709,N_24907,N_25839);
nor U27710 (N_27710,N_25597,N_24558);
and U27711 (N_27711,N_24167,N_25373);
or U27712 (N_27712,N_25486,N_24118);
nor U27713 (N_27713,N_25398,N_24714);
nand U27714 (N_27714,N_25412,N_24198);
or U27715 (N_27715,N_25426,N_24671);
xor U27716 (N_27716,N_24263,N_25791);
nand U27717 (N_27717,N_25770,N_25213);
and U27718 (N_27718,N_24740,N_25861);
or U27719 (N_27719,N_25869,N_25766);
or U27720 (N_27720,N_25248,N_25188);
xor U27721 (N_27721,N_25842,N_25598);
or U27722 (N_27722,N_25545,N_25373);
or U27723 (N_27723,N_24486,N_24177);
nor U27724 (N_27724,N_25597,N_24637);
xnor U27725 (N_27725,N_25210,N_24707);
or U27726 (N_27726,N_25384,N_25867);
or U27727 (N_27727,N_24072,N_24417);
and U27728 (N_27728,N_25838,N_25591);
and U27729 (N_27729,N_24115,N_24143);
and U27730 (N_27730,N_25412,N_25247);
nand U27731 (N_27731,N_24733,N_24034);
nor U27732 (N_27732,N_24445,N_25926);
xnor U27733 (N_27733,N_25735,N_25272);
or U27734 (N_27734,N_25666,N_24175);
or U27735 (N_27735,N_25867,N_24741);
or U27736 (N_27736,N_25849,N_25668);
and U27737 (N_27737,N_24935,N_24100);
and U27738 (N_27738,N_25902,N_25346);
nor U27739 (N_27739,N_24696,N_25363);
or U27740 (N_27740,N_25066,N_24367);
nand U27741 (N_27741,N_24898,N_24147);
nand U27742 (N_27742,N_25787,N_25594);
nor U27743 (N_27743,N_25178,N_24254);
xor U27744 (N_27744,N_25827,N_25973);
xnor U27745 (N_27745,N_25710,N_24965);
and U27746 (N_27746,N_24979,N_25060);
xnor U27747 (N_27747,N_25821,N_25269);
nor U27748 (N_27748,N_25367,N_24964);
nand U27749 (N_27749,N_25580,N_25040);
nor U27750 (N_27750,N_24105,N_24538);
nor U27751 (N_27751,N_25480,N_25315);
xor U27752 (N_27752,N_24370,N_24098);
nor U27753 (N_27753,N_25468,N_25945);
or U27754 (N_27754,N_25668,N_25164);
or U27755 (N_27755,N_24321,N_25835);
nand U27756 (N_27756,N_25754,N_24079);
xor U27757 (N_27757,N_25089,N_24229);
nand U27758 (N_27758,N_24404,N_25061);
nor U27759 (N_27759,N_24790,N_24092);
nand U27760 (N_27760,N_25607,N_24462);
or U27761 (N_27761,N_25464,N_25878);
and U27762 (N_27762,N_25080,N_25634);
and U27763 (N_27763,N_25050,N_24829);
nor U27764 (N_27764,N_25028,N_25603);
and U27765 (N_27765,N_25468,N_24830);
nor U27766 (N_27766,N_24864,N_24304);
or U27767 (N_27767,N_24494,N_24383);
nor U27768 (N_27768,N_24670,N_24938);
and U27769 (N_27769,N_25978,N_24242);
nor U27770 (N_27770,N_25545,N_25597);
nor U27771 (N_27771,N_25305,N_24194);
xnor U27772 (N_27772,N_24269,N_24602);
nand U27773 (N_27773,N_25704,N_25396);
or U27774 (N_27774,N_24324,N_24203);
nand U27775 (N_27775,N_25919,N_25683);
xnor U27776 (N_27776,N_25628,N_24830);
nand U27777 (N_27777,N_25032,N_24956);
and U27778 (N_27778,N_25803,N_24218);
and U27779 (N_27779,N_25478,N_25974);
or U27780 (N_27780,N_24691,N_25538);
xor U27781 (N_27781,N_24490,N_25533);
nor U27782 (N_27782,N_25852,N_25507);
or U27783 (N_27783,N_24641,N_24801);
and U27784 (N_27784,N_24426,N_24206);
nor U27785 (N_27785,N_25276,N_25647);
nand U27786 (N_27786,N_25092,N_24176);
nand U27787 (N_27787,N_25748,N_24766);
xor U27788 (N_27788,N_24668,N_25501);
and U27789 (N_27789,N_24843,N_24393);
nand U27790 (N_27790,N_24542,N_25426);
nand U27791 (N_27791,N_24213,N_25384);
nor U27792 (N_27792,N_24457,N_25148);
nor U27793 (N_27793,N_25875,N_25136);
nor U27794 (N_27794,N_24218,N_24200);
nor U27795 (N_27795,N_24928,N_24323);
or U27796 (N_27796,N_25078,N_24464);
xnor U27797 (N_27797,N_24921,N_25593);
or U27798 (N_27798,N_25082,N_25549);
xor U27799 (N_27799,N_24970,N_25279);
nand U27800 (N_27800,N_25244,N_25060);
xnor U27801 (N_27801,N_25270,N_24572);
xor U27802 (N_27802,N_25622,N_24225);
nor U27803 (N_27803,N_24947,N_24091);
nand U27804 (N_27804,N_25803,N_25203);
nand U27805 (N_27805,N_24727,N_24876);
nor U27806 (N_27806,N_24933,N_24056);
xor U27807 (N_27807,N_24911,N_24466);
nand U27808 (N_27808,N_25358,N_24080);
nand U27809 (N_27809,N_24742,N_25082);
or U27810 (N_27810,N_24228,N_25540);
nor U27811 (N_27811,N_24704,N_25972);
or U27812 (N_27812,N_25625,N_24284);
and U27813 (N_27813,N_24084,N_24473);
nand U27814 (N_27814,N_24778,N_24804);
xor U27815 (N_27815,N_25453,N_25842);
or U27816 (N_27816,N_25366,N_24915);
or U27817 (N_27817,N_25298,N_25503);
nand U27818 (N_27818,N_24237,N_25869);
nand U27819 (N_27819,N_25439,N_25836);
xor U27820 (N_27820,N_24861,N_25822);
nor U27821 (N_27821,N_25709,N_25070);
xor U27822 (N_27822,N_24811,N_24960);
xnor U27823 (N_27823,N_25627,N_24382);
and U27824 (N_27824,N_24857,N_25373);
or U27825 (N_27825,N_25602,N_24740);
xor U27826 (N_27826,N_24703,N_25542);
nor U27827 (N_27827,N_24721,N_24331);
nor U27828 (N_27828,N_25280,N_24249);
nand U27829 (N_27829,N_24413,N_24071);
and U27830 (N_27830,N_24225,N_25797);
nor U27831 (N_27831,N_25429,N_24849);
and U27832 (N_27832,N_25108,N_25813);
and U27833 (N_27833,N_25349,N_25113);
or U27834 (N_27834,N_25008,N_24447);
nor U27835 (N_27835,N_25248,N_24449);
nor U27836 (N_27836,N_24294,N_25470);
xor U27837 (N_27837,N_24766,N_25128);
nand U27838 (N_27838,N_24851,N_25775);
xor U27839 (N_27839,N_25650,N_25174);
and U27840 (N_27840,N_24680,N_24178);
nand U27841 (N_27841,N_25172,N_24910);
nand U27842 (N_27842,N_25209,N_25313);
nand U27843 (N_27843,N_24112,N_25224);
xor U27844 (N_27844,N_25235,N_25835);
nand U27845 (N_27845,N_24480,N_24642);
and U27846 (N_27846,N_24642,N_24921);
and U27847 (N_27847,N_24439,N_24405);
nor U27848 (N_27848,N_24366,N_25273);
and U27849 (N_27849,N_25782,N_24283);
xor U27850 (N_27850,N_24001,N_25830);
or U27851 (N_27851,N_25185,N_24884);
and U27852 (N_27852,N_25765,N_25640);
and U27853 (N_27853,N_24505,N_24293);
and U27854 (N_27854,N_25924,N_24323);
xnor U27855 (N_27855,N_24690,N_25233);
or U27856 (N_27856,N_25098,N_24305);
xnor U27857 (N_27857,N_25235,N_24219);
nor U27858 (N_27858,N_24209,N_25638);
or U27859 (N_27859,N_25375,N_24943);
xor U27860 (N_27860,N_24477,N_24899);
or U27861 (N_27861,N_24936,N_24717);
or U27862 (N_27862,N_25889,N_24196);
and U27863 (N_27863,N_25051,N_25039);
or U27864 (N_27864,N_24523,N_25898);
or U27865 (N_27865,N_25615,N_25459);
or U27866 (N_27866,N_25959,N_25458);
nand U27867 (N_27867,N_24881,N_24156);
xor U27868 (N_27868,N_25113,N_24752);
xnor U27869 (N_27869,N_24344,N_25141);
and U27870 (N_27870,N_24736,N_24682);
or U27871 (N_27871,N_24283,N_25335);
xor U27872 (N_27872,N_25508,N_24978);
nor U27873 (N_27873,N_25642,N_24803);
nor U27874 (N_27874,N_25376,N_24713);
nand U27875 (N_27875,N_25855,N_25980);
nor U27876 (N_27876,N_25728,N_25726);
nor U27877 (N_27877,N_25450,N_25037);
or U27878 (N_27878,N_25217,N_24855);
xnor U27879 (N_27879,N_25712,N_25328);
xnor U27880 (N_27880,N_25750,N_25662);
xnor U27881 (N_27881,N_24086,N_24743);
or U27882 (N_27882,N_25528,N_25273);
xor U27883 (N_27883,N_25105,N_25284);
xor U27884 (N_27884,N_24712,N_24161);
and U27885 (N_27885,N_25339,N_24968);
and U27886 (N_27886,N_24119,N_24821);
and U27887 (N_27887,N_25936,N_25945);
nor U27888 (N_27888,N_25196,N_24639);
nor U27889 (N_27889,N_25228,N_24552);
nor U27890 (N_27890,N_25314,N_24634);
xnor U27891 (N_27891,N_24301,N_25868);
nor U27892 (N_27892,N_24159,N_25815);
nor U27893 (N_27893,N_25896,N_25700);
nand U27894 (N_27894,N_24777,N_25009);
nand U27895 (N_27895,N_24304,N_25203);
xor U27896 (N_27896,N_25928,N_24429);
or U27897 (N_27897,N_24241,N_25349);
xnor U27898 (N_27898,N_24281,N_24901);
xor U27899 (N_27899,N_25676,N_24550);
nor U27900 (N_27900,N_25526,N_24577);
nor U27901 (N_27901,N_25691,N_25323);
nor U27902 (N_27902,N_25295,N_24242);
nor U27903 (N_27903,N_24596,N_24286);
xnor U27904 (N_27904,N_25323,N_25654);
or U27905 (N_27905,N_25166,N_24044);
nor U27906 (N_27906,N_24337,N_25888);
and U27907 (N_27907,N_24866,N_25010);
or U27908 (N_27908,N_24131,N_25181);
xor U27909 (N_27909,N_25030,N_24749);
xor U27910 (N_27910,N_24711,N_25688);
nand U27911 (N_27911,N_24396,N_25728);
nor U27912 (N_27912,N_25191,N_25483);
or U27913 (N_27913,N_24563,N_25657);
nand U27914 (N_27914,N_25044,N_24072);
nor U27915 (N_27915,N_25516,N_25644);
or U27916 (N_27916,N_24201,N_25208);
and U27917 (N_27917,N_25696,N_24622);
xnor U27918 (N_27918,N_24205,N_24877);
nand U27919 (N_27919,N_24297,N_24505);
nor U27920 (N_27920,N_25620,N_24879);
nor U27921 (N_27921,N_25177,N_25671);
nand U27922 (N_27922,N_24192,N_24299);
xor U27923 (N_27923,N_25165,N_25068);
or U27924 (N_27924,N_25547,N_24880);
and U27925 (N_27925,N_25417,N_24462);
xnor U27926 (N_27926,N_25039,N_24147);
xor U27927 (N_27927,N_24477,N_24437);
and U27928 (N_27928,N_24810,N_25291);
or U27929 (N_27929,N_25636,N_25084);
or U27930 (N_27930,N_25467,N_24261);
or U27931 (N_27931,N_24255,N_24457);
xor U27932 (N_27932,N_25450,N_24947);
xor U27933 (N_27933,N_24315,N_25306);
xnor U27934 (N_27934,N_24580,N_25331);
xnor U27935 (N_27935,N_25699,N_25283);
xnor U27936 (N_27936,N_25862,N_24333);
nand U27937 (N_27937,N_24396,N_24606);
nand U27938 (N_27938,N_25918,N_24800);
xor U27939 (N_27939,N_25906,N_25789);
nand U27940 (N_27940,N_24984,N_25677);
or U27941 (N_27941,N_24038,N_24610);
nand U27942 (N_27942,N_24485,N_24298);
and U27943 (N_27943,N_25982,N_25490);
xor U27944 (N_27944,N_25433,N_24585);
nand U27945 (N_27945,N_25025,N_25824);
and U27946 (N_27946,N_25722,N_25879);
nor U27947 (N_27947,N_25724,N_24811);
and U27948 (N_27948,N_24124,N_25771);
nor U27949 (N_27949,N_25318,N_25622);
or U27950 (N_27950,N_24121,N_25872);
nor U27951 (N_27951,N_24822,N_24536);
xnor U27952 (N_27952,N_25835,N_25545);
nor U27953 (N_27953,N_25645,N_24234);
and U27954 (N_27954,N_24040,N_25302);
or U27955 (N_27955,N_24068,N_25290);
nand U27956 (N_27956,N_25070,N_25550);
and U27957 (N_27957,N_24395,N_25462);
or U27958 (N_27958,N_25070,N_25094);
nor U27959 (N_27959,N_24354,N_24372);
and U27960 (N_27960,N_24320,N_24135);
xor U27961 (N_27961,N_25021,N_25857);
and U27962 (N_27962,N_24295,N_25862);
nand U27963 (N_27963,N_24285,N_24959);
xor U27964 (N_27964,N_25712,N_25726);
and U27965 (N_27965,N_25704,N_25329);
nand U27966 (N_27966,N_24691,N_25443);
or U27967 (N_27967,N_24119,N_24142);
or U27968 (N_27968,N_24856,N_25956);
nand U27969 (N_27969,N_25162,N_25147);
or U27970 (N_27970,N_25530,N_25742);
and U27971 (N_27971,N_25527,N_24686);
xnor U27972 (N_27972,N_25207,N_24145);
nor U27973 (N_27973,N_24486,N_24037);
nand U27974 (N_27974,N_24169,N_24233);
or U27975 (N_27975,N_25720,N_25940);
or U27976 (N_27976,N_24821,N_25634);
and U27977 (N_27977,N_25147,N_24282);
or U27978 (N_27978,N_25432,N_24518);
and U27979 (N_27979,N_24444,N_25462);
and U27980 (N_27980,N_25219,N_24941);
nor U27981 (N_27981,N_25939,N_24616);
nand U27982 (N_27982,N_25861,N_25877);
nand U27983 (N_27983,N_25157,N_25926);
nor U27984 (N_27984,N_24833,N_24594);
xnor U27985 (N_27985,N_24959,N_24227);
nor U27986 (N_27986,N_25360,N_25820);
nand U27987 (N_27987,N_25330,N_25158);
or U27988 (N_27988,N_25706,N_24746);
and U27989 (N_27989,N_25847,N_24550);
nor U27990 (N_27990,N_24907,N_25372);
nor U27991 (N_27991,N_25303,N_25753);
or U27992 (N_27992,N_24899,N_24317);
nor U27993 (N_27993,N_24322,N_25357);
nand U27994 (N_27994,N_24160,N_24964);
xnor U27995 (N_27995,N_25632,N_25049);
xor U27996 (N_27996,N_24700,N_24057);
xnor U27997 (N_27997,N_24461,N_25885);
or U27998 (N_27998,N_24332,N_24555);
and U27999 (N_27999,N_25065,N_24856);
nor U28000 (N_28000,N_27928,N_26472);
and U28001 (N_28001,N_27376,N_27372);
and U28002 (N_28002,N_26536,N_27132);
and U28003 (N_28003,N_27649,N_26962);
and U28004 (N_28004,N_26293,N_26414);
and U28005 (N_28005,N_26532,N_26453);
nor U28006 (N_28006,N_26007,N_27872);
and U28007 (N_28007,N_27306,N_26564);
xnor U28008 (N_28008,N_27121,N_26243);
and U28009 (N_28009,N_26753,N_26552);
nand U28010 (N_28010,N_26385,N_26626);
xor U28011 (N_28011,N_26729,N_26415);
nor U28012 (N_28012,N_27340,N_26482);
nand U28013 (N_28013,N_26726,N_26767);
nand U28014 (N_28014,N_26766,N_27887);
xnor U28015 (N_28015,N_27434,N_27144);
and U28016 (N_28016,N_26438,N_27539);
and U28017 (N_28017,N_26092,N_26187);
nand U28018 (N_28018,N_27295,N_27840);
xnor U28019 (N_28019,N_26327,N_27135);
and U28020 (N_28020,N_27666,N_27159);
or U28021 (N_28021,N_26815,N_27604);
nand U28022 (N_28022,N_26288,N_26833);
or U28023 (N_28023,N_27522,N_27425);
nand U28024 (N_28024,N_26731,N_27027);
or U28025 (N_28025,N_27039,N_26356);
xnor U28026 (N_28026,N_26556,N_27967);
or U28027 (N_28027,N_26198,N_26518);
or U28028 (N_28028,N_27163,N_27496);
and U28029 (N_28029,N_27217,N_27919);
or U28030 (N_28030,N_26247,N_26654);
and U28031 (N_28031,N_27782,N_26432);
xnor U28032 (N_28032,N_27056,N_26419);
xnor U28033 (N_28033,N_27102,N_27728);
nand U28034 (N_28034,N_26993,N_27941);
nand U28035 (N_28035,N_27269,N_27738);
nor U28036 (N_28036,N_26969,N_27538);
nor U28037 (N_28037,N_27865,N_26717);
nand U28038 (N_28038,N_27399,N_27473);
xor U28039 (N_28039,N_27282,N_26190);
nor U28040 (N_28040,N_26167,N_26232);
nand U28041 (N_28041,N_27467,N_26876);
and U28042 (N_28042,N_26894,N_27799);
xnor U28043 (N_28043,N_26304,N_27335);
or U28044 (N_28044,N_26347,N_26990);
xnor U28045 (N_28045,N_27612,N_27488);
and U28046 (N_28046,N_26903,N_26761);
nor U28047 (N_28047,N_27515,N_26511);
or U28048 (N_28048,N_26807,N_26269);
nor U28049 (N_28049,N_26774,N_26113);
or U28050 (N_28050,N_27325,N_27686);
and U28051 (N_28051,N_27386,N_26632);
xor U28052 (N_28052,N_27327,N_27851);
nor U28053 (N_28053,N_27007,N_27747);
nand U28054 (N_28054,N_27146,N_27590);
xnor U28055 (N_28055,N_27155,N_26508);
xnor U28056 (N_28056,N_27857,N_26720);
nand U28057 (N_28057,N_26939,N_26219);
xor U28058 (N_28058,N_27959,N_27258);
and U28059 (N_28059,N_26223,N_26871);
nand U28060 (N_28060,N_26644,N_26144);
and U28061 (N_28061,N_26466,N_26320);
xnor U28062 (N_28062,N_27614,N_26989);
or U28063 (N_28063,N_27430,N_26062);
nor U28064 (N_28064,N_26249,N_26209);
xor U28065 (N_28065,N_27384,N_26823);
and U28066 (N_28066,N_27603,N_26836);
xnor U28067 (N_28067,N_27196,N_27804);
nor U28068 (N_28068,N_26631,N_27833);
and U28069 (N_28069,N_27767,N_27518);
nor U28070 (N_28070,N_27288,N_27822);
and U28071 (N_28071,N_27364,N_26839);
or U28072 (N_28072,N_26349,N_26562);
or U28073 (N_28073,N_26695,N_27234);
or U28074 (N_28074,N_27047,N_27647);
nand U28075 (N_28075,N_26315,N_27230);
nand U28076 (N_28076,N_26303,N_27110);
xor U28077 (N_28077,N_27668,N_26423);
and U28078 (N_28078,N_27117,N_27086);
nor U28079 (N_28079,N_26147,N_26373);
nand U28080 (N_28080,N_27888,N_27012);
xnor U28081 (N_28081,N_26862,N_26737);
xnor U28082 (N_28082,N_26809,N_26977);
or U28083 (N_28083,N_27639,N_27861);
and U28084 (N_28084,N_27057,N_26835);
or U28085 (N_28085,N_27030,N_26362);
nor U28086 (N_28086,N_27014,N_27648);
and U28087 (N_28087,N_27800,N_26285);
nor U28088 (N_28088,N_26039,N_26974);
nor U28089 (N_28089,N_26897,N_27720);
nor U28090 (N_28090,N_26802,N_26459);
and U28091 (N_28091,N_26012,N_27633);
xor U28092 (N_28092,N_26988,N_27321);
nand U28093 (N_28093,N_26979,N_27077);
nor U28094 (N_28094,N_26781,N_27341);
nor U28095 (N_28095,N_27354,N_27083);
nor U28096 (N_28096,N_27691,N_27237);
nor U28097 (N_28097,N_27654,N_27715);
and U28098 (N_28098,N_26533,N_26300);
nand U28099 (N_28099,N_26771,N_26843);
xor U28100 (N_28100,N_26528,N_26923);
or U28101 (N_28101,N_26890,N_27271);
and U28102 (N_28102,N_27254,N_26845);
nor U28103 (N_28103,N_26127,N_26649);
and U28104 (N_28104,N_26791,N_26263);
xnor U28105 (N_28105,N_27710,N_27024);
nand U28106 (N_28106,N_26439,N_27148);
and U28107 (N_28107,N_27827,N_27712);
nand U28108 (N_28108,N_27420,N_26653);
xnor U28109 (N_28109,N_27999,N_26768);
or U28110 (N_28110,N_27264,N_27820);
nand U28111 (N_28111,N_27165,N_26081);
xor U28112 (N_28112,N_27629,N_27131);
nand U28113 (N_28113,N_27609,N_26713);
and U28114 (N_28114,N_27916,N_26358);
and U28115 (N_28115,N_26055,N_27022);
nor U28116 (N_28116,N_27737,N_26255);
and U28117 (N_28117,N_27694,N_26191);
and U28118 (N_28118,N_26765,N_27089);
nor U28119 (N_28119,N_26465,N_27255);
and U28120 (N_28120,N_26471,N_26230);
or U28121 (N_28121,N_27331,N_26623);
or U28122 (N_28122,N_26647,N_27699);
and U28123 (N_28123,N_26452,N_26732);
or U28124 (N_28124,N_26367,N_26563);
or U28125 (N_28125,N_26123,N_27808);
xnor U28126 (N_28126,N_27545,N_27523);
xnor U28127 (N_28127,N_26309,N_27220);
and U28128 (N_28128,N_26978,N_27746);
nor U28129 (N_28129,N_27315,N_26294);
xnor U28130 (N_28130,N_27350,N_27279);
or U28131 (N_28131,N_27757,N_26793);
and U28132 (N_28132,N_27011,N_27204);
or U28133 (N_28133,N_26832,N_26698);
xnor U28134 (N_28134,N_27894,N_27546);
or U28135 (N_28135,N_26428,N_26042);
and U28136 (N_28136,N_26566,N_27695);
xor U28137 (N_28137,N_26266,N_27787);
and U28138 (N_28138,N_26301,N_26079);
xnor U28139 (N_28139,N_27931,N_27792);
and U28140 (N_28140,N_27042,N_27316);
nor U28141 (N_28141,N_26818,N_26207);
nor U28142 (N_28142,N_27816,N_27197);
xnor U28143 (N_28143,N_27797,N_26135);
xnor U28144 (N_28144,N_26884,N_26084);
or U28145 (N_28145,N_26467,N_26149);
nand U28146 (N_28146,N_27650,N_26142);
xor U28147 (N_28147,N_26331,N_26251);
and U28148 (N_28148,N_26120,N_27671);
nor U28149 (N_28149,N_26016,N_27417);
nand U28150 (N_28150,N_26455,N_27624);
xor U28151 (N_28151,N_27988,N_27125);
nor U28152 (N_28152,N_27407,N_26277);
nor U28153 (N_28153,N_26248,N_27088);
nor U28154 (N_28154,N_27943,N_26049);
xnor U28155 (N_28155,N_26920,N_27652);
nand U28156 (N_28156,N_27319,N_26093);
or U28157 (N_28157,N_26329,N_27864);
nand U28158 (N_28158,N_27158,N_26476);
xnor U28159 (N_28159,N_27909,N_27463);
nand U28160 (N_28160,N_26867,N_26985);
or U28161 (N_28161,N_26950,N_26316);
nand U28162 (N_28162,N_26214,N_26284);
xor U28163 (N_28163,N_26239,N_27265);
or U28164 (N_28164,N_27889,N_27616);
xor U28165 (N_28165,N_27216,N_26136);
nand U28166 (N_28166,N_27006,N_27210);
xnor U28167 (N_28167,N_27578,N_26422);
or U28168 (N_28168,N_26728,N_27584);
and U28169 (N_28169,N_26549,N_27048);
xnor U28170 (N_28170,N_27651,N_26368);
nand U28171 (N_28171,N_27074,N_27709);
nand U28172 (N_28172,N_27514,N_27934);
xnor U28173 (N_28173,N_26175,N_27563);
nand U28174 (N_28174,N_27577,N_27149);
nor U28175 (N_28175,N_27683,N_27305);
or U28176 (N_28176,N_26256,N_26109);
nand U28177 (N_28177,N_26224,N_27190);
or U28178 (N_28178,N_26283,N_27203);
xor U28179 (N_28179,N_27361,N_26067);
xnor U28180 (N_28180,N_26445,N_26364);
nand U28181 (N_28181,N_26146,N_26576);
nand U28182 (N_28182,N_27280,N_27854);
or U28183 (N_28183,N_26588,N_26208);
nand U28184 (N_28184,N_27530,N_26645);
xor U28185 (N_28185,N_26252,N_27682);
nand U28186 (N_28186,N_27882,N_26826);
or U28187 (N_28187,N_26892,N_27443);
nand U28188 (N_28188,N_26003,N_27892);
and U28189 (N_28189,N_26757,N_27947);
xnor U28190 (N_28190,N_26506,N_26790);
nand U28191 (N_28191,N_26651,N_27107);
and U28192 (N_28192,N_27266,N_26752);
or U28193 (N_28193,N_27094,N_27842);
xnor U28194 (N_28194,N_26088,N_26593);
nand U28195 (N_28195,N_26051,N_27103);
or U28196 (N_28196,N_26888,N_27978);
and U28197 (N_28197,N_26226,N_27655);
or U28198 (N_28198,N_27270,N_27586);
nand U28199 (N_28199,N_26366,N_27613);
and U28200 (N_28200,N_26121,N_27638);
nor U28201 (N_28201,N_27867,N_27708);
nor U28202 (N_28202,N_26868,N_26719);
nor U28203 (N_28203,N_26942,N_27997);
nor U28204 (N_28204,N_26590,N_27465);
nand U28205 (N_28205,N_27895,N_26963);
and U28206 (N_28206,N_26274,N_26205);
or U28207 (N_28207,N_26332,N_27344);
xnor U28208 (N_28208,N_26179,N_26275);
nor U28209 (N_28209,N_27802,N_27940);
nand U28210 (N_28210,N_26748,N_27232);
nor U28211 (N_28211,N_27885,N_26860);
nand U28212 (N_28212,N_27936,N_26642);
nand U28213 (N_28213,N_27451,N_26875);
or U28214 (N_28214,N_27278,N_27949);
nor U28215 (N_28215,N_27557,N_27010);
nor U28216 (N_28216,N_26699,N_26685);
xor U28217 (N_28217,N_27918,N_26795);
or U28218 (N_28218,N_27560,N_27595);
nor U28219 (N_28219,N_26509,N_26499);
nand U28220 (N_28220,N_27718,N_26440);
nand U28221 (N_28221,N_26609,N_26397);
xnor U28222 (N_28222,N_26027,N_27018);
or U28223 (N_28223,N_27771,N_27662);
xnor U28224 (N_28224,N_27847,N_26420);
and U28225 (N_28225,N_27390,N_26424);
nor U28226 (N_28226,N_26053,N_26236);
nor U28227 (N_28227,N_27985,N_26805);
xor U28228 (N_28228,N_26709,N_26145);
nor U28229 (N_28229,N_27445,N_27559);
or U28230 (N_28230,N_26036,N_26234);
nor U28231 (N_28231,N_27824,N_26987);
and U28232 (N_28232,N_27848,N_27664);
nand U28233 (N_28233,N_27766,N_26238);
xor U28234 (N_28234,N_26694,N_26891);
xnor U28235 (N_28235,N_27303,N_26572);
nor U28236 (N_28236,N_27098,N_26662);
nor U28237 (N_28237,N_27636,N_27252);
nor U28238 (N_28238,N_26910,N_26899);
or U28239 (N_28239,N_27469,N_26296);
nand U28240 (N_28240,N_26046,N_27312);
nand U28241 (N_28241,N_27310,N_26106);
nand U28242 (N_28242,N_27675,N_27274);
and U28243 (N_28243,N_27801,N_26825);
or U28244 (N_28244,N_27625,N_27485);
xor U28245 (N_28245,N_26522,N_26025);
or U28246 (N_28246,N_27968,N_27363);
and U28247 (N_28247,N_27351,N_27471);
xnor U28248 (N_28248,N_27605,N_26137);
and U28249 (N_28249,N_26591,N_26189);
and U28250 (N_28250,N_27914,N_27273);
nand U28251 (N_28251,N_27480,N_26480);
xor U28252 (N_28252,N_27549,N_26448);
nand U28253 (N_28253,N_27301,N_26587);
nor U28254 (N_28254,N_26885,N_26715);
and U28255 (N_28255,N_26225,N_27871);
or U28256 (N_28256,N_26363,N_27769);
or U28257 (N_28257,N_26927,N_26583);
and U28258 (N_28258,N_26340,N_27353);
xnor U28259 (N_28259,N_27732,N_26161);
or U28260 (N_28260,N_26534,N_26141);
or U28261 (N_28261,N_27989,N_26325);
xor U28262 (N_28262,N_26352,N_26282);
nand U28263 (N_28263,N_27685,N_26170);
nor U28264 (N_28264,N_26108,N_26741);
and U28265 (N_28265,N_26028,N_27017);
nand U28266 (N_28266,N_27836,N_26210);
xnor U28267 (N_28267,N_26035,N_26160);
nand U28268 (N_28268,N_27565,N_26917);
nor U28269 (N_28269,N_26928,N_26126);
xor U28270 (N_28270,N_27855,N_27926);
and U28271 (N_28271,N_26751,N_26391);
nand U28272 (N_28272,N_27277,N_27287);
nand U28273 (N_28273,N_27778,N_27572);
or U28274 (N_28274,N_26289,N_26722);
nor U28275 (N_28275,N_26607,N_26643);
nor U28276 (N_28276,N_27902,N_26688);
nand U28277 (N_28277,N_26743,N_26931);
nor U28278 (N_28278,N_26272,N_26613);
and U28279 (N_28279,N_26031,N_26865);
and U28280 (N_28280,N_26543,N_26267);
nor U28281 (N_28281,N_26044,N_27908);
and U28282 (N_28282,N_27019,N_26847);
xor U28283 (N_28283,N_27320,N_27189);
nor U28284 (N_28284,N_27368,N_26402);
nand U28285 (N_28285,N_26733,N_26026);
or U28286 (N_28286,N_27140,N_26919);
and U28287 (N_28287,N_27078,N_27065);
and U28288 (N_28288,N_27100,N_26540);
or U28289 (N_28289,N_27725,N_26914);
and U28290 (N_28290,N_27543,N_27831);
nor U28291 (N_28291,N_26004,N_27495);
nand U28292 (N_28292,N_26091,N_27717);
xnor U28293 (N_28293,N_26640,N_27410);
and U28294 (N_28294,N_26032,N_26602);
xor U28295 (N_28295,N_27907,N_26228);
xnor U28296 (N_28296,N_26853,N_27974);
and U28297 (N_28297,N_26433,N_27568);
nor U28298 (N_28298,N_27193,N_27023);
xor U28299 (N_28299,N_26842,N_26451);
or U28300 (N_28300,N_26171,N_27099);
or U28301 (N_28301,N_27194,N_27677);
nand U28302 (N_28302,N_26006,N_27116);
nand U28303 (N_28303,N_26568,N_26059);
and U28304 (N_28304,N_26872,N_26401);
and U28305 (N_28305,N_27336,N_27676);
nor U28306 (N_28306,N_27169,N_27681);
xnor U28307 (N_28307,N_27382,N_26665);
xor U28308 (N_28308,N_26066,N_27329);
xor U28309 (N_28309,N_27900,N_27211);
or U28310 (N_28310,N_27109,N_26199);
and U28311 (N_28311,N_27823,N_27615);
xor U28312 (N_28312,N_26498,N_26041);
xnor U28313 (N_28313,N_26670,N_27793);
xor U28314 (N_28314,N_27753,N_27069);
nor U28315 (N_28315,N_27185,N_26182);
or U28316 (N_28316,N_27423,N_26324);
nor U28317 (N_28317,N_26131,N_26828);
xnor U28318 (N_28318,N_27233,N_26279);
xor U28319 (N_28319,N_26361,N_26378);
xor U28320 (N_28320,N_26298,N_26473);
or U28321 (N_28321,N_27904,N_27242);
and U28322 (N_28322,N_26905,N_27704);
or U28323 (N_28323,N_26968,N_27569);
or U28324 (N_28324,N_27637,N_27644);
nand U28325 (N_28325,N_27810,N_26174);
xnor U28326 (N_28326,N_27528,N_26045);
and U28327 (N_28327,N_26411,N_27945);
or U28328 (N_28328,N_26151,N_27226);
nor U28329 (N_28329,N_26077,N_27172);
or U28330 (N_28330,N_26959,N_26409);
nand U28331 (N_28331,N_27478,N_27874);
and U28332 (N_28332,N_27318,N_26218);
nand U28333 (N_28333,N_26430,N_27182);
and U28334 (N_28334,N_27930,N_26980);
xor U28335 (N_28335,N_26779,N_26525);
and U28336 (N_28336,N_27180,N_27656);
xor U28337 (N_28337,N_27995,N_26904);
and U28338 (N_28338,N_27617,N_27208);
and U28339 (N_28339,N_27119,N_27716);
and U28340 (N_28340,N_27292,N_26738);
or U28341 (N_28341,N_27244,N_27071);
or U28342 (N_28342,N_26196,N_27079);
or U28343 (N_28343,N_27259,N_27005);
nand U28344 (N_28344,N_27238,N_26297);
nor U28345 (N_28345,N_26951,N_27996);
nor U28346 (N_28346,N_27418,N_27573);
or U28347 (N_28347,N_27939,N_27142);
xor U28348 (N_28348,N_26948,N_27973);
nand U28349 (N_28349,N_26050,N_27504);
and U28350 (N_28350,N_26165,N_26947);
or U28351 (N_28351,N_27630,N_27106);
nor U28352 (N_28352,N_27267,N_27598);
xor U28353 (N_28353,N_27791,N_27224);
or U28354 (N_28354,N_26785,N_27524);
and U28355 (N_28355,N_26821,N_27727);
or U28356 (N_28356,N_27670,N_26610);
or U28357 (N_28357,N_27911,N_26940);
nor U28358 (N_28358,N_26803,N_26633);
or U28359 (N_28359,N_27365,N_27853);
nand U28360 (N_28360,N_27108,N_27439);
or U28361 (N_28361,N_27051,N_27923);
and U28362 (N_28362,N_27665,N_27096);
and U28363 (N_28363,N_26128,N_26355);
and U28364 (N_28364,N_26786,N_26787);
and U28365 (N_28365,N_27219,N_26577);
nor U28366 (N_28366,N_26107,N_26510);
or U28367 (N_28367,N_27124,N_26820);
nand U28368 (N_28368,N_26343,N_27186);
nand U28369 (N_28369,N_27877,N_27490);
nor U28370 (N_28370,N_27333,N_27561);
nand U28371 (N_28371,N_26110,N_27356);
xor U28372 (N_28372,N_27123,N_27324);
and U28373 (N_28373,N_26656,N_26002);
or U28374 (N_28374,N_26080,N_27582);
nand U28375 (N_28375,N_27849,N_26663);
and U28376 (N_28376,N_26964,N_27173);
nand U28377 (N_28377,N_27520,N_26176);
xnor U28378 (N_28378,N_27370,N_27832);
or U28379 (N_28379,N_27910,N_26130);
nand U28380 (N_28380,N_27735,N_26851);
nor U28381 (N_28381,N_26557,N_26242);
nand U28382 (N_28382,N_27783,N_27542);
nand U28383 (N_28383,N_27983,N_26558);
xnor U28384 (N_28384,N_27251,N_26442);
or U28385 (N_28385,N_27209,N_27262);
nor U28386 (N_28386,N_26474,N_26701);
nand U28387 (N_28387,N_26554,N_27608);
or U28388 (N_28388,N_26342,N_26104);
xnor U28389 (N_28389,N_26646,N_26392);
or U28390 (N_28390,N_27673,N_27678);
xnor U28391 (N_28391,N_26599,N_26629);
nor U28392 (N_28392,N_27260,N_27897);
nand U28393 (N_28393,N_27075,N_27454);
nor U28394 (N_28394,N_27253,N_26696);
or U28395 (N_28395,N_27393,N_27837);
or U28396 (N_28396,N_26133,N_26960);
nand U28397 (N_28397,N_27736,N_27400);
or U28398 (N_28398,N_27261,N_27516);
nand U28399 (N_28399,N_26736,N_27620);
nand U28400 (N_28400,N_27097,N_26395);
or U28401 (N_28401,N_26734,N_26086);
nand U28402 (N_28402,N_26015,N_27245);
or U28403 (N_28403,N_27763,N_27631);
nand U28404 (N_28404,N_26621,N_26407);
xor U28405 (N_28405,N_27342,N_27413);
xnor U28406 (N_28406,N_26507,N_27241);
nor U28407 (N_28407,N_26898,N_26553);
nor U28408 (N_28408,N_26068,N_26548);
xor U28409 (N_28409,N_27689,N_26431);
xnor U28410 (N_28410,N_26856,N_27153);
nor U28411 (N_28411,N_27986,N_27713);
nor U28412 (N_28412,N_27366,N_27764);
nor U28413 (N_28413,N_26604,N_27028);
nor U28414 (N_28414,N_27362,N_26838);
nand U28415 (N_28415,N_26981,N_27749);
and U28416 (N_28416,N_27517,N_26611);
xnor U28417 (N_28417,N_26911,N_27811);
nor U28418 (N_28418,N_27070,N_27690);
and U28419 (N_28419,N_26155,N_26813);
and U28420 (N_28420,N_27765,N_27427);
or U28421 (N_28421,N_27601,N_27201);
or U28422 (N_28422,N_26233,N_26620);
xor U28423 (N_28423,N_27272,N_26551);
xnor U28424 (N_28424,N_27484,N_27925);
nand U28425 (N_28425,N_26215,N_27537);
and U28426 (N_28426,N_27049,N_27345);
nand U28427 (N_28427,N_26789,N_27134);
or U28428 (N_28428,N_26530,N_27404);
or U28429 (N_28429,N_27429,N_27164);
or U28430 (N_28430,N_26258,N_27195);
and U28431 (N_28431,N_26417,N_26973);
and U28432 (N_28432,N_26018,N_27391);
and U28433 (N_28433,N_26241,N_26716);
xor U28434 (N_28434,N_27571,N_26357);
nand U28435 (N_28435,N_27268,N_26461);
xor U28436 (N_28436,N_27389,N_27453);
and U28437 (N_28437,N_26866,N_26319);
and U28438 (N_28438,N_27510,N_27760);
nor U28439 (N_28439,N_26405,N_27761);
nand U28440 (N_28440,N_26038,N_26011);
or U28441 (N_28441,N_26264,N_26339);
or U28442 (N_28442,N_26485,N_27038);
nor U28443 (N_28443,N_26099,N_26094);
nand U28444 (N_28444,N_26180,N_27846);
nor U28445 (N_28445,N_27845,N_27576);
xor U28446 (N_28446,N_26481,N_27296);
xnor U28447 (N_28447,N_27055,N_26021);
xnor U28448 (N_28448,N_27029,N_27016);
xnor U28449 (N_28449,N_26090,N_26998);
xor U28450 (N_28450,N_26360,N_26527);
or U28451 (N_28451,N_26961,N_26801);
and U28452 (N_28452,N_26908,N_27772);
nand U28453 (N_28453,N_26310,N_26323);
nand U28454 (N_28454,N_27745,N_27085);
nor U28455 (N_28455,N_26883,N_27206);
nand U28456 (N_28456,N_26639,N_26056);
or U28457 (N_28457,N_26075,N_27472);
nand U28458 (N_28458,N_27981,N_26125);
or U28459 (N_28459,N_27001,N_26203);
nand U28460 (N_28460,N_27293,N_27064);
or U28461 (N_28461,N_27618,N_26195);
xnor U28462 (N_28462,N_26115,N_26796);
or U28463 (N_28463,N_27133,N_26353);
xor U28464 (N_28464,N_27143,N_27235);
and U28465 (N_28465,N_26703,N_27969);
and U28466 (N_28466,N_27550,N_27183);
or U28467 (N_28467,N_26777,N_27036);
nand U28468 (N_28468,N_26725,N_27441);
xnor U28469 (N_28469,N_26560,N_26902);
and U28470 (N_28470,N_27229,N_26354);
xnor U28471 (N_28471,N_26671,N_27700);
or U28472 (N_28472,N_26916,N_26048);
xnor U28473 (N_28473,N_26672,N_26907);
nand U28474 (N_28474,N_27138,N_27147);
nand U28475 (N_28475,N_27416,N_27917);
xnor U28476 (N_28476,N_26386,N_26956);
and U28477 (N_28477,N_27574,N_27076);
xor U28478 (N_28478,N_26618,N_26061);
and U28479 (N_28479,N_27236,N_26584);
and U28480 (N_28480,N_26008,N_26287);
nor U28481 (N_28481,N_26922,N_26389);
nor U28482 (N_28482,N_26307,N_27168);
nor U28483 (N_28483,N_26222,N_27788);
or U28484 (N_28484,N_27157,N_27751);
and U28485 (N_28485,N_26449,N_26398);
and U28486 (N_28486,N_27346,N_27663);
and U28487 (N_28487,N_26877,N_27026);
and U28488 (N_28488,N_27977,N_27432);
or U28489 (N_28489,N_26597,N_26776);
nand U28490 (N_28490,N_27095,N_26889);
nor U28491 (N_28491,N_27156,N_26886);
and U28492 (N_28492,N_26484,N_26814);
or U28493 (N_28493,N_27205,N_27322);
and U28494 (N_28494,N_27726,N_27946);
xor U28495 (N_28495,N_27369,N_27397);
nor U28496 (N_28496,N_27246,N_26478);
xor U28497 (N_28497,N_26570,N_27773);
or U28498 (N_28498,N_26864,N_27120);
and U28499 (N_28499,N_27748,N_26070);
and U28500 (N_28500,N_27723,N_27890);
or U28501 (N_28501,N_27875,N_26259);
nand U28502 (N_28502,N_27314,N_26755);
xnor U28503 (N_28503,N_26906,N_26930);
nand U28504 (N_28504,N_26996,N_26966);
or U28505 (N_28505,N_27289,N_26271);
nand U28506 (N_28506,N_27355,N_26706);
or U28507 (N_28507,N_26116,N_26235);
xnor U28508 (N_28508,N_27062,N_26435);
nand U28509 (N_28509,N_27308,N_27583);
and U28510 (N_28510,N_27435,N_26739);
or U28511 (N_28511,N_27881,N_26487);
or U28512 (N_28512,N_27009,N_26336);
xnor U28513 (N_28513,N_27581,N_26521);
or U28514 (N_28514,N_27175,N_27396);
and U28515 (N_28515,N_27597,N_27971);
and U28516 (N_28516,N_26514,N_27489);
nand U28517 (N_28517,N_27426,N_27858);
xor U28518 (N_28518,N_26901,N_27533);
nor U28519 (N_28519,N_26257,N_26896);
and U28520 (N_28520,N_26335,N_27729);
xnor U28521 (N_28521,N_26488,N_27795);
nand U28522 (N_28522,N_26879,N_27456);
nand U28523 (N_28523,N_26058,N_27461);
nand U28524 (N_28524,N_27058,N_26381);
and U28525 (N_28525,N_27352,N_26773);
nand U28526 (N_28526,N_26437,N_27477);
xnor U28527 (N_28527,N_27114,N_27869);
xnor U28528 (N_28528,N_27419,N_27452);
nor U28529 (N_28529,N_26971,N_26657);
and U28530 (N_28530,N_27927,N_27679);
and U28531 (N_28531,N_26955,N_26163);
and U28532 (N_28532,N_26124,N_27415);
and U28533 (N_28533,N_26069,N_27141);
and U28534 (N_28534,N_26469,N_26772);
and U28535 (N_28535,N_27807,N_26129);
nor U28536 (N_28536,N_27798,N_27247);
or U28537 (N_28537,N_26416,N_26636);
or U28538 (N_28538,N_26747,N_27527);
or U28539 (N_28539,N_27509,N_27311);
nor U28540 (N_28540,N_26150,N_27841);
and U28541 (N_28541,N_27965,N_27081);
and U28542 (N_28542,N_26929,N_27044);
and U28543 (N_28543,N_26496,N_26668);
and U28544 (N_28544,N_27170,N_27992);
nor U28545 (N_28545,N_27750,N_27998);
nor U28546 (N_28546,N_26427,N_26759);
nand U28547 (N_28547,N_27722,N_27313);
or U28548 (N_28548,N_26531,N_26965);
and U28549 (N_28549,N_27377,N_26312);
nand U28550 (N_28550,N_27896,N_26505);
and U28551 (N_28551,N_27066,N_26995);
nor U28552 (N_28552,N_27781,N_27606);
nor U28553 (N_28553,N_26087,N_27460);
and U28554 (N_28554,N_26986,N_26667);
xnor U28555 (N_28555,N_27444,N_27130);
nor U28556 (N_28556,N_26060,N_26596);
nand U28557 (N_28557,N_27588,N_26111);
or U28558 (N_28558,N_26200,N_26660);
and U28559 (N_28559,N_26569,N_27046);
and U28560 (N_28560,N_26375,N_26513);
and U28561 (N_28561,N_26714,N_27623);
nor U28562 (N_28562,N_26921,N_26512);
and U28563 (N_28563,N_27291,N_27915);
nor U28564 (N_28564,N_26278,N_26834);
or U28565 (N_28565,N_26935,N_27499);
nor U28566 (N_28566,N_27768,N_27214);
xor U28567 (N_28567,N_27374,N_26290);
nand U28568 (N_28568,N_27790,N_27486);
nand U28569 (N_28569,N_26425,N_27068);
nand U28570 (N_28570,N_27008,N_27448);
nand U28571 (N_28571,N_27375,N_26302);
or U28572 (N_28572,N_26827,N_26273);
nor U28573 (N_28573,N_26158,N_27503);
nand U28574 (N_28574,N_27944,N_26013);
nand U28575 (N_28575,N_27412,N_26043);
xor U28576 (N_28576,N_27526,N_27405);
nand U28577 (N_28577,N_27043,N_26497);
xnor U28578 (N_28578,N_26192,N_27178);
nor U28579 (N_28579,N_27498,N_26983);
nand U28580 (N_28580,N_27087,N_27385);
xor U28581 (N_28581,N_26140,N_26542);
nand U28582 (N_28582,N_26254,N_27886);
xnor U28583 (N_28583,N_27762,N_27326);
nand U28584 (N_28584,N_27693,N_26806);
and U28585 (N_28585,N_27160,N_27529);
nor U28586 (N_28586,N_27596,N_26348);
nand U28587 (N_28587,N_26486,N_27591);
nor U28588 (N_28588,N_27562,N_27589);
and U28589 (N_28589,N_27658,N_26627);
or U28590 (N_28590,N_27428,N_26139);
xor U28591 (N_28591,N_27541,N_27828);
xnor U28592 (N_28592,N_26792,N_26664);
nor U28593 (N_28593,N_26262,N_27249);
and U28594 (N_28594,N_27139,N_26844);
and U28595 (N_28595,N_27703,N_27786);
xnor U28596 (N_28596,N_27493,N_26040);
or U28597 (N_28597,N_26762,N_27740);
nand U28598 (N_28598,N_26341,N_27883);
xnor U28599 (N_28599,N_26516,N_27421);
or U28600 (N_28600,N_26318,N_26691);
or U28601 (N_28601,N_26870,N_26684);
and U28602 (N_28602,N_26970,N_27015);
nor U28603 (N_28603,N_27187,N_26692);
nand U28604 (N_28604,N_26166,N_27304);
nor U28605 (N_28605,N_27646,N_26313);
or U28606 (N_28606,N_27052,N_27813);
and U28607 (N_28607,N_26280,N_26539);
and U28608 (N_28608,N_26764,N_27830);
nor U28609 (N_28609,N_27343,N_26000);
and U28610 (N_28610,N_26387,N_26064);
nor U28611 (N_28611,N_27334,N_27034);
nor U28612 (N_28612,N_27775,N_27337);
or U28613 (N_28613,N_27806,N_26666);
or U28614 (N_28614,N_27993,N_26260);
nor U28615 (N_28615,N_27218,N_26470);
or U28616 (N_28616,N_26648,N_26157);
and U28617 (N_28617,N_26817,N_26641);
and U28618 (N_28618,N_26537,N_26334);
nand U28619 (N_28619,N_27972,N_26918);
nor U28620 (N_28620,N_26601,N_27330);
nand U28621 (N_28621,N_27789,N_26365);
nand U28622 (N_28622,N_27491,N_26658);
nand U28623 (N_28623,N_27129,N_27136);
or U28624 (N_28624,N_27357,N_27544);
and U28625 (N_28625,N_26850,N_26804);
or U28626 (N_28626,N_27228,N_26612);
or U28627 (N_28627,N_26811,N_27373);
nor U28628 (N_28628,N_26383,N_27843);
nand U28629 (N_28629,N_27092,N_26408);
xnor U28630 (N_28630,N_27627,N_26418);
nand U28631 (N_28631,N_26193,N_27150);
xnor U28632 (N_28632,N_26529,N_26984);
and U28633 (N_28633,N_27739,N_26561);
nor U28634 (N_28634,N_27101,N_26143);
nand U28635 (N_28635,N_26456,N_26295);
xor U28636 (N_28636,N_26581,N_26874);
or U28637 (N_28637,N_27579,N_27755);
and U28638 (N_28638,N_26413,N_26893);
and U28639 (N_28639,N_26848,N_27688);
nor U28640 (N_28640,N_27844,N_26211);
xnor U28641 (N_28641,N_26637,N_26909);
and U28642 (N_28642,N_27730,N_26078);
and U28643 (N_28643,N_26686,N_26750);
nand U28644 (N_28644,N_26954,N_26412);
or U28645 (N_28645,N_27093,N_27701);
nand U28646 (N_28646,N_27387,N_26547);
and U28647 (N_28647,N_27770,N_26005);
xnor U28648 (N_28648,N_27021,N_27411);
xor U28649 (N_28649,N_26746,N_27179);
xor U28650 (N_28650,N_27285,N_26479);
nand U28651 (N_28651,N_26925,N_27803);
nand U28652 (N_28652,N_26204,N_27587);
or U28653 (N_28653,N_27963,N_26550);
or U28654 (N_28654,N_27970,N_27711);
xnor U28655 (N_28655,N_27073,N_27174);
xnor U28656 (N_28656,N_26052,N_26708);
xnor U28657 (N_28657,N_27126,N_26669);
nand U28658 (N_28658,N_26689,N_26852);
xor U28659 (N_28659,N_27906,N_27669);
nand U28660 (N_28660,N_27105,N_27276);
nor U28661 (N_28661,N_27899,N_26994);
or U28662 (N_28662,N_26100,N_26376);
xor U28663 (N_28663,N_26798,N_26047);
nor U28664 (N_28664,N_27721,N_26097);
or U28665 (N_28665,N_27383,N_26134);
and U28666 (N_28666,N_27487,N_26429);
and U28667 (N_28667,N_27990,N_26819);
nor U28668 (N_28668,N_26592,N_27567);
xor U28669 (N_28669,N_27935,N_26841);
xnor U28670 (N_28670,N_26338,N_27225);
xor U28671 (N_28671,N_26101,N_26723);
or U28672 (N_28672,N_26541,N_27815);
or U28673 (N_28673,N_27050,N_26679);
nand U28674 (N_28674,N_27905,N_26390);
nand U28675 (N_28675,N_27961,N_27475);
nor U28676 (N_28676,N_26678,N_27113);
nor U28677 (N_28677,N_26846,N_27634);
and U28678 (N_28678,N_26598,N_26579);
or U28679 (N_28679,N_26468,N_27653);
xor U28680 (N_28680,N_26350,N_27424);
nor U28681 (N_28681,N_26936,N_27812);
or U28682 (N_28682,N_27447,N_27884);
nand U28683 (N_28683,N_27555,N_27002);
and U28684 (N_28684,N_26394,N_27367);
nand U28685 (N_28685,N_27580,N_26159);
nand U28686 (N_28686,N_26212,N_26895);
and U28687 (N_28687,N_27891,N_26718);
nor U28688 (N_28688,N_27481,N_27464);
or U28689 (N_28689,N_27659,N_27446);
and U28690 (N_28690,N_27300,N_26083);
nand U28691 (N_28691,N_26403,N_27433);
nand U28692 (N_28692,N_26837,N_26724);
nand U28693 (N_28693,N_27741,N_27564);
nor U28694 (N_28694,N_26869,N_26756);
nor U28695 (N_28695,N_27394,N_27199);
xnor U28696 (N_28696,N_27222,N_27000);
xor U28697 (N_28697,N_27774,N_27924);
nand U28698 (N_28698,N_26578,N_27176);
nor U28699 (N_28699,N_26638,N_27118);
or U28700 (N_28700,N_27408,N_26710);
xor U28701 (N_28701,N_26778,N_27500);
nand U28702 (N_28702,N_27758,N_27553);
and U28703 (N_28703,N_27692,N_26745);
xnor U28704 (N_28704,N_26754,N_26221);
or U28705 (N_28705,N_26220,N_27298);
nor U28706 (N_28706,N_27198,N_27302);
nor U28707 (N_28707,N_26992,N_26464);
xnor U28708 (N_28708,N_26816,N_27231);
nand U28709 (N_28709,N_27257,N_26103);
xnor U28710 (N_28710,N_26102,N_26926);
nor U28711 (N_28711,N_26913,N_27166);
or U28712 (N_28712,N_27628,N_26369);
and U28713 (N_28713,N_26585,N_26410);
and U28714 (N_28714,N_26881,N_26404);
nor U28715 (N_28715,N_27275,N_26625);
xnor U28716 (N_28716,N_26517,N_26524);
nand U28717 (N_28717,N_26628,N_27863);
and U28718 (N_28718,N_26500,N_26337);
nor U28719 (N_28719,N_26526,N_27809);
or U28720 (N_28720,N_27954,N_27743);
or U28721 (N_28721,N_27779,N_26460);
and U28722 (N_28722,N_27060,N_26010);
xnor U28723 (N_28723,N_27672,N_27756);
xor U28724 (N_28724,N_27570,N_26020);
and U28725 (N_28725,N_26682,N_26831);
xor U28726 (N_28726,N_26675,N_26953);
xnor U28727 (N_28727,N_27921,N_26861);
nand U28728 (N_28728,N_26168,N_27674);
nand U28729 (N_28729,N_27643,N_27744);
and U28730 (N_28730,N_27912,N_26074);
nor U28731 (N_28731,N_26085,N_27548);
nor U28732 (N_28732,N_27388,N_27512);
nor U28733 (N_28733,N_26680,N_27040);
nor U28734 (N_28734,N_26436,N_26321);
and U28735 (N_28735,N_26188,N_26800);
or U28736 (N_28736,N_27839,N_26999);
or U28737 (N_28737,N_26808,N_27640);
nor U28738 (N_28738,N_26197,N_27913);
nand U28739 (N_28739,N_26065,N_26001);
nor U28740 (N_28740,N_26702,N_27955);
nand U28741 (N_28741,N_26565,N_27317);
nand U28742 (N_28742,N_27938,N_27061);
nor U28743 (N_28743,N_27436,N_27457);
xor U28744 (N_28744,N_27521,N_27585);
nor U28745 (N_28745,N_27250,N_26494);
xor U28746 (N_28746,N_27212,N_27003);
or U28747 (N_28747,N_26573,N_26555);
or U28748 (N_28748,N_27348,N_26712);
nand U28749 (N_28749,N_27920,N_27979);
xnor U28750 (N_28750,N_26421,N_26545);
or U28751 (N_28751,N_27984,N_26306);
or U28752 (N_28752,N_27513,N_27115);
nor U28753 (N_28753,N_27035,N_26721);
and U28754 (N_28754,N_26119,N_26326);
nor U28755 (N_28755,N_26089,N_26024);
nor U28756 (N_28756,N_26788,N_27450);
and U28757 (N_28757,N_26270,N_27080);
xnor U28758 (N_28758,N_27657,N_27184);
or U28759 (N_28759,N_26617,N_27536);
and U28760 (N_28760,N_27975,N_26949);
and U28761 (N_28761,N_26674,N_26346);
xor U28762 (N_28762,N_27850,N_26393);
xor U28763 (N_28763,N_27987,N_27223);
or U28764 (N_28764,N_26616,N_26172);
and U28765 (N_28765,N_26444,N_27494);
nor U28766 (N_28766,N_26595,N_27734);
nand U28767 (N_28767,N_27128,N_27950);
xnor U28768 (N_28768,N_27826,N_26181);
nand U28769 (N_28769,N_26661,N_27328);
or U28770 (N_28770,N_26794,N_27339);
or U28771 (N_28771,N_26372,N_27084);
and U28772 (N_28772,N_27667,N_27380);
nor U28773 (N_28773,N_26380,N_26034);
or U28774 (N_28774,N_26177,N_26345);
xnor U28775 (N_28775,N_26855,N_27215);
and U28776 (N_28776,N_26250,N_26882);
nand U28777 (N_28777,N_26824,N_27256);
or U28778 (N_28778,N_27566,N_26690);
nand U28779 (N_28779,N_26344,N_27414);
xor U28780 (N_28780,N_27592,N_27594);
nand U28781 (N_28781,N_27025,N_26328);
nor U28782 (N_28782,N_26033,N_26122);
xor U28783 (N_28783,N_27880,N_27552);
nor U28784 (N_28784,N_26237,N_27535);
and U28785 (N_28785,N_26700,N_27004);
and U28786 (N_28786,N_26253,N_27856);
nand U28787 (N_28787,N_27359,N_27202);
nor U28788 (N_28788,N_27299,N_26887);
nand U28789 (N_28789,N_26740,N_27054);
nor U28790 (N_28790,N_27777,N_27281);
nor U28791 (N_28791,N_27661,N_26268);
nor U28792 (N_28792,N_27879,N_27401);
nor U28793 (N_28793,N_27714,N_26178);
nor U28794 (N_28794,N_27167,N_27171);
xor U28795 (N_28795,N_26265,N_27937);
nor U28796 (N_28796,N_27829,N_27962);
and U28797 (N_28797,N_26676,N_26519);
nand U28798 (N_28798,N_26216,N_27593);
and U28799 (N_28799,N_27776,N_26933);
nand U28800 (N_28800,N_26707,N_27151);
xor U28801 (N_28801,N_26492,N_27459);
or U28802 (N_28802,N_27680,N_27466);
xor U28803 (N_28803,N_26359,N_26017);
or U28804 (N_28804,N_27622,N_26932);
or U28805 (N_28805,N_27531,N_26742);
or U28806 (N_28806,N_27707,N_26105);
xnor U28807 (N_28807,N_27759,N_26314);
and U28808 (N_28808,N_27632,N_26370);
nand U28809 (N_28809,N_26374,N_26677);
and U28810 (N_28810,N_26305,N_26063);
and U28811 (N_28811,N_26744,N_26504);
nor U28812 (N_28812,N_26014,N_27705);
nand U28813 (N_28813,N_27127,N_27878);
xor U28814 (N_28814,N_26477,N_27817);
and U28815 (N_28815,N_27525,N_27742);
nand U28816 (N_28816,N_27860,N_26673);
or U28817 (N_28817,N_27645,N_26784);
nand U28818 (N_28818,N_27162,N_27893);
or U28819 (N_28819,N_26538,N_26575);
and U28820 (N_28820,N_27440,N_27403);
xnor U28821 (N_28821,N_26799,N_27032);
and U28822 (N_28822,N_27072,N_26544);
xor U28823 (N_28823,N_27619,N_27398);
or U28824 (N_28824,N_27090,N_26281);
xor U28825 (N_28825,N_26946,N_26333);
or U28826 (N_28826,N_27953,N_27122);
xor U28827 (N_28827,N_26217,N_26501);
and U28828 (N_28828,N_26023,N_26493);
and U28829 (N_28829,N_26458,N_27284);
nand U28830 (N_28830,N_27952,N_26148);
xor U28831 (N_28831,N_27754,N_27455);
and U28832 (N_28832,N_27177,N_27497);
or U28833 (N_28833,N_27371,N_27731);
xor U28834 (N_28834,N_26857,N_27479);
xnor U28835 (N_28835,N_27033,N_27449);
nor U28836 (N_28836,N_27283,N_27506);
and U28837 (N_28837,N_26600,N_27870);
or U28838 (N_28838,N_26118,N_27474);
or U28839 (N_28839,N_27462,N_26261);
nor U28840 (N_28840,N_26938,N_27642);
nor U28841 (N_28841,N_26944,N_27626);
or U28842 (N_28842,N_26924,N_26152);
xor U28843 (N_28843,N_27360,N_27903);
and U28844 (N_28844,N_26117,N_27957);
or U28845 (N_28845,N_26880,N_27794);
nor U28846 (N_28846,N_26606,N_26830);
nor U28847 (N_28847,N_26164,N_27966);
or U28848 (N_28848,N_27192,N_27145);
nand U28849 (N_28849,N_27994,N_26878);
nand U28850 (N_28850,N_26515,N_26317);
nor U28851 (N_28851,N_26571,N_26912);
nand U28852 (N_28852,N_26206,N_26483);
or U28853 (N_28853,N_26608,N_26169);
or U28854 (N_28854,N_26687,N_27991);
nand U28855 (N_28855,N_27602,N_26245);
xnor U28856 (N_28856,N_27821,N_27191);
or U28857 (N_28857,N_26630,N_26434);
or U28858 (N_28858,N_26943,N_26727);
nand U28859 (N_28859,N_26291,N_26184);
xor U28860 (N_28860,N_27635,N_27901);
xnor U28861 (N_28861,N_26286,N_26783);
nand U28862 (N_28862,N_26900,N_26489);
or U28863 (N_28863,N_27951,N_27519);
or U28864 (N_28864,N_27381,N_26782);
or U28865 (N_28865,N_26201,N_27422);
nor U28866 (N_28866,N_27702,N_27112);
or U28867 (N_28867,N_26443,N_27053);
xnor U28868 (N_28868,N_27933,N_27248);
nand U28869 (N_28869,N_27227,N_27263);
nand U28870 (N_28870,N_27200,N_26659);
xnor U28871 (N_28871,N_27876,N_26967);
xor U28872 (N_28872,N_26730,N_26603);
or U28873 (N_28873,N_26490,N_26112);
nor U28874 (N_28874,N_26574,N_26246);
xor U28875 (N_28875,N_26634,N_27600);
nor U28876 (N_28876,N_26941,N_26829);
and U28877 (N_28877,N_26406,N_27825);
and U28878 (N_28878,N_27575,N_26057);
nor U28879 (N_28879,N_26711,N_26863);
nand U28880 (N_28880,N_27378,N_26096);
xor U28881 (N_28881,N_26240,N_27805);
and U28882 (N_28882,N_26934,N_26559);
nand U28883 (N_28883,N_26019,N_27508);
xnor U28884 (N_28884,N_26454,N_27045);
xor U28885 (N_28885,N_27402,N_27780);
or U28886 (N_28886,N_27243,N_26582);
or U28887 (N_28887,N_26945,N_26185);
xnor U28888 (N_28888,N_26071,N_26311);
nor U28889 (N_28889,N_26379,N_27980);
nor U28890 (N_28890,N_26854,N_27610);
or U28891 (N_28891,N_26635,N_26503);
nand U28892 (N_28892,N_27964,N_26213);
and U28893 (N_28893,N_27752,N_27501);
and U28894 (N_28894,N_26073,N_27297);
nor U28895 (N_28895,N_26972,N_27482);
or U28896 (N_28896,N_27838,N_27492);
xnor U28897 (N_28897,N_27307,N_26351);
nand U28898 (N_28898,N_26162,N_26735);
or U28899 (N_28899,N_26991,N_27431);
or U28900 (N_28900,N_27834,N_26450);
xor U28901 (N_28901,N_27082,N_27976);
and U28902 (N_28902,N_27358,N_26655);
xor U28903 (N_28903,N_26399,N_26330);
xnor U28904 (N_28904,N_27239,N_27922);
xnor U28905 (N_28905,N_26153,N_27031);
nand U28906 (N_28906,N_26957,N_27719);
nand U28907 (N_28907,N_26054,N_27558);
and U28908 (N_28908,N_27013,N_27458);
or U28909 (N_28909,N_26447,N_27091);
or U28910 (N_28910,N_27733,N_27309);
xnor U28911 (N_28911,N_27599,N_26589);
xor U28912 (N_28912,N_26705,N_27379);
nand U28913 (N_28913,N_27534,N_26958);
and U28914 (N_28914,N_26915,N_26441);
nand U28915 (N_28915,N_27724,N_27932);
nand U28916 (N_28916,N_27706,N_26586);
nor U28917 (N_28917,N_27392,N_26276);
xnor U28918 (N_28918,N_26976,N_27063);
nand U28919 (N_28919,N_26997,N_26173);
xnor U28920 (N_28920,N_27873,N_26030);
or U28921 (N_28921,N_26194,N_26982);
or U28922 (N_28922,N_26426,N_27502);
nand U28923 (N_28923,N_27409,N_26749);
and U28924 (N_28924,N_26400,N_27556);
or U28925 (N_28925,N_26114,N_26605);
nor U28926 (N_28926,N_26594,N_27684);
or U28927 (N_28927,N_27611,N_27859);
or U28928 (N_28928,N_27294,N_26758);
nor U28929 (N_28929,N_26384,N_26769);
or U28930 (N_28930,N_27476,N_26382);
and U28931 (N_28931,N_27037,N_26009);
or U28932 (N_28932,N_27161,N_27852);
nand U28933 (N_28933,N_26797,N_26546);
or U28934 (N_28934,N_27154,N_27213);
or U28935 (N_28935,N_26614,N_26652);
and U28936 (N_28936,N_26937,N_26770);
nor U28937 (N_28937,N_26780,N_27819);
xnor U28938 (N_28938,N_26760,N_27660);
nor U28939 (N_28939,N_27554,N_27818);
xor U28940 (N_28940,N_26446,N_26377);
and U28941 (N_28941,N_26858,N_26873);
nor U28942 (N_28942,N_27468,N_26183);
nor U28943 (N_28943,N_26308,N_26495);
nand U28944 (N_28944,N_26082,N_27240);
and U28945 (N_28945,N_27207,N_26491);
nand U28946 (N_28946,N_26244,N_26156);
and U28947 (N_28947,N_27785,N_26029);
or U28948 (N_28948,N_27687,N_27696);
or U28949 (N_28949,N_26371,N_26098);
and U28950 (N_28950,N_26388,N_26202);
and U28951 (N_28951,N_27898,N_27323);
nand U28952 (N_28952,N_26227,N_26697);
nand U28953 (N_28953,N_27929,N_27784);
nor U28954 (N_28954,N_26523,N_26763);
and U28955 (N_28955,N_27540,N_27532);
nor U28956 (N_28956,N_26840,N_27507);
nor U28957 (N_28957,N_26975,N_26812);
nor U28958 (N_28958,N_27059,N_27188);
xnor U28959 (N_28959,N_27221,N_26810);
or U28960 (N_28960,N_27942,N_26138);
or U28961 (N_28961,N_26535,N_27338);
nor U28962 (N_28962,N_26520,N_26229);
nor U28963 (N_28963,N_27020,N_26396);
and U28964 (N_28964,N_26622,N_26775);
nor U28965 (N_28965,N_26462,N_26037);
nand U28966 (N_28966,N_27960,N_27505);
and U28967 (N_28967,N_27862,N_26095);
or U28968 (N_28968,N_26822,N_27395);
xor U28969 (N_28969,N_27796,N_27958);
and U28970 (N_28970,N_26683,N_26849);
or U28971 (N_28971,N_26072,N_26022);
or U28972 (N_28972,N_27104,N_26475);
and U28973 (N_28973,N_26952,N_27698);
nor U28974 (N_28974,N_27470,N_26463);
or U28975 (N_28975,N_26619,N_26502);
nand U28976 (N_28976,N_26580,N_26615);
or U28977 (N_28977,N_27286,N_27551);
and U28978 (N_28978,N_26567,N_26322);
and U28979 (N_28979,N_27547,N_26231);
or U28980 (N_28980,N_27349,N_27621);
nor U28981 (N_28981,N_27868,N_27982);
and U28982 (N_28982,N_26704,N_26132);
or U28983 (N_28983,N_27442,N_26693);
nor U28984 (N_28984,N_26859,N_26681);
nand U28985 (N_28985,N_26076,N_26292);
nand U28986 (N_28986,N_27181,N_27814);
nand U28987 (N_28987,N_27483,N_27067);
nor U28988 (N_28988,N_27641,N_26186);
or U28989 (N_28989,N_27835,N_27697);
nor U28990 (N_28990,N_27437,N_27332);
nand U28991 (N_28991,N_27041,N_27511);
nor U28992 (N_28992,N_27438,N_27152);
and U28993 (N_28993,N_27111,N_27607);
or U28994 (N_28994,N_27948,N_26624);
nand U28995 (N_28995,N_26299,N_27866);
nor U28996 (N_28996,N_27137,N_27347);
nor U28997 (N_28997,N_27406,N_27290);
xnor U28998 (N_28998,N_26457,N_26650);
and U28999 (N_28999,N_27956,N_26154);
nor U29000 (N_29000,N_27539,N_26394);
xnor U29001 (N_29001,N_26269,N_27714);
xnor U29002 (N_29002,N_26902,N_27108);
xor U29003 (N_29003,N_26953,N_27254);
xor U29004 (N_29004,N_26927,N_26090);
nor U29005 (N_29005,N_26757,N_27168);
nor U29006 (N_29006,N_26226,N_26309);
and U29007 (N_29007,N_27557,N_27973);
xnor U29008 (N_29008,N_26795,N_26107);
nand U29009 (N_29009,N_26627,N_27528);
or U29010 (N_29010,N_27322,N_26899);
xor U29011 (N_29011,N_27520,N_27867);
nor U29012 (N_29012,N_27103,N_27818);
nor U29013 (N_29013,N_26239,N_26526);
nor U29014 (N_29014,N_27111,N_27680);
and U29015 (N_29015,N_26617,N_27739);
and U29016 (N_29016,N_26646,N_26115);
and U29017 (N_29017,N_27549,N_26901);
nor U29018 (N_29018,N_26846,N_26126);
or U29019 (N_29019,N_27177,N_27436);
nand U29020 (N_29020,N_26822,N_26236);
or U29021 (N_29021,N_26003,N_27912);
xnor U29022 (N_29022,N_26400,N_26408);
and U29023 (N_29023,N_27915,N_27576);
or U29024 (N_29024,N_27745,N_26977);
nand U29025 (N_29025,N_27677,N_27381);
and U29026 (N_29026,N_27989,N_26242);
xnor U29027 (N_29027,N_26391,N_26928);
or U29028 (N_29028,N_27911,N_27311);
or U29029 (N_29029,N_26090,N_27576);
xor U29030 (N_29030,N_27368,N_26813);
nor U29031 (N_29031,N_26926,N_27978);
and U29032 (N_29032,N_27909,N_27730);
or U29033 (N_29033,N_26580,N_26963);
xnor U29034 (N_29034,N_26925,N_26944);
xor U29035 (N_29035,N_27315,N_26267);
nor U29036 (N_29036,N_26959,N_27405);
nor U29037 (N_29037,N_26672,N_26106);
nor U29038 (N_29038,N_26862,N_27847);
xnor U29039 (N_29039,N_26946,N_26731);
nor U29040 (N_29040,N_26091,N_26637);
or U29041 (N_29041,N_26958,N_26021);
nand U29042 (N_29042,N_27548,N_26917);
xor U29043 (N_29043,N_26415,N_27635);
nand U29044 (N_29044,N_26597,N_27422);
nand U29045 (N_29045,N_27769,N_27756);
nand U29046 (N_29046,N_27869,N_26875);
xnor U29047 (N_29047,N_27355,N_27977);
xnor U29048 (N_29048,N_26327,N_26584);
nand U29049 (N_29049,N_26933,N_26670);
nor U29050 (N_29050,N_26629,N_27107);
nand U29051 (N_29051,N_26327,N_27418);
xor U29052 (N_29052,N_26060,N_27076);
xnor U29053 (N_29053,N_27460,N_27754);
xnor U29054 (N_29054,N_26367,N_26599);
nand U29055 (N_29055,N_27907,N_27642);
xor U29056 (N_29056,N_26656,N_27600);
nand U29057 (N_29057,N_27369,N_26931);
xor U29058 (N_29058,N_27276,N_26549);
xor U29059 (N_29059,N_26293,N_26864);
or U29060 (N_29060,N_27557,N_27790);
and U29061 (N_29061,N_27134,N_26398);
nor U29062 (N_29062,N_27935,N_26897);
and U29063 (N_29063,N_26757,N_26540);
or U29064 (N_29064,N_26894,N_26196);
xnor U29065 (N_29065,N_26604,N_27983);
nor U29066 (N_29066,N_26123,N_26951);
nor U29067 (N_29067,N_26805,N_27379);
nor U29068 (N_29068,N_26904,N_27581);
and U29069 (N_29069,N_27129,N_27985);
xnor U29070 (N_29070,N_26762,N_27252);
nand U29071 (N_29071,N_27609,N_26078);
nor U29072 (N_29072,N_27908,N_26082);
or U29073 (N_29073,N_26528,N_27213);
nor U29074 (N_29074,N_27920,N_27137);
xor U29075 (N_29075,N_27832,N_27552);
or U29076 (N_29076,N_26036,N_26868);
xor U29077 (N_29077,N_27639,N_26264);
nor U29078 (N_29078,N_26196,N_27829);
or U29079 (N_29079,N_26858,N_27016);
or U29080 (N_29080,N_26076,N_26808);
xor U29081 (N_29081,N_26058,N_27675);
nand U29082 (N_29082,N_26560,N_26653);
and U29083 (N_29083,N_27883,N_27982);
or U29084 (N_29084,N_27303,N_26807);
or U29085 (N_29085,N_27978,N_27932);
nor U29086 (N_29086,N_26759,N_26790);
or U29087 (N_29087,N_26765,N_26987);
or U29088 (N_29088,N_26502,N_27684);
and U29089 (N_29089,N_26944,N_27217);
or U29090 (N_29090,N_26954,N_26994);
nand U29091 (N_29091,N_26048,N_27321);
nand U29092 (N_29092,N_27591,N_26565);
xor U29093 (N_29093,N_27127,N_27259);
and U29094 (N_29094,N_26638,N_27246);
nor U29095 (N_29095,N_27564,N_27384);
nand U29096 (N_29096,N_27376,N_26462);
nor U29097 (N_29097,N_27601,N_26426);
nand U29098 (N_29098,N_26218,N_26735);
nor U29099 (N_29099,N_26599,N_26325);
nor U29100 (N_29100,N_26247,N_27859);
and U29101 (N_29101,N_26895,N_27525);
xor U29102 (N_29102,N_26662,N_26141);
and U29103 (N_29103,N_27919,N_26971);
or U29104 (N_29104,N_26260,N_27128);
nor U29105 (N_29105,N_27984,N_27884);
or U29106 (N_29106,N_27382,N_27658);
nand U29107 (N_29107,N_26210,N_27977);
and U29108 (N_29108,N_26309,N_27771);
or U29109 (N_29109,N_26458,N_27504);
and U29110 (N_29110,N_26695,N_26444);
and U29111 (N_29111,N_26351,N_27699);
nand U29112 (N_29112,N_27682,N_26417);
and U29113 (N_29113,N_27258,N_26692);
xor U29114 (N_29114,N_27392,N_27989);
nor U29115 (N_29115,N_27878,N_27519);
xnor U29116 (N_29116,N_26777,N_27054);
or U29117 (N_29117,N_26110,N_27906);
and U29118 (N_29118,N_27188,N_27119);
xnor U29119 (N_29119,N_26967,N_27623);
nor U29120 (N_29120,N_26204,N_26486);
nor U29121 (N_29121,N_27904,N_26397);
nor U29122 (N_29122,N_26476,N_27045);
or U29123 (N_29123,N_26808,N_26687);
nor U29124 (N_29124,N_26266,N_27253);
nor U29125 (N_29125,N_27845,N_26135);
nand U29126 (N_29126,N_27858,N_27122);
or U29127 (N_29127,N_26907,N_26896);
xor U29128 (N_29128,N_26561,N_26307);
xor U29129 (N_29129,N_26286,N_26776);
nand U29130 (N_29130,N_26622,N_26534);
nor U29131 (N_29131,N_27709,N_26716);
or U29132 (N_29132,N_26459,N_27333);
nand U29133 (N_29133,N_27879,N_27306);
xnor U29134 (N_29134,N_27729,N_27859);
nor U29135 (N_29135,N_27107,N_27497);
nor U29136 (N_29136,N_27374,N_26797);
and U29137 (N_29137,N_26371,N_26122);
or U29138 (N_29138,N_27263,N_27874);
nor U29139 (N_29139,N_27445,N_26483);
xnor U29140 (N_29140,N_26789,N_27011);
and U29141 (N_29141,N_27218,N_27124);
nand U29142 (N_29142,N_26460,N_27749);
xor U29143 (N_29143,N_27477,N_26175);
nand U29144 (N_29144,N_27979,N_26996);
nand U29145 (N_29145,N_26848,N_27299);
nor U29146 (N_29146,N_27964,N_26996);
nor U29147 (N_29147,N_26037,N_27585);
or U29148 (N_29148,N_27336,N_26427);
or U29149 (N_29149,N_26902,N_27122);
nor U29150 (N_29150,N_26941,N_27973);
nand U29151 (N_29151,N_27936,N_26013);
nor U29152 (N_29152,N_26449,N_26055);
nand U29153 (N_29153,N_27933,N_27461);
nand U29154 (N_29154,N_27974,N_26503);
xor U29155 (N_29155,N_27265,N_27591);
and U29156 (N_29156,N_27105,N_27024);
or U29157 (N_29157,N_27591,N_26682);
and U29158 (N_29158,N_26479,N_26689);
nand U29159 (N_29159,N_26479,N_26883);
nand U29160 (N_29160,N_27083,N_26529);
xor U29161 (N_29161,N_26163,N_26306);
xor U29162 (N_29162,N_27729,N_26063);
and U29163 (N_29163,N_27011,N_27148);
nor U29164 (N_29164,N_27747,N_27099);
xor U29165 (N_29165,N_26367,N_27870);
and U29166 (N_29166,N_26821,N_26536);
nor U29167 (N_29167,N_27047,N_26276);
or U29168 (N_29168,N_27578,N_26710);
nand U29169 (N_29169,N_26713,N_26378);
xor U29170 (N_29170,N_27791,N_27834);
nand U29171 (N_29171,N_27261,N_26112);
or U29172 (N_29172,N_26586,N_26555);
nand U29173 (N_29173,N_26256,N_26731);
nor U29174 (N_29174,N_27058,N_26390);
or U29175 (N_29175,N_26317,N_27428);
and U29176 (N_29176,N_26976,N_26628);
and U29177 (N_29177,N_27391,N_26055);
nand U29178 (N_29178,N_27313,N_26073);
xor U29179 (N_29179,N_26477,N_27037);
xnor U29180 (N_29180,N_27352,N_26400);
or U29181 (N_29181,N_26473,N_27251);
xor U29182 (N_29182,N_27240,N_27217);
nor U29183 (N_29183,N_26838,N_26926);
or U29184 (N_29184,N_27891,N_27539);
nand U29185 (N_29185,N_26650,N_27224);
nand U29186 (N_29186,N_27095,N_26498);
xor U29187 (N_29187,N_27974,N_26079);
nor U29188 (N_29188,N_26421,N_26870);
nor U29189 (N_29189,N_27625,N_26887);
nor U29190 (N_29190,N_27350,N_27039);
nor U29191 (N_29191,N_26629,N_27335);
or U29192 (N_29192,N_26123,N_27163);
nand U29193 (N_29193,N_26445,N_27505);
xor U29194 (N_29194,N_26197,N_26112);
and U29195 (N_29195,N_26318,N_26941);
xor U29196 (N_29196,N_26276,N_26953);
nor U29197 (N_29197,N_26265,N_27195);
xnor U29198 (N_29198,N_26156,N_26020);
xor U29199 (N_29199,N_27932,N_26590);
nand U29200 (N_29200,N_26441,N_27887);
nor U29201 (N_29201,N_26280,N_27696);
or U29202 (N_29202,N_26528,N_26288);
nand U29203 (N_29203,N_27222,N_26220);
nand U29204 (N_29204,N_26265,N_26123);
or U29205 (N_29205,N_27491,N_26089);
xnor U29206 (N_29206,N_27370,N_27382);
xnor U29207 (N_29207,N_27753,N_27896);
xor U29208 (N_29208,N_27825,N_26727);
nor U29209 (N_29209,N_26720,N_26458);
xor U29210 (N_29210,N_27419,N_27875);
nor U29211 (N_29211,N_27502,N_27592);
nor U29212 (N_29212,N_27581,N_26495);
nand U29213 (N_29213,N_26570,N_27020);
and U29214 (N_29214,N_26896,N_26940);
nor U29215 (N_29215,N_27194,N_26547);
xor U29216 (N_29216,N_27606,N_27183);
nor U29217 (N_29217,N_26741,N_27984);
nor U29218 (N_29218,N_27308,N_26254);
nand U29219 (N_29219,N_27746,N_27360);
xor U29220 (N_29220,N_27794,N_27240);
xnor U29221 (N_29221,N_26911,N_26112);
nand U29222 (N_29222,N_27489,N_26290);
or U29223 (N_29223,N_27878,N_27211);
nand U29224 (N_29224,N_27534,N_27760);
xor U29225 (N_29225,N_26978,N_26340);
nand U29226 (N_29226,N_27453,N_26338);
xnor U29227 (N_29227,N_26584,N_27989);
xor U29228 (N_29228,N_26585,N_27791);
or U29229 (N_29229,N_27099,N_27425);
nand U29230 (N_29230,N_26947,N_26986);
nand U29231 (N_29231,N_26531,N_26875);
or U29232 (N_29232,N_27441,N_27496);
and U29233 (N_29233,N_27572,N_26763);
nand U29234 (N_29234,N_26491,N_26050);
nor U29235 (N_29235,N_27784,N_27316);
nor U29236 (N_29236,N_26413,N_26762);
nor U29237 (N_29237,N_26098,N_27647);
nor U29238 (N_29238,N_26790,N_27162);
nand U29239 (N_29239,N_27316,N_27797);
or U29240 (N_29240,N_26342,N_27860);
nor U29241 (N_29241,N_27938,N_26988);
or U29242 (N_29242,N_27937,N_26165);
and U29243 (N_29243,N_27686,N_26493);
nand U29244 (N_29244,N_26414,N_26054);
or U29245 (N_29245,N_26267,N_26569);
or U29246 (N_29246,N_26195,N_26077);
or U29247 (N_29247,N_26880,N_27951);
and U29248 (N_29248,N_27281,N_27635);
or U29249 (N_29249,N_27435,N_27751);
or U29250 (N_29250,N_27517,N_26517);
or U29251 (N_29251,N_26242,N_27953);
nor U29252 (N_29252,N_27264,N_27559);
nor U29253 (N_29253,N_26995,N_26423);
nand U29254 (N_29254,N_26741,N_26674);
and U29255 (N_29255,N_27897,N_26740);
or U29256 (N_29256,N_27636,N_27844);
and U29257 (N_29257,N_27976,N_26804);
nor U29258 (N_29258,N_26289,N_27322);
xor U29259 (N_29259,N_26440,N_26074);
and U29260 (N_29260,N_26107,N_27528);
and U29261 (N_29261,N_27529,N_26007);
nor U29262 (N_29262,N_26141,N_26594);
and U29263 (N_29263,N_26141,N_27539);
xor U29264 (N_29264,N_26698,N_27406);
nand U29265 (N_29265,N_27452,N_26719);
and U29266 (N_29266,N_26115,N_27063);
nor U29267 (N_29267,N_26809,N_27403);
nor U29268 (N_29268,N_27016,N_26970);
nand U29269 (N_29269,N_26298,N_27789);
nand U29270 (N_29270,N_26831,N_26963);
nand U29271 (N_29271,N_26129,N_26544);
or U29272 (N_29272,N_27943,N_27403);
and U29273 (N_29273,N_26941,N_26614);
nor U29274 (N_29274,N_26076,N_27355);
or U29275 (N_29275,N_27300,N_26901);
or U29276 (N_29276,N_26959,N_27591);
or U29277 (N_29277,N_27795,N_27315);
nand U29278 (N_29278,N_27165,N_27941);
nor U29279 (N_29279,N_26541,N_27932);
xor U29280 (N_29280,N_27222,N_27605);
or U29281 (N_29281,N_27582,N_26328);
xnor U29282 (N_29282,N_26907,N_26092);
and U29283 (N_29283,N_27082,N_27774);
or U29284 (N_29284,N_27735,N_27056);
nand U29285 (N_29285,N_26606,N_26204);
nor U29286 (N_29286,N_27689,N_26436);
or U29287 (N_29287,N_27192,N_27469);
xor U29288 (N_29288,N_26896,N_27507);
xor U29289 (N_29289,N_26361,N_26452);
xnor U29290 (N_29290,N_26766,N_26778);
and U29291 (N_29291,N_26886,N_27684);
or U29292 (N_29292,N_26856,N_27638);
and U29293 (N_29293,N_27582,N_27723);
and U29294 (N_29294,N_27283,N_26182);
or U29295 (N_29295,N_26991,N_26072);
or U29296 (N_29296,N_27984,N_26362);
nand U29297 (N_29297,N_26462,N_26461);
xor U29298 (N_29298,N_26192,N_27501);
and U29299 (N_29299,N_27283,N_26860);
xnor U29300 (N_29300,N_26929,N_26326);
or U29301 (N_29301,N_27090,N_27167);
nand U29302 (N_29302,N_27457,N_26180);
xnor U29303 (N_29303,N_26996,N_27601);
xnor U29304 (N_29304,N_26128,N_27065);
nand U29305 (N_29305,N_26957,N_27415);
nand U29306 (N_29306,N_26027,N_27323);
xnor U29307 (N_29307,N_27576,N_27619);
nor U29308 (N_29308,N_26042,N_26276);
or U29309 (N_29309,N_26773,N_26677);
or U29310 (N_29310,N_27729,N_27582);
or U29311 (N_29311,N_27673,N_27902);
nand U29312 (N_29312,N_27810,N_26091);
or U29313 (N_29313,N_27322,N_27631);
or U29314 (N_29314,N_26906,N_26839);
nor U29315 (N_29315,N_26360,N_26880);
xnor U29316 (N_29316,N_26423,N_26316);
and U29317 (N_29317,N_26697,N_27283);
or U29318 (N_29318,N_27155,N_26912);
and U29319 (N_29319,N_26746,N_26358);
or U29320 (N_29320,N_26582,N_26556);
or U29321 (N_29321,N_26837,N_26112);
nand U29322 (N_29322,N_26147,N_26161);
and U29323 (N_29323,N_26904,N_27468);
or U29324 (N_29324,N_27967,N_27175);
and U29325 (N_29325,N_26124,N_26232);
or U29326 (N_29326,N_27160,N_27095);
nand U29327 (N_29327,N_26778,N_26896);
nand U29328 (N_29328,N_26159,N_27880);
nor U29329 (N_29329,N_26180,N_27805);
or U29330 (N_29330,N_26563,N_26362);
nor U29331 (N_29331,N_27841,N_27570);
or U29332 (N_29332,N_27543,N_26881);
or U29333 (N_29333,N_27277,N_26672);
or U29334 (N_29334,N_27536,N_26445);
or U29335 (N_29335,N_26402,N_27022);
or U29336 (N_29336,N_26686,N_26605);
nand U29337 (N_29337,N_26001,N_27522);
nor U29338 (N_29338,N_26138,N_27071);
xor U29339 (N_29339,N_27613,N_27643);
nand U29340 (N_29340,N_26903,N_27825);
nor U29341 (N_29341,N_27197,N_26770);
or U29342 (N_29342,N_27694,N_27297);
nand U29343 (N_29343,N_26711,N_26171);
or U29344 (N_29344,N_26789,N_27588);
or U29345 (N_29345,N_27700,N_26940);
xnor U29346 (N_29346,N_27683,N_26031);
and U29347 (N_29347,N_26973,N_26707);
nand U29348 (N_29348,N_27082,N_27501);
nor U29349 (N_29349,N_26048,N_27634);
xnor U29350 (N_29350,N_26839,N_27754);
and U29351 (N_29351,N_27291,N_27204);
xnor U29352 (N_29352,N_26851,N_26750);
nand U29353 (N_29353,N_26645,N_26234);
and U29354 (N_29354,N_27310,N_27022);
nor U29355 (N_29355,N_26961,N_27195);
xnor U29356 (N_29356,N_27380,N_26931);
and U29357 (N_29357,N_26374,N_27812);
nor U29358 (N_29358,N_26688,N_27254);
nor U29359 (N_29359,N_26537,N_26809);
nand U29360 (N_29360,N_26751,N_27248);
and U29361 (N_29361,N_26834,N_27422);
nand U29362 (N_29362,N_27471,N_27755);
xor U29363 (N_29363,N_27536,N_27198);
xor U29364 (N_29364,N_27773,N_26685);
xnor U29365 (N_29365,N_26450,N_27005);
and U29366 (N_29366,N_27259,N_27894);
xor U29367 (N_29367,N_26945,N_27205);
nand U29368 (N_29368,N_27138,N_27360);
and U29369 (N_29369,N_26296,N_26561);
and U29370 (N_29370,N_27595,N_27364);
nor U29371 (N_29371,N_27303,N_26785);
nor U29372 (N_29372,N_27694,N_26429);
nand U29373 (N_29373,N_27103,N_27212);
and U29374 (N_29374,N_27072,N_27832);
or U29375 (N_29375,N_27194,N_26778);
nor U29376 (N_29376,N_26807,N_26279);
nand U29377 (N_29377,N_27472,N_26627);
or U29378 (N_29378,N_27744,N_26745);
nand U29379 (N_29379,N_26321,N_26689);
and U29380 (N_29380,N_26177,N_26129);
or U29381 (N_29381,N_27484,N_27788);
nand U29382 (N_29382,N_26364,N_27216);
and U29383 (N_29383,N_27095,N_27010);
nor U29384 (N_29384,N_26476,N_26972);
or U29385 (N_29385,N_26054,N_27449);
or U29386 (N_29386,N_27750,N_26636);
and U29387 (N_29387,N_26875,N_26880);
and U29388 (N_29388,N_26932,N_26099);
nor U29389 (N_29389,N_26767,N_26375);
nor U29390 (N_29390,N_26065,N_26574);
and U29391 (N_29391,N_27725,N_26574);
or U29392 (N_29392,N_26214,N_27150);
xor U29393 (N_29393,N_27407,N_26225);
or U29394 (N_29394,N_26323,N_27234);
nor U29395 (N_29395,N_27931,N_27104);
and U29396 (N_29396,N_26736,N_26658);
and U29397 (N_29397,N_27116,N_27336);
xor U29398 (N_29398,N_26410,N_27434);
or U29399 (N_29399,N_27892,N_26584);
or U29400 (N_29400,N_26299,N_26684);
xnor U29401 (N_29401,N_26102,N_27569);
and U29402 (N_29402,N_26918,N_27434);
or U29403 (N_29403,N_27698,N_27919);
nand U29404 (N_29404,N_27484,N_27717);
xor U29405 (N_29405,N_27314,N_26412);
or U29406 (N_29406,N_26242,N_26723);
and U29407 (N_29407,N_27349,N_26592);
xor U29408 (N_29408,N_26594,N_27787);
and U29409 (N_29409,N_27921,N_27178);
nand U29410 (N_29410,N_26483,N_27233);
and U29411 (N_29411,N_27115,N_26481);
or U29412 (N_29412,N_26281,N_27283);
or U29413 (N_29413,N_27450,N_27645);
or U29414 (N_29414,N_26549,N_27659);
nand U29415 (N_29415,N_27997,N_27799);
xnor U29416 (N_29416,N_26300,N_26041);
nand U29417 (N_29417,N_27750,N_26536);
or U29418 (N_29418,N_26122,N_27750);
nor U29419 (N_29419,N_27661,N_26504);
and U29420 (N_29420,N_26042,N_26866);
and U29421 (N_29421,N_27001,N_26207);
and U29422 (N_29422,N_27677,N_26991);
or U29423 (N_29423,N_26016,N_27550);
nor U29424 (N_29424,N_26991,N_26796);
xnor U29425 (N_29425,N_27876,N_26878);
nor U29426 (N_29426,N_26163,N_27695);
xor U29427 (N_29427,N_27621,N_26973);
nand U29428 (N_29428,N_27727,N_26800);
nor U29429 (N_29429,N_26206,N_27366);
xor U29430 (N_29430,N_27713,N_26140);
and U29431 (N_29431,N_26680,N_27260);
nand U29432 (N_29432,N_27405,N_27978);
nor U29433 (N_29433,N_26056,N_26618);
nor U29434 (N_29434,N_27076,N_26192);
and U29435 (N_29435,N_27511,N_27628);
nor U29436 (N_29436,N_27506,N_27198);
or U29437 (N_29437,N_26341,N_26903);
or U29438 (N_29438,N_26462,N_26478);
xnor U29439 (N_29439,N_27155,N_26211);
xnor U29440 (N_29440,N_26369,N_27907);
nand U29441 (N_29441,N_27620,N_27079);
and U29442 (N_29442,N_26886,N_27785);
nor U29443 (N_29443,N_27946,N_27999);
and U29444 (N_29444,N_26789,N_27837);
and U29445 (N_29445,N_27530,N_27697);
nor U29446 (N_29446,N_26060,N_26008);
nor U29447 (N_29447,N_27471,N_26859);
and U29448 (N_29448,N_26773,N_27152);
nor U29449 (N_29449,N_27129,N_27823);
nand U29450 (N_29450,N_27189,N_26201);
or U29451 (N_29451,N_27787,N_27235);
nor U29452 (N_29452,N_27838,N_26376);
nor U29453 (N_29453,N_27946,N_27208);
nor U29454 (N_29454,N_26378,N_26647);
xnor U29455 (N_29455,N_27184,N_26781);
and U29456 (N_29456,N_27375,N_26509);
xnor U29457 (N_29457,N_26428,N_27757);
or U29458 (N_29458,N_27128,N_27511);
nand U29459 (N_29459,N_27266,N_26906);
xnor U29460 (N_29460,N_26512,N_26932);
or U29461 (N_29461,N_26659,N_27268);
xnor U29462 (N_29462,N_26761,N_26207);
xnor U29463 (N_29463,N_26485,N_26352);
and U29464 (N_29464,N_26182,N_26401);
nor U29465 (N_29465,N_27000,N_26187);
nor U29466 (N_29466,N_26292,N_26904);
or U29467 (N_29467,N_27360,N_27989);
nand U29468 (N_29468,N_26740,N_26338);
and U29469 (N_29469,N_26416,N_27822);
nor U29470 (N_29470,N_26821,N_26322);
nor U29471 (N_29471,N_26255,N_27790);
xor U29472 (N_29472,N_26024,N_26297);
nand U29473 (N_29473,N_26863,N_27964);
nand U29474 (N_29474,N_26362,N_27886);
nand U29475 (N_29475,N_27656,N_27405);
or U29476 (N_29476,N_26774,N_27420);
nor U29477 (N_29477,N_26060,N_27775);
and U29478 (N_29478,N_27982,N_26150);
and U29479 (N_29479,N_26629,N_27057);
nand U29480 (N_29480,N_26091,N_26015);
nor U29481 (N_29481,N_26730,N_27252);
or U29482 (N_29482,N_27786,N_26631);
and U29483 (N_29483,N_26064,N_26345);
or U29484 (N_29484,N_26740,N_27511);
xor U29485 (N_29485,N_26035,N_26545);
and U29486 (N_29486,N_26694,N_27146);
nand U29487 (N_29487,N_27688,N_26406);
and U29488 (N_29488,N_27699,N_27931);
nand U29489 (N_29489,N_27661,N_27141);
and U29490 (N_29490,N_26737,N_26569);
nand U29491 (N_29491,N_27028,N_26457);
and U29492 (N_29492,N_27920,N_26397);
or U29493 (N_29493,N_27876,N_26778);
nor U29494 (N_29494,N_26637,N_27095);
xor U29495 (N_29495,N_27086,N_26061);
nand U29496 (N_29496,N_27255,N_26682);
xnor U29497 (N_29497,N_26425,N_26040);
or U29498 (N_29498,N_26719,N_26800);
xor U29499 (N_29499,N_26004,N_27528);
xor U29500 (N_29500,N_27688,N_27615);
nor U29501 (N_29501,N_27726,N_27673);
xor U29502 (N_29502,N_26839,N_27917);
xor U29503 (N_29503,N_27417,N_27770);
xnor U29504 (N_29504,N_27096,N_26091);
nor U29505 (N_29505,N_27983,N_26336);
nand U29506 (N_29506,N_26747,N_26708);
or U29507 (N_29507,N_26843,N_27277);
or U29508 (N_29508,N_26850,N_26259);
or U29509 (N_29509,N_27179,N_26352);
nand U29510 (N_29510,N_26834,N_27464);
nor U29511 (N_29511,N_26272,N_27669);
and U29512 (N_29512,N_27560,N_27038);
xor U29513 (N_29513,N_27679,N_27706);
xnor U29514 (N_29514,N_27489,N_26716);
xor U29515 (N_29515,N_26224,N_26388);
and U29516 (N_29516,N_26745,N_27475);
xnor U29517 (N_29517,N_26004,N_27125);
and U29518 (N_29518,N_26275,N_26353);
or U29519 (N_29519,N_26923,N_26531);
nand U29520 (N_29520,N_26395,N_26151);
nand U29521 (N_29521,N_27873,N_27260);
nor U29522 (N_29522,N_27238,N_26275);
or U29523 (N_29523,N_27680,N_27269);
nand U29524 (N_29524,N_27396,N_26047);
nand U29525 (N_29525,N_27227,N_26593);
or U29526 (N_29526,N_27015,N_27464);
nand U29527 (N_29527,N_26422,N_27774);
or U29528 (N_29528,N_27988,N_26328);
or U29529 (N_29529,N_27930,N_26680);
nor U29530 (N_29530,N_26791,N_27689);
nand U29531 (N_29531,N_27906,N_27646);
and U29532 (N_29532,N_26905,N_26663);
or U29533 (N_29533,N_26770,N_27334);
nor U29534 (N_29534,N_26520,N_26967);
nor U29535 (N_29535,N_27852,N_27482);
or U29536 (N_29536,N_26208,N_27165);
nor U29537 (N_29537,N_27722,N_27590);
or U29538 (N_29538,N_27634,N_26216);
and U29539 (N_29539,N_26754,N_27671);
xor U29540 (N_29540,N_26796,N_27345);
nand U29541 (N_29541,N_27864,N_26117);
nor U29542 (N_29542,N_26395,N_27297);
or U29543 (N_29543,N_27830,N_26552);
nand U29544 (N_29544,N_27533,N_26286);
nand U29545 (N_29545,N_27830,N_26567);
nor U29546 (N_29546,N_27106,N_26371);
nand U29547 (N_29547,N_26300,N_26953);
xor U29548 (N_29548,N_27212,N_26923);
xor U29549 (N_29549,N_26109,N_26276);
nor U29550 (N_29550,N_26864,N_26221);
nor U29551 (N_29551,N_27125,N_27355);
nor U29552 (N_29552,N_26006,N_27102);
xnor U29553 (N_29553,N_27304,N_26472);
nand U29554 (N_29554,N_27037,N_27745);
nand U29555 (N_29555,N_26367,N_27556);
or U29556 (N_29556,N_26475,N_27323);
or U29557 (N_29557,N_27924,N_27629);
and U29558 (N_29558,N_27604,N_26057);
nand U29559 (N_29559,N_26292,N_26549);
and U29560 (N_29560,N_26682,N_27187);
xor U29561 (N_29561,N_27895,N_27602);
and U29562 (N_29562,N_26089,N_26118);
xor U29563 (N_29563,N_27140,N_26090);
nand U29564 (N_29564,N_27346,N_26102);
xnor U29565 (N_29565,N_27476,N_27595);
nand U29566 (N_29566,N_27783,N_27983);
nand U29567 (N_29567,N_26738,N_26853);
and U29568 (N_29568,N_27676,N_27816);
and U29569 (N_29569,N_26458,N_27963);
xor U29570 (N_29570,N_26391,N_27689);
nand U29571 (N_29571,N_27541,N_26167);
or U29572 (N_29572,N_26355,N_27672);
or U29573 (N_29573,N_27914,N_27733);
xnor U29574 (N_29574,N_26654,N_27783);
or U29575 (N_29575,N_27984,N_26593);
or U29576 (N_29576,N_27380,N_26201);
or U29577 (N_29577,N_27784,N_27524);
or U29578 (N_29578,N_27604,N_26567);
nand U29579 (N_29579,N_26398,N_26183);
or U29580 (N_29580,N_26259,N_27454);
nor U29581 (N_29581,N_27160,N_26917);
xnor U29582 (N_29582,N_26537,N_27288);
and U29583 (N_29583,N_26971,N_27853);
nor U29584 (N_29584,N_27091,N_27096);
and U29585 (N_29585,N_26615,N_27203);
and U29586 (N_29586,N_27716,N_27485);
nor U29587 (N_29587,N_26772,N_26038);
xnor U29588 (N_29588,N_27278,N_26602);
nor U29589 (N_29589,N_26831,N_26656);
and U29590 (N_29590,N_27637,N_27529);
or U29591 (N_29591,N_27385,N_26625);
and U29592 (N_29592,N_26198,N_26364);
and U29593 (N_29593,N_27601,N_26473);
xor U29594 (N_29594,N_27577,N_26658);
and U29595 (N_29595,N_26025,N_27958);
nand U29596 (N_29596,N_27593,N_26092);
nand U29597 (N_29597,N_26411,N_27721);
or U29598 (N_29598,N_26386,N_27973);
or U29599 (N_29599,N_26003,N_26270);
and U29600 (N_29600,N_26535,N_26362);
nand U29601 (N_29601,N_26014,N_27093);
nand U29602 (N_29602,N_27826,N_26810);
and U29603 (N_29603,N_27776,N_27107);
nor U29604 (N_29604,N_26713,N_26233);
or U29605 (N_29605,N_26444,N_27151);
xor U29606 (N_29606,N_26858,N_27408);
and U29607 (N_29607,N_26055,N_26672);
xnor U29608 (N_29608,N_26365,N_26540);
nor U29609 (N_29609,N_26858,N_27015);
or U29610 (N_29610,N_26327,N_27702);
xnor U29611 (N_29611,N_26618,N_26858);
nor U29612 (N_29612,N_26060,N_26169);
or U29613 (N_29613,N_27651,N_26103);
nor U29614 (N_29614,N_27509,N_26508);
and U29615 (N_29615,N_27807,N_27630);
nor U29616 (N_29616,N_27291,N_27209);
nand U29617 (N_29617,N_27607,N_26659);
or U29618 (N_29618,N_27127,N_26818);
nand U29619 (N_29619,N_27510,N_26121);
and U29620 (N_29620,N_27362,N_27192);
and U29621 (N_29621,N_27841,N_26733);
or U29622 (N_29622,N_27820,N_27266);
xor U29623 (N_29623,N_27610,N_27310);
nor U29624 (N_29624,N_27392,N_26554);
and U29625 (N_29625,N_26764,N_27714);
or U29626 (N_29626,N_27819,N_26265);
nor U29627 (N_29627,N_27743,N_26875);
or U29628 (N_29628,N_26163,N_26332);
nor U29629 (N_29629,N_27590,N_27682);
or U29630 (N_29630,N_27313,N_27641);
or U29631 (N_29631,N_27545,N_27632);
xor U29632 (N_29632,N_26137,N_26823);
or U29633 (N_29633,N_27445,N_27157);
nand U29634 (N_29634,N_27079,N_27759);
nand U29635 (N_29635,N_27666,N_26952);
nand U29636 (N_29636,N_27414,N_26073);
and U29637 (N_29637,N_27383,N_27832);
nand U29638 (N_29638,N_26837,N_27159);
xor U29639 (N_29639,N_26791,N_27341);
nor U29640 (N_29640,N_26380,N_27939);
xor U29641 (N_29641,N_27179,N_27818);
xnor U29642 (N_29642,N_27821,N_27338);
and U29643 (N_29643,N_27903,N_27730);
nor U29644 (N_29644,N_26415,N_26991);
or U29645 (N_29645,N_26629,N_26460);
nor U29646 (N_29646,N_26499,N_27430);
or U29647 (N_29647,N_27696,N_27430);
nand U29648 (N_29648,N_26850,N_27849);
or U29649 (N_29649,N_27883,N_26742);
xnor U29650 (N_29650,N_27285,N_27609);
xor U29651 (N_29651,N_27289,N_26705);
and U29652 (N_29652,N_26937,N_27594);
and U29653 (N_29653,N_26364,N_26233);
nand U29654 (N_29654,N_26677,N_26760);
and U29655 (N_29655,N_26235,N_27049);
xnor U29656 (N_29656,N_27067,N_27273);
xnor U29657 (N_29657,N_27947,N_27781);
or U29658 (N_29658,N_27385,N_27429);
nand U29659 (N_29659,N_27434,N_26449);
and U29660 (N_29660,N_26977,N_26725);
or U29661 (N_29661,N_27363,N_27025);
xor U29662 (N_29662,N_26504,N_27578);
nand U29663 (N_29663,N_27738,N_27464);
xor U29664 (N_29664,N_27798,N_26854);
or U29665 (N_29665,N_27383,N_27009);
and U29666 (N_29666,N_27347,N_27179);
nand U29667 (N_29667,N_26459,N_26480);
and U29668 (N_29668,N_27001,N_27572);
xor U29669 (N_29669,N_27346,N_26030);
nor U29670 (N_29670,N_26556,N_27768);
nor U29671 (N_29671,N_27277,N_27155);
or U29672 (N_29672,N_26111,N_26185);
nand U29673 (N_29673,N_27262,N_26582);
nor U29674 (N_29674,N_27935,N_27774);
and U29675 (N_29675,N_26581,N_27194);
xor U29676 (N_29676,N_26331,N_26181);
or U29677 (N_29677,N_27977,N_27212);
nand U29678 (N_29678,N_27060,N_26735);
and U29679 (N_29679,N_27934,N_27587);
or U29680 (N_29680,N_26430,N_26263);
xor U29681 (N_29681,N_27462,N_27909);
nand U29682 (N_29682,N_27996,N_26172);
nor U29683 (N_29683,N_27920,N_27157);
nand U29684 (N_29684,N_27642,N_26009);
nand U29685 (N_29685,N_26780,N_26966);
or U29686 (N_29686,N_27901,N_27086);
nor U29687 (N_29687,N_27777,N_26849);
or U29688 (N_29688,N_26041,N_26258);
nor U29689 (N_29689,N_27187,N_26941);
xor U29690 (N_29690,N_26434,N_27568);
nand U29691 (N_29691,N_27835,N_27072);
nor U29692 (N_29692,N_26649,N_27325);
nand U29693 (N_29693,N_27128,N_27423);
nor U29694 (N_29694,N_27668,N_27976);
nand U29695 (N_29695,N_27890,N_27640);
or U29696 (N_29696,N_27418,N_26713);
and U29697 (N_29697,N_27235,N_27525);
nand U29698 (N_29698,N_26164,N_26022);
and U29699 (N_29699,N_26119,N_27166);
nand U29700 (N_29700,N_26410,N_27702);
xnor U29701 (N_29701,N_26829,N_26180);
xnor U29702 (N_29702,N_26034,N_27944);
xor U29703 (N_29703,N_26366,N_26908);
nor U29704 (N_29704,N_26754,N_26778);
xnor U29705 (N_29705,N_27414,N_26036);
or U29706 (N_29706,N_27659,N_27043);
or U29707 (N_29707,N_27189,N_27282);
nand U29708 (N_29708,N_26519,N_26951);
nor U29709 (N_29709,N_26133,N_26484);
nor U29710 (N_29710,N_27756,N_27951);
nor U29711 (N_29711,N_26080,N_27055);
nor U29712 (N_29712,N_26045,N_26240);
and U29713 (N_29713,N_27660,N_26043);
or U29714 (N_29714,N_26086,N_27997);
nor U29715 (N_29715,N_26915,N_27273);
nand U29716 (N_29716,N_26136,N_27655);
nor U29717 (N_29717,N_26349,N_27563);
nand U29718 (N_29718,N_27111,N_27929);
nor U29719 (N_29719,N_27909,N_27996);
nand U29720 (N_29720,N_27903,N_26609);
nor U29721 (N_29721,N_26781,N_26158);
or U29722 (N_29722,N_26830,N_26660);
xor U29723 (N_29723,N_27425,N_27003);
and U29724 (N_29724,N_27769,N_27080);
xnor U29725 (N_29725,N_26598,N_27078);
nor U29726 (N_29726,N_27058,N_27503);
nor U29727 (N_29727,N_26252,N_26925);
nor U29728 (N_29728,N_27692,N_26524);
nor U29729 (N_29729,N_26270,N_27217);
and U29730 (N_29730,N_26700,N_27926);
xnor U29731 (N_29731,N_27568,N_26925);
nand U29732 (N_29732,N_26978,N_27424);
and U29733 (N_29733,N_26169,N_26587);
xor U29734 (N_29734,N_26292,N_26932);
and U29735 (N_29735,N_27838,N_26151);
xor U29736 (N_29736,N_26875,N_27504);
and U29737 (N_29737,N_27309,N_26740);
nor U29738 (N_29738,N_26866,N_26732);
xor U29739 (N_29739,N_27830,N_26252);
nor U29740 (N_29740,N_26918,N_26266);
or U29741 (N_29741,N_26039,N_27121);
nand U29742 (N_29742,N_26755,N_26442);
nand U29743 (N_29743,N_27242,N_26057);
nor U29744 (N_29744,N_27225,N_27720);
nor U29745 (N_29745,N_26191,N_26676);
nor U29746 (N_29746,N_26437,N_26818);
and U29747 (N_29747,N_27961,N_26562);
nor U29748 (N_29748,N_27591,N_26125);
or U29749 (N_29749,N_27622,N_26297);
xor U29750 (N_29750,N_26713,N_27940);
or U29751 (N_29751,N_26040,N_26452);
xnor U29752 (N_29752,N_27705,N_27585);
nand U29753 (N_29753,N_26851,N_27722);
nand U29754 (N_29754,N_27513,N_26800);
and U29755 (N_29755,N_27586,N_26625);
nor U29756 (N_29756,N_27956,N_27122);
nor U29757 (N_29757,N_26184,N_26540);
and U29758 (N_29758,N_27858,N_27495);
and U29759 (N_29759,N_27281,N_27832);
xnor U29760 (N_29760,N_26258,N_27856);
nor U29761 (N_29761,N_26281,N_27669);
or U29762 (N_29762,N_27470,N_26586);
nand U29763 (N_29763,N_26014,N_26760);
nor U29764 (N_29764,N_27938,N_26970);
or U29765 (N_29765,N_26883,N_27934);
xor U29766 (N_29766,N_27143,N_26768);
xor U29767 (N_29767,N_27868,N_26392);
or U29768 (N_29768,N_26704,N_27334);
nand U29769 (N_29769,N_26846,N_27312);
nand U29770 (N_29770,N_27216,N_27118);
xor U29771 (N_29771,N_27284,N_27200);
xnor U29772 (N_29772,N_26022,N_27727);
xor U29773 (N_29773,N_27614,N_27861);
or U29774 (N_29774,N_26195,N_27577);
nand U29775 (N_29775,N_26384,N_26940);
or U29776 (N_29776,N_26388,N_26859);
or U29777 (N_29777,N_26938,N_27141);
nand U29778 (N_29778,N_26010,N_27081);
xnor U29779 (N_29779,N_26376,N_27878);
nand U29780 (N_29780,N_26038,N_27611);
and U29781 (N_29781,N_26040,N_27853);
nand U29782 (N_29782,N_27517,N_27671);
or U29783 (N_29783,N_27605,N_26486);
or U29784 (N_29784,N_27430,N_26010);
xor U29785 (N_29785,N_27912,N_26301);
nor U29786 (N_29786,N_27453,N_26646);
and U29787 (N_29787,N_26174,N_27876);
and U29788 (N_29788,N_27515,N_26713);
nor U29789 (N_29789,N_27427,N_27808);
xor U29790 (N_29790,N_27889,N_27697);
or U29791 (N_29791,N_26729,N_26558);
or U29792 (N_29792,N_26570,N_26027);
nand U29793 (N_29793,N_27163,N_26395);
and U29794 (N_29794,N_27910,N_27877);
nor U29795 (N_29795,N_27982,N_27887);
nor U29796 (N_29796,N_27033,N_26388);
nand U29797 (N_29797,N_27102,N_27021);
nand U29798 (N_29798,N_27174,N_26920);
or U29799 (N_29799,N_27210,N_27311);
or U29800 (N_29800,N_27560,N_27787);
and U29801 (N_29801,N_27363,N_26043);
nor U29802 (N_29802,N_27294,N_27180);
or U29803 (N_29803,N_27432,N_27755);
or U29804 (N_29804,N_26452,N_26956);
and U29805 (N_29805,N_27430,N_26999);
or U29806 (N_29806,N_26120,N_26550);
nor U29807 (N_29807,N_26614,N_27400);
and U29808 (N_29808,N_26022,N_27616);
and U29809 (N_29809,N_27664,N_27268);
nand U29810 (N_29810,N_27875,N_27734);
or U29811 (N_29811,N_26099,N_27170);
nand U29812 (N_29812,N_27212,N_27620);
or U29813 (N_29813,N_27869,N_26972);
nand U29814 (N_29814,N_26795,N_26163);
nor U29815 (N_29815,N_27200,N_27588);
nand U29816 (N_29816,N_27325,N_27914);
xor U29817 (N_29817,N_27438,N_26117);
or U29818 (N_29818,N_27919,N_27346);
or U29819 (N_29819,N_27664,N_26720);
nor U29820 (N_29820,N_27138,N_26309);
nand U29821 (N_29821,N_27795,N_26760);
nand U29822 (N_29822,N_27043,N_27141);
and U29823 (N_29823,N_27815,N_27200);
nor U29824 (N_29824,N_26980,N_27348);
nand U29825 (N_29825,N_27630,N_26411);
nand U29826 (N_29826,N_27490,N_26721);
nand U29827 (N_29827,N_27616,N_27308);
nand U29828 (N_29828,N_26212,N_26480);
nor U29829 (N_29829,N_26839,N_26159);
nand U29830 (N_29830,N_27108,N_26655);
xnor U29831 (N_29831,N_26459,N_26574);
nand U29832 (N_29832,N_27155,N_27529);
and U29833 (N_29833,N_26530,N_26438);
nor U29834 (N_29834,N_27170,N_27896);
and U29835 (N_29835,N_27195,N_27283);
xnor U29836 (N_29836,N_27896,N_27116);
nand U29837 (N_29837,N_27088,N_27971);
nand U29838 (N_29838,N_27568,N_26732);
or U29839 (N_29839,N_26691,N_27351);
xnor U29840 (N_29840,N_27163,N_26482);
nor U29841 (N_29841,N_27077,N_26901);
nand U29842 (N_29842,N_26880,N_26400);
or U29843 (N_29843,N_27816,N_26982);
and U29844 (N_29844,N_27540,N_27636);
and U29845 (N_29845,N_27695,N_26957);
and U29846 (N_29846,N_27372,N_26769);
and U29847 (N_29847,N_27536,N_27912);
or U29848 (N_29848,N_27194,N_26845);
and U29849 (N_29849,N_27615,N_26246);
xnor U29850 (N_29850,N_26697,N_27960);
and U29851 (N_29851,N_26941,N_27821);
nor U29852 (N_29852,N_27633,N_26283);
xnor U29853 (N_29853,N_27944,N_27221);
or U29854 (N_29854,N_26995,N_26886);
nor U29855 (N_29855,N_26001,N_26399);
or U29856 (N_29856,N_27928,N_26247);
and U29857 (N_29857,N_27522,N_27254);
xnor U29858 (N_29858,N_26803,N_27021);
or U29859 (N_29859,N_27928,N_27129);
or U29860 (N_29860,N_26629,N_26736);
or U29861 (N_29861,N_27038,N_26536);
nand U29862 (N_29862,N_27402,N_27666);
nor U29863 (N_29863,N_26711,N_27192);
nor U29864 (N_29864,N_27967,N_26921);
nand U29865 (N_29865,N_26685,N_26566);
or U29866 (N_29866,N_27101,N_26680);
nor U29867 (N_29867,N_27075,N_26566);
and U29868 (N_29868,N_27174,N_27455);
or U29869 (N_29869,N_27271,N_26451);
or U29870 (N_29870,N_27081,N_27849);
nand U29871 (N_29871,N_27392,N_26173);
nand U29872 (N_29872,N_26982,N_27379);
xnor U29873 (N_29873,N_26029,N_27580);
or U29874 (N_29874,N_26381,N_27175);
and U29875 (N_29875,N_27913,N_26457);
xor U29876 (N_29876,N_27910,N_26125);
nor U29877 (N_29877,N_26801,N_27338);
nor U29878 (N_29878,N_27596,N_26880);
nor U29879 (N_29879,N_27379,N_26149);
nor U29880 (N_29880,N_26898,N_27708);
xor U29881 (N_29881,N_27680,N_26859);
and U29882 (N_29882,N_26305,N_26937);
nand U29883 (N_29883,N_26423,N_26143);
and U29884 (N_29884,N_27212,N_26340);
xnor U29885 (N_29885,N_27181,N_26165);
and U29886 (N_29886,N_26520,N_27336);
nor U29887 (N_29887,N_27474,N_26973);
and U29888 (N_29888,N_26649,N_26903);
nand U29889 (N_29889,N_27165,N_27790);
and U29890 (N_29890,N_27305,N_26627);
nand U29891 (N_29891,N_27383,N_26669);
nor U29892 (N_29892,N_27048,N_27468);
and U29893 (N_29893,N_27966,N_26829);
nand U29894 (N_29894,N_27691,N_27085);
and U29895 (N_29895,N_26185,N_27921);
nand U29896 (N_29896,N_26824,N_26868);
nor U29897 (N_29897,N_26481,N_26224);
nand U29898 (N_29898,N_27689,N_26921);
nand U29899 (N_29899,N_26029,N_27523);
and U29900 (N_29900,N_26008,N_26406);
xnor U29901 (N_29901,N_27828,N_27225);
or U29902 (N_29902,N_27361,N_27989);
nand U29903 (N_29903,N_27898,N_27202);
nand U29904 (N_29904,N_26060,N_26371);
or U29905 (N_29905,N_26350,N_26542);
or U29906 (N_29906,N_26416,N_27026);
or U29907 (N_29907,N_27688,N_26135);
and U29908 (N_29908,N_26543,N_27919);
nor U29909 (N_29909,N_27141,N_27653);
or U29910 (N_29910,N_27059,N_26892);
or U29911 (N_29911,N_27935,N_26410);
or U29912 (N_29912,N_26232,N_26003);
nand U29913 (N_29913,N_27992,N_27709);
and U29914 (N_29914,N_27692,N_27572);
xnor U29915 (N_29915,N_27221,N_27117);
xnor U29916 (N_29916,N_26281,N_26806);
and U29917 (N_29917,N_27217,N_26449);
or U29918 (N_29918,N_26203,N_27811);
xnor U29919 (N_29919,N_26533,N_27509);
xor U29920 (N_29920,N_27152,N_26449);
nor U29921 (N_29921,N_26436,N_26536);
xor U29922 (N_29922,N_26848,N_26203);
nor U29923 (N_29923,N_26802,N_26435);
and U29924 (N_29924,N_27570,N_27923);
nand U29925 (N_29925,N_27483,N_27125);
xnor U29926 (N_29926,N_26450,N_26697);
xnor U29927 (N_29927,N_26481,N_26660);
and U29928 (N_29928,N_27099,N_27786);
and U29929 (N_29929,N_27067,N_27308);
and U29930 (N_29930,N_26445,N_26197);
nand U29931 (N_29931,N_27132,N_26992);
and U29932 (N_29932,N_27885,N_27645);
nand U29933 (N_29933,N_27512,N_26440);
or U29934 (N_29934,N_26966,N_27594);
or U29935 (N_29935,N_26595,N_27295);
xor U29936 (N_29936,N_26922,N_26337);
nand U29937 (N_29937,N_27134,N_26689);
nand U29938 (N_29938,N_26866,N_27470);
xnor U29939 (N_29939,N_26456,N_26671);
nand U29940 (N_29940,N_27360,N_27580);
xnor U29941 (N_29941,N_27589,N_27450);
nor U29942 (N_29942,N_26203,N_27760);
or U29943 (N_29943,N_26125,N_26746);
xor U29944 (N_29944,N_26650,N_26278);
nor U29945 (N_29945,N_26105,N_27105);
nand U29946 (N_29946,N_26844,N_27646);
nand U29947 (N_29947,N_27260,N_26181);
xnor U29948 (N_29948,N_26339,N_27676);
nor U29949 (N_29949,N_26919,N_26802);
or U29950 (N_29950,N_27952,N_26942);
xor U29951 (N_29951,N_26963,N_27357);
xor U29952 (N_29952,N_26220,N_27490);
xnor U29953 (N_29953,N_26231,N_27767);
xor U29954 (N_29954,N_26801,N_26532);
xor U29955 (N_29955,N_27662,N_26849);
xnor U29956 (N_29956,N_26970,N_27261);
nand U29957 (N_29957,N_26389,N_27245);
nor U29958 (N_29958,N_26191,N_26907);
nand U29959 (N_29959,N_27586,N_26242);
and U29960 (N_29960,N_27848,N_26911);
or U29961 (N_29961,N_26972,N_27161);
and U29962 (N_29962,N_27048,N_26584);
xor U29963 (N_29963,N_26377,N_26721);
nor U29964 (N_29964,N_26245,N_27442);
xor U29965 (N_29965,N_27747,N_26141);
and U29966 (N_29966,N_27037,N_27605);
and U29967 (N_29967,N_27384,N_26553);
nor U29968 (N_29968,N_26485,N_27065);
and U29969 (N_29969,N_26643,N_27727);
and U29970 (N_29970,N_26505,N_26665);
nand U29971 (N_29971,N_26730,N_27587);
and U29972 (N_29972,N_26287,N_27561);
and U29973 (N_29973,N_26967,N_27530);
or U29974 (N_29974,N_26544,N_26459);
or U29975 (N_29975,N_27519,N_26697);
nor U29976 (N_29976,N_26123,N_26289);
nand U29977 (N_29977,N_26226,N_26842);
and U29978 (N_29978,N_27748,N_27440);
and U29979 (N_29979,N_27222,N_27847);
or U29980 (N_29980,N_27453,N_26683);
or U29981 (N_29981,N_27946,N_27122);
xnor U29982 (N_29982,N_27518,N_27395);
xor U29983 (N_29983,N_27942,N_26704);
nor U29984 (N_29984,N_26014,N_26684);
nand U29985 (N_29985,N_26416,N_26622);
or U29986 (N_29986,N_27397,N_26767);
nor U29987 (N_29987,N_27772,N_27357);
and U29988 (N_29988,N_27326,N_27776);
nor U29989 (N_29989,N_27514,N_27019);
xnor U29990 (N_29990,N_27747,N_27332);
or U29991 (N_29991,N_27196,N_27468);
nand U29992 (N_29992,N_26838,N_26605);
xnor U29993 (N_29993,N_27974,N_27194);
or U29994 (N_29994,N_27260,N_26608);
or U29995 (N_29995,N_26069,N_27611);
and U29996 (N_29996,N_26286,N_27756);
nand U29997 (N_29997,N_26301,N_27646);
or U29998 (N_29998,N_26463,N_26052);
or U29999 (N_29999,N_26945,N_26130);
or UO_0 (O_0,N_29042,N_29863);
nand UO_1 (O_1,N_29309,N_28291);
and UO_2 (O_2,N_29348,N_29623);
nand UO_3 (O_3,N_28327,N_28395);
or UO_4 (O_4,N_29407,N_29932);
or UO_5 (O_5,N_29525,N_28744);
or UO_6 (O_6,N_28606,N_29218);
xnor UO_7 (O_7,N_29220,N_28272);
nor UO_8 (O_8,N_29609,N_28556);
xnor UO_9 (O_9,N_29402,N_29311);
or UO_10 (O_10,N_28234,N_29334);
nand UO_11 (O_11,N_29454,N_28906);
xor UO_12 (O_12,N_29619,N_29360);
nand UO_13 (O_13,N_29099,N_29600);
and UO_14 (O_14,N_29235,N_28146);
and UO_15 (O_15,N_29301,N_29253);
xnor UO_16 (O_16,N_28440,N_28367);
nand UO_17 (O_17,N_29079,N_29989);
nor UO_18 (O_18,N_28654,N_29162);
nor UO_19 (O_19,N_28853,N_28666);
and UO_20 (O_20,N_29438,N_29929);
xnor UO_21 (O_21,N_29138,N_29886);
nand UO_22 (O_22,N_29605,N_28967);
and UO_23 (O_23,N_29261,N_29539);
xnor UO_24 (O_24,N_28060,N_28695);
and UO_25 (O_25,N_28171,N_28577);
and UO_26 (O_26,N_28610,N_28691);
nand UO_27 (O_27,N_29003,N_28715);
nand UO_28 (O_28,N_28878,N_29474);
and UO_29 (O_29,N_29283,N_28549);
nor UO_30 (O_30,N_29233,N_29685);
nor UO_31 (O_31,N_29792,N_29439);
nor UO_32 (O_32,N_29849,N_29114);
nor UO_33 (O_33,N_29538,N_29287);
nor UO_34 (O_34,N_29636,N_29833);
xnor UO_35 (O_35,N_29319,N_28867);
and UO_36 (O_36,N_29304,N_29017);
and UO_37 (O_37,N_29865,N_29071);
or UO_38 (O_38,N_29503,N_28780);
or UO_39 (O_39,N_29483,N_29491);
nand UO_40 (O_40,N_28337,N_28326);
nor UO_41 (O_41,N_29928,N_28576);
nor UO_42 (O_42,N_28965,N_28316);
or UO_43 (O_43,N_28244,N_29655);
xor UO_44 (O_44,N_28584,N_29588);
and UO_45 (O_45,N_29735,N_28685);
or UO_46 (O_46,N_28893,N_28059);
nor UO_47 (O_47,N_29930,N_29453);
and UO_48 (O_48,N_28618,N_28852);
xnor UO_49 (O_49,N_29077,N_28387);
nor UO_50 (O_50,N_28844,N_29761);
or UO_51 (O_51,N_28714,N_28295);
nand UO_52 (O_52,N_28551,N_29194);
and UO_53 (O_53,N_28513,N_28541);
nor UO_54 (O_54,N_29780,N_28493);
and UO_55 (O_55,N_28707,N_29583);
xor UO_56 (O_56,N_29797,N_28939);
and UO_57 (O_57,N_28704,N_28479);
nor UO_58 (O_58,N_28243,N_29812);
nand UO_59 (O_59,N_28616,N_28290);
xor UO_60 (O_60,N_28473,N_29729);
or UO_61 (O_61,N_29034,N_29472);
nor UO_62 (O_62,N_29284,N_29589);
or UO_63 (O_63,N_29405,N_28419);
or UO_64 (O_64,N_29557,N_28001);
or UO_65 (O_65,N_28914,N_28813);
and UO_66 (O_66,N_28548,N_28930);
nand UO_67 (O_67,N_29087,N_28904);
nand UO_68 (O_68,N_29031,N_29744);
nand UO_69 (O_69,N_29248,N_29966);
xnor UO_70 (O_70,N_28846,N_29526);
nand UO_71 (O_71,N_28603,N_29144);
nor UO_72 (O_72,N_28294,N_28038);
xor UO_73 (O_73,N_28518,N_28223);
nor UO_74 (O_74,N_29475,N_28500);
xnor UO_75 (O_75,N_29913,N_28238);
or UO_76 (O_76,N_28094,N_28362);
nor UO_77 (O_77,N_29501,N_29604);
nor UO_78 (O_78,N_29054,N_28894);
xnor UO_79 (O_79,N_28530,N_29924);
and UO_80 (O_80,N_28863,N_29682);
and UO_81 (O_81,N_28206,N_29547);
nor UO_82 (O_82,N_28783,N_29910);
nand UO_83 (O_83,N_29379,N_29452);
xnor UO_84 (O_84,N_29733,N_29070);
or UO_85 (O_85,N_28871,N_29617);
or UO_86 (O_86,N_28035,N_29923);
or UO_87 (O_87,N_28680,N_29393);
nand UO_88 (O_88,N_28850,N_28279);
and UO_89 (O_89,N_29315,N_29188);
nor UO_90 (O_90,N_29982,N_28719);
nor UO_91 (O_91,N_28399,N_28335);
nor UO_92 (O_92,N_28300,N_29414);
or UO_93 (O_93,N_29789,N_28313);
nor UO_94 (O_94,N_29064,N_28683);
nand UO_95 (O_95,N_28127,N_28717);
nand UO_96 (O_96,N_29118,N_29775);
xnor UO_97 (O_97,N_29502,N_28792);
nand UO_98 (O_98,N_28392,N_28420);
nand UO_99 (O_99,N_29081,N_29104);
or UO_100 (O_100,N_29359,N_28946);
or UO_101 (O_101,N_29717,N_28263);
xnor UO_102 (O_102,N_28995,N_28463);
xor UO_103 (O_103,N_28023,N_29920);
nor UO_104 (O_104,N_28802,N_28608);
nor UO_105 (O_105,N_28948,N_28079);
or UO_106 (O_106,N_29339,N_29592);
and UO_107 (O_107,N_28648,N_28653);
and UO_108 (O_108,N_28028,N_29146);
nand UO_109 (O_109,N_28298,N_28321);
xnor UO_110 (O_110,N_28989,N_29460);
and UO_111 (O_111,N_28017,N_29430);
and UO_112 (O_112,N_28828,N_28582);
xor UO_113 (O_113,N_28305,N_29508);
nor UO_114 (O_114,N_28033,N_28255);
nand UO_115 (O_115,N_29317,N_28143);
xor UO_116 (O_116,N_28532,N_28343);
nand UO_117 (O_117,N_28346,N_28815);
or UO_118 (O_118,N_28961,N_28676);
or UO_119 (O_119,N_28614,N_28428);
nand UO_120 (O_120,N_28782,N_29962);
nand UO_121 (O_121,N_28555,N_29570);
xor UO_122 (O_122,N_29521,N_29979);
or UO_123 (O_123,N_29625,N_28120);
or UO_124 (O_124,N_28879,N_29074);
xor UO_125 (O_125,N_28734,N_28843);
xnor UO_126 (O_126,N_29224,N_29116);
xnor UO_127 (O_127,N_28613,N_29613);
nand UO_128 (O_128,N_28988,N_29648);
xor UO_129 (O_129,N_28612,N_29760);
xor UO_130 (O_130,N_28663,N_28916);
xnor UO_131 (O_131,N_29132,N_28202);
nor UO_132 (O_132,N_29062,N_28786);
xnor UO_133 (O_133,N_29545,N_28667);
and UO_134 (O_134,N_28406,N_28553);
xor UO_135 (O_135,N_29963,N_28424);
xor UO_136 (O_136,N_29432,N_28881);
nor UO_137 (O_137,N_29747,N_29773);
or UO_138 (O_138,N_28623,N_28550);
xor UO_139 (O_139,N_29106,N_28566);
or UO_140 (O_140,N_29515,N_28093);
nand UO_141 (O_141,N_28830,N_28960);
xor UO_142 (O_142,N_28086,N_29350);
and UO_143 (O_143,N_28911,N_29902);
nand UO_144 (O_144,N_29927,N_28469);
and UO_145 (O_145,N_29291,N_29415);
xnor UO_146 (O_146,N_28048,N_28776);
xnor UO_147 (O_147,N_28328,N_29282);
or UO_148 (O_148,N_28148,N_28505);
and UO_149 (O_149,N_28250,N_28594);
and UO_150 (O_150,N_29726,N_28448);
xnor UO_151 (O_151,N_29205,N_29170);
nand UO_152 (O_152,N_29462,N_29958);
nand UO_153 (O_153,N_28464,N_28642);
nand UO_154 (O_154,N_28408,N_28798);
xor UO_155 (O_155,N_28465,N_29310);
xnor UO_156 (O_156,N_29043,N_28491);
nor UO_157 (O_157,N_29709,N_28251);
nor UO_158 (O_158,N_28467,N_28742);
xor UO_159 (O_159,N_28753,N_28955);
nor UO_160 (O_160,N_29347,N_28817);
nor UO_161 (O_161,N_28958,N_28882);
xnor UO_162 (O_162,N_28015,N_29829);
nor UO_163 (O_163,N_28746,N_28708);
and UO_164 (O_164,N_28197,N_29548);
nand UO_165 (O_165,N_28103,N_28104);
nor UO_166 (O_166,N_29264,N_29469);
xnor UO_167 (O_167,N_29933,N_29196);
or UO_168 (O_168,N_29791,N_28385);
nor UO_169 (O_169,N_29375,N_28267);
nor UO_170 (O_170,N_28432,N_29703);
nand UO_171 (O_171,N_29968,N_29499);
or UO_172 (O_172,N_28147,N_28884);
nor UO_173 (O_173,N_29954,N_29945);
and UO_174 (O_174,N_29922,N_28917);
xor UO_175 (O_175,N_28745,N_29230);
nor UO_176 (O_176,N_28334,N_28189);
xor UO_177 (O_177,N_28565,N_29739);
nand UO_178 (O_178,N_28230,N_28800);
nor UO_179 (O_179,N_29119,N_29641);
and UO_180 (O_180,N_29399,N_29978);
nor UO_181 (O_181,N_29892,N_29102);
or UO_182 (O_182,N_29243,N_29766);
and UO_183 (O_183,N_29293,N_29810);
nor UO_184 (O_184,N_28311,N_28398);
nand UO_185 (O_185,N_29355,N_28065);
xnor UO_186 (O_186,N_29149,N_29492);
nand UO_187 (O_187,N_29977,N_29326);
and UO_188 (O_188,N_28731,N_28693);
nor UO_189 (O_189,N_28952,N_28055);
xor UO_190 (O_190,N_29630,N_29808);
or UO_191 (O_191,N_29478,N_29436);
nor UO_192 (O_192,N_28677,N_29357);
or UO_193 (O_193,N_29060,N_29518);
or UO_194 (O_194,N_28370,N_29343);
xor UO_195 (O_195,N_28258,N_29671);
or UO_196 (O_196,N_28981,N_28354);
or UO_197 (O_197,N_29085,N_29662);
xor UO_198 (O_198,N_29634,N_29371);
nand UO_199 (O_199,N_29133,N_29616);
nor UO_200 (O_200,N_29562,N_28196);
nor UO_201 (O_201,N_29377,N_28615);
nor UO_202 (O_202,N_29073,N_28456);
nand UO_203 (O_203,N_28444,N_28595);
xor UO_204 (O_204,N_29455,N_28378);
and UO_205 (O_205,N_29909,N_28063);
or UO_206 (O_206,N_29842,N_28322);
xor UO_207 (O_207,N_29160,N_29252);
xnor UO_208 (O_208,N_29354,N_29514);
xnor UO_209 (O_209,N_28159,N_29335);
nor UO_210 (O_210,N_29778,N_29174);
nand UO_211 (O_211,N_29225,N_28791);
nand UO_212 (O_212,N_29649,N_29578);
nand UO_213 (O_213,N_28098,N_29827);
and UO_214 (O_214,N_28301,N_29689);
nor UO_215 (O_215,N_28839,N_28194);
nor UO_216 (O_216,N_29826,N_28203);
nand UO_217 (O_217,N_28052,N_28621);
nor UO_218 (O_218,N_28533,N_29758);
or UO_219 (O_219,N_28212,N_28759);
xor UO_220 (O_220,N_29022,N_29271);
or UO_221 (O_221,N_29496,N_28265);
nand UO_222 (O_222,N_28507,N_28005);
xor UO_223 (O_223,N_29653,N_28178);
nand UO_224 (O_224,N_28993,N_29805);
or UO_225 (O_225,N_29660,N_29896);
nor UO_226 (O_226,N_28087,N_29919);
xnor UO_227 (O_227,N_29900,N_28542);
or UO_228 (O_228,N_29867,N_28716);
nand UO_229 (O_229,N_29782,N_28994);
or UO_230 (O_230,N_29743,N_29516);
and UO_231 (O_231,N_29215,N_28232);
nor UO_232 (O_232,N_28462,N_28264);
nor UO_233 (O_233,N_28150,N_28471);
xnor UO_234 (O_234,N_28942,N_29839);
and UO_235 (O_235,N_29049,N_29723);
or UO_236 (O_236,N_29273,N_28351);
nor UO_237 (O_237,N_29506,N_28635);
nand UO_238 (O_238,N_29051,N_29602);
or UO_239 (O_239,N_29165,N_29817);
xnor UO_240 (O_240,N_29286,N_28389);
nor UO_241 (O_241,N_28137,N_29796);
and UO_242 (O_242,N_28520,N_28587);
or UO_243 (O_243,N_29367,N_29669);
or UO_244 (O_244,N_28900,N_29136);
or UO_245 (O_245,N_29244,N_28283);
nor UO_246 (O_246,N_29100,N_29695);
nand UO_247 (O_247,N_28578,N_29952);
nor UO_248 (O_248,N_28138,N_28651);
and UO_249 (O_249,N_28201,N_28325);
or UO_250 (O_250,N_28669,N_28932);
nor UO_251 (O_251,N_29152,N_28941);
nor UO_252 (O_252,N_28732,N_29524);
nand UO_253 (O_253,N_29195,N_29401);
nor UO_254 (O_254,N_29824,N_28521);
and UO_255 (O_255,N_29258,N_28306);
xor UO_256 (O_256,N_28224,N_28617);
nand UO_257 (O_257,N_29755,N_28276);
or UO_258 (O_258,N_28388,N_29763);
or UO_259 (O_259,N_29056,N_28044);
and UO_260 (O_260,N_28657,N_29332);
nor UO_261 (O_261,N_29970,N_29554);
or UO_262 (O_262,N_29363,N_28278);
xor UO_263 (O_263,N_28236,N_28643);
xnor UO_264 (O_264,N_29127,N_29825);
nand UO_265 (O_265,N_28067,N_29754);
and UO_266 (O_266,N_28910,N_28401);
nand UO_267 (O_267,N_28740,N_29573);
xnor UO_268 (O_268,N_28874,N_29831);
nor UO_269 (O_269,N_28650,N_29096);
xnor UO_270 (O_270,N_29404,N_29358);
and UO_271 (O_271,N_28897,N_29523);
xor UO_272 (O_272,N_29013,N_28253);
or UO_273 (O_273,N_29873,N_28207);
nor UO_274 (O_274,N_28080,N_29765);
and UO_275 (O_275,N_28413,N_29505);
or UO_276 (O_276,N_28484,N_29126);
xor UO_277 (O_277,N_29394,N_28877);
nor UO_278 (O_278,N_28176,N_28849);
nor UO_279 (O_279,N_28811,N_28710);
nor UO_280 (O_280,N_28887,N_29254);
nor UO_281 (O_281,N_29192,N_29059);
xor UO_282 (O_282,N_28854,N_28997);
or UO_283 (O_283,N_28966,N_28826);
nand UO_284 (O_284,N_28356,N_28812);
xor UO_285 (O_285,N_29389,N_29321);
nand UO_286 (O_286,N_29585,N_28105);
nand UO_287 (O_287,N_29352,N_28713);
and UO_288 (O_288,N_28106,N_28488);
nor UO_289 (O_289,N_28240,N_28725);
xor UO_290 (O_290,N_29504,N_28452);
nor UO_291 (O_291,N_29576,N_29659);
and UO_292 (O_292,N_29529,N_28652);
or UO_293 (O_293,N_28135,N_29727);
nor UO_294 (O_294,N_28801,N_29193);
nand UO_295 (O_295,N_29024,N_28529);
nand UO_296 (O_296,N_28115,N_29590);
xor UO_297 (O_297,N_28396,N_28242);
xnor UO_298 (O_298,N_28885,N_29620);
and UO_299 (O_299,N_29901,N_29872);
xor UO_300 (O_300,N_29637,N_28245);
nand UO_301 (O_301,N_28841,N_29877);
xor UO_302 (O_302,N_29214,N_28528);
nor UO_303 (O_303,N_28933,N_29684);
xor UO_304 (O_304,N_29490,N_29368);
xor UO_305 (O_305,N_29058,N_28784);
xnor UO_306 (O_306,N_29818,N_29299);
nor UO_307 (O_307,N_29596,N_28423);
or UO_308 (O_308,N_28282,N_29105);
or UO_309 (O_309,N_29644,N_28477);
or UO_310 (O_310,N_29776,N_28775);
or UO_311 (O_311,N_29316,N_28054);
nand UO_312 (O_312,N_28192,N_28991);
xnor UO_313 (O_313,N_29540,N_28561);
nor UO_314 (O_314,N_28825,N_28547);
or UO_315 (O_315,N_28198,N_28678);
nor UO_316 (O_316,N_28363,N_28156);
or UO_317 (O_317,N_28531,N_28344);
nand UO_318 (O_318,N_29458,N_28002);
nor UO_319 (O_319,N_28437,N_28848);
nor UO_320 (O_320,N_29470,N_28671);
and UO_321 (O_321,N_29388,N_29823);
xnor UO_322 (O_322,N_29172,N_29484);
and UO_323 (O_323,N_29337,N_28497);
or UO_324 (O_324,N_28117,N_28043);
or UO_325 (O_325,N_28478,N_28199);
and UO_326 (O_326,N_28690,N_28050);
or UO_327 (O_327,N_29240,N_28053);
and UO_328 (O_328,N_28524,N_29026);
and UO_329 (O_329,N_29038,N_29510);
nand UO_330 (O_330,N_29365,N_28414);
and UO_331 (O_331,N_28797,N_28233);
xor UO_332 (O_332,N_28943,N_28366);
nor UO_333 (O_333,N_29300,N_29779);
and UO_334 (O_334,N_28774,N_29467);
nand UO_335 (O_335,N_28768,N_28987);
and UO_336 (O_336,N_28949,N_28831);
and UO_337 (O_337,N_28645,N_29292);
or UO_338 (O_338,N_28140,N_28624);
nand UO_339 (O_339,N_28758,N_29719);
nor UO_340 (O_340,N_29822,N_29772);
and UO_341 (O_341,N_28472,N_28421);
or UO_342 (O_342,N_29075,N_28358);
nand UO_343 (O_343,N_28636,N_29323);
nand UO_344 (O_344,N_29905,N_29040);
xor UO_345 (O_345,N_29612,N_29687);
nand UO_346 (O_346,N_28673,N_29329);
nand UO_347 (O_347,N_29028,N_28959);
or UO_348 (O_348,N_28284,N_28110);
nand UO_349 (O_349,N_28903,N_29686);
nor UO_350 (O_350,N_28229,N_28163);
xor UO_351 (O_351,N_29956,N_29520);
or UO_352 (O_352,N_29180,N_28922);
and UO_353 (O_353,N_28186,N_29171);
xnor UO_354 (O_354,N_28173,N_29771);
or UO_355 (O_355,N_28286,N_28895);
and UO_356 (O_356,N_29567,N_29880);
or UO_357 (O_357,N_29495,N_29147);
or UO_358 (O_358,N_29848,N_28179);
and UO_359 (O_359,N_28345,N_29800);
xor UO_360 (O_360,N_28803,N_29851);
or UO_361 (O_361,N_28963,N_28633);
nor UO_362 (O_362,N_29306,N_28468);
xor UO_363 (O_363,N_29429,N_28701);
and UO_364 (O_364,N_28056,N_29876);
nor UO_365 (O_365,N_28976,N_28481);
nand UO_366 (O_366,N_28751,N_28489);
nor UO_367 (O_367,N_28220,N_29698);
and UO_368 (O_368,N_29883,N_28969);
xnor UO_369 (O_369,N_28409,N_28495);
xor UO_370 (O_370,N_28888,N_28076);
xnor UO_371 (O_371,N_28402,N_28269);
nand UO_372 (O_372,N_28304,N_28332);
nand UO_373 (O_373,N_29092,N_29904);
nor UO_374 (O_374,N_28482,N_29450);
or UO_375 (O_375,N_29611,N_28604);
and UO_376 (O_376,N_29618,N_29858);
and UO_377 (O_377,N_28747,N_28441);
and UO_378 (O_378,N_28376,N_28307);
xnor UO_379 (O_379,N_29471,N_28915);
or UO_380 (O_380,N_28560,N_29298);
and UO_381 (O_381,N_29015,N_29084);
xor UO_382 (O_382,N_29097,N_28934);
or UO_383 (O_383,N_29094,N_28051);
nor UO_384 (O_384,N_29090,N_28902);
or UO_385 (O_385,N_29276,N_29652);
or UO_386 (O_386,N_28563,N_29181);
or UO_387 (O_387,N_28804,N_29445);
xor UO_388 (O_388,N_28384,N_29221);
or UO_389 (O_389,N_29828,N_29639);
nand UO_390 (O_390,N_28552,N_28905);
or UO_391 (O_391,N_29724,N_29236);
nor UO_392 (O_392,N_29312,N_29112);
nand UO_393 (O_393,N_29738,N_29005);
xor UO_394 (O_394,N_28820,N_28501);
xnor UO_395 (O_395,N_28208,N_28318);
and UO_396 (O_396,N_28217,N_28866);
xor UO_397 (O_397,N_29037,N_29362);
xor UO_398 (O_398,N_28235,N_29860);
xnor UO_399 (O_399,N_28296,N_29908);
xor UO_400 (O_400,N_29869,N_28446);
and UO_401 (O_401,N_28891,N_28091);
or UO_402 (O_402,N_29658,N_28085);
or UO_403 (O_403,N_29121,N_28153);
nor UO_404 (O_404,N_29412,N_28703);
nand UO_405 (O_405,N_28601,N_29678);
xor UO_406 (O_406,N_28656,N_28368);
nand UO_407 (O_407,N_29535,N_28090);
nor UO_408 (O_408,N_28697,N_28040);
xnor UO_409 (O_409,N_28779,N_29597);
nand UO_410 (O_410,N_29663,N_28570);
nor UO_411 (O_411,N_28069,N_28084);
nor UO_412 (O_412,N_29210,N_29615);
xnor UO_413 (O_413,N_29995,N_29036);
xor UO_414 (O_414,N_28686,N_28899);
or UO_415 (O_415,N_28840,N_28749);
nor UO_416 (O_416,N_29400,N_29975);
nor UO_417 (O_417,N_29798,N_28664);
xnor UO_418 (O_418,N_28324,N_28730);
nand UO_419 (O_419,N_29342,N_29030);
nand UO_420 (O_420,N_29866,N_28720);
and UO_421 (O_421,N_28634,N_29461);
or UO_422 (O_422,N_29943,N_29307);
nand UO_423 (O_423,N_29333,N_28241);
nand UO_424 (O_424,N_28519,N_28609);
nand UO_425 (O_425,N_28918,N_29448);
or UO_426 (O_426,N_28036,N_29594);
nand UO_427 (O_427,N_28757,N_29941);
or UO_428 (O_428,N_29198,N_28886);
nand UO_429 (O_429,N_28277,N_28761);
or UO_430 (O_430,N_28246,N_28266);
and UO_431 (O_431,N_29980,N_28750);
and UO_432 (O_432,N_28926,N_29318);
or UO_433 (O_433,N_29891,N_28107);
nand UO_434 (O_434,N_28458,N_29476);
nor UO_435 (O_435,N_29785,N_28502);
or UO_436 (O_436,N_29178,N_28858);
xor UO_437 (O_437,N_29790,N_29753);
and UO_438 (O_438,N_29752,N_29341);
or UO_439 (O_439,N_28169,N_29008);
xnor UO_440 (O_440,N_29878,N_29494);
xor UO_441 (O_441,N_28436,N_28485);
and UO_442 (O_442,N_28131,N_28130);
xnor UO_443 (O_443,N_29057,N_29257);
or UO_444 (O_444,N_28573,N_29991);
nor UO_445 (O_445,N_28598,N_28494);
nor UO_446 (O_446,N_29123,N_28681);
or UO_447 (O_447,N_29420,N_28487);
or UO_448 (O_448,N_29561,N_29821);
xor UO_449 (O_449,N_29314,N_29629);
and UO_450 (O_450,N_28517,N_28581);
xnor UO_451 (O_451,N_29964,N_28861);
or UO_452 (O_452,N_29973,N_29706);
xor UO_453 (O_453,N_28962,N_28509);
nor UO_454 (O_454,N_29632,N_29794);
nand UO_455 (O_455,N_29227,N_29921);
nor UO_456 (O_456,N_28834,N_28459);
nand UO_457 (O_457,N_29732,N_28213);
xor UO_458 (O_458,N_28205,N_28661);
xor UO_459 (O_459,N_29546,N_28836);
nor UO_460 (O_460,N_29197,N_29640);
nor UO_461 (O_461,N_28096,N_29199);
xnor UO_462 (O_462,N_29907,N_28214);
and UO_463 (O_463,N_28360,N_29345);
or UO_464 (O_464,N_29251,N_29606);
nor UO_465 (O_465,N_29571,N_28964);
and UO_466 (O_466,N_29131,N_29338);
xnor UO_467 (O_467,N_28257,N_29937);
and UO_468 (O_468,N_28544,N_28929);
and UO_469 (O_469,N_29696,N_28134);
nor UO_470 (O_470,N_29422,N_29534);
xor UO_471 (O_471,N_28030,N_29841);
and UO_472 (O_472,N_28377,N_28559);
nor UO_473 (O_473,N_29113,N_28694);
nand UO_474 (O_474,N_29736,N_29268);
or UO_475 (O_475,N_28219,N_28927);
nor UO_476 (O_476,N_29558,N_29093);
or UO_477 (O_477,N_29107,N_28514);
or UO_478 (O_478,N_29710,N_29801);
nor UO_479 (O_479,N_28386,N_28416);
nand UO_480 (O_480,N_28496,N_28262);
xnor UO_481 (O_481,N_28992,N_28014);
and UO_482 (O_482,N_29544,N_29497);
nor UO_483 (O_483,N_29322,N_29574);
nor UO_484 (O_484,N_28457,N_29053);
or UO_485 (O_485,N_29527,N_28515);
nor UO_486 (O_486,N_28350,N_28215);
nand UO_487 (O_487,N_29289,N_28029);
and UO_488 (O_488,N_28429,N_29681);
nor UO_489 (O_489,N_28543,N_29018);
xor UO_490 (O_490,N_29173,N_28193);
nor UO_491 (O_491,N_28764,N_29898);
xor UO_492 (O_492,N_29418,N_29917);
nor UO_493 (O_493,N_28270,N_28799);
and UO_494 (O_494,N_28047,N_29346);
or UO_495 (O_495,N_28081,N_29382);
nand UO_496 (O_496,N_28151,N_29482);
and UO_497 (O_497,N_28982,N_29938);
and UO_498 (O_498,N_28089,N_28600);
and UO_499 (O_499,N_28728,N_28268);
xor UO_500 (O_500,N_28870,N_29749);
or UO_501 (O_501,N_29269,N_28102);
xnor UO_502 (O_502,N_29517,N_28032);
xnor UO_503 (O_503,N_28736,N_29331);
and UO_504 (O_504,N_29325,N_28928);
nor UO_505 (O_505,N_28699,N_29656);
or UO_506 (O_506,N_29751,N_28170);
nor UO_507 (O_507,N_29349,N_28859);
or UO_508 (O_508,N_29434,N_29320);
nand UO_509 (O_509,N_28718,N_29239);
nand UO_510 (O_510,N_28596,N_29950);
or UO_511 (O_511,N_29485,N_28639);
and UO_512 (O_512,N_29313,N_28415);
or UO_513 (O_513,N_29156,N_29683);
xor UO_514 (O_514,N_29290,N_28188);
nor UO_515 (O_515,N_28508,N_29881);
or UO_516 (O_516,N_28185,N_28068);
nand UO_517 (O_517,N_29522,N_29627);
xnor UO_518 (O_518,N_28455,N_29039);
and UO_519 (O_519,N_28302,N_28944);
and UO_520 (O_520,N_28380,N_29598);
and UO_521 (O_521,N_29409,N_29232);
nand UO_522 (O_522,N_29046,N_29427);
xor UO_523 (O_523,N_29424,N_29072);
nand UO_524 (O_524,N_28591,N_29167);
and UO_525 (O_525,N_29820,N_28810);
nor UO_526 (O_526,N_29993,N_29575);
xnor UO_527 (O_527,N_29512,N_28074);
and UO_528 (O_528,N_29294,N_28097);
and UO_529 (O_529,N_29128,N_29076);
xor UO_530 (O_530,N_29871,N_28034);
nand UO_531 (O_531,N_29148,N_29774);
or UO_532 (O_532,N_29741,N_28675);
and UO_533 (O_533,N_28752,N_29542);
or UO_534 (O_534,N_28696,N_28195);
xnor UO_535 (O_535,N_28923,N_29721);
or UO_536 (O_536,N_28778,N_28771);
xnor UO_537 (O_537,N_29874,N_28862);
xor UO_538 (O_538,N_28453,N_29050);
xnor UO_539 (O_539,N_28644,N_29120);
xor UO_540 (O_540,N_28114,N_29944);
and UO_541 (O_541,N_28795,N_28312);
or UO_542 (O_542,N_29440,N_29177);
and UO_543 (O_543,N_28748,N_29336);
nand UO_544 (O_544,N_29700,N_28788);
nand UO_545 (O_545,N_28909,N_28516);
and UO_546 (O_546,N_28379,N_28041);
and UO_547 (O_547,N_29925,N_28483);
nor UO_548 (O_548,N_28249,N_28020);
and UO_549 (O_549,N_29125,N_28434);
or UO_550 (O_550,N_28222,N_29456);
and UO_551 (O_551,N_29748,N_28504);
nand UO_552 (O_552,N_29137,N_29708);
nor UO_553 (O_553,N_28709,N_28141);
and UO_554 (O_554,N_28200,N_29643);
xor UO_555 (O_555,N_28892,N_28510);
or UO_556 (O_556,N_29940,N_29552);
nand UO_557 (O_557,N_28355,N_28924);
and UO_558 (O_558,N_28721,N_28239);
nor UO_559 (O_559,N_29553,N_29903);
nor UO_560 (O_560,N_29231,N_29155);
xor UO_561 (O_561,N_28738,N_29403);
and UO_562 (O_562,N_28225,N_28338);
nand UO_563 (O_563,N_28535,N_29443);
nand UO_564 (O_564,N_28308,N_28772);
nand UO_565 (O_565,N_28474,N_28781);
nand UO_566 (O_566,N_29946,N_28299);
xnor UO_567 (O_567,N_29324,N_29151);
and UO_568 (O_568,N_29117,N_29895);
and UO_569 (O_569,N_28564,N_28129);
nor UO_570 (O_570,N_29651,N_29396);
nor UO_571 (O_571,N_28004,N_28095);
xor UO_572 (O_572,N_29182,N_29089);
xor UO_573 (O_573,N_28537,N_28625);
xnor UO_574 (O_574,N_29124,N_29530);
nand UO_575 (O_575,N_29209,N_28297);
nand UO_576 (O_576,N_28058,N_29769);
and UO_577 (O_577,N_29260,N_28637);
xor UO_578 (O_578,N_28540,N_29280);
nor UO_579 (O_579,N_29983,N_28756);
nor UO_580 (O_580,N_29032,N_29158);
nand UO_581 (O_581,N_29041,N_28273);
or UO_582 (O_582,N_29387,N_28412);
nand UO_583 (O_583,N_28818,N_29002);
nor UO_584 (O_584,N_28369,N_29985);
and UO_585 (O_585,N_29247,N_28868);
nand UO_586 (O_586,N_29098,N_29931);
xor UO_587 (O_587,N_28741,N_29212);
xor UO_588 (O_588,N_29433,N_28417);
xor UO_589 (O_589,N_29654,N_29384);
and UO_590 (O_590,N_29163,N_29411);
nor UO_591 (O_591,N_28875,N_28160);
nor UO_592 (O_592,N_28972,N_29000);
and UO_593 (O_593,N_29463,N_29237);
nor UO_594 (O_594,N_28340,N_29447);
nand UO_595 (O_595,N_28777,N_29423);
nand UO_596 (O_596,N_29421,N_29560);
xnor UO_597 (O_597,N_28706,N_28228);
xor UO_598 (O_598,N_28954,N_28364);
and UO_599 (O_599,N_29374,N_28733);
nor UO_600 (O_600,N_28218,N_28702);
xor UO_601 (O_601,N_28352,N_29067);
xnor UO_602 (O_602,N_28737,N_29555);
or UO_603 (O_603,N_29713,N_28021);
nand UO_604 (O_604,N_28400,N_29513);
nand UO_605 (O_605,N_29216,N_29419);
nor UO_606 (O_606,N_28816,N_28983);
or UO_607 (O_607,N_29226,N_29249);
nand UO_608 (O_608,N_29836,N_28790);
nand UO_609 (O_609,N_29303,N_29256);
nor UO_610 (O_610,N_28789,N_28630);
or UO_611 (O_611,N_29777,N_29795);
and UO_612 (O_612,N_29672,N_29272);
and UO_613 (O_613,N_29595,N_29971);
nor UO_614 (O_614,N_29489,N_29912);
and UO_615 (O_615,N_29987,N_29122);
nor UO_616 (O_616,N_28599,N_29859);
and UO_617 (O_617,N_29001,N_28018);
nand UO_618 (O_618,N_28167,N_29330);
and UO_619 (O_619,N_29431,N_29211);
xor UO_620 (O_620,N_29045,N_28546);
nand UO_621 (O_621,N_29016,N_28970);
nor UO_622 (O_622,N_28700,N_29020);
nand UO_623 (O_623,N_29705,N_29788);
nor UO_624 (O_624,N_29819,N_29141);
xnor UO_625 (O_625,N_28342,N_28112);
and UO_626 (O_626,N_29187,N_29459);
and UO_627 (O_627,N_29191,N_28128);
and UO_628 (O_628,N_28088,N_28373);
xor UO_629 (O_629,N_29014,N_29756);
or UO_630 (O_630,N_29697,N_28712);
or UO_631 (O_631,N_28427,N_29241);
nand UO_632 (O_632,N_28449,N_28289);
or UO_633 (O_633,N_28330,N_28631);
or UO_634 (O_634,N_29340,N_29111);
or UO_635 (O_635,N_29386,N_28049);
nor UO_636 (O_636,N_29278,N_29480);
xor UO_637 (O_637,N_28123,N_29894);
xor UO_638 (O_638,N_28442,N_28064);
nand UO_639 (O_639,N_28980,N_28288);
nand UO_640 (O_640,N_29392,N_28433);
nor UO_641 (O_641,N_28026,N_29992);
and UO_642 (O_642,N_28211,N_29897);
and UO_643 (O_643,N_29101,N_28259);
or UO_644 (O_644,N_29444,N_29843);
and UO_645 (O_645,N_28315,N_28209);
and UO_646 (O_646,N_29887,N_29487);
nor UO_647 (O_647,N_28538,N_28628);
xor UO_648 (O_648,N_29250,N_29029);
xnor UO_649 (O_649,N_28814,N_28957);
xnor UO_650 (O_650,N_29296,N_29972);
or UO_651 (O_651,N_29129,N_29961);
xnor UO_652 (O_652,N_29899,N_29864);
xnor UO_653 (O_653,N_29569,N_28860);
and UO_654 (O_654,N_29680,N_28216);
xor UO_655 (O_655,N_28506,N_29376);
or UO_656 (O_656,N_29219,N_29228);
or UO_657 (O_657,N_28357,N_29862);
or UO_658 (O_658,N_28498,N_29203);
and UO_659 (O_659,N_28646,N_29047);
nand UO_660 (O_660,N_29344,N_29457);
nand UO_661 (O_661,N_28951,N_29308);
nor UO_662 (O_662,N_28404,N_29691);
or UO_663 (O_663,N_28808,N_28118);
and UO_664 (O_664,N_28375,N_28365);
nand UO_665 (O_665,N_29500,N_28231);
nand UO_666 (O_666,N_29677,N_29066);
xor UO_667 (O_667,N_29807,N_28883);
or UO_668 (O_668,N_29638,N_28562);
or UO_669 (O_669,N_28760,N_28641);
or UO_670 (O_670,N_29890,N_28793);
nand UO_671 (O_671,N_29201,N_28727);
nand UO_672 (O_672,N_29591,N_28705);
and UO_673 (O_673,N_29665,N_28688);
xor UO_674 (O_674,N_28066,N_28499);
nor UO_675 (O_675,N_29157,N_29061);
or UO_676 (O_676,N_28381,N_28592);
nor UO_677 (O_677,N_28953,N_28590);
and UO_678 (O_678,N_29728,N_29302);
and UO_679 (O_679,N_28602,N_29486);
or UO_680 (O_680,N_29647,N_28027);
nand UO_681 (O_681,N_29607,N_29207);
nor UO_682 (O_682,N_28142,N_28136);
nand UO_683 (O_683,N_29981,N_29095);
nand UO_684 (O_684,N_28461,N_28687);
or UO_685 (O_685,N_28374,N_29327);
nand UO_686 (O_686,N_28431,N_29217);
xnor UO_687 (O_687,N_29531,N_29185);
nand UO_688 (O_688,N_29134,N_28925);
nand UO_689 (O_689,N_29926,N_29670);
or UO_690 (O_690,N_28122,N_29949);
or UO_691 (O_691,N_28568,N_29441);
nor UO_692 (O_692,N_28372,N_29145);
nand UO_693 (O_693,N_28155,N_29953);
nand UO_694 (O_694,N_29911,N_29245);
or UO_695 (O_695,N_28190,N_28013);
nor UO_696 (O_696,N_29783,N_29850);
nor UO_697 (O_697,N_28046,N_29498);
xor UO_698 (O_698,N_28674,N_28287);
xnor UO_699 (O_699,N_29614,N_29857);
xnor UO_700 (O_700,N_28682,N_28523);
and UO_701 (O_701,N_28672,N_28796);
nand UO_702 (O_702,N_28016,N_28739);
or UO_703 (O_703,N_28006,N_29947);
xor UO_704 (O_704,N_29395,N_29391);
xnor UO_705 (O_705,N_28348,N_29222);
xnor UO_706 (O_706,N_28670,N_28985);
nand UO_707 (O_707,N_28938,N_29610);
and UO_708 (O_708,N_29229,N_28397);
nand UO_709 (O_709,N_29955,N_28503);
nand UO_710 (O_710,N_28655,N_29601);
nand UO_711 (O_711,N_28293,N_29835);
or UO_712 (O_712,N_28785,N_29110);
and UO_713 (O_713,N_29803,N_29563);
and UO_714 (O_714,N_28856,N_28567);
nand UO_715 (O_715,N_29711,N_29010);
nor UO_716 (O_716,N_29238,N_29369);
or UO_717 (O_717,N_29967,N_29948);
and UO_718 (O_718,N_29200,N_29666);
and UO_719 (O_719,N_29275,N_28165);
xor UO_720 (O_720,N_28154,N_29168);
and UO_721 (O_721,N_29694,N_28100);
and UO_722 (O_722,N_29661,N_28443);
xnor UO_723 (O_723,N_28658,N_29701);
and UO_724 (O_724,N_29577,N_28445);
and UO_725 (O_725,N_28569,N_28583);
nand UO_726 (O_726,N_28574,N_29572);
xnor UO_727 (O_727,N_28124,N_29628);
and UO_728 (O_728,N_29852,N_28057);
or UO_729 (O_729,N_28755,N_29715);
and UO_730 (O_730,N_28937,N_28629);
nand UO_731 (O_731,N_29740,N_29465);
xor UO_732 (O_732,N_28986,N_28640);
and UO_733 (O_733,N_28931,N_29893);
or UO_734 (O_734,N_28857,N_28113);
xnor UO_735 (O_735,N_28945,N_29398);
nand UO_736 (O_736,N_29650,N_29550);
xor UO_737 (O_737,N_28184,N_28724);
or UO_738 (O_738,N_29288,N_29722);
xor UO_739 (O_739,N_28492,N_28025);
or UO_740 (O_740,N_28126,N_29426);
nor UO_741 (O_741,N_28072,N_29135);
and UO_742 (O_742,N_28835,N_29048);
or UO_743 (O_743,N_28075,N_28323);
or UO_744 (O_744,N_29668,N_29608);
nand UO_745 (O_745,N_28261,N_29673);
xnor UO_746 (O_746,N_29731,N_29078);
or UO_747 (O_747,N_29587,N_28580);
nor UO_748 (O_748,N_29762,N_29781);
nor UO_749 (O_749,N_29861,N_28872);
nor UO_750 (O_750,N_28019,N_29080);
nor UO_751 (O_751,N_28158,N_29556);
nand UO_752 (O_752,N_28558,N_28766);
xor UO_753 (O_753,N_29353,N_28605);
and UO_754 (O_754,N_29383,N_28070);
and UO_755 (O_755,N_28947,N_29366);
and UO_756 (O_756,N_28393,N_28331);
and UO_757 (O_757,N_28990,N_28806);
xor UO_758 (O_758,N_28082,N_29477);
xor UO_759 (O_759,N_28319,N_28144);
nand UO_760 (O_760,N_29488,N_28407);
or UO_761 (O_761,N_29270,N_28936);
and UO_762 (O_762,N_29809,N_29184);
and UO_763 (O_763,N_29543,N_28819);
xnor UO_764 (O_764,N_28394,N_29186);
nand UO_765 (O_765,N_29208,N_29768);
nor UO_766 (O_766,N_29759,N_28092);
xor UO_767 (O_767,N_29885,N_28317);
xor UO_768 (O_768,N_28978,N_28274);
or UO_769 (O_769,N_28554,N_28626);
xor UO_770 (O_770,N_28827,N_29990);
and UO_771 (O_771,N_29868,N_28480);
xnor UO_772 (O_772,N_29568,N_28638);
or UO_773 (O_773,N_28078,N_28765);
xnor UO_774 (O_774,N_28837,N_28008);
or UO_775 (O_775,N_28204,N_29918);
or UO_776 (O_776,N_29297,N_28622);
xor UO_777 (O_777,N_29770,N_29541);
xor UO_778 (O_778,N_28526,N_29044);
or UO_779 (O_779,N_29951,N_29579);
and UO_780 (O_780,N_28182,N_29664);
or UO_781 (O_781,N_29875,N_29816);
xor UO_782 (O_782,N_28743,N_29844);
nand UO_783 (O_783,N_28009,N_28042);
or UO_784 (O_784,N_29380,N_29939);
nor UO_785 (O_785,N_28996,N_28898);
or UO_786 (O_786,N_29266,N_28157);
nand UO_787 (O_787,N_29473,N_29787);
xnor UO_788 (O_788,N_29262,N_29166);
or UO_789 (O_789,N_28347,N_29027);
xnor UO_790 (O_790,N_28794,N_29830);
or UO_791 (O_791,N_28698,N_29468);
and UO_792 (O_792,N_28821,N_28175);
nand UO_793 (O_793,N_29140,N_29784);
or UO_794 (O_794,N_29507,N_29870);
or UO_795 (O_795,N_29802,N_29189);
nand UO_796 (O_796,N_28907,N_28121);
nor UO_797 (O_797,N_28833,N_28876);
xnor UO_798 (O_798,N_28773,N_28227);
nor UO_799 (O_799,N_29511,N_28956);
or UO_800 (O_800,N_28486,N_29631);
and UO_801 (O_801,N_29793,N_29159);
nor UO_802 (O_802,N_29882,N_29692);
or UO_803 (O_803,N_28162,N_28024);
nor UO_804 (O_804,N_29328,N_29957);
nor UO_805 (O_805,N_29969,N_29019);
xnor UO_806 (O_806,N_29464,N_28039);
and UO_807 (O_807,N_28588,N_29372);
nor UO_808 (O_808,N_28285,N_28940);
nor UO_809 (O_809,N_28083,N_29718);
nand UO_810 (O_810,N_29734,N_28252);
xor UO_811 (O_811,N_29856,N_28684);
and UO_812 (O_812,N_28534,N_29451);
or UO_813 (O_813,N_29549,N_28998);
and UO_814 (O_814,N_29764,N_28880);
nand UO_815 (O_815,N_28139,N_28984);
nand UO_816 (O_816,N_28585,N_29914);
xor UO_817 (O_817,N_29139,N_29234);
and UO_818 (O_818,N_29804,N_29626);
nand UO_819 (O_819,N_29581,N_29091);
nor UO_820 (O_820,N_29811,N_28770);
or UO_821 (O_821,N_29679,N_28527);
nor UO_822 (O_822,N_29410,N_29437);
nor UO_823 (O_823,N_28896,N_28061);
nor UO_824 (O_824,N_28168,N_28425);
or UO_825 (O_825,N_28133,N_29767);
xnor UO_826 (O_826,N_29378,N_29425);
or UO_827 (O_827,N_29150,N_28280);
xor UO_828 (O_828,N_29088,N_28062);
nor UO_829 (O_829,N_28460,N_28571);
nor UO_830 (O_830,N_28920,N_28807);
and UO_831 (O_831,N_28116,N_29737);
nor UO_832 (O_832,N_28586,N_28824);
nand UO_833 (O_833,N_29675,N_28271);
or UO_834 (O_834,N_29063,N_29645);
xor UO_835 (O_835,N_28383,N_28627);
xor UO_836 (O_836,N_29202,N_29559);
and UO_837 (O_837,N_28426,N_28405);
or UO_838 (O_838,N_29204,N_29255);
nand UO_839 (O_839,N_28226,N_28152);
nand UO_840 (O_840,N_29279,N_29840);
nor UO_841 (O_841,N_28187,N_29052);
and UO_842 (O_842,N_29274,N_28303);
and UO_843 (O_843,N_29988,N_28979);
and UO_844 (O_844,N_28975,N_29190);
or UO_845 (O_845,N_29730,N_29974);
or UO_846 (O_846,N_29888,N_29381);
and UO_847 (O_847,N_29164,N_28172);
nand UO_848 (O_848,N_28132,N_29033);
nand UO_849 (O_849,N_29479,N_29536);
nor UO_850 (O_850,N_28145,N_29021);
nor UO_851 (O_851,N_29693,N_29942);
xor UO_852 (O_852,N_29621,N_29109);
nand UO_853 (O_853,N_28829,N_29667);
nor UO_854 (O_854,N_29725,N_29082);
nand UO_855 (O_855,N_28281,N_29277);
or UO_856 (O_856,N_29707,N_28901);
nor UO_857 (O_857,N_28973,N_28855);
nand UO_858 (O_858,N_28071,N_29532);
nand UO_859 (O_859,N_29845,N_29069);
nor UO_860 (O_860,N_28254,N_28000);
and UO_861 (O_861,N_28908,N_29356);
or UO_862 (O_862,N_29175,N_29806);
or UO_863 (O_863,N_29011,N_29757);
and UO_864 (O_864,N_28912,N_28310);
nand UO_865 (O_865,N_29103,N_28632);
nand UO_866 (O_866,N_28403,N_28525);
xor UO_867 (O_867,N_28762,N_29086);
nand UO_868 (O_868,N_28692,N_28919);
nand UO_869 (O_869,N_29712,N_28099);
nor UO_870 (O_870,N_29259,N_28309);
nand UO_871 (O_871,N_28247,N_29143);
and UO_872 (O_872,N_29242,N_28864);
nor UO_873 (O_873,N_28805,N_29603);
xor UO_874 (O_874,N_29565,N_29936);
nor UO_875 (O_875,N_28575,N_28022);
nor UO_876 (O_876,N_29832,N_28177);
nand UO_877 (O_877,N_29361,N_29390);
nor UO_878 (O_878,N_29976,N_29994);
xor UO_879 (O_879,N_28611,N_28689);
nor UO_880 (O_880,N_28410,N_29004);
nand UO_881 (O_881,N_28557,N_29704);
or UO_882 (O_882,N_29142,N_28823);
or UO_883 (O_883,N_29959,N_29635);
nor UO_884 (O_884,N_29622,N_29179);
or UO_885 (O_885,N_28256,N_29012);
and UO_886 (O_886,N_28191,N_29223);
and UO_887 (O_887,N_29351,N_28111);
xor UO_888 (O_888,N_29714,N_29646);
xnor UO_889 (O_889,N_29023,N_28522);
xor UO_890 (O_890,N_29566,N_28977);
xnor UO_891 (O_891,N_28422,N_29688);
xnor UO_892 (O_892,N_29035,N_28619);
and UO_893 (O_893,N_28769,N_29385);
nand UO_894 (O_894,N_28174,N_28073);
or UO_895 (O_895,N_28735,N_29584);
nand UO_896 (O_896,N_28660,N_28974);
xor UO_897 (O_897,N_28418,N_29847);
and UO_898 (O_898,N_28649,N_29624);
xor UO_899 (O_899,N_28320,N_28314);
or UO_900 (O_900,N_28722,N_28662);
or UO_901 (O_901,N_29906,N_28339);
xor UO_902 (O_902,N_29593,N_29493);
xnor UO_903 (O_903,N_28037,N_28999);
or UO_904 (O_904,N_28822,N_29884);
and UO_905 (O_905,N_29206,N_29986);
or UO_906 (O_906,N_28729,N_28371);
or UO_907 (O_907,N_28869,N_29855);
xnor UO_908 (O_908,N_29853,N_29481);
nor UO_909 (O_909,N_29537,N_28971);
or UO_910 (O_910,N_28329,N_29055);
and UO_911 (O_911,N_28435,N_29373);
and UO_912 (O_912,N_28545,N_28851);
nand UO_913 (O_913,N_29998,N_28210);
or UO_914 (O_914,N_28164,N_29997);
xor UO_915 (O_915,N_28361,N_28010);
xor UO_916 (O_916,N_28767,N_29154);
or UO_917 (O_917,N_29633,N_28838);
or UO_918 (O_918,N_29934,N_28382);
nor UO_919 (O_919,N_28447,N_28101);
or UO_920 (O_920,N_28031,N_28607);
nor UO_921 (O_921,N_28349,N_29213);
and UO_922 (O_922,N_29996,N_28183);
and UO_923 (O_923,N_29449,N_29176);
xor UO_924 (O_924,N_28511,N_28539);
xor UO_925 (O_925,N_28333,N_28475);
or UO_926 (O_926,N_28572,N_29674);
or UO_927 (O_927,N_28390,N_28873);
nor UO_928 (O_928,N_29435,N_29813);
xor UO_929 (O_929,N_28921,N_29406);
nor UO_930 (O_930,N_29295,N_28754);
xnor UO_931 (O_931,N_29551,N_28221);
and UO_932 (O_932,N_28620,N_29364);
nand UO_933 (O_933,N_28012,N_28470);
or UO_934 (O_934,N_29130,N_29281);
and UO_935 (O_935,N_28353,N_28341);
xor UO_936 (O_936,N_29786,N_29657);
and UO_937 (O_937,N_28476,N_28439);
and UO_938 (O_938,N_29442,N_29580);
or UO_939 (O_939,N_29564,N_28275);
and UO_940 (O_940,N_28890,N_28125);
xor UO_941 (O_941,N_28411,N_28149);
and UO_942 (O_942,N_28119,N_28007);
or UO_943 (O_943,N_28166,N_29838);
nand UO_944 (O_944,N_28336,N_29446);
nor UO_945 (O_945,N_29416,N_29984);
nand UO_946 (O_946,N_29676,N_29916);
and UO_947 (O_947,N_29509,N_29879);
nor UO_948 (O_948,N_29417,N_29750);
nand UO_949 (O_949,N_28787,N_28809);
nor UO_950 (O_950,N_29115,N_28248);
xor UO_951 (O_951,N_28536,N_28593);
xor UO_952 (O_952,N_28391,N_29746);
xnor UO_953 (O_953,N_29169,N_29742);
nor UO_954 (O_954,N_29702,N_29533);
xor UO_955 (O_955,N_28109,N_28597);
xnor UO_956 (O_956,N_28832,N_29161);
nand UO_957 (O_957,N_28045,N_29068);
and UO_958 (O_958,N_29413,N_28450);
or UO_959 (O_959,N_29599,N_29246);
or UO_960 (O_960,N_28108,N_28430);
xor UO_961 (O_961,N_28451,N_29799);
nor UO_962 (O_962,N_29083,N_28847);
and UO_963 (O_963,N_28668,N_29837);
nor UO_964 (O_964,N_28842,N_28726);
and UO_965 (O_965,N_28579,N_29889);
nor UO_966 (O_966,N_28935,N_29960);
nand UO_967 (O_967,N_28659,N_29935);
or UO_968 (O_968,N_29999,N_29267);
or UO_969 (O_969,N_29690,N_28260);
and UO_970 (O_970,N_28003,N_28889);
xor UO_971 (O_971,N_28180,N_29834);
and UO_972 (O_972,N_29915,N_29519);
nor UO_973 (O_973,N_28589,N_28950);
xnor UO_974 (O_974,N_29263,N_29466);
or UO_975 (O_975,N_28865,N_29699);
nor UO_976 (O_976,N_29108,N_28011);
xor UO_977 (O_977,N_29716,N_28647);
nand UO_978 (O_978,N_29965,N_28913);
nand UO_979 (O_979,N_28490,N_29397);
nand UO_980 (O_980,N_28723,N_29025);
or UO_981 (O_981,N_28763,N_29183);
nor UO_982 (O_982,N_28968,N_29009);
nor UO_983 (O_983,N_28512,N_28845);
nand UO_984 (O_984,N_28181,N_29153);
and UO_985 (O_985,N_29720,N_29586);
nand UO_986 (O_986,N_28711,N_29642);
xor UO_987 (O_987,N_29814,N_29815);
nand UO_988 (O_988,N_29305,N_28454);
nor UO_989 (O_989,N_28237,N_29428);
nand UO_990 (O_990,N_29846,N_29006);
and UO_991 (O_991,N_28438,N_28665);
and UO_992 (O_992,N_29854,N_29745);
nor UO_993 (O_993,N_29265,N_29065);
nor UO_994 (O_994,N_28466,N_28077);
and UO_995 (O_995,N_28161,N_28292);
and UO_996 (O_996,N_29408,N_29285);
nand UO_997 (O_997,N_29007,N_28679);
and UO_998 (O_998,N_29370,N_28359);
xor UO_999 (O_999,N_29528,N_29582);
or UO_1000 (O_1000,N_28182,N_28757);
nor UO_1001 (O_1001,N_28407,N_29399);
nor UO_1002 (O_1002,N_28109,N_28552);
or UO_1003 (O_1003,N_29849,N_28498);
xor UO_1004 (O_1004,N_28278,N_28125);
and UO_1005 (O_1005,N_29060,N_28660);
xor UO_1006 (O_1006,N_28984,N_29562);
nor UO_1007 (O_1007,N_28618,N_28496);
and UO_1008 (O_1008,N_28013,N_29842);
xor UO_1009 (O_1009,N_29160,N_28972);
and UO_1010 (O_1010,N_29893,N_28676);
or UO_1011 (O_1011,N_29563,N_28419);
xor UO_1012 (O_1012,N_29473,N_28651);
nand UO_1013 (O_1013,N_28714,N_28023);
or UO_1014 (O_1014,N_29601,N_28045);
nand UO_1015 (O_1015,N_29959,N_29561);
xnor UO_1016 (O_1016,N_29274,N_28108);
nor UO_1017 (O_1017,N_28078,N_29202);
nand UO_1018 (O_1018,N_29795,N_29194);
xnor UO_1019 (O_1019,N_28756,N_29659);
and UO_1020 (O_1020,N_29294,N_28231);
and UO_1021 (O_1021,N_28379,N_28754);
or UO_1022 (O_1022,N_29601,N_29825);
or UO_1023 (O_1023,N_28850,N_28005);
xor UO_1024 (O_1024,N_28970,N_29522);
nor UO_1025 (O_1025,N_28190,N_28167);
and UO_1026 (O_1026,N_29837,N_29430);
nand UO_1027 (O_1027,N_29324,N_28844);
nor UO_1028 (O_1028,N_28187,N_29236);
or UO_1029 (O_1029,N_29581,N_28557);
or UO_1030 (O_1030,N_29102,N_28014);
and UO_1031 (O_1031,N_28993,N_29794);
nand UO_1032 (O_1032,N_28461,N_28684);
xor UO_1033 (O_1033,N_29196,N_29469);
nor UO_1034 (O_1034,N_29670,N_28161);
or UO_1035 (O_1035,N_29570,N_29116);
or UO_1036 (O_1036,N_28474,N_29022);
nand UO_1037 (O_1037,N_28881,N_29509);
nor UO_1038 (O_1038,N_29502,N_28327);
and UO_1039 (O_1039,N_28315,N_29929);
and UO_1040 (O_1040,N_29431,N_29171);
nor UO_1041 (O_1041,N_29393,N_29902);
or UO_1042 (O_1042,N_28874,N_28193);
and UO_1043 (O_1043,N_28196,N_29198);
nor UO_1044 (O_1044,N_28564,N_28577);
nand UO_1045 (O_1045,N_29929,N_28276);
nand UO_1046 (O_1046,N_29769,N_28523);
nor UO_1047 (O_1047,N_28146,N_29875);
and UO_1048 (O_1048,N_28757,N_28401);
nand UO_1049 (O_1049,N_29132,N_28605);
nor UO_1050 (O_1050,N_28917,N_28244);
nand UO_1051 (O_1051,N_28309,N_29297);
and UO_1052 (O_1052,N_28777,N_28754);
nand UO_1053 (O_1053,N_28825,N_29417);
nor UO_1054 (O_1054,N_28840,N_29503);
and UO_1055 (O_1055,N_29779,N_29231);
nand UO_1056 (O_1056,N_28967,N_28115);
and UO_1057 (O_1057,N_28825,N_28743);
nand UO_1058 (O_1058,N_29166,N_29088);
or UO_1059 (O_1059,N_29565,N_29852);
nor UO_1060 (O_1060,N_28210,N_28867);
nand UO_1061 (O_1061,N_29210,N_28178);
and UO_1062 (O_1062,N_29113,N_29194);
xnor UO_1063 (O_1063,N_29805,N_28724);
nor UO_1064 (O_1064,N_29000,N_28338);
nand UO_1065 (O_1065,N_28806,N_28509);
nand UO_1066 (O_1066,N_29591,N_28653);
nor UO_1067 (O_1067,N_29135,N_29492);
or UO_1068 (O_1068,N_28177,N_28157);
xnor UO_1069 (O_1069,N_28594,N_29073);
and UO_1070 (O_1070,N_29513,N_29841);
nor UO_1071 (O_1071,N_28893,N_29310);
and UO_1072 (O_1072,N_29998,N_29262);
and UO_1073 (O_1073,N_28348,N_28626);
nand UO_1074 (O_1074,N_29237,N_29792);
nor UO_1075 (O_1075,N_29986,N_29449);
nor UO_1076 (O_1076,N_28100,N_28352);
or UO_1077 (O_1077,N_29079,N_29539);
and UO_1078 (O_1078,N_28220,N_28769);
xnor UO_1079 (O_1079,N_29325,N_29003);
nor UO_1080 (O_1080,N_28234,N_29380);
or UO_1081 (O_1081,N_29587,N_29523);
xor UO_1082 (O_1082,N_29739,N_29585);
nor UO_1083 (O_1083,N_29900,N_28558);
or UO_1084 (O_1084,N_28051,N_28413);
or UO_1085 (O_1085,N_28800,N_29654);
or UO_1086 (O_1086,N_28825,N_29600);
and UO_1087 (O_1087,N_29679,N_28690);
nor UO_1088 (O_1088,N_29304,N_28345);
nor UO_1089 (O_1089,N_28410,N_28950);
or UO_1090 (O_1090,N_28024,N_28305);
xor UO_1091 (O_1091,N_29329,N_28757);
nor UO_1092 (O_1092,N_28123,N_28420);
nand UO_1093 (O_1093,N_29532,N_29267);
or UO_1094 (O_1094,N_28459,N_28702);
and UO_1095 (O_1095,N_29596,N_29493);
or UO_1096 (O_1096,N_29613,N_29850);
nor UO_1097 (O_1097,N_28718,N_29198);
or UO_1098 (O_1098,N_29468,N_29704);
nor UO_1099 (O_1099,N_29848,N_28145);
xor UO_1100 (O_1100,N_29592,N_28804);
or UO_1101 (O_1101,N_28432,N_29917);
xnor UO_1102 (O_1102,N_29791,N_29440);
or UO_1103 (O_1103,N_29652,N_29385);
and UO_1104 (O_1104,N_29582,N_28962);
nand UO_1105 (O_1105,N_29438,N_28795);
or UO_1106 (O_1106,N_29149,N_28498);
nor UO_1107 (O_1107,N_29608,N_28820);
nand UO_1108 (O_1108,N_28837,N_29177);
and UO_1109 (O_1109,N_29687,N_29581);
nor UO_1110 (O_1110,N_29408,N_29412);
or UO_1111 (O_1111,N_29441,N_29848);
and UO_1112 (O_1112,N_28587,N_29852);
nand UO_1113 (O_1113,N_29290,N_29044);
nand UO_1114 (O_1114,N_28244,N_28094);
nand UO_1115 (O_1115,N_29920,N_28367);
xnor UO_1116 (O_1116,N_28765,N_29947);
xnor UO_1117 (O_1117,N_28015,N_29272);
nor UO_1118 (O_1118,N_29009,N_28200);
xor UO_1119 (O_1119,N_29716,N_29718);
nand UO_1120 (O_1120,N_29603,N_29397);
nand UO_1121 (O_1121,N_28189,N_29971);
nand UO_1122 (O_1122,N_29890,N_29171);
nand UO_1123 (O_1123,N_29824,N_29454);
nand UO_1124 (O_1124,N_29663,N_29892);
nand UO_1125 (O_1125,N_28962,N_28154);
or UO_1126 (O_1126,N_28858,N_28341);
or UO_1127 (O_1127,N_29423,N_29373);
nor UO_1128 (O_1128,N_29657,N_29828);
nand UO_1129 (O_1129,N_28818,N_29945);
xor UO_1130 (O_1130,N_29296,N_29607);
or UO_1131 (O_1131,N_28316,N_28346);
or UO_1132 (O_1132,N_29905,N_28822);
nor UO_1133 (O_1133,N_28046,N_29489);
and UO_1134 (O_1134,N_29637,N_29184);
xnor UO_1135 (O_1135,N_29510,N_28396);
or UO_1136 (O_1136,N_29777,N_29485);
nand UO_1137 (O_1137,N_28269,N_29135);
nor UO_1138 (O_1138,N_29574,N_28859);
and UO_1139 (O_1139,N_28414,N_28942);
xnor UO_1140 (O_1140,N_28508,N_29505);
or UO_1141 (O_1141,N_28356,N_29375);
and UO_1142 (O_1142,N_29673,N_28385);
and UO_1143 (O_1143,N_29646,N_29213);
xnor UO_1144 (O_1144,N_29792,N_29846);
nand UO_1145 (O_1145,N_29435,N_29891);
and UO_1146 (O_1146,N_29157,N_28458);
nand UO_1147 (O_1147,N_28758,N_28234);
nor UO_1148 (O_1148,N_29178,N_29042);
nand UO_1149 (O_1149,N_28901,N_29839);
and UO_1150 (O_1150,N_28870,N_28781);
nand UO_1151 (O_1151,N_29189,N_29370);
and UO_1152 (O_1152,N_29607,N_29539);
nand UO_1153 (O_1153,N_29931,N_29644);
xor UO_1154 (O_1154,N_29439,N_28452);
xor UO_1155 (O_1155,N_29862,N_29898);
xnor UO_1156 (O_1156,N_28754,N_29861);
or UO_1157 (O_1157,N_29663,N_28438);
xor UO_1158 (O_1158,N_28377,N_29005);
nor UO_1159 (O_1159,N_28786,N_29162);
xor UO_1160 (O_1160,N_29659,N_28193);
or UO_1161 (O_1161,N_28774,N_28237);
or UO_1162 (O_1162,N_28275,N_29027);
xnor UO_1163 (O_1163,N_28626,N_28291);
xnor UO_1164 (O_1164,N_29692,N_28498);
nor UO_1165 (O_1165,N_28543,N_29545);
or UO_1166 (O_1166,N_29924,N_28556);
and UO_1167 (O_1167,N_29882,N_29753);
or UO_1168 (O_1168,N_29075,N_28264);
nor UO_1169 (O_1169,N_29070,N_28230);
or UO_1170 (O_1170,N_28717,N_28910);
nand UO_1171 (O_1171,N_29950,N_29854);
and UO_1172 (O_1172,N_29011,N_29945);
nor UO_1173 (O_1173,N_28057,N_28417);
nand UO_1174 (O_1174,N_28379,N_28868);
nor UO_1175 (O_1175,N_28998,N_28670);
or UO_1176 (O_1176,N_28584,N_28237);
or UO_1177 (O_1177,N_29201,N_28402);
nor UO_1178 (O_1178,N_29776,N_28611);
and UO_1179 (O_1179,N_28649,N_29277);
or UO_1180 (O_1180,N_29932,N_28499);
nand UO_1181 (O_1181,N_28032,N_29266);
and UO_1182 (O_1182,N_29419,N_28210);
or UO_1183 (O_1183,N_29804,N_28723);
xnor UO_1184 (O_1184,N_28874,N_29328);
xnor UO_1185 (O_1185,N_29813,N_28584);
or UO_1186 (O_1186,N_29670,N_29239);
nand UO_1187 (O_1187,N_29796,N_29579);
or UO_1188 (O_1188,N_28334,N_28483);
nand UO_1189 (O_1189,N_29267,N_28167);
and UO_1190 (O_1190,N_28544,N_29332);
xnor UO_1191 (O_1191,N_28909,N_29528);
and UO_1192 (O_1192,N_29986,N_29519);
nor UO_1193 (O_1193,N_29806,N_29471);
or UO_1194 (O_1194,N_28560,N_28282);
nand UO_1195 (O_1195,N_29086,N_28318);
xnor UO_1196 (O_1196,N_29654,N_28759);
xnor UO_1197 (O_1197,N_29984,N_28902);
nor UO_1198 (O_1198,N_29862,N_28673);
or UO_1199 (O_1199,N_29369,N_29746);
or UO_1200 (O_1200,N_28142,N_28810);
nor UO_1201 (O_1201,N_29884,N_28244);
nor UO_1202 (O_1202,N_29898,N_29524);
nor UO_1203 (O_1203,N_29042,N_29389);
nand UO_1204 (O_1204,N_28231,N_29062);
nand UO_1205 (O_1205,N_28667,N_29774);
xnor UO_1206 (O_1206,N_29666,N_28183);
or UO_1207 (O_1207,N_28784,N_28837);
or UO_1208 (O_1208,N_28409,N_28537);
xnor UO_1209 (O_1209,N_29418,N_28725);
and UO_1210 (O_1210,N_29738,N_28058);
xor UO_1211 (O_1211,N_28224,N_29524);
nor UO_1212 (O_1212,N_28858,N_28386);
and UO_1213 (O_1213,N_29656,N_29778);
nand UO_1214 (O_1214,N_29663,N_28264);
xnor UO_1215 (O_1215,N_29109,N_29239);
nor UO_1216 (O_1216,N_28925,N_28977);
and UO_1217 (O_1217,N_28282,N_28620);
nor UO_1218 (O_1218,N_29172,N_29938);
nand UO_1219 (O_1219,N_29547,N_28002);
xnor UO_1220 (O_1220,N_28324,N_28528);
nand UO_1221 (O_1221,N_29143,N_28165);
nor UO_1222 (O_1222,N_28478,N_29870);
or UO_1223 (O_1223,N_28682,N_28760);
nor UO_1224 (O_1224,N_29032,N_29744);
nor UO_1225 (O_1225,N_29331,N_28301);
nor UO_1226 (O_1226,N_28054,N_28326);
nand UO_1227 (O_1227,N_28997,N_28182);
and UO_1228 (O_1228,N_28977,N_28015);
or UO_1229 (O_1229,N_29824,N_29785);
xor UO_1230 (O_1230,N_28691,N_29222);
or UO_1231 (O_1231,N_28952,N_28784);
or UO_1232 (O_1232,N_28304,N_28828);
nor UO_1233 (O_1233,N_28607,N_29634);
and UO_1234 (O_1234,N_28050,N_29375);
xnor UO_1235 (O_1235,N_29384,N_28313);
or UO_1236 (O_1236,N_29732,N_28798);
or UO_1237 (O_1237,N_28435,N_29198);
or UO_1238 (O_1238,N_29136,N_28745);
xnor UO_1239 (O_1239,N_29637,N_28381);
and UO_1240 (O_1240,N_29516,N_28443);
and UO_1241 (O_1241,N_29928,N_28222);
and UO_1242 (O_1242,N_29870,N_29911);
or UO_1243 (O_1243,N_29710,N_28565);
xnor UO_1244 (O_1244,N_29734,N_29075);
nor UO_1245 (O_1245,N_28351,N_28879);
or UO_1246 (O_1246,N_28196,N_29599);
nor UO_1247 (O_1247,N_28760,N_29705);
nand UO_1248 (O_1248,N_28361,N_29306);
xnor UO_1249 (O_1249,N_28693,N_28920);
and UO_1250 (O_1250,N_28254,N_29167);
xor UO_1251 (O_1251,N_28443,N_28323);
xor UO_1252 (O_1252,N_28399,N_28766);
nor UO_1253 (O_1253,N_29876,N_28414);
or UO_1254 (O_1254,N_29930,N_28793);
and UO_1255 (O_1255,N_29152,N_29343);
nor UO_1256 (O_1256,N_28437,N_29258);
nand UO_1257 (O_1257,N_28379,N_28560);
and UO_1258 (O_1258,N_28221,N_28825);
nand UO_1259 (O_1259,N_28314,N_29790);
nor UO_1260 (O_1260,N_29278,N_29018);
and UO_1261 (O_1261,N_28716,N_29474);
nand UO_1262 (O_1262,N_29181,N_28936);
xor UO_1263 (O_1263,N_29395,N_28725);
or UO_1264 (O_1264,N_28439,N_28208);
nand UO_1265 (O_1265,N_28171,N_29883);
nand UO_1266 (O_1266,N_28181,N_28681);
and UO_1267 (O_1267,N_29383,N_28685);
and UO_1268 (O_1268,N_29277,N_29589);
xnor UO_1269 (O_1269,N_28366,N_28899);
xor UO_1270 (O_1270,N_29932,N_29408);
nor UO_1271 (O_1271,N_28344,N_28145);
nand UO_1272 (O_1272,N_28664,N_29258);
or UO_1273 (O_1273,N_28874,N_28602);
nand UO_1274 (O_1274,N_29921,N_28058);
nor UO_1275 (O_1275,N_29291,N_29224);
xnor UO_1276 (O_1276,N_29690,N_29724);
or UO_1277 (O_1277,N_28798,N_28278);
or UO_1278 (O_1278,N_29737,N_28228);
and UO_1279 (O_1279,N_28876,N_28008);
and UO_1280 (O_1280,N_28198,N_28861);
and UO_1281 (O_1281,N_28063,N_29826);
or UO_1282 (O_1282,N_28384,N_28976);
nand UO_1283 (O_1283,N_29921,N_28981);
nor UO_1284 (O_1284,N_29965,N_29052);
xor UO_1285 (O_1285,N_29426,N_29098);
nor UO_1286 (O_1286,N_29987,N_28567);
xor UO_1287 (O_1287,N_29765,N_28038);
and UO_1288 (O_1288,N_29165,N_29948);
nand UO_1289 (O_1289,N_29407,N_28154);
xnor UO_1290 (O_1290,N_28867,N_29801);
or UO_1291 (O_1291,N_28273,N_28251);
and UO_1292 (O_1292,N_28726,N_29549);
or UO_1293 (O_1293,N_29891,N_29532);
nand UO_1294 (O_1294,N_28344,N_29646);
xor UO_1295 (O_1295,N_28991,N_28078);
and UO_1296 (O_1296,N_28894,N_28826);
nor UO_1297 (O_1297,N_28967,N_29101);
xnor UO_1298 (O_1298,N_28791,N_29270);
and UO_1299 (O_1299,N_28092,N_28260);
nor UO_1300 (O_1300,N_29286,N_29604);
nand UO_1301 (O_1301,N_29667,N_28924);
or UO_1302 (O_1302,N_28392,N_29507);
and UO_1303 (O_1303,N_28481,N_28867);
nor UO_1304 (O_1304,N_28405,N_28756);
and UO_1305 (O_1305,N_29933,N_28331);
xor UO_1306 (O_1306,N_29087,N_29634);
and UO_1307 (O_1307,N_29426,N_29774);
nor UO_1308 (O_1308,N_29271,N_28624);
nand UO_1309 (O_1309,N_28509,N_29873);
or UO_1310 (O_1310,N_29391,N_29029);
or UO_1311 (O_1311,N_28572,N_28211);
nor UO_1312 (O_1312,N_28195,N_28105);
or UO_1313 (O_1313,N_28779,N_29433);
or UO_1314 (O_1314,N_29293,N_28756);
or UO_1315 (O_1315,N_28295,N_29931);
nor UO_1316 (O_1316,N_28750,N_29947);
or UO_1317 (O_1317,N_28759,N_29174);
xor UO_1318 (O_1318,N_29852,N_29372);
nor UO_1319 (O_1319,N_29985,N_29015);
nand UO_1320 (O_1320,N_28457,N_28085);
and UO_1321 (O_1321,N_29018,N_29727);
nor UO_1322 (O_1322,N_29991,N_29301);
or UO_1323 (O_1323,N_29289,N_29805);
and UO_1324 (O_1324,N_29945,N_29997);
nand UO_1325 (O_1325,N_28356,N_29496);
or UO_1326 (O_1326,N_29238,N_29595);
and UO_1327 (O_1327,N_28308,N_29931);
nor UO_1328 (O_1328,N_28189,N_29923);
nand UO_1329 (O_1329,N_29924,N_29096);
or UO_1330 (O_1330,N_28024,N_28425);
and UO_1331 (O_1331,N_29138,N_28708);
and UO_1332 (O_1332,N_28807,N_29369);
and UO_1333 (O_1333,N_29880,N_28189);
nor UO_1334 (O_1334,N_29432,N_29049);
xor UO_1335 (O_1335,N_28322,N_29661);
nand UO_1336 (O_1336,N_29992,N_28883);
xor UO_1337 (O_1337,N_29856,N_29767);
xnor UO_1338 (O_1338,N_28458,N_28049);
nor UO_1339 (O_1339,N_28784,N_28551);
and UO_1340 (O_1340,N_29567,N_28554);
xnor UO_1341 (O_1341,N_29387,N_28843);
or UO_1342 (O_1342,N_28247,N_28235);
nor UO_1343 (O_1343,N_28316,N_29127);
nor UO_1344 (O_1344,N_29799,N_29499);
xor UO_1345 (O_1345,N_29783,N_28773);
or UO_1346 (O_1346,N_28568,N_28946);
and UO_1347 (O_1347,N_29538,N_28125);
nand UO_1348 (O_1348,N_28074,N_28013);
and UO_1349 (O_1349,N_29704,N_28870);
nand UO_1350 (O_1350,N_29574,N_29326);
nor UO_1351 (O_1351,N_29858,N_28834);
and UO_1352 (O_1352,N_28241,N_29709);
xor UO_1353 (O_1353,N_28815,N_29830);
xnor UO_1354 (O_1354,N_29904,N_28659);
nor UO_1355 (O_1355,N_29807,N_28751);
xnor UO_1356 (O_1356,N_28190,N_29219);
xor UO_1357 (O_1357,N_29950,N_28721);
nand UO_1358 (O_1358,N_28626,N_29502);
xor UO_1359 (O_1359,N_28616,N_29074);
nor UO_1360 (O_1360,N_29180,N_28900);
nor UO_1361 (O_1361,N_29276,N_28196);
xnor UO_1362 (O_1362,N_29491,N_28473);
nand UO_1363 (O_1363,N_29292,N_28455);
or UO_1364 (O_1364,N_28590,N_29755);
or UO_1365 (O_1365,N_29267,N_29411);
or UO_1366 (O_1366,N_28341,N_29525);
nor UO_1367 (O_1367,N_29250,N_28880);
nor UO_1368 (O_1368,N_29073,N_28475);
and UO_1369 (O_1369,N_29948,N_28298);
xnor UO_1370 (O_1370,N_29802,N_28580);
nand UO_1371 (O_1371,N_28881,N_29007);
xor UO_1372 (O_1372,N_28017,N_29339);
nand UO_1373 (O_1373,N_28841,N_29066);
nor UO_1374 (O_1374,N_29981,N_29531);
and UO_1375 (O_1375,N_28251,N_28970);
and UO_1376 (O_1376,N_28413,N_29389);
nor UO_1377 (O_1377,N_29717,N_28215);
xor UO_1378 (O_1378,N_29839,N_29358);
nor UO_1379 (O_1379,N_29673,N_28324);
nand UO_1380 (O_1380,N_28100,N_28676);
xor UO_1381 (O_1381,N_28980,N_28930);
nand UO_1382 (O_1382,N_29816,N_29053);
xnor UO_1383 (O_1383,N_29785,N_28797);
nand UO_1384 (O_1384,N_29289,N_28863);
or UO_1385 (O_1385,N_28912,N_29802);
nand UO_1386 (O_1386,N_29939,N_28462);
xor UO_1387 (O_1387,N_29227,N_28315);
nand UO_1388 (O_1388,N_28970,N_29864);
nor UO_1389 (O_1389,N_28840,N_29422);
nand UO_1390 (O_1390,N_28960,N_28164);
nand UO_1391 (O_1391,N_28163,N_29925);
nor UO_1392 (O_1392,N_29001,N_28130);
or UO_1393 (O_1393,N_28641,N_29150);
or UO_1394 (O_1394,N_29070,N_28830);
nand UO_1395 (O_1395,N_28171,N_28368);
xor UO_1396 (O_1396,N_28736,N_29705);
or UO_1397 (O_1397,N_28585,N_28376);
nor UO_1398 (O_1398,N_28852,N_28931);
or UO_1399 (O_1399,N_28080,N_28634);
xor UO_1400 (O_1400,N_28243,N_29175);
nor UO_1401 (O_1401,N_28663,N_29318);
xor UO_1402 (O_1402,N_28234,N_29441);
and UO_1403 (O_1403,N_29300,N_28961);
nand UO_1404 (O_1404,N_29266,N_29461);
nand UO_1405 (O_1405,N_29496,N_28173);
or UO_1406 (O_1406,N_29741,N_28316);
nand UO_1407 (O_1407,N_28396,N_29689);
and UO_1408 (O_1408,N_29831,N_29225);
and UO_1409 (O_1409,N_28477,N_29769);
nand UO_1410 (O_1410,N_29826,N_28955);
xor UO_1411 (O_1411,N_28875,N_28980);
and UO_1412 (O_1412,N_28269,N_29514);
and UO_1413 (O_1413,N_29904,N_29587);
xnor UO_1414 (O_1414,N_28059,N_28977);
xnor UO_1415 (O_1415,N_29120,N_28513);
or UO_1416 (O_1416,N_29171,N_29312);
nor UO_1417 (O_1417,N_28223,N_29711);
nand UO_1418 (O_1418,N_28407,N_29543);
and UO_1419 (O_1419,N_28348,N_28792);
and UO_1420 (O_1420,N_29892,N_29960);
nand UO_1421 (O_1421,N_29171,N_29159);
xnor UO_1422 (O_1422,N_28096,N_28703);
xnor UO_1423 (O_1423,N_29682,N_29341);
or UO_1424 (O_1424,N_28269,N_29027);
xnor UO_1425 (O_1425,N_28734,N_28228);
nor UO_1426 (O_1426,N_29147,N_28197);
and UO_1427 (O_1427,N_29335,N_29146);
nor UO_1428 (O_1428,N_28523,N_29864);
and UO_1429 (O_1429,N_29229,N_28761);
nand UO_1430 (O_1430,N_29608,N_28527);
and UO_1431 (O_1431,N_28180,N_28578);
nor UO_1432 (O_1432,N_28633,N_28734);
or UO_1433 (O_1433,N_29839,N_28455);
nand UO_1434 (O_1434,N_29377,N_29824);
nor UO_1435 (O_1435,N_29798,N_29869);
nand UO_1436 (O_1436,N_28934,N_29719);
nand UO_1437 (O_1437,N_29095,N_29416);
xor UO_1438 (O_1438,N_28009,N_28966);
nand UO_1439 (O_1439,N_28990,N_29681);
and UO_1440 (O_1440,N_29880,N_28871);
and UO_1441 (O_1441,N_29236,N_28060);
nand UO_1442 (O_1442,N_29169,N_28211);
xnor UO_1443 (O_1443,N_28832,N_28348);
xnor UO_1444 (O_1444,N_28872,N_29400);
or UO_1445 (O_1445,N_29434,N_29978);
nor UO_1446 (O_1446,N_29936,N_28728);
nor UO_1447 (O_1447,N_29327,N_28858);
xnor UO_1448 (O_1448,N_29553,N_28086);
nor UO_1449 (O_1449,N_28329,N_28223);
and UO_1450 (O_1450,N_28002,N_28352);
and UO_1451 (O_1451,N_29751,N_29363);
nand UO_1452 (O_1452,N_29388,N_28938);
nand UO_1453 (O_1453,N_29338,N_28298);
or UO_1454 (O_1454,N_28259,N_28023);
or UO_1455 (O_1455,N_28256,N_29709);
nor UO_1456 (O_1456,N_28927,N_28838);
xnor UO_1457 (O_1457,N_29541,N_28656);
xor UO_1458 (O_1458,N_29450,N_28883);
xor UO_1459 (O_1459,N_28281,N_29548);
xnor UO_1460 (O_1460,N_28244,N_28896);
or UO_1461 (O_1461,N_29601,N_28343);
nor UO_1462 (O_1462,N_29256,N_29013);
and UO_1463 (O_1463,N_28217,N_28752);
or UO_1464 (O_1464,N_28853,N_29978);
nand UO_1465 (O_1465,N_28542,N_29835);
or UO_1466 (O_1466,N_28838,N_28680);
nor UO_1467 (O_1467,N_28956,N_28346);
xor UO_1468 (O_1468,N_29839,N_28350);
nand UO_1469 (O_1469,N_29559,N_28101);
xnor UO_1470 (O_1470,N_28619,N_29637);
or UO_1471 (O_1471,N_28929,N_28973);
and UO_1472 (O_1472,N_28271,N_28054);
xor UO_1473 (O_1473,N_28351,N_28923);
and UO_1474 (O_1474,N_29046,N_29587);
nor UO_1475 (O_1475,N_29328,N_28539);
xor UO_1476 (O_1476,N_28479,N_28437);
nand UO_1477 (O_1477,N_28380,N_29923);
nand UO_1478 (O_1478,N_28342,N_29154);
xor UO_1479 (O_1479,N_29000,N_29401);
and UO_1480 (O_1480,N_28576,N_28012);
or UO_1481 (O_1481,N_28139,N_28330);
nand UO_1482 (O_1482,N_29650,N_28710);
and UO_1483 (O_1483,N_28587,N_29942);
xor UO_1484 (O_1484,N_29753,N_28853);
xnor UO_1485 (O_1485,N_29509,N_29323);
and UO_1486 (O_1486,N_28661,N_29340);
and UO_1487 (O_1487,N_28834,N_28440);
nor UO_1488 (O_1488,N_28323,N_29846);
or UO_1489 (O_1489,N_28990,N_28420);
and UO_1490 (O_1490,N_28662,N_28484);
xnor UO_1491 (O_1491,N_29286,N_29522);
or UO_1492 (O_1492,N_29073,N_29383);
and UO_1493 (O_1493,N_28247,N_29245);
and UO_1494 (O_1494,N_29027,N_29938);
nor UO_1495 (O_1495,N_29851,N_29484);
or UO_1496 (O_1496,N_28832,N_29255);
nor UO_1497 (O_1497,N_29104,N_29743);
nand UO_1498 (O_1498,N_28464,N_29405);
and UO_1499 (O_1499,N_28371,N_29726);
xnor UO_1500 (O_1500,N_29421,N_28177);
nor UO_1501 (O_1501,N_29116,N_29222);
or UO_1502 (O_1502,N_29975,N_28871);
or UO_1503 (O_1503,N_29047,N_28403);
nor UO_1504 (O_1504,N_28184,N_29838);
or UO_1505 (O_1505,N_28674,N_28435);
nor UO_1506 (O_1506,N_29801,N_28082);
nand UO_1507 (O_1507,N_29142,N_28058);
or UO_1508 (O_1508,N_29155,N_28483);
and UO_1509 (O_1509,N_29583,N_28849);
xnor UO_1510 (O_1510,N_29566,N_28395);
nor UO_1511 (O_1511,N_29964,N_29458);
xnor UO_1512 (O_1512,N_29908,N_29071);
nor UO_1513 (O_1513,N_28257,N_28246);
or UO_1514 (O_1514,N_28671,N_29614);
and UO_1515 (O_1515,N_29894,N_29879);
and UO_1516 (O_1516,N_28790,N_29539);
nand UO_1517 (O_1517,N_28775,N_28174);
nor UO_1518 (O_1518,N_28569,N_29767);
nor UO_1519 (O_1519,N_29150,N_29737);
xor UO_1520 (O_1520,N_28680,N_29666);
nor UO_1521 (O_1521,N_29128,N_28382);
or UO_1522 (O_1522,N_28144,N_28404);
nor UO_1523 (O_1523,N_29203,N_28398);
nor UO_1524 (O_1524,N_29507,N_28003);
xnor UO_1525 (O_1525,N_29737,N_29724);
or UO_1526 (O_1526,N_28884,N_29187);
nand UO_1527 (O_1527,N_28598,N_29424);
xnor UO_1528 (O_1528,N_29964,N_29571);
nand UO_1529 (O_1529,N_28123,N_28943);
nand UO_1530 (O_1530,N_28805,N_28635);
nor UO_1531 (O_1531,N_28945,N_28578);
and UO_1532 (O_1532,N_29437,N_29439);
nor UO_1533 (O_1533,N_29922,N_29221);
and UO_1534 (O_1534,N_29542,N_28956);
xor UO_1535 (O_1535,N_29104,N_28801);
nor UO_1536 (O_1536,N_28778,N_29867);
nand UO_1537 (O_1537,N_28881,N_28909);
or UO_1538 (O_1538,N_29041,N_29345);
nand UO_1539 (O_1539,N_29197,N_28409);
or UO_1540 (O_1540,N_28183,N_29437);
nand UO_1541 (O_1541,N_28884,N_29494);
nor UO_1542 (O_1542,N_28280,N_29419);
or UO_1543 (O_1543,N_29141,N_28892);
and UO_1544 (O_1544,N_29385,N_28195);
nor UO_1545 (O_1545,N_28271,N_29589);
and UO_1546 (O_1546,N_29009,N_28264);
and UO_1547 (O_1547,N_29599,N_28612);
xnor UO_1548 (O_1548,N_29865,N_29384);
or UO_1549 (O_1549,N_29573,N_29832);
nor UO_1550 (O_1550,N_28820,N_28376);
nand UO_1551 (O_1551,N_29569,N_29541);
xnor UO_1552 (O_1552,N_29966,N_28314);
xnor UO_1553 (O_1553,N_29259,N_29014);
nor UO_1554 (O_1554,N_28908,N_29192);
and UO_1555 (O_1555,N_29845,N_29024);
nor UO_1556 (O_1556,N_28069,N_29399);
nor UO_1557 (O_1557,N_28094,N_29592);
nand UO_1558 (O_1558,N_29465,N_28642);
or UO_1559 (O_1559,N_28850,N_28380);
and UO_1560 (O_1560,N_28819,N_28052);
nor UO_1561 (O_1561,N_29480,N_29626);
nand UO_1562 (O_1562,N_28167,N_28566);
nand UO_1563 (O_1563,N_28532,N_28859);
nand UO_1564 (O_1564,N_28619,N_28576);
and UO_1565 (O_1565,N_29777,N_29198);
or UO_1566 (O_1566,N_28722,N_29504);
and UO_1567 (O_1567,N_28187,N_29573);
nand UO_1568 (O_1568,N_29860,N_28451);
xnor UO_1569 (O_1569,N_29355,N_29459);
nor UO_1570 (O_1570,N_28850,N_28637);
or UO_1571 (O_1571,N_29146,N_29678);
and UO_1572 (O_1572,N_29584,N_29655);
and UO_1573 (O_1573,N_29638,N_28407);
xor UO_1574 (O_1574,N_28553,N_28979);
nand UO_1575 (O_1575,N_29781,N_29410);
or UO_1576 (O_1576,N_28777,N_29746);
nand UO_1577 (O_1577,N_29538,N_29559);
and UO_1578 (O_1578,N_28915,N_28351);
nand UO_1579 (O_1579,N_29296,N_29012);
and UO_1580 (O_1580,N_29199,N_28276);
nor UO_1581 (O_1581,N_29878,N_28872);
and UO_1582 (O_1582,N_28164,N_29829);
nor UO_1583 (O_1583,N_29236,N_29076);
or UO_1584 (O_1584,N_28801,N_28892);
and UO_1585 (O_1585,N_28066,N_28338);
nor UO_1586 (O_1586,N_29694,N_28159);
and UO_1587 (O_1587,N_29794,N_29400);
xnor UO_1588 (O_1588,N_28249,N_28401);
and UO_1589 (O_1589,N_29089,N_28496);
nand UO_1590 (O_1590,N_29278,N_28724);
nand UO_1591 (O_1591,N_28944,N_29528);
or UO_1592 (O_1592,N_29830,N_29916);
and UO_1593 (O_1593,N_29886,N_28732);
xor UO_1594 (O_1594,N_29662,N_29082);
or UO_1595 (O_1595,N_28048,N_28039);
and UO_1596 (O_1596,N_28988,N_28603);
nor UO_1597 (O_1597,N_29760,N_29822);
and UO_1598 (O_1598,N_28771,N_29887);
and UO_1599 (O_1599,N_29990,N_29373);
and UO_1600 (O_1600,N_29216,N_29389);
xor UO_1601 (O_1601,N_28238,N_28500);
nor UO_1602 (O_1602,N_29782,N_29270);
or UO_1603 (O_1603,N_29579,N_28466);
nand UO_1604 (O_1604,N_28710,N_28877);
nand UO_1605 (O_1605,N_29585,N_28905);
or UO_1606 (O_1606,N_29325,N_29396);
and UO_1607 (O_1607,N_28655,N_28764);
and UO_1608 (O_1608,N_28368,N_28139);
and UO_1609 (O_1609,N_28001,N_28990);
nand UO_1610 (O_1610,N_28454,N_29873);
xor UO_1611 (O_1611,N_28295,N_28796);
nor UO_1612 (O_1612,N_28970,N_29915);
nor UO_1613 (O_1613,N_28999,N_29693);
or UO_1614 (O_1614,N_29184,N_29128);
or UO_1615 (O_1615,N_28287,N_28054);
or UO_1616 (O_1616,N_28842,N_29597);
nand UO_1617 (O_1617,N_28613,N_28735);
xnor UO_1618 (O_1618,N_29530,N_29691);
or UO_1619 (O_1619,N_29989,N_28121);
or UO_1620 (O_1620,N_29482,N_28159);
xnor UO_1621 (O_1621,N_28725,N_29414);
nor UO_1622 (O_1622,N_29477,N_29328);
nand UO_1623 (O_1623,N_28944,N_29603);
or UO_1624 (O_1624,N_28492,N_29229);
nor UO_1625 (O_1625,N_28680,N_28907);
xor UO_1626 (O_1626,N_29917,N_28136);
nor UO_1627 (O_1627,N_29416,N_28388);
nor UO_1628 (O_1628,N_29393,N_29227);
or UO_1629 (O_1629,N_28690,N_29767);
xor UO_1630 (O_1630,N_29841,N_28229);
and UO_1631 (O_1631,N_28592,N_28393);
xnor UO_1632 (O_1632,N_28971,N_28011);
nor UO_1633 (O_1633,N_29848,N_28521);
nand UO_1634 (O_1634,N_29867,N_28603);
and UO_1635 (O_1635,N_28673,N_29649);
nor UO_1636 (O_1636,N_28867,N_28044);
nand UO_1637 (O_1637,N_28677,N_28679);
or UO_1638 (O_1638,N_29891,N_29007);
and UO_1639 (O_1639,N_28914,N_29209);
or UO_1640 (O_1640,N_28104,N_28060);
nand UO_1641 (O_1641,N_28689,N_29379);
nor UO_1642 (O_1642,N_29921,N_29258);
and UO_1643 (O_1643,N_28486,N_28234);
nand UO_1644 (O_1644,N_29784,N_29814);
nor UO_1645 (O_1645,N_28907,N_29232);
and UO_1646 (O_1646,N_29450,N_28854);
and UO_1647 (O_1647,N_28709,N_28207);
and UO_1648 (O_1648,N_29464,N_29010);
xor UO_1649 (O_1649,N_29680,N_29311);
nor UO_1650 (O_1650,N_29369,N_28158);
or UO_1651 (O_1651,N_29168,N_28717);
nor UO_1652 (O_1652,N_29108,N_29113);
nand UO_1653 (O_1653,N_29489,N_29518);
nor UO_1654 (O_1654,N_28588,N_28717);
xor UO_1655 (O_1655,N_28923,N_29459);
or UO_1656 (O_1656,N_29823,N_29951);
nor UO_1657 (O_1657,N_28885,N_29343);
nor UO_1658 (O_1658,N_28432,N_29839);
xnor UO_1659 (O_1659,N_28160,N_28717);
xor UO_1660 (O_1660,N_28429,N_29539);
and UO_1661 (O_1661,N_29014,N_29619);
or UO_1662 (O_1662,N_28113,N_28806);
nand UO_1663 (O_1663,N_29847,N_29678);
nor UO_1664 (O_1664,N_28810,N_28879);
or UO_1665 (O_1665,N_29392,N_29123);
or UO_1666 (O_1666,N_29147,N_29877);
xnor UO_1667 (O_1667,N_28789,N_28882);
and UO_1668 (O_1668,N_29007,N_29698);
and UO_1669 (O_1669,N_29902,N_28934);
nor UO_1670 (O_1670,N_28463,N_28808);
or UO_1671 (O_1671,N_28553,N_28323);
nor UO_1672 (O_1672,N_29638,N_28932);
and UO_1673 (O_1673,N_29008,N_28105);
nor UO_1674 (O_1674,N_29262,N_28028);
or UO_1675 (O_1675,N_29977,N_28254);
xor UO_1676 (O_1676,N_29294,N_29354);
and UO_1677 (O_1677,N_29324,N_29972);
xnor UO_1678 (O_1678,N_29585,N_28850);
xor UO_1679 (O_1679,N_28852,N_28664);
nor UO_1680 (O_1680,N_28362,N_28096);
nand UO_1681 (O_1681,N_28609,N_29454);
xor UO_1682 (O_1682,N_28490,N_28324);
and UO_1683 (O_1683,N_29009,N_29133);
or UO_1684 (O_1684,N_28979,N_29738);
and UO_1685 (O_1685,N_29175,N_28914);
xor UO_1686 (O_1686,N_28122,N_28241);
nand UO_1687 (O_1687,N_28945,N_28217);
or UO_1688 (O_1688,N_28851,N_29081);
and UO_1689 (O_1689,N_29604,N_29927);
nand UO_1690 (O_1690,N_28560,N_29141);
nor UO_1691 (O_1691,N_29263,N_29786);
nand UO_1692 (O_1692,N_28268,N_28411);
and UO_1693 (O_1693,N_29365,N_29317);
and UO_1694 (O_1694,N_29748,N_28977);
and UO_1695 (O_1695,N_28335,N_28003);
and UO_1696 (O_1696,N_29639,N_29373);
nand UO_1697 (O_1697,N_28720,N_29830);
and UO_1698 (O_1698,N_28265,N_29336);
and UO_1699 (O_1699,N_29004,N_28650);
or UO_1700 (O_1700,N_29873,N_28227);
nand UO_1701 (O_1701,N_28557,N_28775);
nor UO_1702 (O_1702,N_28994,N_28795);
and UO_1703 (O_1703,N_29868,N_28142);
or UO_1704 (O_1704,N_28238,N_28223);
and UO_1705 (O_1705,N_29202,N_28519);
and UO_1706 (O_1706,N_28637,N_29276);
xor UO_1707 (O_1707,N_29206,N_29315);
and UO_1708 (O_1708,N_29419,N_29115);
nand UO_1709 (O_1709,N_29306,N_29377);
and UO_1710 (O_1710,N_29550,N_29589);
nand UO_1711 (O_1711,N_29193,N_29493);
or UO_1712 (O_1712,N_29879,N_29605);
xor UO_1713 (O_1713,N_28522,N_28255);
xor UO_1714 (O_1714,N_29259,N_29614);
nand UO_1715 (O_1715,N_28254,N_28413);
nand UO_1716 (O_1716,N_28075,N_29785);
and UO_1717 (O_1717,N_28526,N_28414);
or UO_1718 (O_1718,N_28059,N_29348);
and UO_1719 (O_1719,N_29410,N_29342);
and UO_1720 (O_1720,N_28626,N_28775);
nor UO_1721 (O_1721,N_29872,N_29652);
nand UO_1722 (O_1722,N_28887,N_28623);
and UO_1723 (O_1723,N_28283,N_29115);
nand UO_1724 (O_1724,N_29238,N_28040);
xnor UO_1725 (O_1725,N_29261,N_29239);
xnor UO_1726 (O_1726,N_28089,N_28612);
and UO_1727 (O_1727,N_28263,N_29840);
nor UO_1728 (O_1728,N_28679,N_29282);
and UO_1729 (O_1729,N_28262,N_28799);
nand UO_1730 (O_1730,N_29731,N_28802);
nand UO_1731 (O_1731,N_28573,N_28129);
or UO_1732 (O_1732,N_29493,N_28777);
or UO_1733 (O_1733,N_28056,N_28325);
and UO_1734 (O_1734,N_28043,N_29864);
and UO_1735 (O_1735,N_28946,N_28601);
xnor UO_1736 (O_1736,N_28335,N_28661);
nor UO_1737 (O_1737,N_29279,N_28544);
or UO_1738 (O_1738,N_28944,N_29108);
or UO_1739 (O_1739,N_29674,N_29215);
xnor UO_1740 (O_1740,N_28002,N_28108);
and UO_1741 (O_1741,N_29922,N_29378);
or UO_1742 (O_1742,N_29985,N_29014);
xnor UO_1743 (O_1743,N_28187,N_28531);
nand UO_1744 (O_1744,N_29530,N_28517);
nand UO_1745 (O_1745,N_28822,N_28204);
nor UO_1746 (O_1746,N_28783,N_29559);
xor UO_1747 (O_1747,N_29148,N_28934);
and UO_1748 (O_1748,N_28475,N_28485);
nand UO_1749 (O_1749,N_29141,N_28969);
nand UO_1750 (O_1750,N_28515,N_28976);
or UO_1751 (O_1751,N_29166,N_28582);
xor UO_1752 (O_1752,N_28318,N_28428);
or UO_1753 (O_1753,N_29008,N_28466);
nand UO_1754 (O_1754,N_29622,N_29014);
nand UO_1755 (O_1755,N_28265,N_28950);
or UO_1756 (O_1756,N_29704,N_29994);
and UO_1757 (O_1757,N_28520,N_29897);
or UO_1758 (O_1758,N_28973,N_29597);
or UO_1759 (O_1759,N_28015,N_29074);
and UO_1760 (O_1760,N_29520,N_29530);
nand UO_1761 (O_1761,N_29307,N_29499);
nor UO_1762 (O_1762,N_28324,N_28566);
and UO_1763 (O_1763,N_29582,N_28602);
and UO_1764 (O_1764,N_29745,N_28391);
xnor UO_1765 (O_1765,N_28193,N_28953);
or UO_1766 (O_1766,N_28519,N_28852);
nand UO_1767 (O_1767,N_28381,N_29068);
nand UO_1768 (O_1768,N_28910,N_29002);
xor UO_1769 (O_1769,N_29489,N_29231);
or UO_1770 (O_1770,N_28805,N_29037);
xor UO_1771 (O_1771,N_29446,N_28086);
nor UO_1772 (O_1772,N_28059,N_28153);
nor UO_1773 (O_1773,N_28359,N_29507);
nor UO_1774 (O_1774,N_28919,N_28656);
and UO_1775 (O_1775,N_29911,N_29788);
xor UO_1776 (O_1776,N_29721,N_28033);
and UO_1777 (O_1777,N_28871,N_29291);
nand UO_1778 (O_1778,N_28105,N_29868);
nor UO_1779 (O_1779,N_28831,N_29744);
and UO_1780 (O_1780,N_29770,N_29601);
xnor UO_1781 (O_1781,N_29545,N_28918);
or UO_1782 (O_1782,N_28906,N_29678);
xnor UO_1783 (O_1783,N_28306,N_29968);
and UO_1784 (O_1784,N_28817,N_28854);
nor UO_1785 (O_1785,N_28429,N_28624);
nand UO_1786 (O_1786,N_29710,N_29186);
nor UO_1787 (O_1787,N_29186,N_29286);
or UO_1788 (O_1788,N_28031,N_28651);
xnor UO_1789 (O_1789,N_28066,N_29913);
nor UO_1790 (O_1790,N_28022,N_28071);
and UO_1791 (O_1791,N_29538,N_28001);
and UO_1792 (O_1792,N_29946,N_29806);
xor UO_1793 (O_1793,N_29318,N_29270);
and UO_1794 (O_1794,N_29526,N_28329);
xnor UO_1795 (O_1795,N_29838,N_28687);
and UO_1796 (O_1796,N_28552,N_29882);
nor UO_1797 (O_1797,N_28344,N_29469);
or UO_1798 (O_1798,N_29916,N_28299);
or UO_1799 (O_1799,N_29343,N_28798);
xor UO_1800 (O_1800,N_28321,N_29724);
nor UO_1801 (O_1801,N_28244,N_29455);
xnor UO_1802 (O_1802,N_29302,N_29487);
nor UO_1803 (O_1803,N_28620,N_28530);
or UO_1804 (O_1804,N_28277,N_28963);
nand UO_1805 (O_1805,N_28457,N_29757);
or UO_1806 (O_1806,N_28014,N_29676);
or UO_1807 (O_1807,N_28782,N_28228);
xnor UO_1808 (O_1808,N_29234,N_28706);
or UO_1809 (O_1809,N_28097,N_29618);
and UO_1810 (O_1810,N_29041,N_29577);
nand UO_1811 (O_1811,N_29742,N_29070);
or UO_1812 (O_1812,N_29142,N_29510);
nand UO_1813 (O_1813,N_28216,N_28644);
nand UO_1814 (O_1814,N_28692,N_28306);
or UO_1815 (O_1815,N_28459,N_28662);
nor UO_1816 (O_1816,N_29658,N_29976);
nor UO_1817 (O_1817,N_28642,N_29126);
and UO_1818 (O_1818,N_29580,N_29526);
nand UO_1819 (O_1819,N_28199,N_29195);
nand UO_1820 (O_1820,N_28236,N_29400);
or UO_1821 (O_1821,N_28355,N_29275);
xor UO_1822 (O_1822,N_28993,N_29381);
and UO_1823 (O_1823,N_28580,N_28714);
or UO_1824 (O_1824,N_29189,N_28789);
or UO_1825 (O_1825,N_29369,N_28766);
nor UO_1826 (O_1826,N_28491,N_29467);
xnor UO_1827 (O_1827,N_29935,N_29775);
nand UO_1828 (O_1828,N_29330,N_28433);
nor UO_1829 (O_1829,N_28107,N_28605);
nand UO_1830 (O_1830,N_29925,N_29734);
xor UO_1831 (O_1831,N_28966,N_29703);
and UO_1832 (O_1832,N_29933,N_29208);
nor UO_1833 (O_1833,N_29212,N_28099);
and UO_1834 (O_1834,N_28854,N_28818);
and UO_1835 (O_1835,N_28719,N_29889);
and UO_1836 (O_1836,N_28502,N_28876);
and UO_1837 (O_1837,N_28318,N_28463);
nand UO_1838 (O_1838,N_29563,N_28054);
or UO_1839 (O_1839,N_28056,N_29499);
or UO_1840 (O_1840,N_29107,N_29559);
nor UO_1841 (O_1841,N_28406,N_28635);
nor UO_1842 (O_1842,N_29727,N_29162);
nand UO_1843 (O_1843,N_28282,N_28211);
and UO_1844 (O_1844,N_28934,N_28044);
or UO_1845 (O_1845,N_28546,N_29077);
and UO_1846 (O_1846,N_28740,N_29102);
or UO_1847 (O_1847,N_29522,N_29159);
xnor UO_1848 (O_1848,N_29360,N_29079);
nand UO_1849 (O_1849,N_29425,N_28938);
nand UO_1850 (O_1850,N_28923,N_28660);
nor UO_1851 (O_1851,N_28158,N_28499);
or UO_1852 (O_1852,N_29684,N_29149);
or UO_1853 (O_1853,N_29995,N_28644);
and UO_1854 (O_1854,N_29854,N_28210);
and UO_1855 (O_1855,N_29626,N_28974);
xor UO_1856 (O_1856,N_28135,N_29532);
xnor UO_1857 (O_1857,N_28387,N_28869);
or UO_1858 (O_1858,N_29102,N_29767);
and UO_1859 (O_1859,N_29640,N_29222);
nand UO_1860 (O_1860,N_28927,N_29091);
nor UO_1861 (O_1861,N_29215,N_28674);
nor UO_1862 (O_1862,N_28997,N_29407);
nor UO_1863 (O_1863,N_29501,N_29668);
xnor UO_1864 (O_1864,N_29424,N_29975);
nor UO_1865 (O_1865,N_29887,N_29979);
and UO_1866 (O_1866,N_29864,N_28614);
or UO_1867 (O_1867,N_29028,N_29432);
and UO_1868 (O_1868,N_29424,N_28597);
xor UO_1869 (O_1869,N_28110,N_29393);
nand UO_1870 (O_1870,N_29136,N_28485);
or UO_1871 (O_1871,N_29404,N_28151);
and UO_1872 (O_1872,N_28390,N_28866);
or UO_1873 (O_1873,N_29291,N_28600);
or UO_1874 (O_1874,N_28852,N_29222);
and UO_1875 (O_1875,N_28487,N_28820);
xor UO_1876 (O_1876,N_29636,N_29405);
and UO_1877 (O_1877,N_29305,N_28463);
xnor UO_1878 (O_1878,N_29720,N_29046);
or UO_1879 (O_1879,N_28747,N_28433);
xor UO_1880 (O_1880,N_29687,N_29780);
xnor UO_1881 (O_1881,N_29603,N_28505);
and UO_1882 (O_1882,N_29976,N_29775);
and UO_1883 (O_1883,N_28911,N_29608);
xnor UO_1884 (O_1884,N_28057,N_28589);
xor UO_1885 (O_1885,N_29815,N_28894);
nor UO_1886 (O_1886,N_28631,N_29848);
or UO_1887 (O_1887,N_28402,N_28623);
and UO_1888 (O_1888,N_29030,N_28884);
and UO_1889 (O_1889,N_28528,N_29919);
or UO_1890 (O_1890,N_28898,N_28755);
or UO_1891 (O_1891,N_29104,N_28276);
nor UO_1892 (O_1892,N_28492,N_28849);
nor UO_1893 (O_1893,N_28160,N_29792);
and UO_1894 (O_1894,N_29967,N_29509);
xor UO_1895 (O_1895,N_29297,N_28845);
xor UO_1896 (O_1896,N_29430,N_29044);
or UO_1897 (O_1897,N_29463,N_28109);
nor UO_1898 (O_1898,N_29511,N_28065);
and UO_1899 (O_1899,N_28782,N_29501);
nor UO_1900 (O_1900,N_29625,N_28232);
nor UO_1901 (O_1901,N_28608,N_28032);
nor UO_1902 (O_1902,N_29866,N_29077);
nor UO_1903 (O_1903,N_28412,N_29665);
nor UO_1904 (O_1904,N_28324,N_29611);
xor UO_1905 (O_1905,N_28362,N_29525);
nor UO_1906 (O_1906,N_29624,N_28268);
nand UO_1907 (O_1907,N_28495,N_28523);
xor UO_1908 (O_1908,N_28944,N_28129);
xnor UO_1909 (O_1909,N_29000,N_28614);
xnor UO_1910 (O_1910,N_29887,N_28545);
and UO_1911 (O_1911,N_28966,N_29849);
xor UO_1912 (O_1912,N_28815,N_28436);
and UO_1913 (O_1913,N_29574,N_28943);
or UO_1914 (O_1914,N_28364,N_29987);
or UO_1915 (O_1915,N_29215,N_28147);
nand UO_1916 (O_1916,N_29207,N_29811);
nand UO_1917 (O_1917,N_28271,N_29563);
or UO_1918 (O_1918,N_29061,N_29435);
xnor UO_1919 (O_1919,N_28384,N_28503);
xnor UO_1920 (O_1920,N_28402,N_28938);
nand UO_1921 (O_1921,N_29854,N_29995);
nor UO_1922 (O_1922,N_29245,N_28288);
xor UO_1923 (O_1923,N_29102,N_29743);
nor UO_1924 (O_1924,N_28392,N_29998);
nor UO_1925 (O_1925,N_29503,N_29130);
nand UO_1926 (O_1926,N_29716,N_28894);
or UO_1927 (O_1927,N_29089,N_28203);
nor UO_1928 (O_1928,N_29799,N_29862);
nand UO_1929 (O_1929,N_28563,N_29789);
nor UO_1930 (O_1930,N_29545,N_29230);
xnor UO_1931 (O_1931,N_29863,N_29552);
and UO_1932 (O_1932,N_29527,N_28251);
xnor UO_1933 (O_1933,N_29017,N_29168);
or UO_1934 (O_1934,N_29449,N_29967);
and UO_1935 (O_1935,N_28346,N_29547);
or UO_1936 (O_1936,N_28806,N_28691);
and UO_1937 (O_1937,N_28599,N_29007);
or UO_1938 (O_1938,N_29390,N_29148);
or UO_1939 (O_1939,N_28348,N_29618);
or UO_1940 (O_1940,N_29781,N_29042);
nand UO_1941 (O_1941,N_29509,N_29328);
or UO_1942 (O_1942,N_29916,N_29458);
nor UO_1943 (O_1943,N_29076,N_29808);
xnor UO_1944 (O_1944,N_28603,N_28762);
nor UO_1945 (O_1945,N_28368,N_28427);
nor UO_1946 (O_1946,N_28680,N_28821);
nand UO_1947 (O_1947,N_28242,N_29596);
and UO_1948 (O_1948,N_28826,N_29259);
and UO_1949 (O_1949,N_28859,N_29206);
or UO_1950 (O_1950,N_29420,N_28683);
or UO_1951 (O_1951,N_29633,N_28290);
or UO_1952 (O_1952,N_29043,N_29619);
nor UO_1953 (O_1953,N_29753,N_29496);
nor UO_1954 (O_1954,N_28743,N_29131);
nor UO_1955 (O_1955,N_29612,N_28415);
xnor UO_1956 (O_1956,N_29645,N_28397);
xnor UO_1957 (O_1957,N_28941,N_29171);
and UO_1958 (O_1958,N_29376,N_29457);
or UO_1959 (O_1959,N_28101,N_28145);
xnor UO_1960 (O_1960,N_28360,N_28141);
xor UO_1961 (O_1961,N_28695,N_28783);
nor UO_1962 (O_1962,N_29074,N_28650);
and UO_1963 (O_1963,N_28599,N_28008);
and UO_1964 (O_1964,N_29021,N_29894);
or UO_1965 (O_1965,N_29213,N_28532);
or UO_1966 (O_1966,N_29007,N_28083);
nand UO_1967 (O_1967,N_28191,N_29172);
xor UO_1968 (O_1968,N_28677,N_28278);
xnor UO_1969 (O_1969,N_28877,N_28617);
xnor UO_1970 (O_1970,N_29958,N_29367);
nor UO_1971 (O_1971,N_29011,N_28197);
xor UO_1972 (O_1972,N_29412,N_29831);
or UO_1973 (O_1973,N_29707,N_28103);
xor UO_1974 (O_1974,N_28249,N_29983);
nor UO_1975 (O_1975,N_28371,N_28498);
and UO_1976 (O_1976,N_29447,N_28821);
or UO_1977 (O_1977,N_28692,N_29816);
or UO_1978 (O_1978,N_28885,N_29528);
nand UO_1979 (O_1979,N_28539,N_29089);
xor UO_1980 (O_1980,N_28787,N_29553);
and UO_1981 (O_1981,N_29087,N_29196);
or UO_1982 (O_1982,N_29957,N_28925);
or UO_1983 (O_1983,N_29372,N_28765);
xor UO_1984 (O_1984,N_28792,N_29108);
xnor UO_1985 (O_1985,N_29008,N_29714);
and UO_1986 (O_1986,N_29665,N_28295);
nor UO_1987 (O_1987,N_29337,N_29972);
and UO_1988 (O_1988,N_29598,N_28320);
xnor UO_1989 (O_1989,N_28067,N_29553);
xor UO_1990 (O_1990,N_28883,N_29697);
or UO_1991 (O_1991,N_28550,N_29838);
nor UO_1992 (O_1992,N_29671,N_28591);
nor UO_1993 (O_1993,N_28034,N_28120);
and UO_1994 (O_1994,N_28293,N_29951);
and UO_1995 (O_1995,N_29436,N_28917);
nand UO_1996 (O_1996,N_28294,N_29287);
nor UO_1997 (O_1997,N_29905,N_29046);
or UO_1998 (O_1998,N_28512,N_29757);
or UO_1999 (O_1999,N_28018,N_29897);
and UO_2000 (O_2000,N_29977,N_28801);
nor UO_2001 (O_2001,N_29838,N_28667);
and UO_2002 (O_2002,N_29624,N_29076);
nand UO_2003 (O_2003,N_29246,N_28392);
xnor UO_2004 (O_2004,N_29397,N_28275);
and UO_2005 (O_2005,N_28974,N_28260);
nor UO_2006 (O_2006,N_29401,N_29553);
or UO_2007 (O_2007,N_28881,N_29930);
and UO_2008 (O_2008,N_29108,N_28000);
and UO_2009 (O_2009,N_29717,N_29063);
or UO_2010 (O_2010,N_28408,N_28845);
nor UO_2011 (O_2011,N_29534,N_29535);
nand UO_2012 (O_2012,N_28555,N_29663);
and UO_2013 (O_2013,N_28940,N_28847);
nand UO_2014 (O_2014,N_29346,N_28086);
xnor UO_2015 (O_2015,N_28318,N_29382);
nand UO_2016 (O_2016,N_28117,N_28479);
or UO_2017 (O_2017,N_29814,N_29496);
xor UO_2018 (O_2018,N_28954,N_28309);
xor UO_2019 (O_2019,N_28441,N_28978);
nand UO_2020 (O_2020,N_29308,N_28036);
or UO_2021 (O_2021,N_28917,N_28213);
xnor UO_2022 (O_2022,N_28712,N_28032);
nor UO_2023 (O_2023,N_29620,N_29171);
or UO_2024 (O_2024,N_29895,N_29651);
xor UO_2025 (O_2025,N_28816,N_29803);
nand UO_2026 (O_2026,N_29505,N_28429);
and UO_2027 (O_2027,N_29981,N_29437);
nor UO_2028 (O_2028,N_28991,N_28828);
or UO_2029 (O_2029,N_28823,N_29864);
nand UO_2030 (O_2030,N_28835,N_28346);
nand UO_2031 (O_2031,N_28621,N_29525);
xnor UO_2032 (O_2032,N_28278,N_28365);
and UO_2033 (O_2033,N_28088,N_29317);
nand UO_2034 (O_2034,N_28734,N_29858);
or UO_2035 (O_2035,N_28704,N_29291);
and UO_2036 (O_2036,N_29608,N_28353);
or UO_2037 (O_2037,N_29136,N_28905);
and UO_2038 (O_2038,N_28798,N_29074);
nor UO_2039 (O_2039,N_29232,N_28563);
nor UO_2040 (O_2040,N_29678,N_28550);
or UO_2041 (O_2041,N_28970,N_29842);
or UO_2042 (O_2042,N_28205,N_28440);
xnor UO_2043 (O_2043,N_29064,N_28029);
xor UO_2044 (O_2044,N_29298,N_28043);
nor UO_2045 (O_2045,N_28929,N_28774);
nor UO_2046 (O_2046,N_28614,N_28801);
nor UO_2047 (O_2047,N_29042,N_29151);
xnor UO_2048 (O_2048,N_29287,N_28004);
xnor UO_2049 (O_2049,N_28138,N_29246);
nand UO_2050 (O_2050,N_29258,N_28522);
nand UO_2051 (O_2051,N_28677,N_28043);
xor UO_2052 (O_2052,N_28768,N_28631);
xnor UO_2053 (O_2053,N_28717,N_29994);
nor UO_2054 (O_2054,N_28985,N_28711);
or UO_2055 (O_2055,N_28783,N_28605);
xor UO_2056 (O_2056,N_28666,N_29672);
nor UO_2057 (O_2057,N_29026,N_28336);
and UO_2058 (O_2058,N_28091,N_28530);
nand UO_2059 (O_2059,N_28835,N_29449);
nand UO_2060 (O_2060,N_28403,N_28391);
nor UO_2061 (O_2061,N_29871,N_28090);
xor UO_2062 (O_2062,N_29700,N_29452);
nor UO_2063 (O_2063,N_28093,N_28467);
or UO_2064 (O_2064,N_29739,N_28310);
nand UO_2065 (O_2065,N_28008,N_28755);
and UO_2066 (O_2066,N_29458,N_29677);
or UO_2067 (O_2067,N_28694,N_29945);
and UO_2068 (O_2068,N_29096,N_29363);
or UO_2069 (O_2069,N_28234,N_29091);
xor UO_2070 (O_2070,N_29243,N_28024);
nor UO_2071 (O_2071,N_29340,N_29971);
or UO_2072 (O_2072,N_28007,N_29204);
xor UO_2073 (O_2073,N_29010,N_29955);
nor UO_2074 (O_2074,N_29554,N_28762);
or UO_2075 (O_2075,N_28970,N_28287);
xor UO_2076 (O_2076,N_28642,N_28596);
or UO_2077 (O_2077,N_28748,N_29354);
nor UO_2078 (O_2078,N_28243,N_28824);
xnor UO_2079 (O_2079,N_29018,N_29816);
and UO_2080 (O_2080,N_29718,N_28484);
and UO_2081 (O_2081,N_28825,N_28849);
and UO_2082 (O_2082,N_28702,N_29897);
nor UO_2083 (O_2083,N_29218,N_29107);
and UO_2084 (O_2084,N_28645,N_28936);
nor UO_2085 (O_2085,N_29754,N_29513);
and UO_2086 (O_2086,N_28721,N_29456);
and UO_2087 (O_2087,N_29047,N_28158);
nor UO_2088 (O_2088,N_29917,N_28213);
xnor UO_2089 (O_2089,N_28091,N_29920);
xor UO_2090 (O_2090,N_29970,N_28162);
nor UO_2091 (O_2091,N_28663,N_29222);
or UO_2092 (O_2092,N_28836,N_29221);
and UO_2093 (O_2093,N_28461,N_29190);
nand UO_2094 (O_2094,N_28821,N_29778);
nand UO_2095 (O_2095,N_29037,N_29394);
nor UO_2096 (O_2096,N_29766,N_28846);
nand UO_2097 (O_2097,N_28387,N_28940);
xor UO_2098 (O_2098,N_29117,N_28252);
or UO_2099 (O_2099,N_29766,N_28180);
and UO_2100 (O_2100,N_28640,N_28524);
xnor UO_2101 (O_2101,N_28547,N_28974);
nor UO_2102 (O_2102,N_29626,N_29672);
nor UO_2103 (O_2103,N_28523,N_28437);
nor UO_2104 (O_2104,N_29349,N_29171);
nand UO_2105 (O_2105,N_29178,N_29146);
or UO_2106 (O_2106,N_29635,N_29535);
nand UO_2107 (O_2107,N_28837,N_29617);
xor UO_2108 (O_2108,N_29372,N_29530);
xor UO_2109 (O_2109,N_29691,N_29017);
and UO_2110 (O_2110,N_29268,N_29233);
nor UO_2111 (O_2111,N_28571,N_29196);
xnor UO_2112 (O_2112,N_28644,N_28866);
xor UO_2113 (O_2113,N_28958,N_28133);
xnor UO_2114 (O_2114,N_28201,N_28813);
nor UO_2115 (O_2115,N_29067,N_28682);
or UO_2116 (O_2116,N_28479,N_28259);
or UO_2117 (O_2117,N_29113,N_28814);
and UO_2118 (O_2118,N_29818,N_28742);
xnor UO_2119 (O_2119,N_29314,N_29063);
and UO_2120 (O_2120,N_28569,N_29831);
xor UO_2121 (O_2121,N_28835,N_29804);
nand UO_2122 (O_2122,N_29689,N_29272);
or UO_2123 (O_2123,N_29713,N_29608);
xor UO_2124 (O_2124,N_28337,N_28453);
and UO_2125 (O_2125,N_29746,N_29751);
nand UO_2126 (O_2126,N_28505,N_28549);
and UO_2127 (O_2127,N_29038,N_28614);
and UO_2128 (O_2128,N_28330,N_29295);
and UO_2129 (O_2129,N_29844,N_29328);
and UO_2130 (O_2130,N_28474,N_29575);
nand UO_2131 (O_2131,N_28219,N_29644);
and UO_2132 (O_2132,N_28790,N_29752);
or UO_2133 (O_2133,N_28469,N_28835);
nor UO_2134 (O_2134,N_28491,N_29465);
xor UO_2135 (O_2135,N_28211,N_29983);
nor UO_2136 (O_2136,N_29046,N_28309);
or UO_2137 (O_2137,N_29397,N_28324);
xnor UO_2138 (O_2138,N_28223,N_29504);
or UO_2139 (O_2139,N_28905,N_29259);
nor UO_2140 (O_2140,N_29222,N_29280);
and UO_2141 (O_2141,N_28570,N_29424);
nor UO_2142 (O_2142,N_28247,N_29739);
or UO_2143 (O_2143,N_29282,N_29064);
xnor UO_2144 (O_2144,N_28421,N_28384);
nand UO_2145 (O_2145,N_29892,N_28553);
and UO_2146 (O_2146,N_29151,N_28593);
and UO_2147 (O_2147,N_28183,N_29921);
or UO_2148 (O_2148,N_28388,N_29856);
nand UO_2149 (O_2149,N_28153,N_29835);
nand UO_2150 (O_2150,N_29636,N_29866);
xnor UO_2151 (O_2151,N_29200,N_29601);
nand UO_2152 (O_2152,N_28176,N_28881);
nor UO_2153 (O_2153,N_28905,N_29483);
and UO_2154 (O_2154,N_29827,N_29569);
or UO_2155 (O_2155,N_29837,N_29499);
xor UO_2156 (O_2156,N_28560,N_29263);
or UO_2157 (O_2157,N_28179,N_29590);
or UO_2158 (O_2158,N_29846,N_29328);
xor UO_2159 (O_2159,N_28268,N_29279);
nor UO_2160 (O_2160,N_28475,N_29048);
or UO_2161 (O_2161,N_29765,N_29912);
or UO_2162 (O_2162,N_29462,N_28181);
or UO_2163 (O_2163,N_28221,N_29668);
xor UO_2164 (O_2164,N_28994,N_29787);
nor UO_2165 (O_2165,N_28957,N_28843);
nor UO_2166 (O_2166,N_29073,N_28665);
xor UO_2167 (O_2167,N_28792,N_28737);
or UO_2168 (O_2168,N_29726,N_29527);
or UO_2169 (O_2169,N_28982,N_29671);
nand UO_2170 (O_2170,N_28876,N_28828);
nor UO_2171 (O_2171,N_29572,N_29061);
nand UO_2172 (O_2172,N_28000,N_28100);
nand UO_2173 (O_2173,N_29321,N_28747);
xnor UO_2174 (O_2174,N_29381,N_29339);
nor UO_2175 (O_2175,N_28866,N_29105);
and UO_2176 (O_2176,N_28584,N_29469);
and UO_2177 (O_2177,N_28511,N_29317);
nor UO_2178 (O_2178,N_28036,N_29743);
and UO_2179 (O_2179,N_29748,N_29707);
nor UO_2180 (O_2180,N_29714,N_29643);
nor UO_2181 (O_2181,N_28128,N_28583);
nor UO_2182 (O_2182,N_28422,N_29869);
nor UO_2183 (O_2183,N_28897,N_29445);
nor UO_2184 (O_2184,N_29770,N_28880);
and UO_2185 (O_2185,N_28797,N_29887);
and UO_2186 (O_2186,N_28313,N_29473);
nand UO_2187 (O_2187,N_28872,N_28097);
nand UO_2188 (O_2188,N_29320,N_29178);
or UO_2189 (O_2189,N_28804,N_28469);
nor UO_2190 (O_2190,N_29915,N_29035);
xor UO_2191 (O_2191,N_29045,N_28613);
and UO_2192 (O_2192,N_28036,N_29087);
nor UO_2193 (O_2193,N_29564,N_29071);
or UO_2194 (O_2194,N_28315,N_29689);
nor UO_2195 (O_2195,N_29756,N_29795);
nor UO_2196 (O_2196,N_29231,N_29175);
nand UO_2197 (O_2197,N_29747,N_29658);
nand UO_2198 (O_2198,N_29585,N_29847);
nand UO_2199 (O_2199,N_28230,N_28931);
nand UO_2200 (O_2200,N_29908,N_28493);
nor UO_2201 (O_2201,N_28575,N_29169);
nand UO_2202 (O_2202,N_28437,N_28529);
xor UO_2203 (O_2203,N_28366,N_28774);
nor UO_2204 (O_2204,N_29285,N_29571);
xnor UO_2205 (O_2205,N_29769,N_29126);
and UO_2206 (O_2206,N_29025,N_28930);
nor UO_2207 (O_2207,N_29603,N_29293);
nor UO_2208 (O_2208,N_28648,N_29244);
xor UO_2209 (O_2209,N_29038,N_29147);
or UO_2210 (O_2210,N_29384,N_28025);
nor UO_2211 (O_2211,N_29683,N_29311);
or UO_2212 (O_2212,N_28194,N_28948);
nor UO_2213 (O_2213,N_28476,N_28988);
nand UO_2214 (O_2214,N_28612,N_29226);
xnor UO_2215 (O_2215,N_28665,N_28042);
xnor UO_2216 (O_2216,N_28915,N_28881);
and UO_2217 (O_2217,N_28397,N_28265);
xor UO_2218 (O_2218,N_28179,N_29622);
or UO_2219 (O_2219,N_29647,N_28016);
xor UO_2220 (O_2220,N_29656,N_28021);
nand UO_2221 (O_2221,N_28829,N_28803);
and UO_2222 (O_2222,N_28246,N_29617);
nand UO_2223 (O_2223,N_29840,N_29719);
nor UO_2224 (O_2224,N_28830,N_29591);
xor UO_2225 (O_2225,N_29958,N_29400);
or UO_2226 (O_2226,N_29162,N_28977);
xnor UO_2227 (O_2227,N_29982,N_29816);
or UO_2228 (O_2228,N_29995,N_28507);
xnor UO_2229 (O_2229,N_29264,N_29140);
or UO_2230 (O_2230,N_29304,N_29395);
and UO_2231 (O_2231,N_28048,N_29579);
nand UO_2232 (O_2232,N_28538,N_28417);
and UO_2233 (O_2233,N_29794,N_28338);
nand UO_2234 (O_2234,N_28914,N_29002);
and UO_2235 (O_2235,N_29145,N_28850);
or UO_2236 (O_2236,N_28446,N_29950);
nand UO_2237 (O_2237,N_29521,N_28133);
nand UO_2238 (O_2238,N_28605,N_28550);
nand UO_2239 (O_2239,N_29554,N_29424);
or UO_2240 (O_2240,N_29112,N_29990);
and UO_2241 (O_2241,N_29000,N_28330);
or UO_2242 (O_2242,N_29119,N_29204);
nor UO_2243 (O_2243,N_29842,N_28373);
nor UO_2244 (O_2244,N_28346,N_28971);
nor UO_2245 (O_2245,N_29983,N_28943);
nand UO_2246 (O_2246,N_29935,N_28872);
xor UO_2247 (O_2247,N_29686,N_29620);
nor UO_2248 (O_2248,N_29421,N_29081);
nor UO_2249 (O_2249,N_28709,N_29863);
nand UO_2250 (O_2250,N_29757,N_29327);
nor UO_2251 (O_2251,N_28611,N_28389);
or UO_2252 (O_2252,N_29213,N_28705);
or UO_2253 (O_2253,N_29266,N_29004);
nand UO_2254 (O_2254,N_28809,N_29904);
xnor UO_2255 (O_2255,N_29484,N_28424);
or UO_2256 (O_2256,N_28597,N_28489);
nand UO_2257 (O_2257,N_29980,N_29446);
xor UO_2258 (O_2258,N_29910,N_28589);
or UO_2259 (O_2259,N_29336,N_28710);
xor UO_2260 (O_2260,N_29702,N_29399);
nand UO_2261 (O_2261,N_28271,N_29241);
xor UO_2262 (O_2262,N_29154,N_28330);
xor UO_2263 (O_2263,N_29891,N_28470);
nor UO_2264 (O_2264,N_29111,N_28962);
xnor UO_2265 (O_2265,N_29216,N_29983);
xor UO_2266 (O_2266,N_29626,N_28850);
nor UO_2267 (O_2267,N_29379,N_28606);
or UO_2268 (O_2268,N_28503,N_28714);
xor UO_2269 (O_2269,N_28385,N_29709);
and UO_2270 (O_2270,N_29866,N_29281);
xnor UO_2271 (O_2271,N_28965,N_28578);
and UO_2272 (O_2272,N_29564,N_28992);
nand UO_2273 (O_2273,N_28757,N_28093);
xor UO_2274 (O_2274,N_28201,N_29115);
and UO_2275 (O_2275,N_29090,N_29484);
nor UO_2276 (O_2276,N_29715,N_28438);
or UO_2277 (O_2277,N_28554,N_28601);
and UO_2278 (O_2278,N_28650,N_29587);
xor UO_2279 (O_2279,N_28632,N_28558);
or UO_2280 (O_2280,N_28972,N_29107);
xnor UO_2281 (O_2281,N_28150,N_29413);
or UO_2282 (O_2282,N_29896,N_29575);
nand UO_2283 (O_2283,N_29667,N_29255);
xor UO_2284 (O_2284,N_29861,N_29702);
or UO_2285 (O_2285,N_29727,N_28334);
xnor UO_2286 (O_2286,N_28498,N_28564);
nor UO_2287 (O_2287,N_28983,N_28210);
nor UO_2288 (O_2288,N_28879,N_28616);
nor UO_2289 (O_2289,N_28091,N_29227);
nor UO_2290 (O_2290,N_29504,N_28570);
and UO_2291 (O_2291,N_28790,N_28450);
or UO_2292 (O_2292,N_28981,N_29788);
nor UO_2293 (O_2293,N_29726,N_29789);
nand UO_2294 (O_2294,N_29346,N_29216);
and UO_2295 (O_2295,N_29271,N_29622);
and UO_2296 (O_2296,N_28886,N_28585);
or UO_2297 (O_2297,N_28752,N_28388);
nor UO_2298 (O_2298,N_28236,N_28753);
xnor UO_2299 (O_2299,N_29692,N_28767);
and UO_2300 (O_2300,N_29353,N_29383);
xor UO_2301 (O_2301,N_29413,N_29158);
nor UO_2302 (O_2302,N_29778,N_28359);
nand UO_2303 (O_2303,N_29425,N_28158);
xnor UO_2304 (O_2304,N_29565,N_28435);
and UO_2305 (O_2305,N_28405,N_28069);
nand UO_2306 (O_2306,N_28346,N_28556);
and UO_2307 (O_2307,N_29225,N_28681);
or UO_2308 (O_2308,N_28438,N_29588);
nor UO_2309 (O_2309,N_29080,N_29890);
xnor UO_2310 (O_2310,N_29469,N_29173);
or UO_2311 (O_2311,N_28920,N_28917);
nand UO_2312 (O_2312,N_29860,N_29968);
or UO_2313 (O_2313,N_29208,N_29033);
or UO_2314 (O_2314,N_28540,N_29248);
nand UO_2315 (O_2315,N_29879,N_28182);
nand UO_2316 (O_2316,N_29190,N_28170);
nor UO_2317 (O_2317,N_28024,N_28087);
nor UO_2318 (O_2318,N_29239,N_29736);
nand UO_2319 (O_2319,N_29508,N_29555);
and UO_2320 (O_2320,N_28969,N_29467);
xor UO_2321 (O_2321,N_28229,N_29853);
and UO_2322 (O_2322,N_28353,N_28297);
nor UO_2323 (O_2323,N_29049,N_29374);
xnor UO_2324 (O_2324,N_28413,N_28914);
xor UO_2325 (O_2325,N_28684,N_29263);
and UO_2326 (O_2326,N_28085,N_28527);
nand UO_2327 (O_2327,N_28559,N_28457);
and UO_2328 (O_2328,N_29189,N_29990);
xnor UO_2329 (O_2329,N_28324,N_28575);
xnor UO_2330 (O_2330,N_28115,N_28031);
or UO_2331 (O_2331,N_29249,N_29481);
nand UO_2332 (O_2332,N_29373,N_28289);
nor UO_2333 (O_2333,N_28872,N_28145);
and UO_2334 (O_2334,N_29789,N_28817);
nand UO_2335 (O_2335,N_28741,N_29446);
or UO_2336 (O_2336,N_28159,N_29973);
and UO_2337 (O_2337,N_29738,N_28998);
or UO_2338 (O_2338,N_29868,N_28058);
and UO_2339 (O_2339,N_29202,N_28530);
or UO_2340 (O_2340,N_29527,N_29368);
or UO_2341 (O_2341,N_28370,N_29751);
and UO_2342 (O_2342,N_28942,N_29093);
xor UO_2343 (O_2343,N_29113,N_29185);
nand UO_2344 (O_2344,N_28187,N_28712);
xor UO_2345 (O_2345,N_29597,N_29055);
xor UO_2346 (O_2346,N_29638,N_29251);
nor UO_2347 (O_2347,N_29325,N_28462);
or UO_2348 (O_2348,N_29083,N_29765);
xnor UO_2349 (O_2349,N_28054,N_29879);
and UO_2350 (O_2350,N_29691,N_29463);
or UO_2351 (O_2351,N_28716,N_28864);
nand UO_2352 (O_2352,N_28147,N_29401);
nor UO_2353 (O_2353,N_29967,N_29866);
and UO_2354 (O_2354,N_29943,N_29406);
and UO_2355 (O_2355,N_28687,N_28110);
nor UO_2356 (O_2356,N_29009,N_29325);
xor UO_2357 (O_2357,N_29547,N_29356);
xor UO_2358 (O_2358,N_29500,N_28651);
nand UO_2359 (O_2359,N_28141,N_28934);
nor UO_2360 (O_2360,N_29726,N_29934);
nand UO_2361 (O_2361,N_28375,N_29918);
nand UO_2362 (O_2362,N_28508,N_29435);
nor UO_2363 (O_2363,N_28735,N_28374);
xor UO_2364 (O_2364,N_29246,N_29609);
and UO_2365 (O_2365,N_28985,N_29642);
or UO_2366 (O_2366,N_28958,N_28139);
and UO_2367 (O_2367,N_29225,N_29769);
nor UO_2368 (O_2368,N_29182,N_28427);
and UO_2369 (O_2369,N_28830,N_29385);
or UO_2370 (O_2370,N_28179,N_28957);
nor UO_2371 (O_2371,N_29172,N_29595);
nor UO_2372 (O_2372,N_29320,N_29824);
or UO_2373 (O_2373,N_28131,N_28027);
and UO_2374 (O_2374,N_29257,N_28278);
nor UO_2375 (O_2375,N_29935,N_29623);
or UO_2376 (O_2376,N_29899,N_29382);
or UO_2377 (O_2377,N_29707,N_29899);
nand UO_2378 (O_2378,N_29736,N_29184);
nor UO_2379 (O_2379,N_29099,N_28421);
or UO_2380 (O_2380,N_28029,N_28188);
nor UO_2381 (O_2381,N_29448,N_28451);
nor UO_2382 (O_2382,N_29719,N_28135);
xor UO_2383 (O_2383,N_29204,N_28274);
nand UO_2384 (O_2384,N_28587,N_29617);
nand UO_2385 (O_2385,N_29276,N_28414);
or UO_2386 (O_2386,N_28441,N_29935);
xor UO_2387 (O_2387,N_28506,N_28747);
nor UO_2388 (O_2388,N_29995,N_29368);
and UO_2389 (O_2389,N_28692,N_28094);
nand UO_2390 (O_2390,N_28462,N_28313);
and UO_2391 (O_2391,N_28525,N_29625);
nor UO_2392 (O_2392,N_29845,N_29858);
nand UO_2393 (O_2393,N_28075,N_28992);
nor UO_2394 (O_2394,N_29942,N_28392);
xor UO_2395 (O_2395,N_29449,N_29438);
nor UO_2396 (O_2396,N_29891,N_28551);
or UO_2397 (O_2397,N_29406,N_29224);
xor UO_2398 (O_2398,N_28884,N_28982);
xnor UO_2399 (O_2399,N_29531,N_29359);
nor UO_2400 (O_2400,N_28782,N_28022);
nor UO_2401 (O_2401,N_29733,N_28054);
and UO_2402 (O_2402,N_28577,N_28015);
xnor UO_2403 (O_2403,N_28948,N_28094);
nor UO_2404 (O_2404,N_28901,N_29325);
nand UO_2405 (O_2405,N_29359,N_28327);
xnor UO_2406 (O_2406,N_28386,N_28260);
nand UO_2407 (O_2407,N_28754,N_29126);
nor UO_2408 (O_2408,N_28061,N_28748);
xor UO_2409 (O_2409,N_29989,N_29314);
nor UO_2410 (O_2410,N_28969,N_28525);
nor UO_2411 (O_2411,N_28576,N_28262);
nand UO_2412 (O_2412,N_28270,N_29077);
nand UO_2413 (O_2413,N_29865,N_29784);
and UO_2414 (O_2414,N_28863,N_28709);
nor UO_2415 (O_2415,N_29073,N_28474);
or UO_2416 (O_2416,N_29778,N_28887);
and UO_2417 (O_2417,N_28994,N_29194);
nand UO_2418 (O_2418,N_28945,N_28260);
xnor UO_2419 (O_2419,N_29245,N_29012);
and UO_2420 (O_2420,N_29001,N_29775);
xor UO_2421 (O_2421,N_29724,N_29424);
xnor UO_2422 (O_2422,N_29227,N_29590);
and UO_2423 (O_2423,N_28943,N_28828);
or UO_2424 (O_2424,N_29633,N_29450);
and UO_2425 (O_2425,N_29950,N_28057);
or UO_2426 (O_2426,N_28231,N_29821);
and UO_2427 (O_2427,N_29710,N_28550);
and UO_2428 (O_2428,N_28263,N_28128);
nand UO_2429 (O_2429,N_28788,N_28075);
and UO_2430 (O_2430,N_28698,N_29251);
xnor UO_2431 (O_2431,N_29430,N_28997);
nand UO_2432 (O_2432,N_28312,N_28175);
or UO_2433 (O_2433,N_29219,N_28561);
nor UO_2434 (O_2434,N_28647,N_28122);
nor UO_2435 (O_2435,N_29815,N_29873);
nand UO_2436 (O_2436,N_28328,N_29697);
nor UO_2437 (O_2437,N_28528,N_29327);
nor UO_2438 (O_2438,N_28515,N_28268);
xor UO_2439 (O_2439,N_29352,N_29578);
and UO_2440 (O_2440,N_28823,N_29687);
xnor UO_2441 (O_2441,N_29862,N_28772);
xor UO_2442 (O_2442,N_29964,N_28552);
or UO_2443 (O_2443,N_29461,N_29212);
or UO_2444 (O_2444,N_29331,N_28456);
xor UO_2445 (O_2445,N_29359,N_29566);
nand UO_2446 (O_2446,N_28949,N_29054);
nand UO_2447 (O_2447,N_29894,N_29743);
nand UO_2448 (O_2448,N_28113,N_28728);
xnor UO_2449 (O_2449,N_29758,N_29226);
and UO_2450 (O_2450,N_29596,N_29433);
and UO_2451 (O_2451,N_29324,N_28191);
xor UO_2452 (O_2452,N_28994,N_29300);
or UO_2453 (O_2453,N_29409,N_29210);
and UO_2454 (O_2454,N_29638,N_28402);
or UO_2455 (O_2455,N_29445,N_29906);
or UO_2456 (O_2456,N_29224,N_29540);
or UO_2457 (O_2457,N_28275,N_29507);
or UO_2458 (O_2458,N_28191,N_28470);
or UO_2459 (O_2459,N_28056,N_28205);
nand UO_2460 (O_2460,N_29219,N_29401);
xnor UO_2461 (O_2461,N_28851,N_28765);
or UO_2462 (O_2462,N_29957,N_28073);
or UO_2463 (O_2463,N_29165,N_28944);
nor UO_2464 (O_2464,N_29586,N_29599);
or UO_2465 (O_2465,N_29522,N_28169);
nand UO_2466 (O_2466,N_28801,N_28293);
nand UO_2467 (O_2467,N_29232,N_28540);
nand UO_2468 (O_2468,N_29826,N_28403);
nor UO_2469 (O_2469,N_29008,N_29391);
nand UO_2470 (O_2470,N_29337,N_29447);
nand UO_2471 (O_2471,N_29921,N_29581);
nand UO_2472 (O_2472,N_28790,N_29269);
nor UO_2473 (O_2473,N_28885,N_28775);
and UO_2474 (O_2474,N_29426,N_29933);
and UO_2475 (O_2475,N_29333,N_28107);
or UO_2476 (O_2476,N_29819,N_29439);
xnor UO_2477 (O_2477,N_29760,N_29342);
nor UO_2478 (O_2478,N_29844,N_28962);
or UO_2479 (O_2479,N_29325,N_28063);
and UO_2480 (O_2480,N_28442,N_29110);
or UO_2481 (O_2481,N_28952,N_28408);
xor UO_2482 (O_2482,N_28154,N_29329);
or UO_2483 (O_2483,N_29940,N_29908);
xnor UO_2484 (O_2484,N_29069,N_29465);
nand UO_2485 (O_2485,N_29193,N_29788);
nand UO_2486 (O_2486,N_28169,N_29660);
nor UO_2487 (O_2487,N_29056,N_28358);
nand UO_2488 (O_2488,N_29690,N_28847);
nand UO_2489 (O_2489,N_29459,N_28706);
nand UO_2490 (O_2490,N_28272,N_28586);
and UO_2491 (O_2491,N_28790,N_29819);
xor UO_2492 (O_2492,N_28553,N_28584);
nor UO_2493 (O_2493,N_28157,N_29761);
or UO_2494 (O_2494,N_28735,N_29442);
and UO_2495 (O_2495,N_29065,N_28026);
nand UO_2496 (O_2496,N_29486,N_28582);
nor UO_2497 (O_2497,N_29492,N_29163);
and UO_2498 (O_2498,N_29965,N_29825);
and UO_2499 (O_2499,N_29188,N_28885);
and UO_2500 (O_2500,N_28628,N_28341);
xnor UO_2501 (O_2501,N_28009,N_29965);
xor UO_2502 (O_2502,N_29934,N_29820);
or UO_2503 (O_2503,N_28747,N_29495);
or UO_2504 (O_2504,N_28606,N_28809);
nor UO_2505 (O_2505,N_29495,N_28228);
or UO_2506 (O_2506,N_28892,N_29724);
nand UO_2507 (O_2507,N_28660,N_29668);
nand UO_2508 (O_2508,N_28762,N_28508);
and UO_2509 (O_2509,N_28861,N_29955);
or UO_2510 (O_2510,N_28644,N_29466);
nand UO_2511 (O_2511,N_28171,N_29818);
nand UO_2512 (O_2512,N_29954,N_29139);
nand UO_2513 (O_2513,N_28371,N_28027);
nand UO_2514 (O_2514,N_29864,N_29748);
or UO_2515 (O_2515,N_29160,N_29720);
and UO_2516 (O_2516,N_28760,N_28964);
and UO_2517 (O_2517,N_28681,N_28207);
nand UO_2518 (O_2518,N_28416,N_29549);
nand UO_2519 (O_2519,N_29800,N_28248);
nand UO_2520 (O_2520,N_28540,N_29348);
xor UO_2521 (O_2521,N_28894,N_29553);
and UO_2522 (O_2522,N_28897,N_28081);
nand UO_2523 (O_2523,N_29994,N_29087);
and UO_2524 (O_2524,N_29646,N_28660);
nor UO_2525 (O_2525,N_28363,N_29593);
or UO_2526 (O_2526,N_29559,N_28841);
or UO_2527 (O_2527,N_29834,N_28882);
nand UO_2528 (O_2528,N_28923,N_28084);
nor UO_2529 (O_2529,N_28245,N_28415);
nand UO_2530 (O_2530,N_28708,N_28833);
and UO_2531 (O_2531,N_28752,N_29065);
xor UO_2532 (O_2532,N_28431,N_29222);
xor UO_2533 (O_2533,N_29276,N_28658);
and UO_2534 (O_2534,N_29361,N_29704);
nand UO_2535 (O_2535,N_28219,N_28210);
nor UO_2536 (O_2536,N_28380,N_29345);
nand UO_2537 (O_2537,N_29277,N_28919);
or UO_2538 (O_2538,N_29754,N_29357);
and UO_2539 (O_2539,N_29973,N_29535);
xnor UO_2540 (O_2540,N_29759,N_29439);
or UO_2541 (O_2541,N_28819,N_29938);
or UO_2542 (O_2542,N_28943,N_29254);
xor UO_2543 (O_2543,N_28033,N_28693);
nor UO_2544 (O_2544,N_29075,N_28690);
nor UO_2545 (O_2545,N_29598,N_29235);
nor UO_2546 (O_2546,N_29563,N_29097);
xnor UO_2547 (O_2547,N_28862,N_28007);
nand UO_2548 (O_2548,N_28039,N_29227);
nor UO_2549 (O_2549,N_28600,N_28931);
xor UO_2550 (O_2550,N_28689,N_28576);
nand UO_2551 (O_2551,N_28314,N_29550);
or UO_2552 (O_2552,N_28519,N_29881);
nor UO_2553 (O_2553,N_28541,N_28711);
nor UO_2554 (O_2554,N_29444,N_29923);
nor UO_2555 (O_2555,N_29620,N_29857);
nand UO_2556 (O_2556,N_29992,N_28823);
xor UO_2557 (O_2557,N_28846,N_28587);
or UO_2558 (O_2558,N_29293,N_29453);
xor UO_2559 (O_2559,N_29648,N_28189);
and UO_2560 (O_2560,N_29007,N_29933);
or UO_2561 (O_2561,N_28297,N_29361);
or UO_2562 (O_2562,N_28873,N_29856);
nor UO_2563 (O_2563,N_28155,N_29129);
and UO_2564 (O_2564,N_29584,N_29808);
or UO_2565 (O_2565,N_29449,N_29338);
nand UO_2566 (O_2566,N_28135,N_28993);
or UO_2567 (O_2567,N_29514,N_28041);
nor UO_2568 (O_2568,N_29002,N_29399);
xor UO_2569 (O_2569,N_28556,N_28596);
nor UO_2570 (O_2570,N_29432,N_28699);
or UO_2571 (O_2571,N_28647,N_29504);
xor UO_2572 (O_2572,N_29515,N_28586);
xor UO_2573 (O_2573,N_28616,N_28032);
xor UO_2574 (O_2574,N_28359,N_29084);
xnor UO_2575 (O_2575,N_28124,N_28356);
nor UO_2576 (O_2576,N_29357,N_29153);
or UO_2577 (O_2577,N_29259,N_29443);
and UO_2578 (O_2578,N_28227,N_28322);
nor UO_2579 (O_2579,N_29783,N_28693);
nor UO_2580 (O_2580,N_28744,N_28235);
nor UO_2581 (O_2581,N_28959,N_28518);
xor UO_2582 (O_2582,N_29458,N_29979);
and UO_2583 (O_2583,N_28187,N_28722);
or UO_2584 (O_2584,N_29655,N_28984);
xnor UO_2585 (O_2585,N_29374,N_29799);
xnor UO_2586 (O_2586,N_29257,N_28995);
xor UO_2587 (O_2587,N_29057,N_29340);
or UO_2588 (O_2588,N_29807,N_29050);
xor UO_2589 (O_2589,N_28859,N_29154);
xnor UO_2590 (O_2590,N_29408,N_28019);
and UO_2591 (O_2591,N_29827,N_29287);
nand UO_2592 (O_2592,N_28322,N_29045);
or UO_2593 (O_2593,N_29785,N_28041);
nand UO_2594 (O_2594,N_28495,N_29590);
nand UO_2595 (O_2595,N_29771,N_28664);
nor UO_2596 (O_2596,N_29017,N_29204);
xnor UO_2597 (O_2597,N_28226,N_29559);
and UO_2598 (O_2598,N_28668,N_29204);
and UO_2599 (O_2599,N_29475,N_29941);
or UO_2600 (O_2600,N_28678,N_28691);
nor UO_2601 (O_2601,N_28875,N_28255);
or UO_2602 (O_2602,N_28795,N_28646);
xnor UO_2603 (O_2603,N_28712,N_29929);
nand UO_2604 (O_2604,N_29421,N_28521);
xnor UO_2605 (O_2605,N_29476,N_28388);
or UO_2606 (O_2606,N_28837,N_29678);
and UO_2607 (O_2607,N_28039,N_28311);
nand UO_2608 (O_2608,N_28337,N_28478);
or UO_2609 (O_2609,N_29570,N_28503);
nor UO_2610 (O_2610,N_28549,N_28474);
xnor UO_2611 (O_2611,N_29771,N_29874);
xor UO_2612 (O_2612,N_28001,N_29683);
nor UO_2613 (O_2613,N_29595,N_28541);
nand UO_2614 (O_2614,N_28942,N_29348);
nor UO_2615 (O_2615,N_29724,N_28675);
and UO_2616 (O_2616,N_28347,N_28425);
or UO_2617 (O_2617,N_28887,N_29109);
xor UO_2618 (O_2618,N_28845,N_28986);
xnor UO_2619 (O_2619,N_29916,N_29317);
or UO_2620 (O_2620,N_29724,N_28541);
or UO_2621 (O_2621,N_29472,N_29321);
and UO_2622 (O_2622,N_29690,N_28967);
nand UO_2623 (O_2623,N_29614,N_28027);
and UO_2624 (O_2624,N_29151,N_29661);
and UO_2625 (O_2625,N_29295,N_28081);
nand UO_2626 (O_2626,N_29016,N_28320);
nand UO_2627 (O_2627,N_28215,N_29221);
or UO_2628 (O_2628,N_28501,N_29158);
nor UO_2629 (O_2629,N_28591,N_28210);
nor UO_2630 (O_2630,N_29796,N_28211);
nor UO_2631 (O_2631,N_29286,N_28225);
nor UO_2632 (O_2632,N_29377,N_29210);
nand UO_2633 (O_2633,N_29029,N_28061);
xnor UO_2634 (O_2634,N_29121,N_28676);
and UO_2635 (O_2635,N_29593,N_28596);
or UO_2636 (O_2636,N_29653,N_28778);
or UO_2637 (O_2637,N_29625,N_29394);
or UO_2638 (O_2638,N_28083,N_28539);
or UO_2639 (O_2639,N_28680,N_28962);
nand UO_2640 (O_2640,N_28528,N_29510);
and UO_2641 (O_2641,N_28649,N_28628);
xnor UO_2642 (O_2642,N_28017,N_28555);
and UO_2643 (O_2643,N_29254,N_29744);
and UO_2644 (O_2644,N_29364,N_29582);
or UO_2645 (O_2645,N_29004,N_29233);
xnor UO_2646 (O_2646,N_29744,N_28931);
nor UO_2647 (O_2647,N_28067,N_29176);
nor UO_2648 (O_2648,N_28445,N_29071);
nand UO_2649 (O_2649,N_29208,N_28711);
or UO_2650 (O_2650,N_29567,N_28972);
nor UO_2651 (O_2651,N_29493,N_28703);
nor UO_2652 (O_2652,N_29046,N_28400);
or UO_2653 (O_2653,N_28738,N_29308);
nand UO_2654 (O_2654,N_29141,N_28110);
nand UO_2655 (O_2655,N_28001,N_29937);
nor UO_2656 (O_2656,N_29000,N_28315);
nand UO_2657 (O_2657,N_29929,N_29768);
nand UO_2658 (O_2658,N_29421,N_28324);
nor UO_2659 (O_2659,N_29513,N_29751);
nand UO_2660 (O_2660,N_28911,N_29121);
xor UO_2661 (O_2661,N_29804,N_28972);
xor UO_2662 (O_2662,N_29719,N_29332);
nand UO_2663 (O_2663,N_29849,N_28963);
nor UO_2664 (O_2664,N_28686,N_28254);
nor UO_2665 (O_2665,N_28932,N_29390);
and UO_2666 (O_2666,N_29189,N_29453);
nor UO_2667 (O_2667,N_29350,N_28423);
nand UO_2668 (O_2668,N_29397,N_29940);
and UO_2669 (O_2669,N_29094,N_29261);
nor UO_2670 (O_2670,N_29878,N_29277);
xnor UO_2671 (O_2671,N_28690,N_29920);
or UO_2672 (O_2672,N_29186,N_29308);
nor UO_2673 (O_2673,N_29837,N_29202);
nand UO_2674 (O_2674,N_29939,N_29296);
xor UO_2675 (O_2675,N_28810,N_28356);
nand UO_2676 (O_2676,N_28148,N_28008);
nand UO_2677 (O_2677,N_29490,N_28125);
and UO_2678 (O_2678,N_28815,N_28439);
or UO_2679 (O_2679,N_28614,N_28750);
xor UO_2680 (O_2680,N_29505,N_29286);
xor UO_2681 (O_2681,N_28849,N_29531);
nand UO_2682 (O_2682,N_29500,N_29710);
and UO_2683 (O_2683,N_29144,N_29008);
nor UO_2684 (O_2684,N_29653,N_28567);
nand UO_2685 (O_2685,N_28831,N_29247);
xor UO_2686 (O_2686,N_29149,N_28130);
and UO_2687 (O_2687,N_29851,N_29396);
nand UO_2688 (O_2688,N_29325,N_28825);
or UO_2689 (O_2689,N_29896,N_29883);
or UO_2690 (O_2690,N_28990,N_28402);
xor UO_2691 (O_2691,N_28682,N_28946);
nand UO_2692 (O_2692,N_29726,N_29746);
nand UO_2693 (O_2693,N_29662,N_28789);
nand UO_2694 (O_2694,N_29154,N_28952);
nor UO_2695 (O_2695,N_28626,N_28383);
or UO_2696 (O_2696,N_29467,N_28689);
nor UO_2697 (O_2697,N_28101,N_28130);
xnor UO_2698 (O_2698,N_29117,N_29558);
or UO_2699 (O_2699,N_28766,N_29601);
xnor UO_2700 (O_2700,N_28957,N_29412);
and UO_2701 (O_2701,N_28383,N_29941);
nor UO_2702 (O_2702,N_29049,N_28098);
nand UO_2703 (O_2703,N_28254,N_29467);
or UO_2704 (O_2704,N_28553,N_28389);
or UO_2705 (O_2705,N_29548,N_29772);
and UO_2706 (O_2706,N_28247,N_28866);
and UO_2707 (O_2707,N_29585,N_28109);
xor UO_2708 (O_2708,N_29216,N_29808);
or UO_2709 (O_2709,N_28647,N_29225);
and UO_2710 (O_2710,N_29602,N_28366);
xor UO_2711 (O_2711,N_28409,N_28582);
nand UO_2712 (O_2712,N_28515,N_28498);
nand UO_2713 (O_2713,N_29374,N_28847);
nand UO_2714 (O_2714,N_28316,N_28933);
nand UO_2715 (O_2715,N_28097,N_28605);
and UO_2716 (O_2716,N_28947,N_29264);
or UO_2717 (O_2717,N_29690,N_28627);
nor UO_2718 (O_2718,N_28877,N_29183);
xnor UO_2719 (O_2719,N_28553,N_29795);
nor UO_2720 (O_2720,N_28412,N_29139);
nand UO_2721 (O_2721,N_29116,N_28086);
and UO_2722 (O_2722,N_28259,N_29026);
nand UO_2723 (O_2723,N_29679,N_29103);
or UO_2724 (O_2724,N_28463,N_29943);
and UO_2725 (O_2725,N_28450,N_28575);
nand UO_2726 (O_2726,N_28689,N_28881);
xor UO_2727 (O_2727,N_28854,N_28252);
xor UO_2728 (O_2728,N_29728,N_29192);
xor UO_2729 (O_2729,N_28559,N_28190);
xor UO_2730 (O_2730,N_29055,N_29957);
nor UO_2731 (O_2731,N_29688,N_28170);
or UO_2732 (O_2732,N_28481,N_28166);
and UO_2733 (O_2733,N_28625,N_28343);
xor UO_2734 (O_2734,N_28735,N_28028);
and UO_2735 (O_2735,N_29007,N_28699);
or UO_2736 (O_2736,N_28335,N_28707);
nand UO_2737 (O_2737,N_29208,N_28739);
nand UO_2738 (O_2738,N_29523,N_28028);
nor UO_2739 (O_2739,N_28269,N_29436);
and UO_2740 (O_2740,N_28335,N_28111);
nor UO_2741 (O_2741,N_29925,N_29000);
and UO_2742 (O_2742,N_28743,N_28403);
nor UO_2743 (O_2743,N_28711,N_28123);
and UO_2744 (O_2744,N_29753,N_28213);
xnor UO_2745 (O_2745,N_29095,N_28015);
or UO_2746 (O_2746,N_29669,N_29321);
nand UO_2747 (O_2747,N_29222,N_29470);
xor UO_2748 (O_2748,N_29924,N_29301);
nand UO_2749 (O_2749,N_28792,N_28525);
nand UO_2750 (O_2750,N_29839,N_29242);
nand UO_2751 (O_2751,N_28665,N_29503);
xnor UO_2752 (O_2752,N_28471,N_29979);
or UO_2753 (O_2753,N_28415,N_29940);
xnor UO_2754 (O_2754,N_28552,N_28587);
xor UO_2755 (O_2755,N_29884,N_29777);
or UO_2756 (O_2756,N_28513,N_29386);
xnor UO_2757 (O_2757,N_28145,N_29620);
and UO_2758 (O_2758,N_29588,N_29464);
nor UO_2759 (O_2759,N_28710,N_28789);
nor UO_2760 (O_2760,N_29403,N_29072);
nor UO_2761 (O_2761,N_28956,N_29890);
xor UO_2762 (O_2762,N_29654,N_29548);
xor UO_2763 (O_2763,N_29737,N_28150);
and UO_2764 (O_2764,N_28869,N_28483);
nand UO_2765 (O_2765,N_28891,N_29965);
nor UO_2766 (O_2766,N_29421,N_29686);
xor UO_2767 (O_2767,N_29204,N_29893);
xor UO_2768 (O_2768,N_29160,N_28247);
nand UO_2769 (O_2769,N_29234,N_29694);
nand UO_2770 (O_2770,N_28865,N_29476);
or UO_2771 (O_2771,N_28283,N_28511);
and UO_2772 (O_2772,N_28109,N_29440);
nor UO_2773 (O_2773,N_29360,N_29994);
and UO_2774 (O_2774,N_28059,N_29314);
or UO_2775 (O_2775,N_28396,N_28856);
xnor UO_2776 (O_2776,N_29814,N_29318);
nor UO_2777 (O_2777,N_28823,N_28995);
xnor UO_2778 (O_2778,N_28502,N_28673);
or UO_2779 (O_2779,N_29609,N_28425);
or UO_2780 (O_2780,N_29382,N_29618);
nor UO_2781 (O_2781,N_28473,N_29520);
nand UO_2782 (O_2782,N_28866,N_29334);
xor UO_2783 (O_2783,N_28169,N_29076);
nand UO_2784 (O_2784,N_28124,N_29344);
and UO_2785 (O_2785,N_28270,N_28345);
nand UO_2786 (O_2786,N_29631,N_29484);
and UO_2787 (O_2787,N_29188,N_29731);
nand UO_2788 (O_2788,N_28130,N_28981);
or UO_2789 (O_2789,N_29458,N_28595);
and UO_2790 (O_2790,N_28679,N_29597);
and UO_2791 (O_2791,N_29725,N_28179);
and UO_2792 (O_2792,N_29609,N_28562);
nor UO_2793 (O_2793,N_29917,N_29979);
nand UO_2794 (O_2794,N_28984,N_29685);
or UO_2795 (O_2795,N_28324,N_28376);
xnor UO_2796 (O_2796,N_28985,N_28257);
xnor UO_2797 (O_2797,N_29832,N_28641);
nand UO_2798 (O_2798,N_28456,N_28957);
and UO_2799 (O_2799,N_29899,N_28200);
nand UO_2800 (O_2800,N_29657,N_29934);
nor UO_2801 (O_2801,N_28224,N_29692);
nand UO_2802 (O_2802,N_29827,N_28658);
or UO_2803 (O_2803,N_29809,N_29624);
and UO_2804 (O_2804,N_29922,N_28189);
nand UO_2805 (O_2805,N_28369,N_29837);
or UO_2806 (O_2806,N_28358,N_28033);
nand UO_2807 (O_2807,N_29964,N_29732);
nand UO_2808 (O_2808,N_29378,N_28839);
nor UO_2809 (O_2809,N_28768,N_29229);
and UO_2810 (O_2810,N_28780,N_28174);
and UO_2811 (O_2811,N_28042,N_28293);
xor UO_2812 (O_2812,N_28270,N_29214);
xnor UO_2813 (O_2813,N_29258,N_29880);
nand UO_2814 (O_2814,N_28857,N_29142);
or UO_2815 (O_2815,N_28606,N_29188);
xor UO_2816 (O_2816,N_28156,N_28885);
or UO_2817 (O_2817,N_28194,N_29644);
xor UO_2818 (O_2818,N_28214,N_29835);
and UO_2819 (O_2819,N_28295,N_28741);
xor UO_2820 (O_2820,N_28171,N_29115);
nor UO_2821 (O_2821,N_28770,N_29158);
nand UO_2822 (O_2822,N_28871,N_28346);
nor UO_2823 (O_2823,N_29827,N_29695);
or UO_2824 (O_2824,N_29722,N_28759);
or UO_2825 (O_2825,N_29954,N_28574);
nand UO_2826 (O_2826,N_28133,N_29020);
or UO_2827 (O_2827,N_29913,N_29263);
nor UO_2828 (O_2828,N_28709,N_29940);
and UO_2829 (O_2829,N_28493,N_28920);
and UO_2830 (O_2830,N_28050,N_28899);
xor UO_2831 (O_2831,N_29212,N_29752);
nand UO_2832 (O_2832,N_29872,N_28690);
xnor UO_2833 (O_2833,N_29338,N_29129);
or UO_2834 (O_2834,N_28521,N_28704);
xor UO_2835 (O_2835,N_28110,N_28156);
nor UO_2836 (O_2836,N_28749,N_28774);
and UO_2837 (O_2837,N_28792,N_29927);
xor UO_2838 (O_2838,N_28621,N_28177);
or UO_2839 (O_2839,N_28525,N_29763);
nand UO_2840 (O_2840,N_29173,N_29442);
or UO_2841 (O_2841,N_29177,N_28009);
nand UO_2842 (O_2842,N_29061,N_29960);
xor UO_2843 (O_2843,N_29967,N_29425);
nand UO_2844 (O_2844,N_28615,N_28418);
xor UO_2845 (O_2845,N_28117,N_28530);
nor UO_2846 (O_2846,N_28889,N_28464);
and UO_2847 (O_2847,N_29203,N_28039);
and UO_2848 (O_2848,N_29656,N_29595);
nor UO_2849 (O_2849,N_28411,N_29176);
nor UO_2850 (O_2850,N_28804,N_29939);
or UO_2851 (O_2851,N_29360,N_29850);
nand UO_2852 (O_2852,N_29477,N_28477);
nor UO_2853 (O_2853,N_28483,N_29960);
nand UO_2854 (O_2854,N_29008,N_29822);
or UO_2855 (O_2855,N_28954,N_29722);
or UO_2856 (O_2856,N_28878,N_29062);
and UO_2857 (O_2857,N_29422,N_29005);
xnor UO_2858 (O_2858,N_28067,N_28140);
or UO_2859 (O_2859,N_29147,N_28812);
or UO_2860 (O_2860,N_29971,N_28672);
nand UO_2861 (O_2861,N_28934,N_29781);
xor UO_2862 (O_2862,N_29934,N_28288);
nand UO_2863 (O_2863,N_28439,N_29525);
or UO_2864 (O_2864,N_29933,N_28912);
nand UO_2865 (O_2865,N_29963,N_29399);
nand UO_2866 (O_2866,N_29656,N_28842);
nor UO_2867 (O_2867,N_29258,N_28357);
and UO_2868 (O_2868,N_28753,N_28102);
nand UO_2869 (O_2869,N_28105,N_29332);
and UO_2870 (O_2870,N_28513,N_28381);
nor UO_2871 (O_2871,N_28885,N_29379);
nand UO_2872 (O_2872,N_28512,N_29498);
nor UO_2873 (O_2873,N_28003,N_28564);
nand UO_2874 (O_2874,N_29477,N_29774);
nor UO_2875 (O_2875,N_28501,N_28277);
or UO_2876 (O_2876,N_29279,N_28165);
nor UO_2877 (O_2877,N_28023,N_28473);
nor UO_2878 (O_2878,N_28819,N_29730);
and UO_2879 (O_2879,N_29148,N_29342);
and UO_2880 (O_2880,N_29501,N_28949);
or UO_2881 (O_2881,N_29561,N_29334);
nand UO_2882 (O_2882,N_29481,N_28397);
nor UO_2883 (O_2883,N_29681,N_29037);
or UO_2884 (O_2884,N_29623,N_29600);
and UO_2885 (O_2885,N_28907,N_29246);
nor UO_2886 (O_2886,N_28147,N_28779);
and UO_2887 (O_2887,N_29492,N_28082);
xnor UO_2888 (O_2888,N_28571,N_28495);
or UO_2889 (O_2889,N_29948,N_28103);
xnor UO_2890 (O_2890,N_28453,N_28165);
xor UO_2891 (O_2891,N_29965,N_29476);
or UO_2892 (O_2892,N_29941,N_29875);
nor UO_2893 (O_2893,N_29780,N_28129);
and UO_2894 (O_2894,N_28587,N_28321);
or UO_2895 (O_2895,N_28418,N_28276);
nand UO_2896 (O_2896,N_29623,N_28864);
nor UO_2897 (O_2897,N_29778,N_29311);
nand UO_2898 (O_2898,N_29889,N_29242);
nor UO_2899 (O_2899,N_29594,N_29343);
and UO_2900 (O_2900,N_28590,N_28389);
or UO_2901 (O_2901,N_28471,N_29014);
or UO_2902 (O_2902,N_28888,N_28268);
and UO_2903 (O_2903,N_28461,N_29853);
nand UO_2904 (O_2904,N_29967,N_28747);
nand UO_2905 (O_2905,N_28101,N_28749);
nor UO_2906 (O_2906,N_29102,N_28807);
nor UO_2907 (O_2907,N_29695,N_28260);
xor UO_2908 (O_2908,N_29946,N_29131);
nor UO_2909 (O_2909,N_29605,N_29575);
nand UO_2910 (O_2910,N_28129,N_29849);
nand UO_2911 (O_2911,N_29547,N_28027);
nor UO_2912 (O_2912,N_29705,N_29965);
xor UO_2913 (O_2913,N_29419,N_28868);
or UO_2914 (O_2914,N_29755,N_29162);
and UO_2915 (O_2915,N_29500,N_28358);
xnor UO_2916 (O_2916,N_29737,N_28372);
and UO_2917 (O_2917,N_29019,N_29501);
and UO_2918 (O_2918,N_28009,N_29499);
nor UO_2919 (O_2919,N_28660,N_29164);
nor UO_2920 (O_2920,N_29754,N_29184);
or UO_2921 (O_2921,N_28410,N_28390);
nand UO_2922 (O_2922,N_29630,N_29026);
xor UO_2923 (O_2923,N_29093,N_29597);
and UO_2924 (O_2924,N_29834,N_28436);
and UO_2925 (O_2925,N_29617,N_28983);
or UO_2926 (O_2926,N_29486,N_28584);
and UO_2927 (O_2927,N_29240,N_28950);
or UO_2928 (O_2928,N_29096,N_29830);
nand UO_2929 (O_2929,N_28414,N_29911);
nor UO_2930 (O_2930,N_28453,N_29818);
nor UO_2931 (O_2931,N_29123,N_29796);
and UO_2932 (O_2932,N_29215,N_28456);
and UO_2933 (O_2933,N_28096,N_29917);
xnor UO_2934 (O_2934,N_28834,N_28201);
nand UO_2935 (O_2935,N_29346,N_28002);
nor UO_2936 (O_2936,N_29249,N_28131);
xnor UO_2937 (O_2937,N_28636,N_29299);
nor UO_2938 (O_2938,N_28022,N_28839);
or UO_2939 (O_2939,N_28357,N_29437);
nand UO_2940 (O_2940,N_29379,N_28967);
and UO_2941 (O_2941,N_29109,N_28171);
nand UO_2942 (O_2942,N_29961,N_29560);
xnor UO_2943 (O_2943,N_28584,N_28438);
or UO_2944 (O_2944,N_28027,N_28458);
or UO_2945 (O_2945,N_29749,N_29279);
nand UO_2946 (O_2946,N_29097,N_28402);
xor UO_2947 (O_2947,N_29308,N_29893);
or UO_2948 (O_2948,N_28996,N_29191);
and UO_2949 (O_2949,N_29735,N_28241);
xnor UO_2950 (O_2950,N_28105,N_28283);
nor UO_2951 (O_2951,N_29314,N_29449);
and UO_2952 (O_2952,N_28865,N_29631);
and UO_2953 (O_2953,N_28464,N_28610);
nor UO_2954 (O_2954,N_29788,N_28638);
xnor UO_2955 (O_2955,N_29121,N_28276);
xnor UO_2956 (O_2956,N_28891,N_29840);
and UO_2957 (O_2957,N_28356,N_28558);
and UO_2958 (O_2958,N_29556,N_29732);
and UO_2959 (O_2959,N_29273,N_29770);
xnor UO_2960 (O_2960,N_29527,N_28779);
or UO_2961 (O_2961,N_28423,N_28705);
nor UO_2962 (O_2962,N_29773,N_28975);
or UO_2963 (O_2963,N_28259,N_28959);
xnor UO_2964 (O_2964,N_29486,N_29347);
or UO_2965 (O_2965,N_29681,N_28025);
nand UO_2966 (O_2966,N_29780,N_28883);
and UO_2967 (O_2967,N_29400,N_29573);
and UO_2968 (O_2968,N_29459,N_29153);
nand UO_2969 (O_2969,N_29174,N_28035);
nor UO_2970 (O_2970,N_29662,N_28186);
and UO_2971 (O_2971,N_28512,N_28026);
nand UO_2972 (O_2972,N_29359,N_28689);
nor UO_2973 (O_2973,N_29516,N_28245);
nor UO_2974 (O_2974,N_28489,N_29621);
nand UO_2975 (O_2975,N_29669,N_28876);
nand UO_2976 (O_2976,N_29112,N_28174);
xor UO_2977 (O_2977,N_28198,N_29016);
nand UO_2978 (O_2978,N_29551,N_29265);
and UO_2979 (O_2979,N_29350,N_28477);
xor UO_2980 (O_2980,N_28090,N_29891);
nand UO_2981 (O_2981,N_28908,N_29391);
nor UO_2982 (O_2982,N_29996,N_29490);
xnor UO_2983 (O_2983,N_28965,N_29232);
and UO_2984 (O_2984,N_28690,N_29747);
or UO_2985 (O_2985,N_29377,N_29739);
nor UO_2986 (O_2986,N_28892,N_28951);
xor UO_2987 (O_2987,N_28229,N_29537);
and UO_2988 (O_2988,N_29845,N_29686);
and UO_2989 (O_2989,N_29589,N_28131);
and UO_2990 (O_2990,N_29999,N_28708);
and UO_2991 (O_2991,N_28774,N_29522);
nand UO_2992 (O_2992,N_29658,N_28326);
nor UO_2993 (O_2993,N_28874,N_29825);
xor UO_2994 (O_2994,N_29643,N_28417);
xnor UO_2995 (O_2995,N_28937,N_29235);
nor UO_2996 (O_2996,N_29738,N_29498);
and UO_2997 (O_2997,N_29227,N_28763);
xor UO_2998 (O_2998,N_29694,N_28101);
and UO_2999 (O_2999,N_28028,N_29192);
xor UO_3000 (O_3000,N_28590,N_28146);
nor UO_3001 (O_3001,N_28846,N_28615);
nor UO_3002 (O_3002,N_28884,N_29155);
or UO_3003 (O_3003,N_28005,N_29306);
nand UO_3004 (O_3004,N_29817,N_28876);
and UO_3005 (O_3005,N_28721,N_29047);
xnor UO_3006 (O_3006,N_28469,N_29438);
and UO_3007 (O_3007,N_28798,N_28124);
nor UO_3008 (O_3008,N_28344,N_29179);
or UO_3009 (O_3009,N_28449,N_29900);
and UO_3010 (O_3010,N_29729,N_29957);
nor UO_3011 (O_3011,N_28695,N_29434);
and UO_3012 (O_3012,N_28911,N_28566);
nor UO_3013 (O_3013,N_29989,N_29673);
and UO_3014 (O_3014,N_29784,N_28007);
and UO_3015 (O_3015,N_29196,N_28759);
xnor UO_3016 (O_3016,N_29756,N_28481);
nand UO_3017 (O_3017,N_29127,N_28931);
nor UO_3018 (O_3018,N_28778,N_28732);
nand UO_3019 (O_3019,N_28655,N_29839);
or UO_3020 (O_3020,N_29737,N_29220);
and UO_3021 (O_3021,N_28915,N_29388);
nand UO_3022 (O_3022,N_29466,N_29992);
nor UO_3023 (O_3023,N_29354,N_28977);
xnor UO_3024 (O_3024,N_28009,N_28730);
nand UO_3025 (O_3025,N_29010,N_29775);
nor UO_3026 (O_3026,N_28096,N_29937);
nand UO_3027 (O_3027,N_29179,N_29635);
or UO_3028 (O_3028,N_28630,N_29407);
nor UO_3029 (O_3029,N_29991,N_28876);
nor UO_3030 (O_3030,N_29797,N_28190);
nor UO_3031 (O_3031,N_28722,N_28342);
nor UO_3032 (O_3032,N_28966,N_28366);
or UO_3033 (O_3033,N_28939,N_29429);
nor UO_3034 (O_3034,N_28877,N_29565);
and UO_3035 (O_3035,N_28852,N_28298);
nand UO_3036 (O_3036,N_28567,N_29057);
xnor UO_3037 (O_3037,N_28845,N_29961);
or UO_3038 (O_3038,N_29873,N_29727);
or UO_3039 (O_3039,N_28308,N_28201);
xnor UO_3040 (O_3040,N_29033,N_29626);
nor UO_3041 (O_3041,N_29666,N_29767);
or UO_3042 (O_3042,N_29499,N_29370);
or UO_3043 (O_3043,N_28993,N_28970);
nor UO_3044 (O_3044,N_29678,N_28123);
nand UO_3045 (O_3045,N_28240,N_28984);
nor UO_3046 (O_3046,N_28919,N_29968);
and UO_3047 (O_3047,N_29803,N_29505);
nor UO_3048 (O_3048,N_28556,N_28150);
nand UO_3049 (O_3049,N_29754,N_29767);
or UO_3050 (O_3050,N_28585,N_28877);
nand UO_3051 (O_3051,N_28036,N_29111);
nor UO_3052 (O_3052,N_28938,N_29001);
xnor UO_3053 (O_3053,N_28581,N_29988);
xor UO_3054 (O_3054,N_28432,N_29358);
nor UO_3055 (O_3055,N_29354,N_29339);
or UO_3056 (O_3056,N_29422,N_29844);
or UO_3057 (O_3057,N_28143,N_29127);
nor UO_3058 (O_3058,N_29539,N_28451);
and UO_3059 (O_3059,N_29478,N_28409);
and UO_3060 (O_3060,N_28020,N_29832);
and UO_3061 (O_3061,N_29560,N_29817);
and UO_3062 (O_3062,N_28966,N_28752);
xor UO_3063 (O_3063,N_28046,N_28945);
or UO_3064 (O_3064,N_28902,N_29105);
xnor UO_3065 (O_3065,N_29299,N_28433);
xor UO_3066 (O_3066,N_29097,N_28687);
or UO_3067 (O_3067,N_28564,N_29395);
xor UO_3068 (O_3068,N_28796,N_28248);
nand UO_3069 (O_3069,N_29453,N_29696);
or UO_3070 (O_3070,N_29002,N_29743);
nor UO_3071 (O_3071,N_29852,N_28523);
xor UO_3072 (O_3072,N_29163,N_28145);
or UO_3073 (O_3073,N_28931,N_28623);
or UO_3074 (O_3074,N_28465,N_28840);
or UO_3075 (O_3075,N_28856,N_29490);
or UO_3076 (O_3076,N_29351,N_28440);
nor UO_3077 (O_3077,N_29243,N_29205);
or UO_3078 (O_3078,N_29922,N_29560);
or UO_3079 (O_3079,N_28356,N_29511);
nand UO_3080 (O_3080,N_28163,N_28476);
xor UO_3081 (O_3081,N_28930,N_28542);
or UO_3082 (O_3082,N_28726,N_29859);
nand UO_3083 (O_3083,N_28094,N_29250);
xnor UO_3084 (O_3084,N_29734,N_29354);
and UO_3085 (O_3085,N_28283,N_29233);
and UO_3086 (O_3086,N_28246,N_28260);
xnor UO_3087 (O_3087,N_28922,N_28243);
nor UO_3088 (O_3088,N_29732,N_28899);
or UO_3089 (O_3089,N_28422,N_28101);
nor UO_3090 (O_3090,N_29277,N_29779);
nor UO_3091 (O_3091,N_28844,N_29822);
nand UO_3092 (O_3092,N_29724,N_28076);
nor UO_3093 (O_3093,N_29267,N_29894);
xnor UO_3094 (O_3094,N_29151,N_29182);
nor UO_3095 (O_3095,N_28931,N_28832);
xnor UO_3096 (O_3096,N_28527,N_28764);
nand UO_3097 (O_3097,N_29710,N_28637);
nand UO_3098 (O_3098,N_28828,N_29289);
nor UO_3099 (O_3099,N_29138,N_29134);
nor UO_3100 (O_3100,N_29879,N_28496);
nor UO_3101 (O_3101,N_29303,N_29762);
and UO_3102 (O_3102,N_29958,N_28589);
nand UO_3103 (O_3103,N_29820,N_29195);
nand UO_3104 (O_3104,N_28490,N_28629);
nor UO_3105 (O_3105,N_28906,N_28604);
xnor UO_3106 (O_3106,N_28382,N_28013);
nor UO_3107 (O_3107,N_29605,N_29701);
nand UO_3108 (O_3108,N_29027,N_28012);
or UO_3109 (O_3109,N_28052,N_28604);
nor UO_3110 (O_3110,N_29394,N_28066);
nor UO_3111 (O_3111,N_29304,N_28788);
and UO_3112 (O_3112,N_29975,N_28559);
or UO_3113 (O_3113,N_29271,N_29479);
xor UO_3114 (O_3114,N_28326,N_29922);
nand UO_3115 (O_3115,N_29064,N_28556);
xor UO_3116 (O_3116,N_28471,N_28010);
xnor UO_3117 (O_3117,N_28026,N_29719);
and UO_3118 (O_3118,N_29043,N_29563);
or UO_3119 (O_3119,N_28650,N_28122);
nand UO_3120 (O_3120,N_28175,N_29472);
nand UO_3121 (O_3121,N_28644,N_29782);
nand UO_3122 (O_3122,N_29739,N_28449);
or UO_3123 (O_3123,N_28602,N_29682);
and UO_3124 (O_3124,N_29098,N_28383);
xnor UO_3125 (O_3125,N_28149,N_28661);
nor UO_3126 (O_3126,N_28221,N_28780);
or UO_3127 (O_3127,N_28139,N_28515);
nor UO_3128 (O_3128,N_28439,N_28650);
and UO_3129 (O_3129,N_29111,N_29594);
xnor UO_3130 (O_3130,N_28217,N_29703);
xor UO_3131 (O_3131,N_29243,N_28760);
or UO_3132 (O_3132,N_28525,N_28711);
or UO_3133 (O_3133,N_29238,N_28267);
nor UO_3134 (O_3134,N_28317,N_28139);
nor UO_3135 (O_3135,N_28091,N_29119);
nor UO_3136 (O_3136,N_28795,N_28558);
or UO_3137 (O_3137,N_28043,N_28460);
and UO_3138 (O_3138,N_28141,N_29122);
and UO_3139 (O_3139,N_28190,N_29460);
or UO_3140 (O_3140,N_29114,N_28453);
or UO_3141 (O_3141,N_29879,N_28516);
nand UO_3142 (O_3142,N_28205,N_28555);
nor UO_3143 (O_3143,N_29572,N_29107);
and UO_3144 (O_3144,N_28663,N_28325);
and UO_3145 (O_3145,N_29259,N_29389);
xnor UO_3146 (O_3146,N_28319,N_28534);
nand UO_3147 (O_3147,N_28489,N_29583);
nand UO_3148 (O_3148,N_28392,N_29738);
nand UO_3149 (O_3149,N_28432,N_28879);
and UO_3150 (O_3150,N_29643,N_28157);
nand UO_3151 (O_3151,N_28016,N_29785);
nor UO_3152 (O_3152,N_28150,N_29282);
xor UO_3153 (O_3153,N_28288,N_28935);
and UO_3154 (O_3154,N_28504,N_28701);
or UO_3155 (O_3155,N_29404,N_29326);
or UO_3156 (O_3156,N_29407,N_28572);
xnor UO_3157 (O_3157,N_28809,N_29169);
and UO_3158 (O_3158,N_28665,N_28173);
xor UO_3159 (O_3159,N_29109,N_28814);
or UO_3160 (O_3160,N_29538,N_29145);
nor UO_3161 (O_3161,N_29054,N_29234);
nor UO_3162 (O_3162,N_28048,N_29903);
nand UO_3163 (O_3163,N_28960,N_29992);
xnor UO_3164 (O_3164,N_29767,N_28007);
or UO_3165 (O_3165,N_29064,N_29691);
nand UO_3166 (O_3166,N_28301,N_28601);
xnor UO_3167 (O_3167,N_28526,N_29256);
xor UO_3168 (O_3168,N_28889,N_29929);
and UO_3169 (O_3169,N_29692,N_28427);
nor UO_3170 (O_3170,N_28478,N_29241);
or UO_3171 (O_3171,N_28244,N_28343);
nand UO_3172 (O_3172,N_28121,N_28950);
and UO_3173 (O_3173,N_29995,N_28550);
and UO_3174 (O_3174,N_29749,N_28105);
nand UO_3175 (O_3175,N_28636,N_28938);
xor UO_3176 (O_3176,N_28926,N_28710);
or UO_3177 (O_3177,N_29544,N_29890);
and UO_3178 (O_3178,N_29250,N_28848);
nor UO_3179 (O_3179,N_28255,N_28998);
or UO_3180 (O_3180,N_28487,N_28706);
xnor UO_3181 (O_3181,N_29662,N_28306);
nor UO_3182 (O_3182,N_28775,N_29669);
or UO_3183 (O_3183,N_29374,N_28534);
nand UO_3184 (O_3184,N_29277,N_29210);
or UO_3185 (O_3185,N_28592,N_29922);
nor UO_3186 (O_3186,N_28635,N_29934);
or UO_3187 (O_3187,N_29482,N_28990);
or UO_3188 (O_3188,N_29920,N_28755);
nand UO_3189 (O_3189,N_29678,N_29791);
nand UO_3190 (O_3190,N_28298,N_28492);
nor UO_3191 (O_3191,N_29993,N_29677);
and UO_3192 (O_3192,N_29008,N_29081);
nor UO_3193 (O_3193,N_28343,N_28819);
xor UO_3194 (O_3194,N_29388,N_28180);
nor UO_3195 (O_3195,N_28138,N_29442);
nor UO_3196 (O_3196,N_28581,N_28725);
and UO_3197 (O_3197,N_28527,N_29764);
and UO_3198 (O_3198,N_29888,N_28845);
and UO_3199 (O_3199,N_28050,N_28449);
nand UO_3200 (O_3200,N_29947,N_28441);
xnor UO_3201 (O_3201,N_29464,N_29815);
nand UO_3202 (O_3202,N_28700,N_28074);
or UO_3203 (O_3203,N_29855,N_29132);
nand UO_3204 (O_3204,N_28557,N_28577);
xor UO_3205 (O_3205,N_29656,N_28497);
nand UO_3206 (O_3206,N_28424,N_29341);
and UO_3207 (O_3207,N_28310,N_28374);
nor UO_3208 (O_3208,N_28111,N_29975);
and UO_3209 (O_3209,N_28069,N_28494);
xnor UO_3210 (O_3210,N_28525,N_28889);
nand UO_3211 (O_3211,N_28749,N_29298);
or UO_3212 (O_3212,N_29660,N_29272);
or UO_3213 (O_3213,N_29369,N_28168);
xor UO_3214 (O_3214,N_29763,N_29587);
and UO_3215 (O_3215,N_28393,N_29466);
nand UO_3216 (O_3216,N_29512,N_28813);
nor UO_3217 (O_3217,N_28340,N_29069);
xnor UO_3218 (O_3218,N_29174,N_29423);
or UO_3219 (O_3219,N_28422,N_28548);
nor UO_3220 (O_3220,N_29967,N_28265);
and UO_3221 (O_3221,N_29334,N_28862);
and UO_3222 (O_3222,N_29284,N_28632);
nand UO_3223 (O_3223,N_29146,N_29386);
nor UO_3224 (O_3224,N_28239,N_28482);
nand UO_3225 (O_3225,N_29292,N_28130);
nand UO_3226 (O_3226,N_29664,N_29047);
or UO_3227 (O_3227,N_29900,N_29654);
xnor UO_3228 (O_3228,N_28092,N_28498);
and UO_3229 (O_3229,N_29849,N_28793);
xnor UO_3230 (O_3230,N_29747,N_28142);
and UO_3231 (O_3231,N_29338,N_29754);
xnor UO_3232 (O_3232,N_29952,N_28046);
and UO_3233 (O_3233,N_29647,N_29749);
or UO_3234 (O_3234,N_28099,N_29837);
or UO_3235 (O_3235,N_29201,N_28109);
and UO_3236 (O_3236,N_29847,N_28327);
xnor UO_3237 (O_3237,N_29130,N_29190);
nor UO_3238 (O_3238,N_28431,N_28960);
nand UO_3239 (O_3239,N_29525,N_28003);
or UO_3240 (O_3240,N_29399,N_29248);
nor UO_3241 (O_3241,N_29655,N_29050);
or UO_3242 (O_3242,N_28688,N_28798);
nor UO_3243 (O_3243,N_29913,N_29458);
nor UO_3244 (O_3244,N_28502,N_29090);
and UO_3245 (O_3245,N_29153,N_28987);
nand UO_3246 (O_3246,N_29836,N_28442);
or UO_3247 (O_3247,N_28613,N_28168);
nor UO_3248 (O_3248,N_29932,N_29162);
nor UO_3249 (O_3249,N_29495,N_29310);
xor UO_3250 (O_3250,N_28513,N_29658);
or UO_3251 (O_3251,N_28585,N_29737);
and UO_3252 (O_3252,N_29625,N_28836);
and UO_3253 (O_3253,N_29605,N_29199);
xor UO_3254 (O_3254,N_29136,N_29878);
or UO_3255 (O_3255,N_28965,N_28687);
nor UO_3256 (O_3256,N_29268,N_28089);
xor UO_3257 (O_3257,N_28859,N_29291);
xor UO_3258 (O_3258,N_28425,N_29191);
and UO_3259 (O_3259,N_28631,N_29766);
and UO_3260 (O_3260,N_29075,N_28275);
nor UO_3261 (O_3261,N_28902,N_29450);
xnor UO_3262 (O_3262,N_28195,N_28588);
nand UO_3263 (O_3263,N_29916,N_29399);
nor UO_3264 (O_3264,N_28914,N_29631);
nand UO_3265 (O_3265,N_29160,N_28404);
nand UO_3266 (O_3266,N_29283,N_28079);
and UO_3267 (O_3267,N_29896,N_28813);
and UO_3268 (O_3268,N_29321,N_29682);
and UO_3269 (O_3269,N_29521,N_28813);
xor UO_3270 (O_3270,N_28236,N_29903);
and UO_3271 (O_3271,N_29319,N_29363);
xnor UO_3272 (O_3272,N_29425,N_29048);
nor UO_3273 (O_3273,N_28616,N_29879);
or UO_3274 (O_3274,N_29699,N_28574);
and UO_3275 (O_3275,N_28448,N_28965);
nor UO_3276 (O_3276,N_28276,N_28302);
or UO_3277 (O_3277,N_29744,N_28443);
xnor UO_3278 (O_3278,N_29958,N_28808);
nand UO_3279 (O_3279,N_29223,N_28266);
or UO_3280 (O_3280,N_29926,N_29893);
or UO_3281 (O_3281,N_28192,N_28273);
or UO_3282 (O_3282,N_29998,N_29356);
and UO_3283 (O_3283,N_28977,N_29369);
nand UO_3284 (O_3284,N_28259,N_29437);
or UO_3285 (O_3285,N_29460,N_29665);
nor UO_3286 (O_3286,N_28536,N_29013);
nor UO_3287 (O_3287,N_28294,N_28768);
nor UO_3288 (O_3288,N_28858,N_29963);
and UO_3289 (O_3289,N_29686,N_28671);
nand UO_3290 (O_3290,N_28155,N_28380);
and UO_3291 (O_3291,N_28784,N_29831);
and UO_3292 (O_3292,N_29337,N_28083);
and UO_3293 (O_3293,N_29483,N_29185);
and UO_3294 (O_3294,N_29961,N_29846);
nand UO_3295 (O_3295,N_29204,N_28948);
nand UO_3296 (O_3296,N_28732,N_28940);
xnor UO_3297 (O_3297,N_29223,N_29240);
nor UO_3298 (O_3298,N_28055,N_28986);
nand UO_3299 (O_3299,N_28917,N_29625);
and UO_3300 (O_3300,N_28475,N_29089);
nand UO_3301 (O_3301,N_29013,N_29079);
nand UO_3302 (O_3302,N_29266,N_28146);
nand UO_3303 (O_3303,N_29943,N_28397);
and UO_3304 (O_3304,N_28196,N_28348);
or UO_3305 (O_3305,N_28385,N_28967);
and UO_3306 (O_3306,N_29343,N_28882);
xnor UO_3307 (O_3307,N_28802,N_28588);
nand UO_3308 (O_3308,N_28556,N_28809);
nand UO_3309 (O_3309,N_29092,N_29629);
and UO_3310 (O_3310,N_29859,N_29722);
and UO_3311 (O_3311,N_28108,N_28061);
and UO_3312 (O_3312,N_28048,N_28021);
nor UO_3313 (O_3313,N_28248,N_28390);
or UO_3314 (O_3314,N_28317,N_29279);
and UO_3315 (O_3315,N_28271,N_28960);
and UO_3316 (O_3316,N_28979,N_29405);
and UO_3317 (O_3317,N_28362,N_28113);
and UO_3318 (O_3318,N_29294,N_29683);
xnor UO_3319 (O_3319,N_28410,N_28437);
xnor UO_3320 (O_3320,N_28509,N_28378);
nand UO_3321 (O_3321,N_29728,N_28031);
nand UO_3322 (O_3322,N_29423,N_29849);
and UO_3323 (O_3323,N_28987,N_29082);
nor UO_3324 (O_3324,N_29170,N_28525);
or UO_3325 (O_3325,N_29581,N_29097);
nand UO_3326 (O_3326,N_28980,N_28387);
xor UO_3327 (O_3327,N_29274,N_28943);
and UO_3328 (O_3328,N_29104,N_28710);
or UO_3329 (O_3329,N_29702,N_29783);
or UO_3330 (O_3330,N_29376,N_29994);
and UO_3331 (O_3331,N_29180,N_28118);
nand UO_3332 (O_3332,N_28008,N_28158);
nor UO_3333 (O_3333,N_29556,N_28856);
xor UO_3334 (O_3334,N_28914,N_28964);
and UO_3335 (O_3335,N_29880,N_28287);
and UO_3336 (O_3336,N_28873,N_29411);
nor UO_3337 (O_3337,N_28705,N_28934);
nor UO_3338 (O_3338,N_28263,N_28769);
or UO_3339 (O_3339,N_29669,N_29138);
nand UO_3340 (O_3340,N_29319,N_28841);
xor UO_3341 (O_3341,N_28275,N_29356);
and UO_3342 (O_3342,N_28728,N_28899);
or UO_3343 (O_3343,N_28333,N_29688);
xor UO_3344 (O_3344,N_29469,N_29672);
nand UO_3345 (O_3345,N_29500,N_29716);
nor UO_3346 (O_3346,N_29178,N_29227);
nand UO_3347 (O_3347,N_29993,N_28700);
nor UO_3348 (O_3348,N_28680,N_28920);
nor UO_3349 (O_3349,N_28623,N_28719);
xor UO_3350 (O_3350,N_28762,N_29218);
nand UO_3351 (O_3351,N_29139,N_29491);
nor UO_3352 (O_3352,N_28931,N_29148);
nand UO_3353 (O_3353,N_28543,N_28875);
xnor UO_3354 (O_3354,N_28185,N_28813);
nor UO_3355 (O_3355,N_28597,N_28910);
xnor UO_3356 (O_3356,N_28226,N_29130);
nor UO_3357 (O_3357,N_28491,N_29333);
and UO_3358 (O_3358,N_29723,N_28572);
nor UO_3359 (O_3359,N_29187,N_29918);
nand UO_3360 (O_3360,N_29793,N_29742);
xnor UO_3361 (O_3361,N_28456,N_29102);
and UO_3362 (O_3362,N_29562,N_29833);
nor UO_3363 (O_3363,N_28107,N_28991);
and UO_3364 (O_3364,N_28714,N_29482);
nand UO_3365 (O_3365,N_28066,N_28371);
nand UO_3366 (O_3366,N_28738,N_29829);
or UO_3367 (O_3367,N_29694,N_28637);
and UO_3368 (O_3368,N_29569,N_28211);
nand UO_3369 (O_3369,N_29578,N_29333);
and UO_3370 (O_3370,N_28096,N_28537);
nand UO_3371 (O_3371,N_29497,N_28851);
nand UO_3372 (O_3372,N_28263,N_28926);
xor UO_3373 (O_3373,N_28986,N_28299);
nand UO_3374 (O_3374,N_29631,N_29627);
or UO_3375 (O_3375,N_28920,N_29597);
nand UO_3376 (O_3376,N_28640,N_28300);
or UO_3377 (O_3377,N_28513,N_29676);
or UO_3378 (O_3378,N_28070,N_28722);
or UO_3379 (O_3379,N_29352,N_29109);
nor UO_3380 (O_3380,N_29846,N_29089);
or UO_3381 (O_3381,N_28866,N_28307);
nand UO_3382 (O_3382,N_28232,N_29880);
and UO_3383 (O_3383,N_29210,N_28187);
or UO_3384 (O_3384,N_28814,N_29312);
nand UO_3385 (O_3385,N_29995,N_28754);
nand UO_3386 (O_3386,N_29170,N_28703);
and UO_3387 (O_3387,N_29639,N_28363);
or UO_3388 (O_3388,N_29619,N_29967);
xor UO_3389 (O_3389,N_28615,N_29984);
or UO_3390 (O_3390,N_28248,N_28526);
nand UO_3391 (O_3391,N_28155,N_28334);
nand UO_3392 (O_3392,N_28821,N_29997);
and UO_3393 (O_3393,N_29605,N_28774);
xnor UO_3394 (O_3394,N_29614,N_28848);
xor UO_3395 (O_3395,N_29260,N_28888);
or UO_3396 (O_3396,N_29862,N_28881);
or UO_3397 (O_3397,N_28517,N_28336);
or UO_3398 (O_3398,N_29642,N_28106);
nor UO_3399 (O_3399,N_29570,N_28565);
nor UO_3400 (O_3400,N_29895,N_29628);
nor UO_3401 (O_3401,N_28092,N_29371);
and UO_3402 (O_3402,N_28230,N_28420);
and UO_3403 (O_3403,N_28638,N_29329);
xnor UO_3404 (O_3404,N_28409,N_29340);
or UO_3405 (O_3405,N_28977,N_28322);
or UO_3406 (O_3406,N_29422,N_29369);
or UO_3407 (O_3407,N_29002,N_29223);
or UO_3408 (O_3408,N_28716,N_29205);
and UO_3409 (O_3409,N_29185,N_28944);
nand UO_3410 (O_3410,N_29633,N_29155);
nand UO_3411 (O_3411,N_28540,N_29052);
nor UO_3412 (O_3412,N_29497,N_29762);
nor UO_3413 (O_3413,N_28432,N_29221);
nor UO_3414 (O_3414,N_29456,N_28040);
nand UO_3415 (O_3415,N_29516,N_28281);
nor UO_3416 (O_3416,N_29288,N_29591);
nor UO_3417 (O_3417,N_28381,N_28824);
and UO_3418 (O_3418,N_28302,N_29822);
xor UO_3419 (O_3419,N_28025,N_28777);
nor UO_3420 (O_3420,N_29953,N_29029);
and UO_3421 (O_3421,N_28472,N_28437);
or UO_3422 (O_3422,N_28606,N_28321);
and UO_3423 (O_3423,N_28380,N_29171);
or UO_3424 (O_3424,N_28723,N_28509);
nor UO_3425 (O_3425,N_29318,N_28788);
nor UO_3426 (O_3426,N_28935,N_28353);
xor UO_3427 (O_3427,N_28119,N_28497);
nand UO_3428 (O_3428,N_29812,N_29146);
and UO_3429 (O_3429,N_28010,N_28131);
and UO_3430 (O_3430,N_28699,N_29566);
or UO_3431 (O_3431,N_29958,N_29557);
nor UO_3432 (O_3432,N_28815,N_29440);
or UO_3433 (O_3433,N_28741,N_29300);
or UO_3434 (O_3434,N_29635,N_28561);
nand UO_3435 (O_3435,N_29193,N_28432);
nor UO_3436 (O_3436,N_28901,N_28290);
nor UO_3437 (O_3437,N_29476,N_29240);
or UO_3438 (O_3438,N_28318,N_29370);
nand UO_3439 (O_3439,N_28202,N_28081);
xor UO_3440 (O_3440,N_29297,N_28069);
nor UO_3441 (O_3441,N_28523,N_29929);
xor UO_3442 (O_3442,N_29724,N_28021);
and UO_3443 (O_3443,N_29052,N_28120);
xnor UO_3444 (O_3444,N_29104,N_28365);
xnor UO_3445 (O_3445,N_29016,N_28107);
nand UO_3446 (O_3446,N_29970,N_29372);
nor UO_3447 (O_3447,N_29208,N_29493);
xnor UO_3448 (O_3448,N_29656,N_29684);
xor UO_3449 (O_3449,N_28588,N_29108);
nor UO_3450 (O_3450,N_29265,N_28045);
nand UO_3451 (O_3451,N_28569,N_29796);
nand UO_3452 (O_3452,N_28915,N_29065);
or UO_3453 (O_3453,N_29267,N_29862);
or UO_3454 (O_3454,N_28932,N_28049);
and UO_3455 (O_3455,N_28185,N_28621);
xor UO_3456 (O_3456,N_28481,N_29142);
xor UO_3457 (O_3457,N_29528,N_29818);
nand UO_3458 (O_3458,N_29930,N_28728);
nand UO_3459 (O_3459,N_28427,N_29818);
and UO_3460 (O_3460,N_29793,N_29639);
xor UO_3461 (O_3461,N_29221,N_28891);
and UO_3462 (O_3462,N_28963,N_28407);
nand UO_3463 (O_3463,N_29026,N_28666);
xor UO_3464 (O_3464,N_28077,N_29456);
nor UO_3465 (O_3465,N_29097,N_29695);
nor UO_3466 (O_3466,N_28873,N_28536);
nor UO_3467 (O_3467,N_28959,N_28578);
nor UO_3468 (O_3468,N_28207,N_29654);
or UO_3469 (O_3469,N_28215,N_29948);
nor UO_3470 (O_3470,N_29934,N_29101);
nand UO_3471 (O_3471,N_28103,N_29951);
xor UO_3472 (O_3472,N_29734,N_29843);
and UO_3473 (O_3473,N_28024,N_28522);
or UO_3474 (O_3474,N_28150,N_29100);
and UO_3475 (O_3475,N_28272,N_29696);
or UO_3476 (O_3476,N_29530,N_29829);
or UO_3477 (O_3477,N_28130,N_29784);
nor UO_3478 (O_3478,N_28608,N_29939);
nor UO_3479 (O_3479,N_28121,N_28580);
nor UO_3480 (O_3480,N_28198,N_28127);
and UO_3481 (O_3481,N_28067,N_28709);
or UO_3482 (O_3482,N_28426,N_29390);
or UO_3483 (O_3483,N_29033,N_29942);
nand UO_3484 (O_3484,N_29261,N_28425);
nor UO_3485 (O_3485,N_28581,N_28848);
nor UO_3486 (O_3486,N_28236,N_29517);
nor UO_3487 (O_3487,N_29535,N_29031);
nand UO_3488 (O_3488,N_29696,N_29374);
and UO_3489 (O_3489,N_28116,N_29343);
nor UO_3490 (O_3490,N_29716,N_28475);
xnor UO_3491 (O_3491,N_28952,N_29665);
or UO_3492 (O_3492,N_28797,N_29443);
xor UO_3493 (O_3493,N_29799,N_28203);
and UO_3494 (O_3494,N_28823,N_28445);
or UO_3495 (O_3495,N_28816,N_28869);
or UO_3496 (O_3496,N_29438,N_29189);
and UO_3497 (O_3497,N_28021,N_28766);
xor UO_3498 (O_3498,N_28217,N_28862);
xor UO_3499 (O_3499,N_29436,N_29645);
endmodule