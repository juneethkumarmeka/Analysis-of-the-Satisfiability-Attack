module basic_1500_15000_2000_15_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1381,In_995);
nand U1 (N_1,In_665,In_537);
or U2 (N_2,In_1335,In_590);
nor U3 (N_3,In_92,In_229);
and U4 (N_4,In_1077,In_831);
nor U5 (N_5,In_425,In_918);
nor U6 (N_6,In_18,In_957);
and U7 (N_7,In_217,In_1113);
and U8 (N_8,In_1477,In_685);
nand U9 (N_9,In_1029,In_1331);
and U10 (N_10,In_1407,In_800);
xnor U11 (N_11,In_90,In_658);
xor U12 (N_12,In_112,In_477);
nand U13 (N_13,In_446,In_505);
nand U14 (N_14,In_78,In_419);
nand U15 (N_15,In_948,In_1124);
xor U16 (N_16,In_579,In_1071);
and U17 (N_17,In_539,In_25);
nand U18 (N_18,In_508,In_258);
nor U19 (N_19,In_1023,In_6);
or U20 (N_20,In_1020,In_306);
and U21 (N_21,In_808,In_615);
nor U22 (N_22,In_281,In_708);
xnor U23 (N_23,In_712,In_432);
or U24 (N_24,In_1248,In_383);
nand U25 (N_25,In_450,In_784);
and U26 (N_26,In_773,In_305);
xor U27 (N_27,In_710,In_749);
nor U28 (N_28,In_558,In_42);
nor U29 (N_29,In_168,In_1024);
or U30 (N_30,In_729,In_1106);
nand U31 (N_31,In_62,In_1281);
or U32 (N_32,In_805,In_1263);
xnor U33 (N_33,In_923,In_673);
and U34 (N_34,In_696,In_101);
nor U35 (N_35,In_719,In_867);
xnor U36 (N_36,In_460,In_843);
nand U37 (N_37,In_1090,In_1069);
nor U38 (N_38,In_1366,In_556);
nor U39 (N_39,In_553,In_1070);
xnor U40 (N_40,In_853,In_69);
and U41 (N_41,In_1437,In_41);
nand U42 (N_42,In_384,In_604);
and U43 (N_43,In_605,In_983);
and U44 (N_44,In_1093,In_565);
nor U45 (N_45,In_294,In_500);
nand U46 (N_46,In_375,In_836);
and U47 (N_47,In_1279,In_1210);
and U48 (N_48,In_1095,In_1296);
or U49 (N_49,In_910,In_531);
xnor U50 (N_50,In_895,In_1190);
and U51 (N_51,In_1392,In_801);
or U52 (N_52,In_1044,In_851);
nand U53 (N_53,In_886,In_462);
and U54 (N_54,In_322,In_880);
and U55 (N_55,In_1158,In_1267);
xnor U56 (N_56,In_23,In_1143);
xor U57 (N_57,In_823,In_405);
xor U58 (N_58,In_730,In_1235);
xor U59 (N_59,In_1048,In_635);
or U60 (N_60,In_1209,In_1138);
and U61 (N_61,In_1183,In_1394);
and U62 (N_62,In_706,In_1205);
nand U63 (N_63,In_1242,In_1174);
or U64 (N_64,In_950,In_1297);
xnor U65 (N_65,In_968,In_630);
or U66 (N_66,In_1012,In_507);
nor U67 (N_67,In_26,In_50);
and U68 (N_68,In_1160,In_793);
or U69 (N_69,In_1412,In_203);
nand U70 (N_70,In_687,In_978);
nor U71 (N_71,In_1232,In_1014);
xnor U72 (N_72,In_1206,In_755);
or U73 (N_73,In_1363,In_602);
and U74 (N_74,In_767,In_1162);
and U75 (N_75,In_1447,In_591);
or U76 (N_76,In_1184,In_1045);
and U77 (N_77,In_1416,In_27);
xnor U78 (N_78,In_574,In_457);
and U79 (N_79,In_702,In_1362);
or U80 (N_80,In_237,In_901);
and U81 (N_81,In_1096,In_1116);
nand U82 (N_82,In_377,In_109);
or U83 (N_83,In_942,In_88);
or U84 (N_84,In_741,In_881);
nor U85 (N_85,In_965,In_1457);
or U86 (N_86,In_796,In_1060);
nand U87 (N_87,In_1390,In_415);
nand U88 (N_88,In_1317,In_249);
nand U89 (N_89,In_699,In_642);
nand U90 (N_90,In_795,In_344);
nor U91 (N_91,In_1323,In_1038);
nand U92 (N_92,In_1130,In_182);
and U93 (N_93,In_1370,In_842);
and U94 (N_94,In_355,In_363);
and U95 (N_95,In_445,In_1291);
xor U96 (N_96,In_745,In_964);
xor U97 (N_97,In_728,In_868);
nor U98 (N_98,In_1334,In_548);
and U99 (N_99,In_386,In_198);
and U100 (N_100,In_94,In_854);
or U101 (N_101,In_1240,In_1223);
or U102 (N_102,In_649,In_1440);
nor U103 (N_103,In_1161,In_282);
xnor U104 (N_104,In_424,In_463);
nor U105 (N_105,In_686,In_739);
xor U106 (N_106,In_40,In_13);
nor U107 (N_107,In_396,In_291);
or U108 (N_108,In_1136,In_1236);
and U109 (N_109,In_85,In_871);
and U110 (N_110,In_847,In_572);
nand U111 (N_111,In_530,In_1298);
or U112 (N_112,In_1135,In_194);
nand U113 (N_113,In_285,In_102);
and U114 (N_114,In_1097,In_583);
nand U115 (N_115,In_212,In_131);
or U116 (N_116,In_1021,In_632);
xor U117 (N_117,In_452,In_1387);
or U118 (N_118,In_1483,In_753);
nor U119 (N_119,In_1204,In_1156);
nor U120 (N_120,In_925,In_533);
or U121 (N_121,In_411,In_916);
or U122 (N_122,In_1153,In_1046);
or U123 (N_123,In_1426,In_0);
or U124 (N_124,In_1377,In_662);
xnor U125 (N_125,In_585,In_147);
nor U126 (N_126,In_139,In_426);
nand U127 (N_127,In_311,In_1389);
and U128 (N_128,In_380,In_179);
nor U129 (N_129,In_1461,In_584);
nand U130 (N_130,In_466,In_276);
nor U131 (N_131,In_716,In_546);
or U132 (N_132,In_1163,In_1451);
xnor U133 (N_133,In_1428,In_1469);
xnor U134 (N_134,In_1121,In_816);
nor U135 (N_135,In_159,In_345);
and U136 (N_136,In_829,In_900);
or U137 (N_137,In_1167,In_811);
or U138 (N_138,In_161,In_905);
and U139 (N_139,In_492,In_813);
or U140 (N_140,In_888,In_87);
nand U141 (N_141,In_550,In_233);
xor U142 (N_142,In_1176,In_164);
xor U143 (N_143,In_664,In_19);
nand U144 (N_144,In_966,In_563);
or U145 (N_145,In_1127,In_731);
xor U146 (N_146,In_1404,In_403);
and U147 (N_147,In_1348,In_20);
or U148 (N_148,In_1122,In_547);
nand U149 (N_149,In_1215,In_652);
nand U150 (N_150,In_1269,In_1364);
nor U151 (N_151,In_732,In_596);
nor U152 (N_152,In_681,In_207);
xnor U153 (N_153,In_191,In_1255);
or U154 (N_154,In_428,In_595);
nand U155 (N_155,In_387,In_837);
or U156 (N_156,In_1256,In_1201);
nand U157 (N_157,In_832,In_1057);
or U158 (N_158,In_1109,In_47);
nor U159 (N_159,In_526,In_586);
or U160 (N_160,In_1119,In_218);
xor U161 (N_161,In_346,In_903);
xnor U162 (N_162,In_35,In_328);
and U163 (N_163,In_354,In_1067);
nor U164 (N_164,In_1139,In_10);
or U165 (N_165,In_296,In_820);
nor U166 (N_166,In_86,In_248);
xor U167 (N_167,In_737,In_520);
xnor U168 (N_168,In_1462,In_1033);
or U169 (N_169,In_789,In_638);
xnor U170 (N_170,In_39,In_1354);
or U171 (N_171,In_1244,In_393);
or U172 (N_172,In_758,In_1011);
xnor U173 (N_173,In_241,In_110);
or U174 (N_174,In_711,In_1349);
or U175 (N_175,In_496,In_1499);
or U176 (N_176,In_442,In_969);
xor U177 (N_177,In_1100,In_1207);
xor U178 (N_178,In_892,In_222);
nor U179 (N_179,In_1101,In_513);
nand U180 (N_180,In_277,In_788);
xnor U181 (N_181,In_83,In_435);
nor U182 (N_182,In_1105,In_1013);
nor U183 (N_183,In_436,In_341);
xor U184 (N_184,In_772,In_1003);
nor U185 (N_185,In_724,In_1233);
and U186 (N_186,In_1487,In_210);
nand U187 (N_187,In_848,In_797);
nor U188 (N_188,In_734,In_613);
nand U189 (N_189,In_742,In_744);
nand U190 (N_190,In_468,In_336);
nor U191 (N_191,In_554,In_709);
xnor U192 (N_192,In_321,In_1353);
and U193 (N_193,In_999,In_756);
or U194 (N_194,In_91,In_1250);
xnor U195 (N_195,In_618,In_1155);
and U196 (N_196,In_348,In_421);
or U197 (N_197,In_984,In_1464);
xnor U198 (N_198,In_482,In_1081);
or U199 (N_199,In_838,In_1166);
or U200 (N_200,In_438,In_799);
and U201 (N_201,In_245,In_389);
xor U202 (N_202,In_822,In_1226);
xor U203 (N_203,In_57,In_1344);
nand U204 (N_204,In_924,In_429);
or U205 (N_205,In_67,In_1102);
xor U206 (N_206,In_691,In_485);
nand U207 (N_207,In_1478,In_295);
xor U208 (N_208,In_1374,In_45);
xnor U209 (N_209,In_859,In_764);
nand U210 (N_210,In_422,In_1063);
nor U211 (N_211,In_1196,In_143);
or U212 (N_212,In_1430,In_1260);
nand U213 (N_213,In_633,In_266);
nor U214 (N_214,In_890,In_236);
and U215 (N_215,In_982,In_1328);
nor U216 (N_216,In_476,In_3);
or U217 (N_217,In_1347,In_524);
nor U218 (N_218,In_1406,In_418);
or U219 (N_219,In_451,In_1025);
nor U220 (N_220,In_358,In_825);
nand U221 (N_221,In_1322,In_184);
nor U222 (N_222,In_571,In_573);
xnor U223 (N_223,In_1006,In_1324);
nand U224 (N_224,In_488,In_1005);
xnor U225 (N_225,In_1141,In_250);
xnor U226 (N_226,In_954,In_1049);
xor U227 (N_227,In_459,In_1403);
nand U228 (N_228,In_48,In_1286);
or U229 (N_229,In_472,In_557);
xnor U230 (N_230,In_1342,In_815);
or U231 (N_231,In_352,In_495);
or U232 (N_232,In_864,In_1150);
nand U233 (N_233,In_1120,In_224);
xor U234 (N_234,In_597,In_1495);
and U235 (N_235,In_1018,In_1327);
nor U236 (N_236,In_576,In_578);
or U237 (N_237,In_1243,In_1287);
nor U238 (N_238,In_270,In_587);
nand U239 (N_239,In_259,In_163);
and U240 (N_240,In_1088,In_944);
nor U241 (N_241,In_891,In_707);
and U242 (N_242,In_1361,In_51);
or U243 (N_243,In_1041,In_621);
and U244 (N_244,In_1089,In_568);
xnor U245 (N_245,In_934,In_975);
nor U246 (N_246,In_132,In_214);
or U247 (N_247,In_819,In_287);
nor U248 (N_248,In_1031,In_5);
nor U249 (N_249,In_59,In_223);
or U250 (N_250,In_126,In_1315);
nor U251 (N_251,In_407,In_105);
nand U252 (N_252,In_804,In_402);
and U253 (N_253,In_1316,In_920);
nand U254 (N_254,In_653,In_200);
nor U255 (N_255,In_499,In_142);
xnor U256 (N_256,In_659,In_521);
nor U257 (N_257,In_661,In_735);
xor U258 (N_258,In_911,In_1200);
or U259 (N_259,In_909,In_1091);
nor U260 (N_260,In_1264,In_412);
xnor U261 (N_261,In_1369,In_1386);
xnor U262 (N_262,In_77,In_378);
and U263 (N_263,In_1072,In_1313);
xnor U264 (N_264,In_1219,In_726);
xnor U265 (N_265,In_157,In_154);
xor U266 (N_266,In_677,In_927);
nor U267 (N_267,In_703,In_283);
xnor U268 (N_268,In_458,In_759);
xnor U269 (N_269,In_951,In_993);
or U270 (N_270,In_398,In_271);
or U271 (N_271,In_1132,In_979);
and U272 (N_272,In_1148,In_1239);
nor U273 (N_273,In_616,In_814);
or U274 (N_274,In_478,In_766);
nand U275 (N_275,In_906,In_1473);
nand U276 (N_276,In_810,In_251);
nor U277 (N_277,In_327,In_1383);
and U278 (N_278,In_360,In_1214);
and U279 (N_279,In_1002,In_185);
nor U280 (N_280,In_350,In_1497);
and U281 (N_281,In_221,In_1492);
xnor U282 (N_282,In_998,In_674);
xor U283 (N_283,In_1360,In_882);
or U284 (N_284,In_146,In_1133);
or U285 (N_285,In_1123,In_44);
nand U286 (N_286,In_382,In_858);
xor U287 (N_287,In_280,In_1418);
nand U288 (N_288,In_1254,In_1217);
nor U289 (N_289,In_1192,In_1458);
and U290 (N_290,In_1427,In_1180);
or U291 (N_291,In_610,In_1465);
or U292 (N_292,In_433,In_970);
nor U293 (N_293,In_1154,In_1227);
nand U294 (N_294,In_444,In_1401);
nor U295 (N_295,In_1482,In_791);
and U296 (N_296,In_809,In_697);
nand U297 (N_297,In_798,In_36);
or U298 (N_298,In_1146,In_73);
or U299 (N_299,In_1409,In_542);
or U300 (N_300,In_896,In_1047);
and U301 (N_301,In_260,In_1218);
nor U302 (N_302,In_971,In_611);
xor U303 (N_303,In_932,In_256);
nand U304 (N_304,In_471,In_834);
nor U305 (N_305,In_30,In_675);
nand U306 (N_306,In_308,In_265);
xnor U307 (N_307,In_1157,In_778);
xor U308 (N_308,In_908,In_64);
or U309 (N_309,In_70,In_512);
or U310 (N_310,In_263,In_700);
nand U311 (N_311,In_1015,In_518);
nand U312 (N_312,In_1149,In_330);
or U313 (N_313,In_125,In_592);
and U314 (N_314,In_409,In_1336);
nor U315 (N_315,In_1452,In_1170);
nand U316 (N_316,In_863,In_643);
and U317 (N_317,In_670,In_1350);
or U318 (N_318,In_4,In_1380);
or U319 (N_319,In_679,In_540);
nor U320 (N_320,In_1134,In_869);
xnor U321 (N_321,In_955,In_37);
and U322 (N_322,In_1125,In_1075);
or U323 (N_323,In_528,In_1026);
or U324 (N_324,In_1491,In_581);
nor U325 (N_325,In_818,In_1356);
nand U326 (N_326,In_988,In_1169);
nand U327 (N_327,In_388,In_987);
and U328 (N_328,In_483,In_253);
nor U329 (N_329,In_128,In_1187);
xnor U330 (N_330,In_449,In_503);
nor U331 (N_331,In_781,In_830);
or U332 (N_332,In_977,In_82);
or U333 (N_333,In_1303,In_666);
nor U334 (N_334,In_430,In_1036);
xor U335 (N_335,In_63,In_274);
nand U336 (N_336,In_371,In_1054);
or U337 (N_337,In_943,In_356);
and U338 (N_338,In_28,In_1388);
xor U339 (N_339,In_588,In_316);
or U340 (N_340,In_608,In_849);
nor U341 (N_341,In_535,In_783);
or U342 (N_342,In_961,In_1073);
xnor U343 (N_343,In_213,In_657);
and U344 (N_344,In_351,In_1490);
nor U345 (N_345,In_1308,In_516);
and U346 (N_346,In_1103,In_522);
or U347 (N_347,In_244,In_401);
nor U348 (N_348,In_567,In_205);
or U349 (N_349,In_1198,In_230);
nor U350 (N_350,In_1142,In_1);
and U351 (N_351,In_31,In_1199);
or U352 (N_352,In_671,In_391);
nor U353 (N_353,In_189,In_1221);
nor U354 (N_354,In_1284,In_115);
nand U355 (N_355,In_416,In_684);
nand U356 (N_356,In_1251,In_678);
nor U357 (N_357,In_1159,In_989);
and U358 (N_358,In_866,In_107);
and U359 (N_359,In_252,In_614);
nand U360 (N_360,In_997,In_770);
or U361 (N_361,In_746,In_510);
and U362 (N_362,In_1410,In_1065);
nand U363 (N_363,In_617,In_1338);
xor U364 (N_364,In_569,In_343);
and U365 (N_365,In_1488,In_1129);
xnor U366 (N_366,In_768,In_1456);
and U367 (N_367,In_1310,In_262);
and U368 (N_368,In_1332,In_1325);
xor U369 (N_369,In_1399,In_307);
xor U370 (N_370,In_1424,In_1266);
nor U371 (N_371,In_698,In_72);
and U372 (N_372,In_129,In_357);
nor U373 (N_373,In_956,In_1280);
or U374 (N_374,In_1337,In_623);
and U375 (N_375,In_1474,In_622);
nor U376 (N_376,In_400,In_137);
nand U377 (N_377,In_779,In_166);
nor U378 (N_378,In_1442,In_440);
nand U379 (N_379,In_181,In_1395);
or U380 (N_380,In_104,In_748);
or U381 (N_381,In_1290,In_55);
nand U382 (N_382,In_1178,In_1016);
xor U383 (N_383,In_74,In_990);
nand U384 (N_384,In_727,In_913);
and U385 (N_385,In_1471,In_195);
or U386 (N_386,In_455,In_1411);
or U387 (N_387,In_963,In_803);
nor U388 (N_388,In_536,In_1402);
nor U389 (N_389,In_193,In_876);
or U390 (N_390,In_566,In_1008);
nand U391 (N_391,In_197,In_760);
nor U392 (N_392,In_1193,In_1445);
or U393 (N_393,In_626,In_2);
nand U394 (N_394,In_1234,In_1268);
xor U395 (N_395,In_845,In_267);
xor U396 (N_396,In_645,In_582);
or U397 (N_397,In_1439,In_1321);
or U398 (N_398,In_1295,In_828);
or U399 (N_399,In_647,In_172);
nor U400 (N_400,In_1400,In_1479);
xnor U401 (N_401,In_169,In_1118);
nor U402 (N_402,In_1448,In_1053);
nor U403 (N_403,In_1068,In_541);
nand U404 (N_404,In_1229,In_723);
and U405 (N_405,In_366,In_339);
or U406 (N_406,In_751,In_1164);
xor U407 (N_407,In_490,In_1340);
and U408 (N_408,In_899,In_694);
xor U409 (N_409,In_314,In_108);
nor U410 (N_410,In_594,In_121);
nor U411 (N_411,In_1294,In_123);
or U412 (N_412,In_634,In_43);
xnor U413 (N_413,In_312,In_949);
xnor U414 (N_414,In_9,In_941);
or U415 (N_415,In_552,In_1319);
nand U416 (N_416,In_1498,In_738);
and U417 (N_417,In_1379,In_1421);
and U418 (N_418,In_1237,In_1034);
or U419 (N_419,In_1433,In_150);
and U420 (N_420,In_857,In_1352);
nor U421 (N_421,In_370,In_414);
nand U422 (N_422,In_1191,In_1432);
and U423 (N_423,In_216,In_273);
xor U424 (N_424,In_878,In_12);
nor U425 (N_425,In_1076,In_1372);
nand U426 (N_426,In_1126,In_1419);
nand U427 (N_427,In_235,In_215);
nor U428 (N_428,In_1151,In_152);
and U429 (N_429,In_668,In_921);
nor U430 (N_430,In_58,In_1165);
xnor U431 (N_431,In_127,In_1476);
xnor U432 (N_432,In_228,In_1066);
xor U433 (N_433,In_1019,In_410);
nor U434 (N_434,In_562,In_1343);
or U435 (N_435,In_437,In_497);
or U436 (N_436,In_279,In_1171);
and U437 (N_437,In_1341,In_757);
nor U438 (N_438,In_494,In_15);
or U439 (N_439,In_417,In_717);
nor U440 (N_440,In_912,In_1262);
or U441 (N_441,In_17,In_874);
nand U442 (N_442,In_824,In_232);
xor U443 (N_443,In_22,In_1289);
nand U444 (N_444,In_93,In_646);
nor U445 (N_445,In_855,In_504);
nand U446 (N_446,In_68,In_332);
or U447 (N_447,In_762,In_1043);
or U448 (N_448,In_1382,In_619);
xor U449 (N_449,In_1450,In_862);
nor U450 (N_450,In_1274,In_1376);
or U451 (N_451,In_376,In_1459);
xor U452 (N_452,In_885,In_175);
xnor U453 (N_453,In_794,In_434);
and U454 (N_454,In_1037,In_1391);
xor U455 (N_455,In_1496,In_329);
xnor U456 (N_456,In_683,In_514);
or U457 (N_457,In_721,In_149);
and U458 (N_458,In_240,In_1117);
nor U459 (N_459,In_821,In_1318);
or U460 (N_460,In_517,In_373);
or U461 (N_461,In_967,In_171);
xnor U462 (N_462,In_113,In_1493);
nor U463 (N_463,In_532,In_538);
xor U464 (N_464,In_158,In_1213);
xor U465 (N_465,In_1001,In_593);
nand U466 (N_466,In_688,In_204);
nand U467 (N_467,In_714,In_1030);
xor U468 (N_468,In_960,In_176);
and U469 (N_469,In_1282,In_850);
nand U470 (N_470,In_1486,In_636);
or U471 (N_471,In_1485,In_144);
and U472 (N_472,In_1004,In_713);
nand U473 (N_473,In_272,In_994);
and U474 (N_474,In_1438,In_269);
xor U475 (N_475,In_359,In_114);
or U476 (N_476,In_715,In_750);
and U477 (N_477,In_1259,In_290);
and U478 (N_478,In_1258,In_682);
nor U479 (N_479,In_861,In_397);
or U480 (N_480,In_420,In_247);
or U481 (N_481,In_1058,In_693);
xnor U482 (N_482,In_1114,In_170);
nor U483 (N_483,In_947,In_1224);
xnor U484 (N_484,In_774,In_511);
nor U485 (N_485,In_173,In_936);
xor U486 (N_486,In_315,In_138);
and U487 (N_487,In_133,In_326);
xor U488 (N_488,In_1357,In_21);
nand U489 (N_489,In_575,In_543);
or U490 (N_490,In_560,In_1228);
or U491 (N_491,In_454,In_225);
nand U492 (N_492,In_928,In_1345);
nor U493 (N_493,In_790,In_525);
nand U494 (N_494,In_612,In_1320);
or U495 (N_495,In_992,In_399);
xor U496 (N_496,In_826,In_206);
xor U497 (N_497,In_1009,In_1351);
and U498 (N_498,In_226,In_549);
nor U499 (N_499,In_211,In_1017);
nand U500 (N_500,In_1056,In_786);
xor U501 (N_501,In_1186,In_802);
and U502 (N_502,In_148,In_1484);
and U503 (N_503,In_733,In_856);
xor U504 (N_504,In_116,In_1252);
and U505 (N_505,In_1415,In_7);
or U506 (N_506,In_487,In_902);
nor U507 (N_507,In_1230,In_1027);
xnor U508 (N_508,In_667,In_1444);
and U509 (N_509,In_769,In_763);
or U510 (N_510,In_1085,In_1082);
nand U511 (N_511,In_1467,In_996);
nor U512 (N_512,In_651,In_1453);
nor U513 (N_513,In_1099,In_564);
nor U514 (N_514,In_718,In_570);
nor U515 (N_515,In_1472,In_381);
nand U516 (N_516,In_441,In_135);
xnor U517 (N_517,In_484,In_243);
and U518 (N_518,In_833,In_1108);
nor U519 (N_519,In_353,In_394);
and U520 (N_520,In_29,In_1197);
or U521 (N_521,In_162,In_1080);
or U522 (N_522,In_1311,In_310);
or U523 (N_523,In_656,In_930);
or U524 (N_524,In_220,In_80);
nor U525 (N_525,In_1249,In_323);
nor U526 (N_526,In_817,In_624);
nand U527 (N_527,In_1212,In_493);
and U528 (N_528,In_374,In_95);
nor U529 (N_529,In_75,In_736);
xnor U530 (N_530,In_1083,In_787);
or U531 (N_531,In_219,In_1115);
nor U532 (N_532,In_1431,In_1359);
and U533 (N_533,In_776,In_334);
and U534 (N_534,In_501,In_938);
or U535 (N_535,In_117,In_54);
nand U536 (N_536,In_1181,In_752);
nand U537 (N_537,In_156,In_14);
and U538 (N_538,In_89,In_1211);
nand U539 (N_539,In_806,In_264);
or U540 (N_540,In_897,In_165);
nor U541 (N_541,In_958,In_1463);
xnor U542 (N_542,In_60,In_309);
and U543 (N_543,In_527,In_475);
nor U544 (N_544,In_84,In_448);
or U545 (N_545,In_695,In_785);
or U546 (N_546,In_1194,In_1074);
xnor U547 (N_547,In_1455,In_96);
or U548 (N_548,In_654,In_1367);
and U549 (N_549,In_973,In_190);
nand U550 (N_550,In_1147,In_1333);
nor U551 (N_551,In_519,In_268);
nand U552 (N_552,In_284,In_406);
xor U553 (N_553,In_1064,In_1062);
nand U554 (N_554,In_1408,In_1481);
xor U555 (N_555,In_46,In_929);
nor U556 (N_556,In_1470,In_1028);
nand U557 (N_557,In_705,In_904);
or U558 (N_558,In_1022,In_1460);
and U559 (N_559,In_187,In_1371);
nand U560 (N_560,In_239,In_1241);
xor U561 (N_561,In_379,In_775);
and U562 (N_562,In_447,In_663);
xor U563 (N_563,In_474,In_1208);
nor U564 (N_564,In_201,In_639);
and U565 (N_565,In_523,In_1378);
nor U566 (N_566,In_640,In_369);
and U567 (N_567,In_1309,In_609);
and U568 (N_568,In_1173,In_1265);
or U569 (N_569,In_561,In_491);
xor U570 (N_570,In_141,In_349);
xor U571 (N_571,In_1288,In_151);
and U572 (N_572,In_986,In_914);
nand U573 (N_573,In_303,In_1112);
or U574 (N_574,In_61,In_1413);
xor U575 (N_575,In_292,In_680);
or U576 (N_576,In_395,In_242);
and U577 (N_577,In_545,In_479);
and U578 (N_578,In_648,In_1285);
nor U579 (N_579,In_1238,In_1189);
xnor U580 (N_580,In_1272,In_907);
or U581 (N_581,In_317,In_32);
xnor U582 (N_582,In_362,In_461);
and U583 (N_583,In_1397,In_1301);
nor U584 (N_584,In_1300,In_607);
nor U585 (N_585,In_506,In_1039);
and U586 (N_586,In_196,In_1446);
nand U587 (N_587,In_1225,In_722);
nand U588 (N_588,In_589,In_841);
and U589 (N_589,In_946,In_1128);
nand U590 (N_590,In_740,In_884);
and U591 (N_591,In_33,In_486);
and U592 (N_592,In_627,In_1436);
nor U593 (N_593,In_620,In_1111);
or U594 (N_594,In_1079,In_606);
or U595 (N_595,In_177,In_1094);
or U596 (N_596,In_972,In_469);
or U597 (N_597,In_1104,In_453);
xor U598 (N_598,In_761,In_780);
nand U599 (N_599,In_660,In_1302);
nand U600 (N_600,In_1307,In_180);
and U601 (N_601,In_246,In_1454);
or U602 (N_602,In_1185,In_875);
and U603 (N_603,In_1202,In_318);
or U604 (N_604,In_1414,In_1299);
xor U605 (N_605,In_883,In_603);
nand U606 (N_606,In_628,In_1231);
nor U607 (N_607,In_893,In_1385);
or U608 (N_608,In_427,In_940);
nand U609 (N_609,In_962,In_1042);
nand U610 (N_610,In_1384,In_34);
nand U611 (N_611,In_481,In_192);
nand U612 (N_612,In_160,In_183);
nand U613 (N_613,In_771,In_1393);
nand U614 (N_614,In_1179,In_765);
xor U615 (N_615,In_782,In_122);
xor U616 (N_616,In_340,In_238);
and U617 (N_617,In_56,In_1175);
and U618 (N_618,In_79,In_257);
nor U619 (N_619,In_1368,In_300);
nand U620 (N_620,In_1168,In_286);
and U621 (N_621,In_140,In_134);
or U622 (N_622,In_392,In_464);
xnor U623 (N_623,In_413,In_655);
nor U624 (N_624,In_11,In_625);
and U625 (N_625,In_8,In_555);
nand U626 (N_626,In_917,In_580);
and U627 (N_627,In_720,In_839);
nor U628 (N_628,In_629,In_985);
or U629 (N_629,In_926,In_976);
nand U630 (N_630,In_777,In_106);
xor U631 (N_631,In_991,In_208);
nor U632 (N_632,In_701,In_1283);
or U633 (N_633,In_840,In_347);
nand U634 (N_634,In_692,In_1087);
xor U635 (N_635,In_1330,In_637);
nor U636 (N_636,In_1188,In_1007);
or U637 (N_637,In_509,In_1365);
nand U638 (N_638,In_404,In_1423);
nand U639 (N_639,In_439,In_390);
nor U640 (N_640,In_945,In_534);
nor U641 (N_641,In_807,In_364);
nor U642 (N_642,In_1422,In_1131);
xor U643 (N_643,In_1086,In_935);
and U644 (N_644,In_600,In_443);
and U645 (N_645,In_1061,In_1172);
and U646 (N_646,In_261,In_1052);
nand U647 (N_647,In_980,In_598);
and U648 (N_648,In_1276,In_1000);
nor U649 (N_649,In_98,In_1441);
nand U650 (N_650,In_293,In_812);
nand U651 (N_651,In_1396,In_342);
nand U652 (N_652,In_118,In_870);
xnor U653 (N_653,In_385,In_465);
xnor U654 (N_654,In_1326,In_337);
nor U655 (N_655,In_1084,In_178);
or U656 (N_656,In_288,In_1059);
nand U657 (N_657,In_873,In_304);
and U658 (N_658,In_1277,In_754);
xnor U659 (N_659,In_704,In_1203);
xnor U660 (N_660,In_1140,In_186);
nand U661 (N_661,In_502,In_959);
nor U662 (N_662,In_320,In_1305);
and U663 (N_663,In_898,In_1055);
or U664 (N_664,In_456,In_1468);
xnor U665 (N_665,In_1253,In_939);
xor U666 (N_666,In_915,In_1293);
nor U667 (N_667,In_298,In_1314);
nor U668 (N_668,In_24,In_227);
xor U669 (N_669,In_1040,In_254);
or U670 (N_670,In_1278,In_1443);
and U671 (N_671,In_601,In_1329);
nor U672 (N_672,In_1247,In_278);
and U673 (N_673,In_1358,In_76);
nor U674 (N_674,In_408,In_65);
xor U675 (N_675,In_299,In_1312);
nand U676 (N_676,In_1107,In_689);
nor U677 (N_677,In_1270,In_1110);
nor U678 (N_678,In_331,In_52);
or U679 (N_679,In_1098,In_690);
and U680 (N_680,In_130,In_1032);
and U681 (N_681,In_887,In_852);
nor U682 (N_682,In_1035,In_365);
and U683 (N_683,In_1306,In_188);
nand U684 (N_684,In_1434,In_1273);
nor U685 (N_685,In_551,In_199);
and U686 (N_686,In_100,In_1425);
or U687 (N_687,In_953,In_301);
or U688 (N_688,In_599,In_97);
or U689 (N_689,In_877,In_872);
or U690 (N_690,In_865,In_1220);
and U691 (N_691,In_631,In_846);
and U692 (N_692,In_489,In_124);
nor U693 (N_693,In_431,In_725);
or U694 (N_694,In_1292,In_1475);
nor U695 (N_695,In_361,In_1152);
or U696 (N_696,In_1466,In_302);
nor U697 (N_697,In_153,In_559);
xnor U698 (N_698,In_641,In_879);
or U699 (N_699,In_99,In_1429);
xor U700 (N_700,In_53,In_167);
nor U701 (N_701,In_672,In_1261);
xor U702 (N_702,In_372,In_669);
nor U703 (N_703,In_577,In_933);
nor U704 (N_704,In_1257,In_49);
and U705 (N_705,In_981,In_1050);
and U706 (N_706,In_792,In_1494);
or U707 (N_707,In_16,In_234);
xor U708 (N_708,In_1182,In_423);
or U709 (N_709,In_275,In_480);
nor U710 (N_710,In_894,In_844);
xnor U711 (N_711,In_1339,In_470);
and U712 (N_712,In_313,In_889);
and U713 (N_713,In_1449,In_136);
and U714 (N_714,In_81,In_289);
nor U715 (N_715,In_145,In_650);
xor U716 (N_716,In_644,In_529);
nand U717 (N_717,In_544,In_297);
nor U718 (N_718,In_860,In_1195);
nand U719 (N_719,In_38,In_333);
nand U720 (N_720,In_319,In_255);
nor U721 (N_721,In_231,In_1246);
nor U722 (N_722,In_937,In_827);
nand U723 (N_723,In_676,In_338);
and U724 (N_724,In_155,In_1398);
nor U725 (N_725,In_335,In_919);
nor U726 (N_726,In_1137,In_835);
xor U727 (N_727,In_1177,In_931);
nor U728 (N_728,In_1346,In_1375);
xor U729 (N_729,In_922,In_1480);
nor U730 (N_730,In_1420,In_120);
nor U731 (N_731,In_1051,In_974);
nor U732 (N_732,In_367,In_1092);
xnor U733 (N_733,In_1417,In_1373);
or U734 (N_734,In_1216,In_71);
or U735 (N_735,In_1405,In_515);
or U736 (N_736,In_1435,In_209);
nand U737 (N_737,In_467,In_498);
nor U738 (N_738,In_1145,In_747);
or U739 (N_739,In_1245,In_1304);
nand U740 (N_740,In_103,In_1489);
or U741 (N_741,In_743,In_1144);
nor U742 (N_742,In_1010,In_66);
nand U743 (N_743,In_1222,In_952);
nor U744 (N_744,In_1355,In_1078);
or U745 (N_745,In_174,In_324);
xor U746 (N_746,In_368,In_111);
nor U747 (N_747,In_1275,In_1271);
and U748 (N_748,In_473,In_119);
nand U749 (N_749,In_202,In_325);
and U750 (N_750,In_657,In_1257);
or U751 (N_751,In_1150,In_1476);
xor U752 (N_752,In_602,In_606);
or U753 (N_753,In_139,In_1390);
or U754 (N_754,In_799,In_1236);
and U755 (N_755,In_872,In_782);
and U756 (N_756,In_55,In_1138);
or U757 (N_757,In_617,In_1212);
xnor U758 (N_758,In_1333,In_574);
nand U759 (N_759,In_706,In_369);
nor U760 (N_760,In_403,In_1477);
and U761 (N_761,In_838,In_813);
nor U762 (N_762,In_1148,In_1488);
xnor U763 (N_763,In_477,In_792);
nor U764 (N_764,In_339,In_963);
nand U765 (N_765,In_93,In_664);
or U766 (N_766,In_1068,In_285);
xnor U767 (N_767,In_221,In_1077);
nand U768 (N_768,In_1095,In_210);
xnor U769 (N_769,In_1197,In_658);
and U770 (N_770,In_1367,In_296);
nor U771 (N_771,In_1357,In_33);
or U772 (N_772,In_1031,In_322);
nand U773 (N_773,In_1246,In_1025);
and U774 (N_774,In_738,In_1365);
and U775 (N_775,In_867,In_210);
nand U776 (N_776,In_1010,In_1253);
nand U777 (N_777,In_1228,In_103);
nor U778 (N_778,In_1329,In_3);
nand U779 (N_779,In_587,In_570);
nor U780 (N_780,In_409,In_787);
xnor U781 (N_781,In_794,In_823);
nor U782 (N_782,In_592,In_92);
xor U783 (N_783,In_179,In_689);
nor U784 (N_784,In_100,In_203);
nor U785 (N_785,In_554,In_846);
and U786 (N_786,In_1047,In_470);
xor U787 (N_787,In_112,In_1129);
and U788 (N_788,In_1276,In_1030);
nor U789 (N_789,In_1334,In_565);
nand U790 (N_790,In_1484,In_1137);
xnor U791 (N_791,In_836,In_1348);
nand U792 (N_792,In_1014,In_235);
or U793 (N_793,In_45,In_807);
or U794 (N_794,In_1325,In_1201);
and U795 (N_795,In_943,In_932);
nand U796 (N_796,In_1481,In_149);
nor U797 (N_797,In_195,In_362);
xor U798 (N_798,In_1303,In_1038);
xnor U799 (N_799,In_541,In_44);
nand U800 (N_800,In_596,In_166);
or U801 (N_801,In_1428,In_1098);
or U802 (N_802,In_717,In_286);
nor U803 (N_803,In_649,In_349);
and U804 (N_804,In_1005,In_540);
and U805 (N_805,In_1129,In_106);
nor U806 (N_806,In_940,In_571);
and U807 (N_807,In_720,In_215);
nor U808 (N_808,In_782,In_1143);
xnor U809 (N_809,In_1288,In_116);
and U810 (N_810,In_1060,In_954);
and U811 (N_811,In_517,In_946);
nor U812 (N_812,In_749,In_1214);
and U813 (N_813,In_1276,In_199);
xor U814 (N_814,In_636,In_222);
or U815 (N_815,In_1294,In_733);
xnor U816 (N_816,In_418,In_47);
or U817 (N_817,In_354,In_71);
or U818 (N_818,In_881,In_518);
xor U819 (N_819,In_1108,In_330);
nand U820 (N_820,In_104,In_730);
nand U821 (N_821,In_779,In_119);
xor U822 (N_822,In_1,In_524);
or U823 (N_823,In_795,In_294);
or U824 (N_824,In_1471,In_251);
nor U825 (N_825,In_732,In_779);
or U826 (N_826,In_784,In_48);
or U827 (N_827,In_1460,In_1083);
xnor U828 (N_828,In_479,In_659);
and U829 (N_829,In_1225,In_1459);
xnor U830 (N_830,In_902,In_618);
nand U831 (N_831,In_1003,In_516);
and U832 (N_832,In_558,In_143);
and U833 (N_833,In_1448,In_833);
nor U834 (N_834,In_811,In_323);
xnor U835 (N_835,In_1017,In_699);
or U836 (N_836,In_1000,In_651);
or U837 (N_837,In_1385,In_1043);
nor U838 (N_838,In_1395,In_1383);
nand U839 (N_839,In_1030,In_936);
nand U840 (N_840,In_928,In_734);
nand U841 (N_841,In_1413,In_383);
nand U842 (N_842,In_801,In_1005);
and U843 (N_843,In_841,In_697);
nor U844 (N_844,In_89,In_967);
or U845 (N_845,In_1214,In_55);
and U846 (N_846,In_115,In_1340);
nand U847 (N_847,In_1237,In_214);
or U848 (N_848,In_455,In_93);
or U849 (N_849,In_613,In_380);
or U850 (N_850,In_811,In_1221);
and U851 (N_851,In_718,In_841);
xnor U852 (N_852,In_647,In_408);
or U853 (N_853,In_453,In_1404);
nand U854 (N_854,In_304,In_324);
and U855 (N_855,In_609,In_1135);
or U856 (N_856,In_87,In_1484);
nor U857 (N_857,In_1132,In_1159);
xnor U858 (N_858,In_1272,In_1288);
xor U859 (N_859,In_1229,In_381);
xnor U860 (N_860,In_868,In_78);
or U861 (N_861,In_1079,In_465);
xnor U862 (N_862,In_125,In_1406);
nor U863 (N_863,In_471,In_733);
and U864 (N_864,In_1476,In_133);
nor U865 (N_865,In_426,In_261);
and U866 (N_866,In_516,In_1186);
nand U867 (N_867,In_202,In_273);
xor U868 (N_868,In_613,In_806);
nand U869 (N_869,In_1403,In_1366);
and U870 (N_870,In_917,In_474);
and U871 (N_871,In_326,In_50);
or U872 (N_872,In_394,In_768);
xnor U873 (N_873,In_48,In_99);
nand U874 (N_874,In_870,In_1317);
nor U875 (N_875,In_227,In_806);
and U876 (N_876,In_1494,In_1384);
nand U877 (N_877,In_718,In_174);
and U878 (N_878,In_836,In_144);
or U879 (N_879,In_742,In_649);
or U880 (N_880,In_16,In_877);
nor U881 (N_881,In_1342,In_560);
nand U882 (N_882,In_700,In_1447);
and U883 (N_883,In_202,In_1219);
nand U884 (N_884,In_676,In_140);
and U885 (N_885,In_754,In_939);
nand U886 (N_886,In_226,In_862);
nor U887 (N_887,In_742,In_528);
or U888 (N_888,In_611,In_376);
nand U889 (N_889,In_252,In_14);
or U890 (N_890,In_80,In_393);
and U891 (N_891,In_820,In_1387);
xnor U892 (N_892,In_1130,In_1103);
or U893 (N_893,In_409,In_373);
xnor U894 (N_894,In_282,In_292);
nor U895 (N_895,In_1155,In_522);
xnor U896 (N_896,In_1494,In_681);
and U897 (N_897,In_1460,In_20);
or U898 (N_898,In_669,In_61);
or U899 (N_899,In_1327,In_1091);
or U900 (N_900,In_170,In_989);
xor U901 (N_901,In_850,In_1350);
or U902 (N_902,In_839,In_809);
or U903 (N_903,In_1052,In_497);
xor U904 (N_904,In_897,In_1088);
and U905 (N_905,In_1036,In_925);
or U906 (N_906,In_282,In_1180);
xor U907 (N_907,In_684,In_1280);
nand U908 (N_908,In_674,In_141);
xnor U909 (N_909,In_1283,In_725);
nor U910 (N_910,In_338,In_1243);
nor U911 (N_911,In_1164,In_8);
nor U912 (N_912,In_1143,In_1452);
xnor U913 (N_913,In_509,In_461);
nand U914 (N_914,In_642,In_767);
nor U915 (N_915,In_1106,In_1128);
and U916 (N_916,In_1414,In_129);
xor U917 (N_917,In_960,In_1419);
and U918 (N_918,In_1106,In_1138);
and U919 (N_919,In_153,In_660);
nand U920 (N_920,In_258,In_1109);
nand U921 (N_921,In_47,In_1193);
nand U922 (N_922,In_1395,In_866);
and U923 (N_923,In_81,In_4);
nand U924 (N_924,In_128,In_842);
and U925 (N_925,In_1417,In_322);
or U926 (N_926,In_902,In_1104);
or U927 (N_927,In_1468,In_881);
nand U928 (N_928,In_1222,In_1089);
nand U929 (N_929,In_595,In_240);
and U930 (N_930,In_745,In_226);
nand U931 (N_931,In_824,In_1291);
nand U932 (N_932,In_1134,In_259);
and U933 (N_933,In_892,In_1256);
xor U934 (N_934,In_24,In_1326);
or U935 (N_935,In_849,In_288);
xnor U936 (N_936,In_91,In_1044);
or U937 (N_937,In_933,In_379);
or U938 (N_938,In_1457,In_988);
or U939 (N_939,In_744,In_477);
nand U940 (N_940,In_664,In_477);
nor U941 (N_941,In_1495,In_865);
nor U942 (N_942,In_966,In_708);
nor U943 (N_943,In_631,In_349);
nand U944 (N_944,In_761,In_810);
and U945 (N_945,In_601,In_822);
and U946 (N_946,In_1431,In_1496);
xor U947 (N_947,In_345,In_761);
or U948 (N_948,In_1363,In_1487);
nor U949 (N_949,In_1106,In_1453);
or U950 (N_950,In_287,In_582);
xor U951 (N_951,In_1424,In_1134);
and U952 (N_952,In_1215,In_666);
and U953 (N_953,In_542,In_436);
nand U954 (N_954,In_209,In_1445);
or U955 (N_955,In_229,In_708);
xor U956 (N_956,In_1380,In_960);
nand U957 (N_957,In_1166,In_965);
and U958 (N_958,In_59,In_330);
nand U959 (N_959,In_621,In_595);
or U960 (N_960,In_1324,In_1297);
or U961 (N_961,In_256,In_29);
nor U962 (N_962,In_468,In_366);
xor U963 (N_963,In_414,In_1164);
xor U964 (N_964,In_932,In_164);
nor U965 (N_965,In_958,In_1219);
nor U966 (N_966,In_1495,In_135);
nand U967 (N_967,In_1412,In_150);
and U968 (N_968,In_546,In_661);
nand U969 (N_969,In_624,In_190);
or U970 (N_970,In_888,In_1188);
or U971 (N_971,In_994,In_1176);
and U972 (N_972,In_1224,In_635);
nand U973 (N_973,In_657,In_1069);
nor U974 (N_974,In_1434,In_1397);
and U975 (N_975,In_314,In_1018);
nor U976 (N_976,In_350,In_384);
nand U977 (N_977,In_646,In_366);
xor U978 (N_978,In_536,In_483);
nor U979 (N_979,In_1383,In_955);
nor U980 (N_980,In_339,In_1327);
xor U981 (N_981,In_399,In_1069);
nand U982 (N_982,In_738,In_348);
xor U983 (N_983,In_262,In_399);
and U984 (N_984,In_1356,In_865);
nand U985 (N_985,In_1302,In_1079);
and U986 (N_986,In_1161,In_739);
and U987 (N_987,In_220,In_177);
nor U988 (N_988,In_47,In_1366);
nand U989 (N_989,In_312,In_462);
or U990 (N_990,In_1453,In_131);
nand U991 (N_991,In_251,In_111);
nand U992 (N_992,In_1006,In_919);
nor U993 (N_993,In_272,In_938);
or U994 (N_994,In_404,In_413);
xnor U995 (N_995,In_1061,In_1080);
nor U996 (N_996,In_894,In_1171);
or U997 (N_997,In_1034,In_1197);
and U998 (N_998,In_162,In_4);
nand U999 (N_999,In_1223,In_442);
nand U1000 (N_1000,N_732,N_32);
xor U1001 (N_1001,N_598,N_859);
nand U1002 (N_1002,N_967,N_460);
xnor U1003 (N_1003,N_861,N_128);
nand U1004 (N_1004,N_139,N_361);
nand U1005 (N_1005,N_433,N_363);
nand U1006 (N_1006,N_971,N_898);
nand U1007 (N_1007,N_317,N_891);
xnor U1008 (N_1008,N_911,N_922);
nand U1009 (N_1009,N_521,N_275);
xor U1010 (N_1010,N_590,N_833);
xor U1011 (N_1011,N_577,N_594);
nand U1012 (N_1012,N_314,N_60);
nor U1013 (N_1013,N_441,N_745);
xor U1014 (N_1014,N_235,N_386);
xnor U1015 (N_1015,N_160,N_855);
nor U1016 (N_1016,N_676,N_737);
and U1017 (N_1017,N_155,N_259);
and U1018 (N_1018,N_831,N_684);
nand U1019 (N_1019,N_338,N_987);
and U1020 (N_1020,N_917,N_455);
nand U1021 (N_1021,N_391,N_184);
or U1022 (N_1022,N_566,N_395);
xnor U1023 (N_1023,N_587,N_932);
xor U1024 (N_1024,N_746,N_269);
xor U1025 (N_1025,N_740,N_758);
nor U1026 (N_1026,N_456,N_557);
nand U1027 (N_1027,N_254,N_309);
nor U1028 (N_1028,N_933,N_935);
xnor U1029 (N_1029,N_171,N_620);
xnor U1030 (N_1030,N_137,N_9);
nand U1031 (N_1031,N_220,N_219);
xor U1032 (N_1032,N_948,N_981);
nand U1033 (N_1033,N_57,N_790);
xor U1034 (N_1034,N_936,N_663);
nor U1035 (N_1035,N_975,N_674);
or U1036 (N_1036,N_697,N_972);
nor U1037 (N_1037,N_628,N_672);
xor U1038 (N_1038,N_79,N_182);
or U1039 (N_1039,N_467,N_290);
and U1040 (N_1040,N_609,N_59);
xnor U1041 (N_1041,N_812,N_471);
or U1042 (N_1042,N_292,N_461);
nand U1043 (N_1043,N_50,N_531);
nor U1044 (N_1044,N_547,N_424);
nor U1045 (N_1045,N_903,N_507);
and U1046 (N_1046,N_869,N_615);
nor U1047 (N_1047,N_366,N_631);
xor U1048 (N_1048,N_454,N_834);
nand U1049 (N_1049,N_358,N_976);
xnor U1050 (N_1050,N_170,N_371);
nand U1051 (N_1051,N_111,N_546);
or U1052 (N_1052,N_736,N_66);
or U1053 (N_1053,N_326,N_670);
nor U1054 (N_1054,N_955,N_823);
nor U1055 (N_1055,N_343,N_478);
nand U1056 (N_1056,N_180,N_192);
nand U1057 (N_1057,N_311,N_19);
xor U1058 (N_1058,N_883,N_263);
nor U1059 (N_1059,N_880,N_801);
xnor U1060 (N_1060,N_305,N_618);
nand U1061 (N_1061,N_996,N_67);
or U1062 (N_1062,N_923,N_156);
xor U1063 (N_1063,N_431,N_350);
xor U1064 (N_1064,N_808,N_444);
nand U1065 (N_1065,N_998,N_256);
nor U1066 (N_1066,N_793,N_864);
nor U1067 (N_1067,N_796,N_76);
nand U1068 (N_1068,N_163,N_608);
nand U1069 (N_1069,N_420,N_261);
and U1070 (N_1070,N_775,N_599);
or U1071 (N_1071,N_501,N_397);
and U1072 (N_1072,N_3,N_567);
or U1073 (N_1073,N_581,N_469);
nand U1074 (N_1074,N_141,N_990);
or U1075 (N_1075,N_525,N_143);
or U1076 (N_1076,N_770,N_465);
or U1077 (N_1077,N_665,N_713);
nor U1078 (N_1078,N_988,N_767);
nor U1079 (N_1079,N_227,N_157);
or U1080 (N_1080,N_502,N_330);
nand U1081 (N_1081,N_225,N_781);
nor U1082 (N_1082,N_828,N_321);
nor U1083 (N_1083,N_778,N_701);
nand U1084 (N_1084,N_822,N_319);
and U1085 (N_1085,N_307,N_33);
xor U1086 (N_1086,N_607,N_191);
and U1087 (N_1087,N_44,N_728);
and U1088 (N_1088,N_532,N_856);
nor U1089 (N_1089,N_222,N_117);
xnor U1090 (N_1090,N_421,N_519);
nand U1091 (N_1091,N_483,N_46);
nor U1092 (N_1092,N_459,N_62);
and U1093 (N_1093,N_84,N_535);
or U1094 (N_1094,N_132,N_591);
and U1095 (N_1095,N_819,N_355);
xor U1096 (N_1096,N_751,N_905);
nand U1097 (N_1097,N_708,N_447);
xor U1098 (N_1098,N_230,N_208);
xnor U1099 (N_1099,N_849,N_681);
and U1100 (N_1100,N_429,N_520);
and U1101 (N_1101,N_492,N_228);
nand U1102 (N_1102,N_413,N_387);
nand U1103 (N_1103,N_584,N_78);
or U1104 (N_1104,N_264,N_87);
and U1105 (N_1105,N_121,N_408);
nand U1106 (N_1106,N_422,N_814);
or U1107 (N_1107,N_244,N_866);
nand U1108 (N_1108,N_85,N_86);
or U1109 (N_1109,N_841,N_640);
or U1110 (N_1110,N_985,N_638);
and U1111 (N_1111,N_937,N_716);
and U1112 (N_1112,N_622,N_16);
and U1113 (N_1113,N_647,N_500);
xor U1114 (N_1114,N_807,N_956);
nand U1115 (N_1115,N_271,N_2);
xnor U1116 (N_1116,N_963,N_876);
or U1117 (N_1117,N_662,N_18);
or U1118 (N_1118,N_53,N_417);
xor U1119 (N_1119,N_154,N_52);
and U1120 (N_1120,N_895,N_616);
or U1121 (N_1121,N_407,N_293);
nor U1122 (N_1122,N_887,N_797);
and U1123 (N_1123,N_938,N_989);
xor U1124 (N_1124,N_415,N_405);
or U1125 (N_1125,N_342,N_692);
or U1126 (N_1126,N_120,N_994);
or U1127 (N_1127,N_301,N_573);
nand U1128 (N_1128,N_639,N_36);
xnor U1129 (N_1129,N_34,N_482);
xor U1130 (N_1130,N_38,N_910);
or U1131 (N_1131,N_485,N_931);
nor U1132 (N_1132,N_352,N_136);
nor U1133 (N_1133,N_439,N_768);
xnor U1134 (N_1134,N_418,N_392);
nor U1135 (N_1135,N_809,N_916);
nand U1136 (N_1136,N_498,N_473);
nand U1137 (N_1137,N_960,N_749);
nand U1138 (N_1138,N_537,N_660);
or U1139 (N_1139,N_29,N_509);
xnor U1140 (N_1140,N_602,N_406);
or U1141 (N_1141,N_97,N_239);
and U1142 (N_1142,N_357,N_627);
xnor U1143 (N_1143,N_695,N_206);
xor U1144 (N_1144,N_724,N_394);
or U1145 (N_1145,N_688,N_106);
or U1146 (N_1146,N_739,N_541);
nor U1147 (N_1147,N_150,N_947);
nand U1148 (N_1148,N_379,N_513);
and U1149 (N_1149,N_879,N_510);
nand U1150 (N_1150,N_419,N_297);
nand U1151 (N_1151,N_772,N_491);
or U1152 (N_1152,N_995,N_28);
or U1153 (N_1153,N_245,N_427);
and U1154 (N_1154,N_284,N_811);
or U1155 (N_1155,N_842,N_738);
nor U1156 (N_1156,N_795,N_318);
nor U1157 (N_1157,N_47,N_747);
or U1158 (N_1158,N_533,N_824);
nor U1159 (N_1159,N_354,N_236);
xnor U1160 (N_1160,N_881,N_780);
nand U1161 (N_1161,N_642,N_659);
nand U1162 (N_1162,N_127,N_138);
xnor U1163 (N_1163,N_197,N_251);
nand U1164 (N_1164,N_497,N_585);
xnor U1165 (N_1165,N_511,N_756);
xnor U1166 (N_1166,N_700,N_709);
nand U1167 (N_1167,N_390,N_798);
nor U1168 (N_1168,N_753,N_452);
and U1169 (N_1169,N_399,N_920);
nand U1170 (N_1170,N_103,N_396);
nand U1171 (N_1171,N_21,N_131);
nor U1172 (N_1172,N_765,N_82);
nand U1173 (N_1173,N_964,N_900);
and U1174 (N_1174,N_635,N_523);
and U1175 (N_1175,N_530,N_327);
or U1176 (N_1176,N_604,N_877);
nand U1177 (N_1177,N_682,N_517);
xor U1178 (N_1178,N_969,N_897);
or U1179 (N_1179,N_630,N_49);
or U1180 (N_1180,N_158,N_94);
and U1181 (N_1181,N_815,N_102);
and U1182 (N_1182,N_324,N_489);
or U1183 (N_1183,N_838,N_636);
nor U1184 (N_1184,N_524,N_65);
xnor U1185 (N_1185,N_445,N_273);
xnor U1186 (N_1186,N_845,N_962);
xnor U1187 (N_1187,N_122,N_777);
nor U1188 (N_1188,N_555,N_204);
and U1189 (N_1189,N_89,N_164);
and U1190 (N_1190,N_691,N_169);
xnor U1191 (N_1191,N_203,N_218);
xnor U1192 (N_1192,N_582,N_458);
nor U1193 (N_1193,N_238,N_830);
nand U1194 (N_1194,N_161,N_888);
and U1195 (N_1195,N_852,N_80);
nor U1196 (N_1196,N_679,N_690);
nand U1197 (N_1197,N_167,N_205);
xnor U1198 (N_1198,N_255,N_943);
and U1199 (N_1199,N_725,N_827);
nor U1200 (N_1200,N_425,N_162);
and U1201 (N_1201,N_748,N_761);
or U1202 (N_1202,N_626,N_915);
or U1203 (N_1203,N_870,N_258);
nand U1204 (N_1204,N_176,N_250);
xnor U1205 (N_1205,N_726,N_580);
xnor U1206 (N_1206,N_862,N_522);
xor U1207 (N_1207,N_508,N_463);
or U1208 (N_1208,N_351,N_596);
and U1209 (N_1209,N_730,N_277);
and U1210 (N_1210,N_704,N_901);
xor U1211 (N_1211,N_331,N_83);
and U1212 (N_1212,N_868,N_705);
nor U1213 (N_1213,N_641,N_110);
xor U1214 (N_1214,N_300,N_526);
nand U1215 (N_1215,N_490,N_872);
xor U1216 (N_1216,N_69,N_744);
nor U1217 (N_1217,N_189,N_806);
nand U1218 (N_1218,N_773,N_643);
or U1219 (N_1219,N_552,N_446);
xor U1220 (N_1220,N_17,N_320);
or U1221 (N_1221,N_899,N_821);
xnor U1222 (N_1222,N_409,N_720);
and U1223 (N_1223,N_241,N_623);
or U1224 (N_1224,N_779,N_614);
and U1225 (N_1225,N_310,N_677);
nand U1226 (N_1226,N_249,N_769);
xor U1227 (N_1227,N_119,N_126);
nor U1228 (N_1228,N_648,N_179);
or U1229 (N_1229,N_123,N_560);
nor U1230 (N_1230,N_484,N_389);
or U1231 (N_1231,N_107,N_805);
xor U1232 (N_1232,N_597,N_341);
and U1233 (N_1233,N_359,N_23);
xor U1234 (N_1234,N_914,N_837);
and U1235 (N_1235,N_952,N_711);
and U1236 (N_1236,N_878,N_875);
and U1237 (N_1237,N_11,N_412);
nor U1238 (N_1238,N_882,N_957);
nand U1239 (N_1239,N_619,N_742);
or U1240 (N_1240,N_857,N_72);
nand U1241 (N_1241,N_430,N_966);
nor U1242 (N_1242,N_918,N_979);
and U1243 (N_1243,N_867,N_142);
or U1244 (N_1244,N_426,N_115);
nand U1245 (N_1245,N_783,N_287);
and U1246 (N_1246,N_764,N_306);
xnor U1247 (N_1247,N_999,N_743);
xor U1248 (N_1248,N_130,N_5);
or U1249 (N_1249,N_265,N_542);
nor U1250 (N_1250,N_221,N_570);
nor U1251 (N_1251,N_216,N_214);
or U1252 (N_1252,N_217,N_982);
xnor U1253 (N_1253,N_734,N_649);
or U1254 (N_1254,N_468,N_496);
and U1255 (N_1255,N_817,N_193);
nor U1256 (N_1256,N_388,N_792);
xnor U1257 (N_1257,N_476,N_810);
xnor U1258 (N_1258,N_88,N_578);
nand U1259 (N_1259,N_505,N_248);
nor U1260 (N_1260,N_718,N_980);
nor U1261 (N_1261,N_632,N_951);
nand U1262 (N_1262,N_257,N_393);
xor U1263 (N_1263,N_921,N_759);
nand U1264 (N_1264,N_516,N_166);
xor U1265 (N_1265,N_104,N_63);
nand U1266 (N_1266,N_81,N_983);
nor U1267 (N_1267,N_763,N_281);
xor U1268 (N_1268,N_410,N_381);
nand U1269 (N_1269,N_159,N_909);
nor U1270 (N_1270,N_315,N_202);
and U1271 (N_1271,N_816,N_907);
or U1272 (N_1272,N_551,N_186);
xor U1273 (N_1273,N_651,N_210);
xor U1274 (N_1274,N_226,N_274);
and U1275 (N_1275,N_144,N_657);
nor U1276 (N_1276,N_475,N_108);
or U1277 (N_1277,N_68,N_586);
xnor U1278 (N_1278,N_453,N_800);
xnor U1279 (N_1279,N_603,N_696);
nor U1280 (N_1280,N_893,N_348);
nor U1281 (N_1281,N_243,N_506);
and U1282 (N_1282,N_435,N_685);
xnor U1283 (N_1283,N_561,N_652);
or U1284 (N_1284,N_634,N_280);
xor U1285 (N_1285,N_527,N_771);
or U1286 (N_1286,N_858,N_70);
nor U1287 (N_1287,N_55,N_149);
and U1288 (N_1288,N_645,N_185);
nor U1289 (N_1289,N_195,N_291);
nor U1290 (N_1290,N_15,N_368);
nand U1291 (N_1291,N_710,N_754);
and U1292 (N_1292,N_24,N_470);
and U1293 (N_1293,N_304,N_847);
or U1294 (N_1294,N_428,N_401);
nand U1295 (N_1295,N_486,N_913);
nor U1296 (N_1296,N_26,N_212);
and U1297 (N_1297,N_750,N_906);
xor U1298 (N_1298,N_403,N_295);
xor U1299 (N_1299,N_91,N_384);
and U1300 (N_1300,N_339,N_949);
nor U1301 (N_1301,N_349,N_188);
nand U1302 (N_1302,N_374,N_650);
or U1303 (N_1303,N_224,N_863);
and U1304 (N_1304,N_984,N_512);
and U1305 (N_1305,N_178,N_977);
xnor U1306 (N_1306,N_125,N_680);
and U1307 (N_1307,N_853,N_312);
and U1308 (N_1308,N_646,N_328);
or U1309 (N_1309,N_246,N_114);
nor U1310 (N_1310,N_873,N_940);
nand U1311 (N_1311,N_353,N_42);
xor U1312 (N_1312,N_364,N_335);
and U1313 (N_1313,N_272,N_965);
or U1314 (N_1314,N_534,N_928);
and U1315 (N_1315,N_825,N_973);
xnor U1316 (N_1316,N_556,N_147);
xnor U1317 (N_1317,N_565,N_653);
nor U1318 (N_1318,N_787,N_481);
nand U1319 (N_1319,N_367,N_958);
nor U1320 (N_1320,N_1,N_707);
and U1321 (N_1321,N_175,N_538);
and U1322 (N_1322,N_934,N_885);
or U1323 (N_1323,N_432,N_198);
xor U1324 (N_1324,N_74,N_440);
nand U1325 (N_1325,N_702,N_360);
and U1326 (N_1326,N_575,N_563);
or U1327 (N_1327,N_14,N_762);
nand U1328 (N_1328,N_518,N_190);
nor U1329 (N_1329,N_487,N_583);
nand U1330 (N_1330,N_978,N_233);
xor U1331 (N_1331,N_959,N_991);
or U1332 (N_1332,N_774,N_100);
or U1333 (N_1333,N_495,N_174);
or U1334 (N_1334,N_474,N_493);
nand U1335 (N_1335,N_151,N_558);
and U1336 (N_1336,N_283,N_892);
and U1337 (N_1337,N_851,N_889);
xnor U1338 (N_1338,N_544,N_347);
or U1339 (N_1339,N_504,N_741);
and U1340 (N_1340,N_322,N_543);
xnor U1341 (N_1341,N_961,N_997);
nand U1342 (N_1342,N_992,N_664);
or U1343 (N_1343,N_884,N_73);
nand U1344 (N_1344,N_832,N_803);
nor U1345 (N_1345,N_438,N_788);
nor U1346 (N_1346,N_35,N_610);
or U1347 (N_1347,N_472,N_633);
or U1348 (N_1348,N_687,N_116);
nand U1349 (N_1349,N_299,N_926);
and U1350 (N_1350,N_133,N_377);
nand U1351 (N_1351,N_229,N_286);
xnor U1352 (N_1352,N_323,N_568);
or U1353 (N_1353,N_369,N_37);
and U1354 (N_1354,N_223,N_942);
nand U1355 (N_1355,N_373,N_276);
and U1356 (N_1356,N_316,N_766);
and U1357 (N_1357,N_30,N_515);
or U1358 (N_1358,N_545,N_536);
nand U1359 (N_1359,N_818,N_242);
xnor U1360 (N_1360,N_564,N_58);
and U1361 (N_1361,N_296,N_904);
nor U1362 (N_1362,N_279,N_715);
xnor U1363 (N_1363,N_378,N_278);
or U1364 (N_1364,N_362,N_950);
or U1365 (N_1365,N_625,N_621);
or U1366 (N_1366,N_48,N_51);
xnor U1367 (N_1367,N_802,N_289);
xor U1368 (N_1368,N_336,N_874);
nor U1369 (N_1369,N_140,N_43);
xor U1370 (N_1370,N_268,N_294);
nand U1371 (N_1371,N_499,N_252);
nand U1372 (N_1372,N_712,N_232);
nor U1373 (N_1373,N_61,N_528);
nand U1374 (N_1374,N_199,N_253);
nor U1375 (N_1375,N_804,N_562);
nand U1376 (N_1376,N_211,N_101);
nor U1377 (N_1377,N_113,N_683);
and U1378 (N_1378,N_168,N_56);
xor U1379 (N_1379,N_954,N_450);
and U1380 (N_1380,N_201,N_550);
xnor U1381 (N_1381,N_267,N_105);
xor U1382 (N_1382,N_668,N_90);
nand U1383 (N_1383,N_514,N_466);
nor U1384 (N_1384,N_826,N_488);
or U1385 (N_1385,N_172,N_376);
or U1386 (N_1386,N_600,N_423);
nor U1387 (N_1387,N_346,N_96);
and U1388 (N_1388,N_706,N_333);
nor U1389 (N_1389,N_173,N_656);
nand U1390 (N_1390,N_605,N_654);
or U1391 (N_1391,N_416,N_22);
and U1392 (N_1392,N_671,N_448);
nor U1393 (N_1393,N_231,N_109);
nand U1394 (N_1394,N_477,N_929);
nand U1395 (N_1395,N_442,N_402);
nand U1396 (N_1396,N_946,N_494);
nand U1397 (N_1397,N_124,N_789);
or U1398 (N_1398,N_303,N_974);
nor U1399 (N_1399,N_675,N_332);
and U1400 (N_1400,N_209,N_719);
nand U1401 (N_1401,N_77,N_644);
or U1402 (N_1402,N_678,N_344);
xnor U1403 (N_1403,N_569,N_247);
xor U1404 (N_1404,N_820,N_93);
and U1405 (N_1405,N_945,N_41);
nand U1406 (N_1406,N_404,N_75);
and U1407 (N_1407,N_0,N_152);
nor U1408 (N_1408,N_177,N_689);
or U1409 (N_1409,N_4,N_592);
and U1410 (N_1410,N_529,N_449);
nand U1411 (N_1411,N_970,N_380);
or U1412 (N_1412,N_71,N_927);
or U1413 (N_1413,N_372,N_673);
or U1414 (N_1414,N_503,N_7);
and U1415 (N_1415,N_757,N_593);
nor U1416 (N_1416,N_345,N_703);
nor U1417 (N_1417,N_993,N_611);
or U1418 (N_1418,N_613,N_365);
xor U1419 (N_1419,N_939,N_146);
xnor U1420 (N_1420,N_576,N_755);
or U1421 (N_1421,N_925,N_554);
nand U1422 (N_1422,N_443,N_601);
nand U1423 (N_1423,N_785,N_727);
nor U1424 (N_1424,N_944,N_574);
xnor U1425 (N_1425,N_571,N_850);
and U1426 (N_1426,N_285,N_20);
nand U1427 (N_1427,N_13,N_840);
xor U1428 (N_1428,N_553,N_207);
and U1429 (N_1429,N_782,N_92);
and U1430 (N_1430,N_148,N_464);
nand U1431 (N_1431,N_839,N_12);
nand U1432 (N_1432,N_722,N_637);
and U1433 (N_1433,N_540,N_382);
nand U1434 (N_1434,N_181,N_579);
or U1435 (N_1435,N_735,N_848);
nor U1436 (N_1436,N_968,N_165);
xnor U1437 (N_1437,N_479,N_729);
nor U1438 (N_1438,N_462,N_865);
nor U1439 (N_1439,N_437,N_617);
nor U1440 (N_1440,N_731,N_559);
or U1441 (N_1441,N_908,N_375);
xor U1442 (N_1442,N_54,N_40);
nand U1443 (N_1443,N_340,N_752);
and U1444 (N_1444,N_924,N_836);
or U1445 (N_1445,N_356,N_200);
or U1446 (N_1446,N_325,N_183);
nor U1447 (N_1447,N_10,N_846);
and U1448 (N_1448,N_694,N_776);
and U1449 (N_1449,N_799,N_786);
or U1450 (N_1450,N_667,N_153);
nor U1451 (N_1451,N_288,N_894);
or U1452 (N_1452,N_398,N_27);
nor U1453 (N_1453,N_194,N_31);
xnor U1454 (N_1454,N_595,N_733);
or U1455 (N_1455,N_539,N_693);
or U1456 (N_1456,N_8,N_118);
or U1457 (N_1457,N_39,N_98);
nand U1458 (N_1458,N_572,N_282);
or U1459 (N_1459,N_890,N_95);
and U1460 (N_1460,N_835,N_25);
or U1461 (N_1461,N_548,N_196);
nor U1462 (N_1462,N_329,N_436);
and U1463 (N_1463,N_699,N_145);
xnor U1464 (N_1464,N_919,N_854);
nand U1465 (N_1465,N_624,N_308);
nor U1466 (N_1466,N_234,N_370);
or U1467 (N_1467,N_135,N_686);
xnor U1468 (N_1468,N_237,N_658);
or U1469 (N_1469,N_723,N_383);
xor U1470 (N_1470,N_99,N_457);
nand U1471 (N_1471,N_871,N_337);
and U1472 (N_1472,N_986,N_213);
or U1473 (N_1473,N_262,N_480);
xor U1474 (N_1474,N_886,N_240);
or U1475 (N_1475,N_843,N_813);
and U1476 (N_1476,N_589,N_612);
and U1477 (N_1477,N_334,N_411);
or U1478 (N_1478,N_655,N_669);
xnor U1479 (N_1479,N_896,N_606);
and U1480 (N_1480,N_588,N_385);
and U1481 (N_1481,N_298,N_941);
and U1482 (N_1482,N_661,N_215);
nand U1483 (N_1483,N_721,N_549);
nand U1484 (N_1484,N_270,N_829);
xor U1485 (N_1485,N_260,N_451);
nand U1486 (N_1486,N_112,N_629);
nor U1487 (N_1487,N_666,N_129);
xor U1488 (N_1488,N_717,N_45);
xor U1489 (N_1489,N_64,N_953);
xor U1490 (N_1490,N_791,N_912);
or U1491 (N_1491,N_902,N_313);
or U1492 (N_1492,N_760,N_794);
nand U1493 (N_1493,N_784,N_844);
or U1494 (N_1494,N_266,N_6);
nand U1495 (N_1495,N_187,N_714);
and U1496 (N_1496,N_414,N_434);
xor U1497 (N_1497,N_302,N_400);
xor U1498 (N_1498,N_134,N_698);
and U1499 (N_1499,N_860,N_930);
xnor U1500 (N_1500,N_191,N_654);
nand U1501 (N_1501,N_147,N_516);
xnor U1502 (N_1502,N_646,N_126);
nor U1503 (N_1503,N_211,N_361);
nand U1504 (N_1504,N_774,N_457);
xnor U1505 (N_1505,N_86,N_987);
or U1506 (N_1506,N_823,N_476);
or U1507 (N_1507,N_218,N_565);
nand U1508 (N_1508,N_46,N_858);
xnor U1509 (N_1509,N_334,N_46);
nor U1510 (N_1510,N_975,N_200);
xor U1511 (N_1511,N_216,N_227);
xor U1512 (N_1512,N_928,N_811);
nor U1513 (N_1513,N_237,N_831);
xnor U1514 (N_1514,N_965,N_739);
nor U1515 (N_1515,N_14,N_391);
or U1516 (N_1516,N_410,N_462);
xnor U1517 (N_1517,N_791,N_459);
nor U1518 (N_1518,N_532,N_398);
nand U1519 (N_1519,N_324,N_648);
xor U1520 (N_1520,N_982,N_26);
nor U1521 (N_1521,N_977,N_962);
and U1522 (N_1522,N_714,N_997);
xnor U1523 (N_1523,N_693,N_843);
nor U1524 (N_1524,N_31,N_467);
or U1525 (N_1525,N_466,N_681);
nand U1526 (N_1526,N_666,N_187);
or U1527 (N_1527,N_662,N_598);
or U1528 (N_1528,N_269,N_943);
xor U1529 (N_1529,N_473,N_558);
nor U1530 (N_1530,N_127,N_51);
nor U1531 (N_1531,N_82,N_45);
or U1532 (N_1532,N_891,N_182);
nand U1533 (N_1533,N_304,N_785);
xor U1534 (N_1534,N_800,N_951);
and U1535 (N_1535,N_146,N_416);
or U1536 (N_1536,N_975,N_643);
or U1537 (N_1537,N_323,N_626);
or U1538 (N_1538,N_543,N_880);
and U1539 (N_1539,N_259,N_512);
and U1540 (N_1540,N_410,N_985);
nand U1541 (N_1541,N_1,N_113);
nand U1542 (N_1542,N_294,N_634);
or U1543 (N_1543,N_651,N_966);
or U1544 (N_1544,N_148,N_801);
or U1545 (N_1545,N_498,N_314);
or U1546 (N_1546,N_75,N_42);
nor U1547 (N_1547,N_17,N_841);
nand U1548 (N_1548,N_583,N_897);
nand U1549 (N_1549,N_495,N_678);
nand U1550 (N_1550,N_863,N_189);
and U1551 (N_1551,N_684,N_182);
and U1552 (N_1552,N_88,N_755);
or U1553 (N_1553,N_242,N_847);
or U1554 (N_1554,N_127,N_183);
xnor U1555 (N_1555,N_50,N_141);
or U1556 (N_1556,N_62,N_467);
nor U1557 (N_1557,N_870,N_802);
and U1558 (N_1558,N_654,N_572);
nor U1559 (N_1559,N_173,N_961);
nor U1560 (N_1560,N_491,N_482);
nor U1561 (N_1561,N_724,N_295);
or U1562 (N_1562,N_804,N_673);
nand U1563 (N_1563,N_907,N_786);
or U1564 (N_1564,N_423,N_773);
nor U1565 (N_1565,N_148,N_877);
or U1566 (N_1566,N_766,N_459);
nand U1567 (N_1567,N_467,N_843);
or U1568 (N_1568,N_460,N_735);
nor U1569 (N_1569,N_379,N_601);
nor U1570 (N_1570,N_472,N_505);
and U1571 (N_1571,N_820,N_338);
xnor U1572 (N_1572,N_639,N_260);
or U1573 (N_1573,N_639,N_491);
nor U1574 (N_1574,N_913,N_354);
nand U1575 (N_1575,N_48,N_781);
and U1576 (N_1576,N_904,N_579);
xnor U1577 (N_1577,N_792,N_922);
or U1578 (N_1578,N_336,N_307);
nand U1579 (N_1579,N_211,N_75);
nand U1580 (N_1580,N_562,N_814);
or U1581 (N_1581,N_843,N_830);
or U1582 (N_1582,N_665,N_396);
and U1583 (N_1583,N_982,N_92);
or U1584 (N_1584,N_766,N_19);
or U1585 (N_1585,N_664,N_509);
and U1586 (N_1586,N_420,N_801);
or U1587 (N_1587,N_866,N_937);
and U1588 (N_1588,N_531,N_38);
nor U1589 (N_1589,N_612,N_6);
nor U1590 (N_1590,N_481,N_35);
nand U1591 (N_1591,N_314,N_823);
nor U1592 (N_1592,N_234,N_480);
nand U1593 (N_1593,N_193,N_914);
nor U1594 (N_1594,N_765,N_594);
and U1595 (N_1595,N_88,N_215);
xnor U1596 (N_1596,N_597,N_425);
nor U1597 (N_1597,N_818,N_573);
or U1598 (N_1598,N_955,N_19);
nor U1599 (N_1599,N_114,N_600);
nand U1600 (N_1600,N_411,N_527);
nand U1601 (N_1601,N_500,N_861);
nand U1602 (N_1602,N_825,N_604);
or U1603 (N_1603,N_956,N_802);
nor U1604 (N_1604,N_407,N_230);
nor U1605 (N_1605,N_306,N_881);
nor U1606 (N_1606,N_46,N_673);
xnor U1607 (N_1607,N_991,N_420);
nand U1608 (N_1608,N_372,N_907);
xnor U1609 (N_1609,N_3,N_299);
and U1610 (N_1610,N_0,N_422);
and U1611 (N_1611,N_830,N_371);
xnor U1612 (N_1612,N_378,N_206);
or U1613 (N_1613,N_818,N_428);
and U1614 (N_1614,N_17,N_481);
or U1615 (N_1615,N_30,N_771);
nor U1616 (N_1616,N_452,N_297);
xor U1617 (N_1617,N_824,N_65);
xnor U1618 (N_1618,N_361,N_755);
and U1619 (N_1619,N_559,N_311);
or U1620 (N_1620,N_184,N_871);
or U1621 (N_1621,N_962,N_42);
or U1622 (N_1622,N_479,N_40);
and U1623 (N_1623,N_873,N_782);
xor U1624 (N_1624,N_974,N_333);
nor U1625 (N_1625,N_264,N_993);
and U1626 (N_1626,N_360,N_370);
nor U1627 (N_1627,N_860,N_565);
xor U1628 (N_1628,N_994,N_621);
or U1629 (N_1629,N_318,N_751);
nand U1630 (N_1630,N_1,N_552);
xor U1631 (N_1631,N_880,N_667);
nor U1632 (N_1632,N_885,N_129);
and U1633 (N_1633,N_223,N_411);
and U1634 (N_1634,N_840,N_629);
and U1635 (N_1635,N_731,N_378);
nor U1636 (N_1636,N_348,N_258);
and U1637 (N_1637,N_306,N_682);
and U1638 (N_1638,N_413,N_808);
and U1639 (N_1639,N_593,N_562);
and U1640 (N_1640,N_236,N_483);
nor U1641 (N_1641,N_934,N_199);
nor U1642 (N_1642,N_560,N_201);
and U1643 (N_1643,N_268,N_866);
nor U1644 (N_1644,N_604,N_116);
and U1645 (N_1645,N_115,N_77);
and U1646 (N_1646,N_521,N_953);
or U1647 (N_1647,N_579,N_531);
nand U1648 (N_1648,N_214,N_303);
and U1649 (N_1649,N_376,N_9);
nor U1650 (N_1650,N_179,N_539);
or U1651 (N_1651,N_37,N_379);
xor U1652 (N_1652,N_250,N_126);
nor U1653 (N_1653,N_963,N_754);
nand U1654 (N_1654,N_966,N_33);
and U1655 (N_1655,N_987,N_978);
xor U1656 (N_1656,N_489,N_144);
and U1657 (N_1657,N_419,N_541);
and U1658 (N_1658,N_743,N_812);
and U1659 (N_1659,N_183,N_933);
nor U1660 (N_1660,N_437,N_195);
nor U1661 (N_1661,N_764,N_191);
nand U1662 (N_1662,N_994,N_379);
and U1663 (N_1663,N_809,N_628);
or U1664 (N_1664,N_448,N_731);
nor U1665 (N_1665,N_159,N_177);
nor U1666 (N_1666,N_25,N_174);
and U1667 (N_1667,N_471,N_213);
xor U1668 (N_1668,N_53,N_192);
nor U1669 (N_1669,N_548,N_504);
nor U1670 (N_1670,N_401,N_597);
nor U1671 (N_1671,N_46,N_880);
nand U1672 (N_1672,N_506,N_99);
nor U1673 (N_1673,N_825,N_422);
and U1674 (N_1674,N_499,N_240);
nand U1675 (N_1675,N_847,N_438);
nand U1676 (N_1676,N_510,N_759);
and U1677 (N_1677,N_142,N_947);
nand U1678 (N_1678,N_335,N_37);
or U1679 (N_1679,N_611,N_895);
and U1680 (N_1680,N_285,N_419);
nor U1681 (N_1681,N_970,N_139);
or U1682 (N_1682,N_32,N_429);
and U1683 (N_1683,N_466,N_316);
xnor U1684 (N_1684,N_255,N_364);
or U1685 (N_1685,N_98,N_427);
nand U1686 (N_1686,N_737,N_882);
nor U1687 (N_1687,N_515,N_792);
xnor U1688 (N_1688,N_933,N_605);
and U1689 (N_1689,N_614,N_367);
xor U1690 (N_1690,N_664,N_994);
and U1691 (N_1691,N_336,N_930);
nor U1692 (N_1692,N_907,N_970);
nor U1693 (N_1693,N_339,N_984);
nand U1694 (N_1694,N_609,N_707);
xor U1695 (N_1695,N_634,N_895);
xor U1696 (N_1696,N_782,N_31);
or U1697 (N_1697,N_415,N_565);
nand U1698 (N_1698,N_939,N_539);
nor U1699 (N_1699,N_960,N_682);
nor U1700 (N_1700,N_255,N_312);
nand U1701 (N_1701,N_934,N_815);
and U1702 (N_1702,N_956,N_447);
nand U1703 (N_1703,N_544,N_251);
or U1704 (N_1704,N_589,N_750);
nand U1705 (N_1705,N_664,N_448);
or U1706 (N_1706,N_147,N_811);
xnor U1707 (N_1707,N_548,N_311);
xnor U1708 (N_1708,N_394,N_541);
or U1709 (N_1709,N_428,N_215);
nand U1710 (N_1710,N_485,N_515);
xor U1711 (N_1711,N_389,N_306);
xor U1712 (N_1712,N_622,N_625);
xor U1713 (N_1713,N_899,N_627);
and U1714 (N_1714,N_498,N_165);
nand U1715 (N_1715,N_255,N_568);
xor U1716 (N_1716,N_808,N_136);
xor U1717 (N_1717,N_253,N_321);
nand U1718 (N_1718,N_859,N_157);
nand U1719 (N_1719,N_98,N_670);
or U1720 (N_1720,N_648,N_724);
and U1721 (N_1721,N_755,N_698);
nor U1722 (N_1722,N_712,N_266);
xnor U1723 (N_1723,N_352,N_786);
nand U1724 (N_1724,N_770,N_834);
nand U1725 (N_1725,N_28,N_498);
nor U1726 (N_1726,N_41,N_162);
nand U1727 (N_1727,N_344,N_316);
and U1728 (N_1728,N_108,N_981);
and U1729 (N_1729,N_506,N_667);
nor U1730 (N_1730,N_858,N_186);
nor U1731 (N_1731,N_391,N_874);
or U1732 (N_1732,N_421,N_636);
or U1733 (N_1733,N_195,N_583);
and U1734 (N_1734,N_565,N_847);
or U1735 (N_1735,N_860,N_896);
nand U1736 (N_1736,N_299,N_828);
nand U1737 (N_1737,N_971,N_419);
and U1738 (N_1738,N_338,N_941);
xnor U1739 (N_1739,N_928,N_199);
and U1740 (N_1740,N_690,N_992);
xnor U1741 (N_1741,N_378,N_987);
xnor U1742 (N_1742,N_183,N_268);
and U1743 (N_1743,N_950,N_66);
or U1744 (N_1744,N_128,N_203);
and U1745 (N_1745,N_630,N_157);
nand U1746 (N_1746,N_504,N_871);
and U1747 (N_1747,N_731,N_976);
xnor U1748 (N_1748,N_590,N_495);
or U1749 (N_1749,N_419,N_429);
or U1750 (N_1750,N_458,N_852);
xor U1751 (N_1751,N_324,N_951);
nor U1752 (N_1752,N_430,N_708);
xnor U1753 (N_1753,N_313,N_546);
or U1754 (N_1754,N_411,N_156);
nand U1755 (N_1755,N_864,N_277);
nand U1756 (N_1756,N_29,N_609);
nand U1757 (N_1757,N_823,N_453);
and U1758 (N_1758,N_557,N_422);
nand U1759 (N_1759,N_524,N_730);
nand U1760 (N_1760,N_641,N_188);
xnor U1761 (N_1761,N_423,N_456);
nand U1762 (N_1762,N_944,N_87);
xnor U1763 (N_1763,N_332,N_3);
and U1764 (N_1764,N_534,N_550);
and U1765 (N_1765,N_40,N_859);
nor U1766 (N_1766,N_192,N_73);
or U1767 (N_1767,N_266,N_450);
nand U1768 (N_1768,N_848,N_103);
xor U1769 (N_1769,N_134,N_537);
xor U1770 (N_1770,N_310,N_9);
and U1771 (N_1771,N_686,N_643);
nor U1772 (N_1772,N_830,N_191);
xor U1773 (N_1773,N_497,N_37);
nand U1774 (N_1774,N_635,N_883);
xnor U1775 (N_1775,N_88,N_843);
nor U1776 (N_1776,N_142,N_21);
nor U1777 (N_1777,N_591,N_942);
xor U1778 (N_1778,N_751,N_504);
nor U1779 (N_1779,N_651,N_232);
and U1780 (N_1780,N_278,N_264);
or U1781 (N_1781,N_3,N_811);
nor U1782 (N_1782,N_106,N_197);
nor U1783 (N_1783,N_368,N_364);
or U1784 (N_1784,N_567,N_442);
xnor U1785 (N_1785,N_71,N_837);
nor U1786 (N_1786,N_820,N_192);
nor U1787 (N_1787,N_782,N_506);
xor U1788 (N_1788,N_748,N_52);
nand U1789 (N_1789,N_598,N_114);
xor U1790 (N_1790,N_663,N_845);
xnor U1791 (N_1791,N_131,N_355);
nand U1792 (N_1792,N_858,N_525);
or U1793 (N_1793,N_304,N_765);
nand U1794 (N_1794,N_69,N_160);
xor U1795 (N_1795,N_23,N_30);
xor U1796 (N_1796,N_794,N_884);
or U1797 (N_1797,N_772,N_651);
xor U1798 (N_1798,N_72,N_997);
and U1799 (N_1799,N_612,N_193);
nor U1800 (N_1800,N_310,N_105);
and U1801 (N_1801,N_770,N_500);
nor U1802 (N_1802,N_842,N_26);
and U1803 (N_1803,N_839,N_476);
nand U1804 (N_1804,N_922,N_545);
xor U1805 (N_1805,N_548,N_870);
or U1806 (N_1806,N_885,N_636);
and U1807 (N_1807,N_486,N_379);
or U1808 (N_1808,N_843,N_715);
xnor U1809 (N_1809,N_953,N_925);
nor U1810 (N_1810,N_256,N_636);
and U1811 (N_1811,N_782,N_375);
and U1812 (N_1812,N_252,N_284);
nand U1813 (N_1813,N_266,N_873);
nor U1814 (N_1814,N_385,N_960);
nand U1815 (N_1815,N_568,N_196);
nand U1816 (N_1816,N_467,N_823);
and U1817 (N_1817,N_340,N_965);
nor U1818 (N_1818,N_827,N_74);
and U1819 (N_1819,N_160,N_347);
or U1820 (N_1820,N_457,N_179);
or U1821 (N_1821,N_260,N_657);
nor U1822 (N_1822,N_904,N_260);
nor U1823 (N_1823,N_322,N_522);
nor U1824 (N_1824,N_950,N_232);
or U1825 (N_1825,N_808,N_543);
and U1826 (N_1826,N_993,N_452);
and U1827 (N_1827,N_276,N_422);
nand U1828 (N_1828,N_74,N_111);
nand U1829 (N_1829,N_968,N_170);
and U1830 (N_1830,N_417,N_547);
xor U1831 (N_1831,N_931,N_128);
or U1832 (N_1832,N_780,N_509);
nor U1833 (N_1833,N_474,N_253);
or U1834 (N_1834,N_571,N_260);
nand U1835 (N_1835,N_123,N_827);
nand U1836 (N_1836,N_582,N_637);
nand U1837 (N_1837,N_910,N_170);
or U1838 (N_1838,N_464,N_608);
and U1839 (N_1839,N_9,N_633);
nor U1840 (N_1840,N_769,N_917);
and U1841 (N_1841,N_9,N_103);
xnor U1842 (N_1842,N_344,N_270);
nand U1843 (N_1843,N_5,N_523);
nand U1844 (N_1844,N_387,N_871);
and U1845 (N_1845,N_379,N_264);
nand U1846 (N_1846,N_843,N_783);
or U1847 (N_1847,N_284,N_278);
nor U1848 (N_1848,N_642,N_981);
nor U1849 (N_1849,N_974,N_413);
nor U1850 (N_1850,N_883,N_877);
nand U1851 (N_1851,N_270,N_981);
nor U1852 (N_1852,N_782,N_242);
or U1853 (N_1853,N_608,N_280);
xnor U1854 (N_1854,N_990,N_989);
nand U1855 (N_1855,N_590,N_72);
xnor U1856 (N_1856,N_904,N_908);
nor U1857 (N_1857,N_373,N_564);
xnor U1858 (N_1858,N_416,N_558);
or U1859 (N_1859,N_303,N_707);
xnor U1860 (N_1860,N_684,N_664);
xor U1861 (N_1861,N_977,N_87);
and U1862 (N_1862,N_264,N_745);
and U1863 (N_1863,N_25,N_548);
and U1864 (N_1864,N_95,N_294);
nor U1865 (N_1865,N_718,N_569);
and U1866 (N_1866,N_769,N_340);
and U1867 (N_1867,N_363,N_864);
nor U1868 (N_1868,N_41,N_949);
or U1869 (N_1869,N_468,N_426);
nor U1870 (N_1870,N_153,N_149);
nor U1871 (N_1871,N_9,N_397);
or U1872 (N_1872,N_684,N_115);
or U1873 (N_1873,N_881,N_539);
nand U1874 (N_1874,N_413,N_261);
nand U1875 (N_1875,N_234,N_489);
and U1876 (N_1876,N_487,N_754);
or U1877 (N_1877,N_711,N_389);
nand U1878 (N_1878,N_300,N_253);
and U1879 (N_1879,N_906,N_58);
or U1880 (N_1880,N_810,N_90);
and U1881 (N_1881,N_672,N_769);
nand U1882 (N_1882,N_883,N_124);
nor U1883 (N_1883,N_605,N_523);
nand U1884 (N_1884,N_705,N_360);
nor U1885 (N_1885,N_408,N_83);
nor U1886 (N_1886,N_670,N_757);
or U1887 (N_1887,N_600,N_24);
xnor U1888 (N_1888,N_707,N_892);
xor U1889 (N_1889,N_813,N_606);
xor U1890 (N_1890,N_581,N_575);
and U1891 (N_1891,N_842,N_739);
nand U1892 (N_1892,N_239,N_365);
xor U1893 (N_1893,N_176,N_169);
nand U1894 (N_1894,N_254,N_438);
nor U1895 (N_1895,N_345,N_388);
nand U1896 (N_1896,N_539,N_253);
xor U1897 (N_1897,N_618,N_904);
nor U1898 (N_1898,N_399,N_127);
and U1899 (N_1899,N_841,N_735);
nor U1900 (N_1900,N_732,N_327);
nand U1901 (N_1901,N_531,N_113);
nand U1902 (N_1902,N_26,N_773);
or U1903 (N_1903,N_0,N_328);
or U1904 (N_1904,N_747,N_476);
xnor U1905 (N_1905,N_628,N_839);
xnor U1906 (N_1906,N_960,N_73);
nor U1907 (N_1907,N_382,N_502);
nor U1908 (N_1908,N_405,N_470);
or U1909 (N_1909,N_907,N_547);
and U1910 (N_1910,N_746,N_130);
and U1911 (N_1911,N_617,N_838);
and U1912 (N_1912,N_332,N_710);
and U1913 (N_1913,N_53,N_617);
nand U1914 (N_1914,N_932,N_810);
nor U1915 (N_1915,N_753,N_102);
or U1916 (N_1916,N_332,N_39);
or U1917 (N_1917,N_654,N_185);
or U1918 (N_1918,N_586,N_826);
or U1919 (N_1919,N_166,N_685);
nor U1920 (N_1920,N_745,N_454);
or U1921 (N_1921,N_884,N_242);
nand U1922 (N_1922,N_759,N_659);
or U1923 (N_1923,N_862,N_141);
nand U1924 (N_1924,N_452,N_618);
nor U1925 (N_1925,N_396,N_630);
nor U1926 (N_1926,N_495,N_508);
or U1927 (N_1927,N_727,N_411);
nor U1928 (N_1928,N_4,N_949);
or U1929 (N_1929,N_174,N_51);
nor U1930 (N_1930,N_593,N_961);
or U1931 (N_1931,N_797,N_943);
or U1932 (N_1932,N_118,N_85);
nand U1933 (N_1933,N_684,N_290);
and U1934 (N_1934,N_63,N_727);
and U1935 (N_1935,N_73,N_563);
and U1936 (N_1936,N_301,N_908);
or U1937 (N_1937,N_618,N_630);
and U1938 (N_1938,N_68,N_919);
and U1939 (N_1939,N_2,N_365);
or U1940 (N_1940,N_747,N_252);
nand U1941 (N_1941,N_850,N_960);
and U1942 (N_1942,N_970,N_455);
and U1943 (N_1943,N_672,N_751);
and U1944 (N_1944,N_861,N_956);
nand U1945 (N_1945,N_679,N_448);
or U1946 (N_1946,N_63,N_510);
nor U1947 (N_1947,N_653,N_737);
nand U1948 (N_1948,N_424,N_499);
nor U1949 (N_1949,N_69,N_560);
nand U1950 (N_1950,N_808,N_687);
nor U1951 (N_1951,N_341,N_661);
and U1952 (N_1952,N_517,N_267);
nand U1953 (N_1953,N_931,N_473);
nand U1954 (N_1954,N_290,N_635);
xor U1955 (N_1955,N_132,N_705);
xor U1956 (N_1956,N_103,N_833);
xor U1957 (N_1957,N_389,N_94);
and U1958 (N_1958,N_633,N_196);
or U1959 (N_1959,N_293,N_777);
xnor U1960 (N_1960,N_487,N_542);
nand U1961 (N_1961,N_647,N_949);
nor U1962 (N_1962,N_385,N_749);
and U1963 (N_1963,N_892,N_864);
xor U1964 (N_1964,N_921,N_687);
nand U1965 (N_1965,N_47,N_383);
nand U1966 (N_1966,N_612,N_925);
nand U1967 (N_1967,N_764,N_89);
and U1968 (N_1968,N_316,N_452);
xnor U1969 (N_1969,N_455,N_953);
and U1970 (N_1970,N_735,N_125);
and U1971 (N_1971,N_503,N_155);
nand U1972 (N_1972,N_90,N_273);
and U1973 (N_1973,N_552,N_241);
xor U1974 (N_1974,N_2,N_534);
or U1975 (N_1975,N_60,N_4);
and U1976 (N_1976,N_177,N_256);
xor U1977 (N_1977,N_525,N_211);
nor U1978 (N_1978,N_816,N_331);
xnor U1979 (N_1979,N_474,N_105);
xnor U1980 (N_1980,N_49,N_260);
nand U1981 (N_1981,N_173,N_619);
nor U1982 (N_1982,N_666,N_662);
nor U1983 (N_1983,N_891,N_388);
nor U1984 (N_1984,N_138,N_891);
or U1985 (N_1985,N_548,N_626);
and U1986 (N_1986,N_850,N_423);
nand U1987 (N_1987,N_627,N_427);
or U1988 (N_1988,N_513,N_303);
xnor U1989 (N_1989,N_86,N_376);
xnor U1990 (N_1990,N_629,N_59);
xnor U1991 (N_1991,N_191,N_293);
nand U1992 (N_1992,N_589,N_597);
nand U1993 (N_1993,N_186,N_120);
nand U1994 (N_1994,N_68,N_92);
nand U1995 (N_1995,N_914,N_181);
or U1996 (N_1996,N_205,N_688);
nor U1997 (N_1997,N_414,N_573);
xnor U1998 (N_1998,N_143,N_322);
nand U1999 (N_1999,N_936,N_182);
xor U2000 (N_2000,N_1023,N_1402);
or U2001 (N_2001,N_1191,N_1911);
or U2002 (N_2002,N_1861,N_1229);
nand U2003 (N_2003,N_1112,N_1493);
or U2004 (N_2004,N_1097,N_1894);
and U2005 (N_2005,N_1615,N_1814);
or U2006 (N_2006,N_1523,N_1371);
xnor U2007 (N_2007,N_1537,N_1723);
and U2008 (N_2008,N_1747,N_1156);
nor U2009 (N_2009,N_1059,N_1483);
and U2010 (N_2010,N_1282,N_1575);
nand U2011 (N_2011,N_1104,N_1953);
nor U2012 (N_2012,N_1708,N_1225);
nand U2013 (N_2013,N_1611,N_1718);
and U2014 (N_2014,N_1734,N_1871);
nand U2015 (N_2015,N_1567,N_1391);
nor U2016 (N_2016,N_1377,N_1100);
nor U2017 (N_2017,N_1548,N_1950);
xnor U2018 (N_2018,N_1613,N_1769);
and U2019 (N_2019,N_1269,N_1686);
and U2020 (N_2020,N_1754,N_1743);
and U2021 (N_2021,N_1499,N_1252);
and U2022 (N_2022,N_1309,N_1710);
or U2023 (N_2023,N_1595,N_1116);
and U2024 (N_2024,N_1141,N_1995);
and U2025 (N_2025,N_1588,N_1698);
xor U2026 (N_2026,N_1713,N_1078);
nor U2027 (N_2027,N_1699,N_1964);
nand U2028 (N_2028,N_1675,N_1832);
nor U2029 (N_2029,N_1153,N_1135);
or U2030 (N_2030,N_1924,N_1621);
nand U2031 (N_2031,N_1159,N_1014);
nor U2032 (N_2032,N_1876,N_1231);
and U2033 (N_2033,N_1981,N_1232);
nor U2034 (N_2034,N_1239,N_1126);
nor U2035 (N_2035,N_1919,N_1898);
nand U2036 (N_2036,N_1749,N_1857);
and U2037 (N_2037,N_1230,N_1323);
or U2038 (N_2038,N_1477,N_1016);
nand U2039 (N_2039,N_1730,N_1461);
nor U2040 (N_2040,N_1865,N_1278);
xor U2041 (N_2041,N_1004,N_1008);
nand U2042 (N_2042,N_1958,N_1322);
nand U2043 (N_2043,N_1934,N_1666);
or U2044 (N_2044,N_1224,N_1353);
or U2045 (N_2045,N_1329,N_1390);
nor U2046 (N_2046,N_1152,N_1201);
or U2047 (N_2047,N_1826,N_1987);
and U2048 (N_2048,N_1733,N_1923);
nand U2049 (N_2049,N_1338,N_1946);
nor U2050 (N_2050,N_1645,N_1512);
and U2051 (N_2051,N_1080,N_1472);
or U2052 (N_2052,N_1728,N_1850);
or U2053 (N_2053,N_1215,N_1418);
nor U2054 (N_2054,N_1770,N_1074);
nor U2055 (N_2055,N_1419,N_1815);
or U2056 (N_2056,N_1572,N_1219);
nand U2057 (N_2057,N_1318,N_1683);
nor U2058 (N_2058,N_1626,N_1562);
nor U2059 (N_2059,N_1476,N_1073);
nand U2060 (N_2060,N_1001,N_1672);
nand U2061 (N_2061,N_1839,N_1695);
xor U2062 (N_2062,N_1556,N_1093);
nand U2063 (N_2063,N_1807,N_1564);
nor U2064 (N_2064,N_1868,N_1380);
and U2065 (N_2065,N_1929,N_1862);
and U2066 (N_2066,N_1714,N_1451);
or U2067 (N_2067,N_1139,N_1196);
or U2068 (N_2068,N_1151,N_1180);
or U2069 (N_2069,N_1211,N_1577);
nand U2070 (N_2070,N_1185,N_1503);
nand U2071 (N_2071,N_1197,N_1400);
xor U2072 (N_2072,N_1550,N_1809);
nand U2073 (N_2073,N_1509,N_1133);
nand U2074 (N_2074,N_1541,N_1762);
and U2075 (N_2075,N_1144,N_1131);
or U2076 (N_2076,N_1337,N_1242);
xnor U2077 (N_2077,N_1971,N_1842);
nor U2078 (N_2078,N_1125,N_1960);
and U2079 (N_2079,N_1557,N_1266);
or U2080 (N_2080,N_1838,N_1887);
and U2081 (N_2081,N_1555,N_1109);
xnor U2082 (N_2082,N_1755,N_1130);
or U2083 (N_2083,N_1386,N_1775);
nand U2084 (N_2084,N_1115,N_1692);
or U2085 (N_2085,N_1018,N_1590);
nor U2086 (N_2086,N_1798,N_1792);
nor U2087 (N_2087,N_1993,N_1333);
nor U2088 (N_2088,N_1384,N_1789);
and U2089 (N_2089,N_1712,N_1988);
nand U2090 (N_2090,N_1768,N_1358);
xnor U2091 (N_2091,N_1538,N_1462);
nand U2092 (N_2092,N_1439,N_1039);
and U2093 (N_2093,N_1817,N_1241);
and U2094 (N_2094,N_1758,N_1157);
nand U2095 (N_2095,N_1441,N_1812);
nand U2096 (N_2096,N_1199,N_1667);
or U2097 (N_2097,N_1020,N_1393);
xnor U2098 (N_2098,N_1081,N_1030);
nor U2099 (N_2099,N_1289,N_1641);
and U2100 (N_2100,N_1580,N_1134);
nor U2101 (N_2101,N_1421,N_1409);
or U2102 (N_2102,N_1951,N_1138);
nor U2103 (N_2103,N_1859,N_1387);
nand U2104 (N_2104,N_1369,N_1473);
and U2105 (N_2105,N_1394,N_1546);
and U2106 (N_2106,N_1610,N_1422);
nand U2107 (N_2107,N_1335,N_1644);
or U2108 (N_2108,N_1584,N_1547);
and U2109 (N_2109,N_1846,N_1956);
or U2110 (N_2110,N_1399,N_1571);
nand U2111 (N_2111,N_1217,N_1293);
nand U2112 (N_2112,N_1277,N_1721);
and U2113 (N_2113,N_1620,N_1527);
nor U2114 (N_2114,N_1200,N_1188);
nand U2115 (N_2115,N_1288,N_1502);
nor U2116 (N_2116,N_1381,N_1107);
or U2117 (N_2117,N_1404,N_1388);
and U2118 (N_2118,N_1583,N_1805);
xnor U2119 (N_2119,N_1326,N_1189);
nand U2120 (N_2120,N_1598,N_1636);
and U2121 (N_2121,N_1592,N_1111);
or U2122 (N_2122,N_1006,N_1905);
and U2123 (N_2123,N_1685,N_1653);
and U2124 (N_2124,N_1468,N_1693);
or U2125 (N_2125,N_1720,N_1938);
nand U2126 (N_2126,N_1656,N_1634);
and U2127 (N_2127,N_1440,N_1715);
xnor U2128 (N_2128,N_1351,N_1825);
and U2129 (N_2129,N_1983,N_1706);
xor U2130 (N_2130,N_1984,N_1478);
and U2131 (N_2131,N_1648,N_1649);
xnor U2132 (N_2132,N_1514,N_1009);
xnor U2133 (N_2133,N_1046,N_1961);
or U2134 (N_2134,N_1246,N_1348);
and U2135 (N_2135,N_1047,N_1629);
and U2136 (N_2136,N_1132,N_1284);
nand U2137 (N_2137,N_1646,N_1797);
nand U2138 (N_2138,N_1013,N_1777);
xnor U2139 (N_2139,N_1704,N_1048);
nand U2140 (N_2140,N_1885,N_1488);
and U2141 (N_2141,N_1467,N_1233);
and U2142 (N_2142,N_1298,N_1517);
and U2143 (N_2143,N_1513,N_1062);
or U2144 (N_2144,N_1883,N_1820);
or U2145 (N_2145,N_1137,N_1935);
nand U2146 (N_2146,N_1250,N_1494);
nand U2147 (N_2147,N_1286,N_1510);
nand U2148 (N_2148,N_1244,N_1785);
and U2149 (N_2149,N_1521,N_1818);
nor U2150 (N_2150,N_1428,N_1623);
and U2151 (N_2151,N_1536,N_1341);
nand U2152 (N_2152,N_1829,N_1896);
or U2153 (N_2153,N_1186,N_1444);
nand U2154 (N_2154,N_1204,N_1819);
and U2155 (N_2155,N_1776,N_1345);
or U2156 (N_2156,N_1314,N_1084);
nand U2157 (N_2157,N_1085,N_1912);
nor U2158 (N_2158,N_1296,N_1102);
nor U2159 (N_2159,N_1560,N_1779);
and U2160 (N_2160,N_1772,N_1851);
and U2161 (N_2161,N_1764,N_1460);
and U2162 (N_2162,N_1978,N_1259);
and U2163 (N_2163,N_1903,N_1945);
nand U2164 (N_2164,N_1670,N_1178);
nand U2165 (N_2165,N_1681,N_1121);
xnor U2166 (N_2166,N_1976,N_1315);
xnor U2167 (N_2167,N_1140,N_1276);
or U2168 (N_2168,N_1203,N_1780);
xnor U2169 (N_2169,N_1379,N_1576);
nor U2170 (N_2170,N_1803,N_1982);
xnor U2171 (N_2171,N_1311,N_1750);
xor U2172 (N_2172,N_1810,N_1587);
nor U2173 (N_2173,N_1928,N_1830);
xnor U2174 (N_2174,N_1396,N_1145);
or U2175 (N_2175,N_1173,N_1553);
or U2176 (N_2176,N_1034,N_1049);
xnor U2177 (N_2177,N_1941,N_1114);
nand U2178 (N_2178,N_1258,N_1700);
and U2179 (N_2179,N_1937,N_1346);
nand U2180 (N_2180,N_1906,N_1821);
xnor U2181 (N_2181,N_1012,N_1058);
xnor U2182 (N_2182,N_1913,N_1535);
and U2183 (N_2183,N_1352,N_1312);
and U2184 (N_2184,N_1454,N_1035);
and U2185 (N_2185,N_1356,N_1927);
xor U2186 (N_2186,N_1471,N_1365);
xnor U2187 (N_2187,N_1302,N_1474);
or U2188 (N_2188,N_1195,N_1465);
nor U2189 (N_2189,N_1375,N_1223);
and U2190 (N_2190,N_1449,N_1852);
nor U2191 (N_2191,N_1989,N_1459);
nor U2192 (N_2192,N_1411,N_1806);
or U2193 (N_2193,N_1783,N_1482);
or U2194 (N_2194,N_1342,N_1528);
or U2195 (N_2195,N_1979,N_1257);
or U2196 (N_2196,N_1870,N_1740);
xnor U2197 (N_2197,N_1736,N_1042);
nor U2198 (N_2198,N_1060,N_1495);
and U2199 (N_2199,N_1781,N_1210);
and U2200 (N_2200,N_1249,N_1726);
nand U2201 (N_2201,N_1811,N_1002);
or U2202 (N_2202,N_1848,N_1824);
and U2203 (N_2203,N_1498,N_1751);
nand U2204 (N_2204,N_1889,N_1642);
or U2205 (N_2205,N_1143,N_1999);
xor U2206 (N_2206,N_1403,N_1243);
nand U2207 (N_2207,N_1307,N_1029);
or U2208 (N_2208,N_1168,N_1000);
nand U2209 (N_2209,N_1586,N_1694);
nor U2210 (N_2210,N_1432,N_1456);
nor U2211 (N_2211,N_1187,N_1605);
nand U2212 (N_2212,N_1110,N_1174);
nor U2213 (N_2213,N_1050,N_1028);
or U2214 (N_2214,N_1319,N_1317);
nand U2215 (N_2215,N_1633,N_1118);
and U2216 (N_2216,N_1866,N_1281);
and U2217 (N_2217,N_1659,N_1585);
xor U2218 (N_2218,N_1164,N_1155);
nor U2219 (N_2219,N_1382,N_1893);
nand U2220 (N_2220,N_1602,N_1136);
nor U2221 (N_2221,N_1414,N_1665);
xor U2222 (N_2222,N_1888,N_1884);
xor U2223 (N_2223,N_1627,N_1652);
nand U2224 (N_2224,N_1321,N_1662);
nor U2225 (N_2225,N_1767,N_1574);
nand U2226 (N_2226,N_1205,N_1603);
xnor U2227 (N_2227,N_1872,N_1362);
nor U2228 (N_2228,N_1183,N_1900);
nor U2229 (N_2229,N_1997,N_1198);
nor U2230 (N_2230,N_1835,N_1032);
or U2231 (N_2231,N_1702,N_1182);
or U2232 (N_2232,N_1455,N_1925);
nand U2233 (N_2233,N_1711,N_1918);
xnor U2234 (N_2234,N_1899,N_1531);
xnor U2235 (N_2235,N_1881,N_1267);
or U2236 (N_2236,N_1447,N_1841);
or U2237 (N_2237,N_1766,N_1354);
nor U2238 (N_2238,N_1606,N_1773);
xnor U2239 (N_2239,N_1823,N_1631);
and U2240 (N_2240,N_1294,N_1607);
nand U2241 (N_2241,N_1745,N_1533);
xor U2242 (N_2242,N_1443,N_1496);
and U2243 (N_2243,N_1735,N_1691);
xor U2244 (N_2244,N_1072,N_1774);
nor U2245 (N_2245,N_1932,N_1882);
nor U2246 (N_2246,N_1742,N_1630);
or U2247 (N_2247,N_1596,N_1914);
or U2248 (N_2248,N_1235,N_1096);
nor U2249 (N_2249,N_1207,N_1328);
and U2250 (N_2250,N_1778,N_1657);
xor U2251 (N_2251,N_1206,N_1367);
or U2252 (N_2252,N_1664,N_1026);
and U2253 (N_2253,N_1962,N_1845);
nor U2254 (N_2254,N_1007,N_1901);
xor U2255 (N_2255,N_1324,N_1690);
or U2256 (N_2256,N_1895,N_1150);
and U2257 (N_2257,N_1113,N_1705);
nor U2258 (N_2258,N_1784,N_1808);
nand U2259 (N_2259,N_1724,N_1942);
nor U2260 (N_2260,N_1725,N_1063);
xor U2261 (N_2261,N_1522,N_1024);
xor U2262 (N_2262,N_1990,N_1669);
or U2263 (N_2263,N_1632,N_1415);
or U2264 (N_2264,N_1996,N_1285);
and U2265 (N_2265,N_1304,N_1480);
or U2266 (N_2266,N_1038,N_1208);
xnor U2267 (N_2267,N_1051,N_1160);
or U2268 (N_2268,N_1619,N_1265);
nand U2269 (N_2269,N_1067,N_1660);
nor U2270 (N_2270,N_1340,N_1616);
nand U2271 (N_2271,N_1332,N_1213);
nor U2272 (N_2272,N_1301,N_1466);
and U2273 (N_2273,N_1065,N_1383);
xnor U2274 (N_2274,N_1628,N_1907);
nor U2275 (N_2275,N_1202,N_1497);
and U2276 (N_2276,N_1782,N_1218);
and U2277 (N_2277,N_1108,N_1920);
and U2278 (N_2278,N_1994,N_1552);
or U2279 (N_2279,N_1417,N_1299);
nand U2280 (N_2280,N_1303,N_1822);
and U2281 (N_2281,N_1300,N_1248);
and U2282 (N_2282,N_1036,N_1308);
nor U2283 (N_2283,N_1663,N_1904);
nand U2284 (N_2284,N_1520,N_1469);
and U2285 (N_2285,N_1696,N_1194);
nand U2286 (N_2286,N_1279,N_1043);
nand U2287 (N_2287,N_1916,N_1647);
or U2288 (N_2288,N_1879,N_1359);
and U2289 (N_2289,N_1076,N_1238);
nand U2290 (N_2290,N_1408,N_1931);
nor U2291 (N_2291,N_1435,N_1947);
and U2292 (N_2292,N_1098,N_1974);
nor U2293 (N_2293,N_1505,N_1668);
nor U2294 (N_2294,N_1212,N_1955);
nor U2295 (N_2295,N_1253,N_1347);
xnor U2296 (N_2296,N_1019,N_1475);
or U2297 (N_2297,N_1917,N_1120);
and U2298 (N_2298,N_1395,N_1273);
xnor U2299 (N_2299,N_1330,N_1457);
nand U2300 (N_2300,N_1325,N_1753);
nor U2301 (N_2301,N_1998,N_1554);
or U2302 (N_2302,N_1529,N_1054);
or U2303 (N_2303,N_1270,N_1260);
xnor U2304 (N_2304,N_1658,N_1123);
or U2305 (N_2305,N_1853,N_1343);
nand U2306 (N_2306,N_1149,N_1334);
or U2307 (N_2307,N_1413,N_1017);
nor U2308 (N_2308,N_1184,N_1245);
xor U2309 (N_2309,N_1492,N_1431);
xnor U2310 (N_2310,N_1117,N_1426);
or U2311 (N_2311,N_1703,N_1816);
nor U2312 (N_2312,N_1970,N_1424);
xor U2313 (N_2313,N_1066,N_1678);
or U2314 (N_2314,N_1331,N_1410);
nor U2315 (N_2315,N_1739,N_1094);
or U2316 (N_2316,N_1310,N_1374);
nor U2317 (N_2317,N_1673,N_1055);
xor U2318 (N_2318,N_1687,N_1524);
xnor U2319 (N_2319,N_1350,N_1701);
xor U2320 (N_2320,N_1487,N_1171);
xnor U2321 (N_2321,N_1570,N_1237);
xnor U2322 (N_2322,N_1129,N_1161);
or U2323 (N_2323,N_1370,N_1902);
and U2324 (N_2324,N_1221,N_1041);
or U2325 (N_2325,N_1122,N_1654);
and U2326 (N_2326,N_1719,N_1729);
nand U2327 (N_2327,N_1716,N_1617);
or U2328 (N_2328,N_1831,N_1061);
or U2329 (N_2329,N_1448,N_1392);
nand U2330 (N_2330,N_1597,N_1291);
nor U2331 (N_2331,N_1939,N_1867);
or U2332 (N_2332,N_1092,N_1127);
or U2333 (N_2333,N_1834,N_1637);
or U2334 (N_2334,N_1275,N_1290);
nand U2335 (N_2335,N_1190,N_1481);
or U2336 (N_2336,N_1869,N_1875);
or U2337 (N_2337,N_1463,N_1599);
and U2338 (N_2338,N_1280,N_1915);
xor U2339 (N_2339,N_1105,N_1589);
xor U2340 (N_2340,N_1837,N_1373);
or U2341 (N_2341,N_1949,N_1873);
and U2342 (N_2342,N_1437,N_1090);
nor U2343 (N_2343,N_1306,N_1760);
and U2344 (N_2344,N_1389,N_1316);
nor U2345 (N_2345,N_1709,N_1433);
nor U2346 (N_2346,N_1697,N_1957);
nor U2347 (N_2347,N_1177,N_1618);
nor U2348 (N_2348,N_1025,N_1858);
nand U2349 (N_2349,N_1559,N_1262);
nand U2350 (N_2350,N_1165,N_1479);
xor U2351 (N_2351,N_1795,N_1794);
nand U2352 (N_2352,N_1401,N_1578);
nor U2353 (N_2353,N_1357,N_1142);
or U2354 (N_2354,N_1470,N_1731);
nand U2355 (N_2355,N_1166,N_1124);
xor U2356 (N_2356,N_1878,N_1453);
xnor U2357 (N_2357,N_1622,N_1682);
xnor U2358 (N_2358,N_1608,N_1813);
and U2359 (N_2359,N_1689,N_1786);
xnor U2360 (N_2360,N_1486,N_1075);
or U2361 (N_2361,N_1748,N_1926);
nor U2362 (N_2362,N_1068,N_1082);
nand U2363 (N_2363,N_1087,N_1506);
nor U2364 (N_2364,N_1052,N_1385);
nor U2365 (N_2365,N_1563,N_1534);
nand U2366 (N_2366,N_1193,N_1936);
and U2367 (N_2367,N_1849,N_1045);
nor U2368 (N_2368,N_1101,N_1565);
xor U2369 (N_2369,N_1398,N_1635);
or U2370 (N_2370,N_1741,N_1793);
nor U2371 (N_2371,N_1801,N_1214);
nor U2372 (N_2372,N_1843,N_1890);
nor U2373 (N_2373,N_1429,N_1056);
nand U2374 (N_2374,N_1349,N_1484);
and U2375 (N_2375,N_1943,N_1015);
or U2376 (N_2376,N_1676,N_1033);
xnor U2377 (N_2377,N_1226,N_1991);
and U2378 (N_2378,N_1167,N_1737);
nor U2379 (N_2379,N_1684,N_1909);
nand U2380 (N_2380,N_1796,N_1880);
xnor U2381 (N_2381,N_1944,N_1376);
nand U2382 (N_2382,N_1146,N_1738);
xnor U2383 (N_2383,N_1625,N_1490);
and U2384 (N_2384,N_1655,N_1847);
or U2385 (N_2385,N_1247,N_1344);
nor U2386 (N_2386,N_1295,N_1254);
nand U2387 (N_2387,N_1727,N_1162);
xor U2388 (N_2388,N_1464,N_1504);
nor U2389 (N_2389,N_1106,N_1763);
nor U2390 (N_2390,N_1256,N_1169);
and U2391 (N_2391,N_1959,N_1922);
nand U2392 (N_2392,N_1368,N_1840);
nor U2393 (N_2393,N_1886,N_1220);
and U2394 (N_2394,N_1671,N_1397);
or U2395 (N_2395,N_1158,N_1119);
and U2396 (N_2396,N_1446,N_1545);
nor U2397 (N_2397,N_1442,N_1021);
nand U2398 (N_2398,N_1091,N_1549);
or U2399 (N_2399,N_1877,N_1089);
nor U2400 (N_2400,N_1327,N_1799);
and U2401 (N_2401,N_1568,N_1854);
or U2402 (N_2402,N_1163,N_1430);
xor U2403 (N_2403,N_1434,N_1975);
nand U2404 (N_2404,N_1305,N_1566);
nor U2405 (N_2405,N_1170,N_1175);
and U2406 (N_2406,N_1010,N_1027);
xnor U2407 (N_2407,N_1176,N_1236);
and U2408 (N_2408,N_1261,N_1591);
and U2409 (N_2409,N_1438,N_1594);
xor U2410 (N_2410,N_1037,N_1746);
or U2411 (N_2411,N_1406,N_1558);
and U2412 (N_2412,N_1707,N_1601);
nand U2413 (N_2413,N_1897,N_1181);
nand U2414 (N_2414,N_1227,N_1952);
nand U2415 (N_2415,N_1500,N_1516);
xnor U2416 (N_2416,N_1057,N_1154);
or U2417 (N_2417,N_1679,N_1372);
and U2418 (N_2418,N_1680,N_1540);
xor U2419 (N_2419,N_1086,N_1968);
or U2420 (N_2420,N_1833,N_1407);
or U2421 (N_2421,N_1844,N_1624);
or U2422 (N_2422,N_1966,N_1542);
xor U2423 (N_2423,N_1079,N_1855);
nand U2424 (N_2424,N_1378,N_1609);
nor U2425 (N_2425,N_1532,N_1283);
and U2426 (N_2426,N_1800,N_1573);
xor U2427 (N_2427,N_1530,N_1507);
and U2428 (N_2428,N_1526,N_1069);
nand U2429 (N_2429,N_1864,N_1525);
nor U2430 (N_2430,N_1539,N_1228);
xor U2431 (N_2431,N_1921,N_1234);
nand U2432 (N_2432,N_1717,N_1489);
xnor U2433 (N_2433,N_1948,N_1364);
nand U2434 (N_2434,N_1071,N_1452);
nor U2435 (N_2435,N_1450,N_1972);
nor U2436 (N_2436,N_1095,N_1003);
nor U2437 (N_2437,N_1423,N_1405);
or U2438 (N_2438,N_1638,N_1569);
nand U2439 (N_2439,N_1360,N_1581);
nor U2440 (N_2440,N_1077,N_1209);
or U2441 (N_2441,N_1765,N_1802);
xnor U2442 (N_2442,N_1579,N_1933);
nor U2443 (N_2443,N_1519,N_1355);
and U2444 (N_2444,N_1420,N_1491);
nand U2445 (N_2445,N_1172,N_1445);
nor U2446 (N_2446,N_1969,N_1860);
xnor U2447 (N_2447,N_1752,N_1910);
and U2448 (N_2448,N_1271,N_1005);
or U2449 (N_2449,N_1674,N_1366);
or U2450 (N_2450,N_1192,N_1083);
xnor U2451 (N_2451,N_1561,N_1518);
nor U2452 (N_2452,N_1600,N_1240);
and U2453 (N_2453,N_1651,N_1954);
nand U2454 (N_2454,N_1501,N_1980);
nor U2455 (N_2455,N_1582,N_1264);
or U2456 (N_2456,N_1031,N_1053);
nand U2457 (N_2457,N_1361,N_1744);
or U2458 (N_2458,N_1614,N_1011);
and U2459 (N_2459,N_1064,N_1458);
nor U2460 (N_2460,N_1863,N_1427);
or U2461 (N_2461,N_1791,N_1732);
and U2462 (N_2462,N_1593,N_1757);
nand U2463 (N_2463,N_1216,N_1892);
nand U2464 (N_2464,N_1363,N_1836);
or U2465 (N_2465,N_1044,N_1639);
or U2466 (N_2466,N_1722,N_1771);
or U2467 (N_2467,N_1643,N_1977);
or U2468 (N_2468,N_1650,N_1930);
nand U2469 (N_2469,N_1436,N_1148);
nor U2470 (N_2470,N_1856,N_1268);
nand U2471 (N_2471,N_1992,N_1287);
and U2472 (N_2472,N_1640,N_1688);
xor U2473 (N_2473,N_1828,N_1416);
nand U2474 (N_2474,N_1511,N_1251);
nor U2475 (N_2475,N_1179,N_1508);
and U2476 (N_2476,N_1973,N_1255);
or U2477 (N_2477,N_1790,N_1891);
or U2478 (N_2478,N_1272,N_1543);
nand U2479 (N_2479,N_1551,N_1908);
and U2480 (N_2480,N_1874,N_1544);
xnor U2481 (N_2481,N_1339,N_1515);
or U2482 (N_2482,N_1222,N_1788);
or U2483 (N_2483,N_1940,N_1756);
xor U2484 (N_2484,N_1827,N_1313);
nor U2485 (N_2485,N_1070,N_1128);
xor U2486 (N_2486,N_1099,N_1292);
and U2487 (N_2487,N_1147,N_1022);
and U2488 (N_2488,N_1985,N_1263);
nor U2489 (N_2489,N_1320,N_1761);
or U2490 (N_2490,N_1965,N_1412);
xnor U2491 (N_2491,N_1274,N_1759);
and U2492 (N_2492,N_1967,N_1103);
nor U2493 (N_2493,N_1040,N_1485);
xor U2494 (N_2494,N_1661,N_1612);
and U2495 (N_2495,N_1804,N_1297);
nor U2496 (N_2496,N_1336,N_1963);
or U2497 (N_2497,N_1425,N_1986);
nor U2498 (N_2498,N_1787,N_1088);
xor U2499 (N_2499,N_1604,N_1677);
nor U2500 (N_2500,N_1860,N_1957);
xnor U2501 (N_2501,N_1888,N_1785);
and U2502 (N_2502,N_1655,N_1161);
xor U2503 (N_2503,N_1838,N_1113);
xor U2504 (N_2504,N_1183,N_1023);
and U2505 (N_2505,N_1932,N_1030);
xor U2506 (N_2506,N_1213,N_1551);
xnor U2507 (N_2507,N_1622,N_1673);
and U2508 (N_2508,N_1769,N_1947);
xor U2509 (N_2509,N_1774,N_1706);
nand U2510 (N_2510,N_1256,N_1195);
xnor U2511 (N_2511,N_1648,N_1071);
nand U2512 (N_2512,N_1405,N_1847);
xnor U2513 (N_2513,N_1788,N_1588);
and U2514 (N_2514,N_1275,N_1955);
nor U2515 (N_2515,N_1666,N_1664);
or U2516 (N_2516,N_1525,N_1931);
nand U2517 (N_2517,N_1869,N_1429);
nand U2518 (N_2518,N_1624,N_1672);
or U2519 (N_2519,N_1311,N_1842);
nor U2520 (N_2520,N_1887,N_1700);
xnor U2521 (N_2521,N_1197,N_1219);
or U2522 (N_2522,N_1800,N_1982);
and U2523 (N_2523,N_1717,N_1243);
nand U2524 (N_2524,N_1077,N_1449);
and U2525 (N_2525,N_1272,N_1758);
and U2526 (N_2526,N_1529,N_1520);
and U2527 (N_2527,N_1113,N_1575);
or U2528 (N_2528,N_1950,N_1491);
nand U2529 (N_2529,N_1926,N_1096);
nand U2530 (N_2530,N_1398,N_1508);
or U2531 (N_2531,N_1925,N_1895);
nor U2532 (N_2532,N_1862,N_1467);
nor U2533 (N_2533,N_1475,N_1288);
nor U2534 (N_2534,N_1210,N_1067);
nor U2535 (N_2535,N_1579,N_1483);
or U2536 (N_2536,N_1437,N_1929);
nand U2537 (N_2537,N_1639,N_1892);
xnor U2538 (N_2538,N_1283,N_1952);
and U2539 (N_2539,N_1380,N_1105);
or U2540 (N_2540,N_1367,N_1691);
xor U2541 (N_2541,N_1288,N_1108);
nand U2542 (N_2542,N_1213,N_1129);
nor U2543 (N_2543,N_1402,N_1067);
and U2544 (N_2544,N_1141,N_1870);
or U2545 (N_2545,N_1434,N_1036);
xnor U2546 (N_2546,N_1856,N_1788);
nor U2547 (N_2547,N_1761,N_1729);
xor U2548 (N_2548,N_1729,N_1483);
nor U2549 (N_2549,N_1772,N_1599);
nand U2550 (N_2550,N_1031,N_1303);
and U2551 (N_2551,N_1715,N_1231);
nor U2552 (N_2552,N_1516,N_1225);
or U2553 (N_2553,N_1411,N_1119);
nand U2554 (N_2554,N_1625,N_1463);
nor U2555 (N_2555,N_1741,N_1138);
nand U2556 (N_2556,N_1593,N_1051);
xor U2557 (N_2557,N_1714,N_1622);
and U2558 (N_2558,N_1248,N_1526);
or U2559 (N_2559,N_1373,N_1732);
nor U2560 (N_2560,N_1911,N_1103);
nand U2561 (N_2561,N_1558,N_1168);
nor U2562 (N_2562,N_1908,N_1575);
or U2563 (N_2563,N_1538,N_1056);
xnor U2564 (N_2564,N_1299,N_1611);
and U2565 (N_2565,N_1776,N_1937);
nand U2566 (N_2566,N_1580,N_1269);
or U2567 (N_2567,N_1225,N_1321);
xor U2568 (N_2568,N_1337,N_1631);
nand U2569 (N_2569,N_1215,N_1466);
xnor U2570 (N_2570,N_1619,N_1202);
nand U2571 (N_2571,N_1383,N_1157);
and U2572 (N_2572,N_1896,N_1161);
and U2573 (N_2573,N_1348,N_1789);
nand U2574 (N_2574,N_1819,N_1222);
or U2575 (N_2575,N_1940,N_1154);
and U2576 (N_2576,N_1217,N_1572);
or U2577 (N_2577,N_1938,N_1173);
nand U2578 (N_2578,N_1432,N_1649);
or U2579 (N_2579,N_1314,N_1829);
xor U2580 (N_2580,N_1953,N_1502);
and U2581 (N_2581,N_1709,N_1837);
nand U2582 (N_2582,N_1708,N_1190);
or U2583 (N_2583,N_1727,N_1369);
nor U2584 (N_2584,N_1086,N_1882);
xnor U2585 (N_2585,N_1235,N_1300);
nor U2586 (N_2586,N_1367,N_1304);
xnor U2587 (N_2587,N_1952,N_1316);
nor U2588 (N_2588,N_1758,N_1436);
and U2589 (N_2589,N_1464,N_1067);
xor U2590 (N_2590,N_1596,N_1915);
nand U2591 (N_2591,N_1275,N_1370);
and U2592 (N_2592,N_1553,N_1134);
or U2593 (N_2593,N_1572,N_1419);
nor U2594 (N_2594,N_1784,N_1463);
nand U2595 (N_2595,N_1028,N_1269);
or U2596 (N_2596,N_1083,N_1583);
and U2597 (N_2597,N_1521,N_1925);
or U2598 (N_2598,N_1894,N_1901);
nor U2599 (N_2599,N_1605,N_1277);
or U2600 (N_2600,N_1231,N_1632);
xor U2601 (N_2601,N_1185,N_1874);
nand U2602 (N_2602,N_1618,N_1026);
nor U2603 (N_2603,N_1089,N_1401);
nand U2604 (N_2604,N_1578,N_1650);
nor U2605 (N_2605,N_1496,N_1830);
nand U2606 (N_2606,N_1686,N_1780);
or U2607 (N_2607,N_1500,N_1102);
xor U2608 (N_2608,N_1097,N_1254);
nand U2609 (N_2609,N_1212,N_1751);
nand U2610 (N_2610,N_1361,N_1460);
and U2611 (N_2611,N_1553,N_1897);
nor U2612 (N_2612,N_1659,N_1394);
and U2613 (N_2613,N_1705,N_1137);
nor U2614 (N_2614,N_1691,N_1124);
nand U2615 (N_2615,N_1939,N_1139);
and U2616 (N_2616,N_1659,N_1460);
xor U2617 (N_2617,N_1138,N_1468);
xor U2618 (N_2618,N_1870,N_1588);
nand U2619 (N_2619,N_1758,N_1082);
and U2620 (N_2620,N_1000,N_1679);
xor U2621 (N_2621,N_1419,N_1456);
nor U2622 (N_2622,N_1903,N_1267);
and U2623 (N_2623,N_1433,N_1423);
xnor U2624 (N_2624,N_1316,N_1640);
nand U2625 (N_2625,N_1422,N_1910);
nand U2626 (N_2626,N_1025,N_1087);
nor U2627 (N_2627,N_1458,N_1115);
or U2628 (N_2628,N_1277,N_1896);
xor U2629 (N_2629,N_1253,N_1450);
xnor U2630 (N_2630,N_1117,N_1072);
xor U2631 (N_2631,N_1802,N_1840);
or U2632 (N_2632,N_1727,N_1959);
nor U2633 (N_2633,N_1845,N_1439);
nand U2634 (N_2634,N_1729,N_1070);
nand U2635 (N_2635,N_1735,N_1979);
or U2636 (N_2636,N_1093,N_1340);
and U2637 (N_2637,N_1970,N_1326);
or U2638 (N_2638,N_1960,N_1326);
nor U2639 (N_2639,N_1412,N_1409);
nor U2640 (N_2640,N_1879,N_1400);
and U2641 (N_2641,N_1398,N_1089);
xnor U2642 (N_2642,N_1964,N_1907);
xor U2643 (N_2643,N_1659,N_1408);
or U2644 (N_2644,N_1332,N_1492);
and U2645 (N_2645,N_1824,N_1504);
and U2646 (N_2646,N_1413,N_1477);
xor U2647 (N_2647,N_1934,N_1096);
and U2648 (N_2648,N_1877,N_1487);
nor U2649 (N_2649,N_1743,N_1965);
nor U2650 (N_2650,N_1131,N_1870);
and U2651 (N_2651,N_1917,N_1405);
nand U2652 (N_2652,N_1958,N_1952);
nor U2653 (N_2653,N_1350,N_1998);
xor U2654 (N_2654,N_1317,N_1662);
nand U2655 (N_2655,N_1231,N_1758);
xor U2656 (N_2656,N_1899,N_1485);
xor U2657 (N_2657,N_1035,N_1414);
xor U2658 (N_2658,N_1313,N_1472);
and U2659 (N_2659,N_1604,N_1135);
and U2660 (N_2660,N_1649,N_1347);
nor U2661 (N_2661,N_1876,N_1819);
nor U2662 (N_2662,N_1583,N_1319);
or U2663 (N_2663,N_1197,N_1435);
nor U2664 (N_2664,N_1503,N_1793);
and U2665 (N_2665,N_1043,N_1098);
and U2666 (N_2666,N_1844,N_1001);
or U2667 (N_2667,N_1417,N_1282);
nand U2668 (N_2668,N_1234,N_1590);
or U2669 (N_2669,N_1870,N_1204);
nor U2670 (N_2670,N_1574,N_1421);
xor U2671 (N_2671,N_1245,N_1437);
nand U2672 (N_2672,N_1895,N_1227);
nor U2673 (N_2673,N_1535,N_1615);
or U2674 (N_2674,N_1810,N_1298);
and U2675 (N_2675,N_1449,N_1952);
or U2676 (N_2676,N_1657,N_1078);
nand U2677 (N_2677,N_1013,N_1836);
or U2678 (N_2678,N_1420,N_1679);
or U2679 (N_2679,N_1896,N_1867);
xor U2680 (N_2680,N_1521,N_1643);
and U2681 (N_2681,N_1312,N_1228);
or U2682 (N_2682,N_1752,N_1722);
xnor U2683 (N_2683,N_1942,N_1591);
nor U2684 (N_2684,N_1271,N_1768);
xnor U2685 (N_2685,N_1801,N_1908);
nand U2686 (N_2686,N_1484,N_1825);
and U2687 (N_2687,N_1267,N_1658);
nor U2688 (N_2688,N_1993,N_1717);
nor U2689 (N_2689,N_1386,N_1837);
nor U2690 (N_2690,N_1393,N_1070);
or U2691 (N_2691,N_1790,N_1009);
xor U2692 (N_2692,N_1430,N_1289);
xor U2693 (N_2693,N_1205,N_1060);
or U2694 (N_2694,N_1965,N_1780);
or U2695 (N_2695,N_1340,N_1815);
xnor U2696 (N_2696,N_1648,N_1807);
nand U2697 (N_2697,N_1458,N_1688);
and U2698 (N_2698,N_1187,N_1019);
nor U2699 (N_2699,N_1514,N_1546);
or U2700 (N_2700,N_1232,N_1056);
or U2701 (N_2701,N_1615,N_1447);
nor U2702 (N_2702,N_1458,N_1285);
xor U2703 (N_2703,N_1168,N_1642);
or U2704 (N_2704,N_1682,N_1370);
nor U2705 (N_2705,N_1737,N_1929);
nand U2706 (N_2706,N_1035,N_1648);
or U2707 (N_2707,N_1708,N_1509);
and U2708 (N_2708,N_1740,N_1441);
and U2709 (N_2709,N_1018,N_1389);
nor U2710 (N_2710,N_1316,N_1152);
nor U2711 (N_2711,N_1713,N_1755);
nand U2712 (N_2712,N_1927,N_1163);
nand U2713 (N_2713,N_1274,N_1745);
xnor U2714 (N_2714,N_1491,N_1377);
nand U2715 (N_2715,N_1075,N_1641);
nor U2716 (N_2716,N_1788,N_1757);
xnor U2717 (N_2717,N_1480,N_1074);
nand U2718 (N_2718,N_1998,N_1414);
nand U2719 (N_2719,N_1346,N_1182);
and U2720 (N_2720,N_1203,N_1746);
or U2721 (N_2721,N_1972,N_1504);
or U2722 (N_2722,N_1072,N_1335);
xor U2723 (N_2723,N_1433,N_1107);
xor U2724 (N_2724,N_1137,N_1275);
xor U2725 (N_2725,N_1265,N_1260);
and U2726 (N_2726,N_1521,N_1321);
nor U2727 (N_2727,N_1521,N_1638);
or U2728 (N_2728,N_1587,N_1474);
nand U2729 (N_2729,N_1263,N_1485);
and U2730 (N_2730,N_1647,N_1912);
and U2731 (N_2731,N_1037,N_1381);
nor U2732 (N_2732,N_1940,N_1348);
nand U2733 (N_2733,N_1456,N_1006);
nor U2734 (N_2734,N_1351,N_1570);
and U2735 (N_2735,N_1892,N_1052);
or U2736 (N_2736,N_1609,N_1642);
and U2737 (N_2737,N_1199,N_1042);
nand U2738 (N_2738,N_1224,N_1341);
and U2739 (N_2739,N_1865,N_1118);
and U2740 (N_2740,N_1544,N_1897);
xor U2741 (N_2741,N_1471,N_1160);
and U2742 (N_2742,N_1541,N_1969);
nor U2743 (N_2743,N_1149,N_1225);
xnor U2744 (N_2744,N_1063,N_1580);
xor U2745 (N_2745,N_1843,N_1084);
or U2746 (N_2746,N_1855,N_1895);
xor U2747 (N_2747,N_1762,N_1188);
or U2748 (N_2748,N_1216,N_1470);
or U2749 (N_2749,N_1946,N_1087);
nor U2750 (N_2750,N_1868,N_1639);
or U2751 (N_2751,N_1933,N_1972);
and U2752 (N_2752,N_1283,N_1169);
or U2753 (N_2753,N_1897,N_1101);
xnor U2754 (N_2754,N_1674,N_1263);
nor U2755 (N_2755,N_1088,N_1045);
xor U2756 (N_2756,N_1995,N_1077);
nand U2757 (N_2757,N_1810,N_1921);
xnor U2758 (N_2758,N_1544,N_1361);
or U2759 (N_2759,N_1055,N_1920);
or U2760 (N_2760,N_1674,N_1754);
nor U2761 (N_2761,N_1050,N_1970);
xor U2762 (N_2762,N_1232,N_1693);
xor U2763 (N_2763,N_1593,N_1477);
xor U2764 (N_2764,N_1169,N_1719);
or U2765 (N_2765,N_1610,N_1829);
nor U2766 (N_2766,N_1522,N_1189);
nor U2767 (N_2767,N_1457,N_1687);
nand U2768 (N_2768,N_1116,N_1111);
and U2769 (N_2769,N_1207,N_1725);
or U2770 (N_2770,N_1444,N_1593);
nor U2771 (N_2771,N_1124,N_1641);
nand U2772 (N_2772,N_1070,N_1637);
xnor U2773 (N_2773,N_1682,N_1528);
nor U2774 (N_2774,N_1771,N_1378);
or U2775 (N_2775,N_1243,N_1477);
or U2776 (N_2776,N_1721,N_1357);
nor U2777 (N_2777,N_1781,N_1864);
nor U2778 (N_2778,N_1480,N_1906);
nand U2779 (N_2779,N_1171,N_1508);
and U2780 (N_2780,N_1426,N_1947);
or U2781 (N_2781,N_1069,N_1638);
or U2782 (N_2782,N_1344,N_1546);
or U2783 (N_2783,N_1994,N_1330);
xor U2784 (N_2784,N_1493,N_1841);
nand U2785 (N_2785,N_1257,N_1661);
nor U2786 (N_2786,N_1386,N_1124);
and U2787 (N_2787,N_1608,N_1086);
or U2788 (N_2788,N_1089,N_1604);
xnor U2789 (N_2789,N_1859,N_1901);
and U2790 (N_2790,N_1168,N_1540);
nand U2791 (N_2791,N_1952,N_1713);
xor U2792 (N_2792,N_1433,N_1447);
nor U2793 (N_2793,N_1287,N_1787);
and U2794 (N_2794,N_1355,N_1695);
xor U2795 (N_2795,N_1923,N_1910);
nand U2796 (N_2796,N_1218,N_1631);
or U2797 (N_2797,N_1512,N_1219);
nor U2798 (N_2798,N_1334,N_1067);
nor U2799 (N_2799,N_1268,N_1496);
xor U2800 (N_2800,N_1235,N_1983);
or U2801 (N_2801,N_1676,N_1797);
nor U2802 (N_2802,N_1115,N_1196);
xnor U2803 (N_2803,N_1319,N_1525);
nand U2804 (N_2804,N_1850,N_1267);
and U2805 (N_2805,N_1646,N_1786);
xnor U2806 (N_2806,N_1151,N_1438);
and U2807 (N_2807,N_1919,N_1385);
and U2808 (N_2808,N_1994,N_1583);
nor U2809 (N_2809,N_1189,N_1011);
and U2810 (N_2810,N_1106,N_1241);
and U2811 (N_2811,N_1439,N_1866);
xnor U2812 (N_2812,N_1480,N_1120);
nor U2813 (N_2813,N_1379,N_1381);
or U2814 (N_2814,N_1281,N_1992);
and U2815 (N_2815,N_1040,N_1845);
and U2816 (N_2816,N_1175,N_1764);
xnor U2817 (N_2817,N_1620,N_1948);
or U2818 (N_2818,N_1359,N_1964);
xor U2819 (N_2819,N_1763,N_1828);
and U2820 (N_2820,N_1734,N_1426);
or U2821 (N_2821,N_1112,N_1698);
and U2822 (N_2822,N_1177,N_1670);
nor U2823 (N_2823,N_1385,N_1367);
nand U2824 (N_2824,N_1766,N_1427);
or U2825 (N_2825,N_1448,N_1202);
and U2826 (N_2826,N_1992,N_1210);
nand U2827 (N_2827,N_1575,N_1727);
or U2828 (N_2828,N_1086,N_1541);
or U2829 (N_2829,N_1703,N_1930);
xnor U2830 (N_2830,N_1978,N_1591);
nor U2831 (N_2831,N_1339,N_1058);
xor U2832 (N_2832,N_1093,N_1996);
nand U2833 (N_2833,N_1340,N_1334);
or U2834 (N_2834,N_1096,N_1500);
and U2835 (N_2835,N_1834,N_1985);
or U2836 (N_2836,N_1297,N_1156);
xnor U2837 (N_2837,N_1002,N_1743);
xor U2838 (N_2838,N_1618,N_1468);
nand U2839 (N_2839,N_1564,N_1673);
xor U2840 (N_2840,N_1523,N_1446);
or U2841 (N_2841,N_1912,N_1051);
nor U2842 (N_2842,N_1243,N_1823);
xor U2843 (N_2843,N_1300,N_1000);
or U2844 (N_2844,N_1252,N_1226);
xor U2845 (N_2845,N_1783,N_1032);
and U2846 (N_2846,N_1596,N_1684);
nand U2847 (N_2847,N_1340,N_1176);
nand U2848 (N_2848,N_1385,N_1897);
xor U2849 (N_2849,N_1415,N_1150);
nand U2850 (N_2850,N_1094,N_1959);
xnor U2851 (N_2851,N_1166,N_1249);
nor U2852 (N_2852,N_1294,N_1374);
or U2853 (N_2853,N_1112,N_1974);
or U2854 (N_2854,N_1505,N_1170);
or U2855 (N_2855,N_1878,N_1325);
or U2856 (N_2856,N_1430,N_1009);
nand U2857 (N_2857,N_1491,N_1433);
nand U2858 (N_2858,N_1505,N_1270);
nand U2859 (N_2859,N_1936,N_1684);
nand U2860 (N_2860,N_1172,N_1542);
and U2861 (N_2861,N_1515,N_1005);
nor U2862 (N_2862,N_1727,N_1067);
nor U2863 (N_2863,N_1396,N_1540);
or U2864 (N_2864,N_1324,N_1148);
nor U2865 (N_2865,N_1456,N_1247);
or U2866 (N_2866,N_1489,N_1210);
xnor U2867 (N_2867,N_1973,N_1055);
and U2868 (N_2868,N_1535,N_1706);
or U2869 (N_2869,N_1283,N_1353);
and U2870 (N_2870,N_1978,N_1834);
or U2871 (N_2871,N_1558,N_1564);
xor U2872 (N_2872,N_1541,N_1898);
nand U2873 (N_2873,N_1566,N_1743);
xor U2874 (N_2874,N_1362,N_1522);
nor U2875 (N_2875,N_1356,N_1174);
and U2876 (N_2876,N_1789,N_1607);
nand U2877 (N_2877,N_1681,N_1186);
xnor U2878 (N_2878,N_1601,N_1161);
nand U2879 (N_2879,N_1534,N_1738);
nand U2880 (N_2880,N_1766,N_1292);
xnor U2881 (N_2881,N_1067,N_1326);
nand U2882 (N_2882,N_1899,N_1343);
nand U2883 (N_2883,N_1789,N_1209);
and U2884 (N_2884,N_1766,N_1305);
xnor U2885 (N_2885,N_1672,N_1974);
nand U2886 (N_2886,N_1478,N_1472);
nor U2887 (N_2887,N_1206,N_1063);
and U2888 (N_2888,N_1669,N_1450);
nor U2889 (N_2889,N_1872,N_1740);
and U2890 (N_2890,N_1510,N_1383);
nor U2891 (N_2891,N_1697,N_1069);
and U2892 (N_2892,N_1445,N_1534);
nand U2893 (N_2893,N_1548,N_1905);
nor U2894 (N_2894,N_1924,N_1791);
or U2895 (N_2895,N_1873,N_1394);
or U2896 (N_2896,N_1360,N_1827);
xnor U2897 (N_2897,N_1034,N_1955);
and U2898 (N_2898,N_1304,N_1953);
nand U2899 (N_2899,N_1362,N_1786);
and U2900 (N_2900,N_1583,N_1498);
nand U2901 (N_2901,N_1009,N_1187);
and U2902 (N_2902,N_1483,N_1813);
xnor U2903 (N_2903,N_1934,N_1821);
or U2904 (N_2904,N_1486,N_1361);
nand U2905 (N_2905,N_1533,N_1256);
xnor U2906 (N_2906,N_1838,N_1282);
or U2907 (N_2907,N_1139,N_1888);
nand U2908 (N_2908,N_1804,N_1381);
nor U2909 (N_2909,N_1713,N_1437);
nor U2910 (N_2910,N_1686,N_1392);
nand U2911 (N_2911,N_1049,N_1653);
nor U2912 (N_2912,N_1376,N_1179);
nor U2913 (N_2913,N_1076,N_1682);
xor U2914 (N_2914,N_1064,N_1516);
xnor U2915 (N_2915,N_1392,N_1905);
and U2916 (N_2916,N_1779,N_1521);
xor U2917 (N_2917,N_1672,N_1018);
nor U2918 (N_2918,N_1567,N_1236);
or U2919 (N_2919,N_1854,N_1358);
xor U2920 (N_2920,N_1748,N_1650);
xnor U2921 (N_2921,N_1921,N_1941);
nand U2922 (N_2922,N_1530,N_1397);
and U2923 (N_2923,N_1878,N_1813);
xnor U2924 (N_2924,N_1064,N_1036);
and U2925 (N_2925,N_1201,N_1330);
nand U2926 (N_2926,N_1624,N_1497);
nor U2927 (N_2927,N_1280,N_1510);
and U2928 (N_2928,N_1481,N_1162);
or U2929 (N_2929,N_1722,N_1035);
or U2930 (N_2930,N_1312,N_1676);
and U2931 (N_2931,N_1749,N_1304);
and U2932 (N_2932,N_1819,N_1267);
nor U2933 (N_2933,N_1315,N_1798);
nand U2934 (N_2934,N_1037,N_1760);
nand U2935 (N_2935,N_1134,N_1828);
xor U2936 (N_2936,N_1456,N_1063);
nand U2937 (N_2937,N_1314,N_1368);
xor U2938 (N_2938,N_1611,N_1885);
and U2939 (N_2939,N_1573,N_1183);
nor U2940 (N_2940,N_1694,N_1120);
nor U2941 (N_2941,N_1373,N_1954);
and U2942 (N_2942,N_1429,N_1197);
nand U2943 (N_2943,N_1539,N_1502);
and U2944 (N_2944,N_1659,N_1948);
and U2945 (N_2945,N_1847,N_1167);
nand U2946 (N_2946,N_1338,N_1023);
or U2947 (N_2947,N_1997,N_1221);
nand U2948 (N_2948,N_1767,N_1026);
and U2949 (N_2949,N_1422,N_1237);
nand U2950 (N_2950,N_1112,N_1789);
nor U2951 (N_2951,N_1149,N_1692);
xnor U2952 (N_2952,N_1874,N_1687);
nand U2953 (N_2953,N_1386,N_1940);
nor U2954 (N_2954,N_1982,N_1675);
xor U2955 (N_2955,N_1392,N_1768);
xnor U2956 (N_2956,N_1564,N_1586);
xnor U2957 (N_2957,N_1126,N_1895);
xor U2958 (N_2958,N_1334,N_1577);
nand U2959 (N_2959,N_1696,N_1150);
nor U2960 (N_2960,N_1588,N_1532);
nor U2961 (N_2961,N_1439,N_1907);
nor U2962 (N_2962,N_1650,N_1546);
nand U2963 (N_2963,N_1352,N_1006);
or U2964 (N_2964,N_1290,N_1450);
or U2965 (N_2965,N_1889,N_1977);
or U2966 (N_2966,N_1795,N_1809);
xnor U2967 (N_2967,N_1607,N_1878);
nor U2968 (N_2968,N_1531,N_1039);
nand U2969 (N_2969,N_1790,N_1392);
or U2970 (N_2970,N_1622,N_1288);
nor U2971 (N_2971,N_1623,N_1140);
xor U2972 (N_2972,N_1709,N_1882);
or U2973 (N_2973,N_1768,N_1119);
or U2974 (N_2974,N_1762,N_1143);
xnor U2975 (N_2975,N_1519,N_1093);
nand U2976 (N_2976,N_1976,N_1953);
and U2977 (N_2977,N_1964,N_1686);
nand U2978 (N_2978,N_1994,N_1435);
or U2979 (N_2979,N_1754,N_1667);
xor U2980 (N_2980,N_1397,N_1550);
nor U2981 (N_2981,N_1764,N_1451);
xnor U2982 (N_2982,N_1244,N_1367);
and U2983 (N_2983,N_1276,N_1154);
nor U2984 (N_2984,N_1163,N_1370);
and U2985 (N_2985,N_1917,N_1582);
nor U2986 (N_2986,N_1247,N_1726);
xnor U2987 (N_2987,N_1410,N_1153);
or U2988 (N_2988,N_1838,N_1102);
and U2989 (N_2989,N_1026,N_1519);
xnor U2990 (N_2990,N_1769,N_1297);
nor U2991 (N_2991,N_1465,N_1731);
xor U2992 (N_2992,N_1019,N_1703);
nand U2993 (N_2993,N_1266,N_1871);
xor U2994 (N_2994,N_1804,N_1187);
nand U2995 (N_2995,N_1046,N_1500);
nand U2996 (N_2996,N_1919,N_1673);
or U2997 (N_2997,N_1486,N_1004);
nand U2998 (N_2998,N_1385,N_1417);
and U2999 (N_2999,N_1905,N_1988);
or U3000 (N_3000,N_2885,N_2997);
xor U3001 (N_3001,N_2332,N_2802);
nand U3002 (N_3002,N_2824,N_2845);
and U3003 (N_3003,N_2543,N_2615);
or U3004 (N_3004,N_2699,N_2320);
or U3005 (N_3005,N_2273,N_2898);
and U3006 (N_3006,N_2105,N_2049);
xnor U3007 (N_3007,N_2361,N_2249);
and U3008 (N_3008,N_2602,N_2648);
and U3009 (N_3009,N_2117,N_2723);
or U3010 (N_3010,N_2402,N_2902);
xnor U3011 (N_3011,N_2920,N_2035);
xnor U3012 (N_3012,N_2005,N_2950);
and U3013 (N_3013,N_2869,N_2224);
xnor U3014 (N_3014,N_2722,N_2422);
xnor U3015 (N_3015,N_2796,N_2962);
nor U3016 (N_3016,N_2265,N_2888);
nor U3017 (N_3017,N_2212,N_2019);
nor U3018 (N_3018,N_2673,N_2551);
xor U3019 (N_3019,N_2496,N_2907);
and U3020 (N_3020,N_2868,N_2376);
xor U3021 (N_3021,N_2952,N_2115);
nand U3022 (N_3022,N_2283,N_2009);
or U3023 (N_3023,N_2524,N_2136);
and U3024 (N_3024,N_2610,N_2667);
nor U3025 (N_3025,N_2291,N_2507);
or U3026 (N_3026,N_2252,N_2965);
and U3027 (N_3027,N_2135,N_2839);
nand U3028 (N_3028,N_2169,N_2742);
xnor U3029 (N_3029,N_2506,N_2387);
nor U3030 (N_3030,N_2852,N_2978);
xor U3031 (N_3031,N_2398,N_2977);
or U3032 (N_3032,N_2934,N_2548);
xnor U3033 (N_3033,N_2143,N_2479);
xor U3034 (N_3034,N_2955,N_2598);
xnor U3035 (N_3035,N_2605,N_2349);
xor U3036 (N_3036,N_2979,N_2038);
or U3037 (N_3037,N_2566,N_2011);
xnor U3038 (N_3038,N_2989,N_2270);
or U3039 (N_3039,N_2938,N_2941);
or U3040 (N_3040,N_2816,N_2284);
xnor U3041 (N_3041,N_2031,N_2980);
xnor U3042 (N_3042,N_2672,N_2683);
nor U3043 (N_3043,N_2963,N_2500);
or U3044 (N_3044,N_2331,N_2485);
or U3045 (N_3045,N_2604,N_2383);
and U3046 (N_3046,N_2037,N_2835);
or U3047 (N_3047,N_2858,N_2318);
nor U3048 (N_3048,N_2828,N_2294);
and U3049 (N_3049,N_2231,N_2581);
and U3050 (N_3050,N_2146,N_2008);
xnor U3051 (N_3051,N_2002,N_2493);
nand U3052 (N_3052,N_2514,N_2185);
and U3053 (N_3053,N_2090,N_2101);
or U3054 (N_3054,N_2083,N_2862);
nor U3055 (N_3055,N_2245,N_2756);
nor U3056 (N_3056,N_2597,N_2201);
xnor U3057 (N_3057,N_2366,N_2119);
or U3058 (N_3058,N_2084,N_2323);
xnor U3059 (N_3059,N_2694,N_2867);
xnor U3060 (N_3060,N_2000,N_2365);
xor U3061 (N_3061,N_2333,N_2933);
and U3062 (N_3062,N_2140,N_2026);
or U3063 (N_3063,N_2822,N_2141);
nor U3064 (N_3064,N_2298,N_2513);
xor U3065 (N_3065,N_2727,N_2385);
and U3066 (N_3066,N_2488,N_2821);
nand U3067 (N_3067,N_2810,N_2209);
and U3068 (N_3068,N_2882,N_2712);
nand U3069 (N_3069,N_2515,N_2290);
xnor U3070 (N_3070,N_2057,N_2906);
xor U3071 (N_3071,N_2794,N_2216);
and U3072 (N_3072,N_2416,N_2181);
nand U3073 (N_3073,N_2919,N_2653);
or U3074 (N_3074,N_2313,N_2658);
nor U3075 (N_3075,N_2188,N_2996);
xnor U3076 (N_3076,N_2519,N_2271);
nor U3077 (N_3077,N_2544,N_2420);
nor U3078 (N_3078,N_2122,N_2295);
nor U3079 (N_3079,N_2655,N_2899);
or U3080 (N_3080,N_2157,N_2912);
or U3081 (N_3081,N_2477,N_2126);
nand U3082 (N_3082,N_2687,N_2556);
or U3083 (N_3083,N_2260,N_2873);
or U3084 (N_3084,N_2628,N_2277);
nor U3085 (N_3085,N_2576,N_2746);
xnor U3086 (N_3086,N_2510,N_2702);
nor U3087 (N_3087,N_2393,N_2749);
or U3088 (N_3088,N_2030,N_2713);
and U3089 (N_3089,N_2395,N_2645);
or U3090 (N_3090,N_2586,N_2879);
or U3091 (N_3091,N_2613,N_2847);
xnor U3092 (N_3092,N_2456,N_2646);
or U3093 (N_3093,N_2161,N_2937);
nand U3094 (N_3094,N_2220,N_2518);
and U3095 (N_3095,N_2511,N_2842);
nand U3096 (N_3096,N_2327,N_2991);
nand U3097 (N_3097,N_2974,N_2164);
xnor U3098 (N_3098,N_2239,N_2109);
nand U3099 (N_3099,N_2244,N_2721);
or U3100 (N_3100,N_2476,N_2329);
nand U3101 (N_3101,N_2995,N_2436);
and U3102 (N_3102,N_2338,N_2235);
nand U3103 (N_3103,N_2959,N_2681);
or U3104 (N_3104,N_2193,N_2582);
and U3105 (N_3105,N_2800,N_2512);
xnor U3106 (N_3106,N_2175,N_2641);
or U3107 (N_3107,N_2584,N_2783);
or U3108 (N_3108,N_2982,N_2106);
nor U3109 (N_3109,N_2182,N_2826);
xnor U3110 (N_3110,N_2324,N_2123);
nor U3111 (N_3111,N_2555,N_2047);
nand U3112 (N_3112,N_2150,N_2368);
xnor U3113 (N_3113,N_2166,N_2677);
or U3114 (N_3114,N_2362,N_2676);
xnor U3115 (N_3115,N_2442,N_2183);
nand U3116 (N_3116,N_2373,N_2369);
nor U3117 (N_3117,N_2798,N_2241);
nor U3118 (N_3118,N_2799,N_2326);
or U3119 (N_3119,N_2056,N_2389);
and U3120 (N_3120,N_2390,N_2179);
or U3121 (N_3121,N_2303,N_2403);
and U3122 (N_3122,N_2599,N_2872);
or U3123 (N_3123,N_2527,N_2480);
xor U3124 (N_3124,N_2767,N_2423);
xnor U3125 (N_3125,N_2027,N_2345);
and U3126 (N_3126,N_2431,N_2944);
or U3127 (N_3127,N_2219,N_2714);
or U3128 (N_3128,N_2081,N_2042);
nand U3129 (N_3129,N_2690,N_2426);
nand U3130 (N_3130,N_2396,N_2595);
nor U3131 (N_3131,N_2116,N_2635);
or U3132 (N_3132,N_2302,N_2987);
nor U3133 (N_3133,N_2846,N_2281);
nand U3134 (N_3134,N_2350,N_2264);
nor U3135 (N_3135,N_2654,N_2675);
xor U3136 (N_3136,N_2204,N_2787);
nand U3137 (N_3137,N_2400,N_2473);
xor U3138 (N_3138,N_2099,N_2454);
and U3139 (N_3139,N_2770,N_2680);
nand U3140 (N_3140,N_2497,N_2730);
and U3141 (N_3141,N_2659,N_2568);
and U3142 (N_3142,N_2399,N_2900);
nor U3143 (N_3143,N_2718,N_2129);
or U3144 (N_3144,N_2625,N_2642);
nand U3145 (N_3145,N_2128,N_2697);
nand U3146 (N_3146,N_2278,N_2177);
nor U3147 (N_3147,N_2428,N_2623);
nand U3148 (N_3148,N_2616,N_2936);
and U3149 (N_3149,N_2768,N_2010);
and U3150 (N_3150,N_2843,N_2939);
or U3151 (N_3151,N_2203,N_2516);
and U3152 (N_3152,N_2620,N_2643);
or U3153 (N_3153,N_2634,N_2779);
nand U3154 (N_3154,N_2296,N_2475);
or U3155 (N_3155,N_2788,N_2577);
or U3156 (N_3156,N_2441,N_2017);
nor U3157 (N_3157,N_2662,N_2619);
nor U3158 (N_3158,N_2703,N_2587);
nand U3159 (N_3159,N_2674,N_2606);
nand U3160 (N_3160,N_2994,N_2924);
nand U3161 (N_3161,N_2469,N_2127);
xnor U3162 (N_3162,N_2927,N_2559);
or U3163 (N_3163,N_2857,N_2525);
nand U3164 (N_3164,N_2227,N_2550);
nand U3165 (N_3165,N_2501,N_2414);
xnor U3166 (N_3166,N_2915,N_2750);
xnor U3167 (N_3167,N_2339,N_2829);
xnor U3168 (N_3168,N_2693,N_2124);
xor U3169 (N_3169,N_2614,N_2021);
nor U3170 (N_3170,N_2992,N_2443);
and U3171 (N_3171,N_2754,N_2744);
xor U3172 (N_3172,N_2347,N_2719);
xnor U3173 (N_3173,N_2063,N_2285);
xor U3174 (N_3174,N_2608,N_2110);
or U3175 (N_3175,N_2528,N_2180);
and U3176 (N_3176,N_2388,N_2863);
and U3177 (N_3177,N_2287,N_2752);
xor U3178 (N_3178,N_2738,N_2158);
xnor U3179 (N_3179,N_2357,N_2808);
nor U3180 (N_3180,N_2904,N_2151);
and U3181 (N_3181,N_2640,N_2553);
and U3182 (N_3182,N_2014,N_2195);
xor U3183 (N_3183,N_2045,N_2751);
and U3184 (N_3184,N_2948,N_2878);
nand U3185 (N_3185,N_2592,N_2541);
nor U3186 (N_3186,N_2272,N_2424);
xnor U3187 (N_3187,N_2459,N_2893);
and U3188 (N_3188,N_2032,N_2044);
or U3189 (N_3189,N_2975,N_2689);
or U3190 (N_3190,N_2538,N_2825);
nand U3191 (N_3191,N_2678,N_2237);
xor U3192 (N_3192,N_2053,N_2375);
and U3193 (N_3193,N_2956,N_2755);
nand U3194 (N_3194,N_2359,N_2916);
nand U3195 (N_3195,N_2665,N_2013);
or U3196 (N_3196,N_2134,N_2757);
nand U3197 (N_3197,N_2760,N_2268);
nand U3198 (N_3198,N_2269,N_2579);
and U3199 (N_3199,N_2957,N_2363);
nor U3200 (N_3200,N_2707,N_2895);
nor U3201 (N_3201,N_2230,N_2133);
or U3202 (N_3202,N_2438,N_2953);
or U3203 (N_3203,N_2671,N_2542);
or U3204 (N_3204,N_2591,N_2552);
or U3205 (N_3205,N_2050,N_2334);
nor U3206 (N_3206,N_2207,N_2095);
nand U3207 (N_3207,N_2897,N_2540);
and U3208 (N_3208,N_2517,N_2322);
nor U3209 (N_3209,N_2004,N_2509);
nand U3210 (N_3210,N_2851,N_2533);
xor U3211 (N_3211,N_2711,N_2132);
nand U3212 (N_3212,N_2205,N_2708);
xor U3213 (N_3213,N_2661,N_2739);
or U3214 (N_3214,N_2728,N_2892);
xnor U3215 (N_3215,N_2998,N_2812);
nand U3216 (N_3216,N_2669,N_2064);
and U3217 (N_3217,N_2918,N_2412);
or U3218 (N_3218,N_2217,N_2404);
nor U3219 (N_3219,N_2173,N_2487);
and U3220 (N_3220,N_2560,N_2776);
and U3221 (N_3221,N_2321,N_2418);
or U3222 (N_3222,N_2870,N_2649);
and U3223 (N_3223,N_2379,N_2214);
nor U3224 (N_3224,N_2815,N_2314);
and U3225 (N_3225,N_2831,N_2240);
or U3226 (N_3226,N_2600,N_2526);
and U3227 (N_3227,N_2360,N_2837);
xnor U3228 (N_3228,N_2999,N_2208);
xnor U3229 (N_3229,N_2494,N_2773);
nand U3230 (N_3230,N_2850,N_2262);
xnor U3231 (N_3231,N_2701,N_2336);
xor U3232 (N_3232,N_2896,N_2905);
nor U3233 (N_3233,N_2710,N_2276);
and U3234 (N_3234,N_2725,N_2142);
nand U3235 (N_3235,N_2621,N_2306);
xnor U3236 (N_3236,N_2356,N_2251);
xnor U3237 (N_3237,N_2853,N_2985);
and U3238 (N_3238,N_2964,N_2622);
or U3239 (N_3239,N_2917,N_2883);
or U3240 (N_3240,N_2753,N_2909);
nand U3241 (N_3241,N_2198,N_2951);
nand U3242 (N_3242,N_2889,N_2585);
nor U3243 (N_3243,N_2624,N_2337);
xnor U3244 (N_3244,N_2946,N_2864);
nand U3245 (N_3245,N_2588,N_2293);
xnor U3246 (N_3246,N_2392,N_2445);
or U3247 (N_3247,N_2068,N_2736);
or U3248 (N_3248,N_2601,N_2886);
nor U3249 (N_3249,N_2297,N_2894);
xor U3250 (N_3250,N_2328,N_2156);
nand U3251 (N_3251,N_2092,N_2644);
xnor U3252 (N_3252,N_2261,N_2930);
xnor U3253 (N_3253,N_2319,N_2256);
xor U3254 (N_3254,N_2351,N_2961);
and U3255 (N_3255,N_2355,N_2374);
nor U3256 (N_3256,N_2700,N_2887);
xnor U3257 (N_3257,N_2534,N_2967);
xor U3258 (N_3258,N_2435,N_2499);
xnor U3259 (N_3259,N_2731,N_2748);
nor U3260 (N_3260,N_2405,N_2343);
xor U3261 (N_3261,N_2455,N_2732);
nand U3262 (N_3262,N_2317,N_2636);
xor U3263 (N_3263,N_2811,N_2429);
nor U3264 (N_3264,N_2949,N_2809);
nand U3265 (N_3265,N_2470,N_2733);
nand U3266 (N_3266,N_2679,N_2263);
nor U3267 (N_3267,N_2472,N_2197);
xnor U3268 (N_3268,N_2187,N_2299);
and U3269 (N_3269,N_2647,N_2073);
xor U3270 (N_3270,N_2639,N_2218);
xnor U3271 (N_3271,N_2066,N_2695);
xnor U3272 (N_3272,N_2759,N_2481);
nand U3273 (N_3273,N_2567,N_2737);
or U3274 (N_3274,N_2311,N_2921);
nand U3275 (N_3275,N_2091,N_2165);
and U3276 (N_3276,N_2108,N_2532);
nor U3277 (N_3277,N_2025,N_2795);
nand U3278 (N_3278,N_2061,N_2451);
nor U3279 (N_3279,N_2280,N_2250);
nor U3280 (N_3280,N_2943,N_2503);
or U3281 (N_3281,N_2765,N_2942);
or U3282 (N_3282,N_2255,N_2861);
or U3283 (N_3283,N_2530,N_2232);
and U3284 (N_3284,N_2401,N_2492);
nand U3285 (N_3285,N_2215,N_2785);
and U3286 (N_3286,N_2908,N_2876);
nand U3287 (N_3287,N_2784,N_2618);
nor U3288 (N_3288,N_2086,N_2705);
and U3289 (N_3289,N_2437,N_2603);
and U3290 (N_3290,N_2419,N_2814);
nand U3291 (N_3291,N_2384,N_2176);
nor U3292 (N_3292,N_2028,N_2935);
and U3293 (N_3293,N_2266,N_2844);
or U3294 (N_3294,N_2397,N_2415);
nor U3295 (N_3295,N_2663,N_2148);
nor U3296 (N_3296,N_2447,N_2570);
xor U3297 (N_3297,N_2929,N_2001);
or U3298 (N_3298,N_2346,N_2801);
nand U3299 (N_3299,N_2305,N_2316);
nor U3300 (N_3300,N_2211,N_2098);
xnor U3301 (N_3301,N_2529,N_2791);
and U3302 (N_3302,N_2370,N_2832);
xnor U3303 (N_3303,N_2743,N_2820);
nor U3304 (N_3304,N_2107,N_2840);
or U3305 (N_3305,N_2594,N_2466);
nor U3306 (N_3306,N_2970,N_2629);
or U3307 (N_3307,N_2039,N_2131);
xnor U3308 (N_3308,N_2471,N_2167);
nand U3309 (N_3309,N_2223,N_2780);
nand U3310 (N_3310,N_2221,N_2981);
xnor U3311 (N_3311,N_2254,N_2609);
or U3312 (N_3312,N_2571,N_2911);
and U3313 (N_3313,N_2782,N_2626);
xor U3314 (N_3314,N_2865,N_2903);
nand U3315 (N_3315,N_2590,N_2386);
or U3316 (N_3316,N_2154,N_2352);
and U3317 (N_3317,N_2856,N_2758);
xnor U3318 (N_3318,N_2309,N_2225);
xor U3319 (N_3319,N_2766,N_2656);
or U3320 (N_3320,N_2194,N_2304);
and U3321 (N_3321,N_2813,N_2015);
nor U3322 (N_3322,N_2666,N_2928);
nand U3323 (N_3323,N_2474,N_2686);
or U3324 (N_3324,N_2046,N_2380);
or U3325 (N_3325,N_2698,N_2724);
or U3326 (N_3326,N_2490,N_2578);
nor U3327 (N_3327,N_2922,N_2267);
or U3328 (N_3328,N_2051,N_2054);
nor U3329 (N_3329,N_2554,N_2682);
nor U3330 (N_3330,N_2461,N_2575);
nor U3331 (N_3331,N_2875,N_2772);
xnor U3332 (N_3332,N_2206,N_2834);
or U3333 (N_3333,N_2781,N_2630);
nor U3334 (N_3334,N_2391,N_2539);
nor U3335 (N_3335,N_2547,N_2657);
nor U3336 (N_3336,N_2972,N_2102);
nand U3337 (N_3337,N_2052,N_2427);
nand U3338 (N_3338,N_2836,N_2914);
or U3339 (N_3339,N_2508,N_2171);
xnor U3340 (N_3340,N_2130,N_2866);
and U3341 (N_3341,N_2411,N_2279);
xor U3342 (N_3342,N_2521,N_2838);
nand U3343 (N_3343,N_2243,N_2762);
or U3344 (N_3344,N_2089,N_2104);
nor U3345 (N_3345,N_2817,N_2716);
nand U3346 (N_3346,N_2200,N_2282);
xnor U3347 (N_3347,N_2377,N_2631);
nand U3348 (N_3348,N_2155,N_2486);
or U3349 (N_3349,N_2463,N_2034);
and U3350 (N_3350,N_2353,N_2855);
xnor U3351 (N_3351,N_2633,N_2777);
nor U3352 (N_3352,N_2531,N_2335);
and U3353 (N_3353,N_2342,N_2112);
xor U3354 (N_3354,N_2545,N_2189);
nor U3355 (N_3355,N_2465,N_2877);
xor U3356 (N_3356,N_2307,N_2096);
xnor U3357 (N_3357,N_2007,N_2163);
nand U3358 (N_3358,N_2596,N_2792);
and U3359 (N_3359,N_2184,N_2274);
nor U3360 (N_3360,N_2706,N_2325);
and U3361 (N_3361,N_2670,N_2890);
nor U3362 (N_3362,N_2704,N_2976);
nor U3363 (N_3363,N_2523,N_2080);
and U3364 (N_3364,N_2988,N_2734);
or U3365 (N_3365,N_2139,N_2823);
nor U3366 (N_3366,N_2522,N_2078);
nand U3367 (N_3367,N_2968,N_2196);
nor U3368 (N_3368,N_2060,N_2036);
and U3369 (N_3369,N_2043,N_2790);
and U3370 (N_3370,N_2969,N_2789);
and U3371 (N_3371,N_2536,N_2315);
or U3372 (N_3372,N_2087,N_2460);
nand U3373 (N_3373,N_2430,N_2312);
or U3374 (N_3374,N_2668,N_2717);
or U3375 (N_3375,N_2583,N_2803);
nand U3376 (N_3376,N_2074,N_2786);
or U3377 (N_3377,N_2881,N_2071);
nand U3378 (N_3378,N_2557,N_2275);
nor U3379 (N_3379,N_2685,N_2288);
nor U3380 (N_3380,N_2040,N_2120);
or U3381 (N_3381,N_2145,N_2072);
or U3382 (N_3382,N_2168,N_2178);
or U3383 (N_3383,N_2213,N_2162);
nand U3384 (N_3384,N_2923,N_2520);
or U3385 (N_3385,N_2449,N_2041);
xor U3386 (N_3386,N_2771,N_2023);
nor U3387 (N_3387,N_2121,N_2382);
xor U3388 (N_3388,N_2286,N_2569);
nand U3389 (N_3389,N_2259,N_2709);
or U3390 (N_3390,N_2637,N_2174);
xnor U3391 (N_3391,N_2495,N_2891);
xor U3392 (N_3392,N_2144,N_2354);
or U3393 (N_3393,N_2300,N_2075);
and U3394 (N_3394,N_2082,N_2925);
nor U3395 (N_3395,N_2229,N_2458);
nand U3396 (N_3396,N_2931,N_2258);
nand U3397 (N_3397,N_2421,N_2372);
nand U3398 (N_3398,N_2993,N_2960);
nand U3399 (N_3399,N_2192,N_2761);
or U3400 (N_3400,N_2448,N_2003);
nand U3401 (N_3401,N_2573,N_2535);
nand U3402 (N_3402,N_2860,N_2880);
and U3403 (N_3403,N_2793,N_2688);
nor U3404 (N_3404,N_2113,N_2806);
nor U3405 (N_3405,N_2100,N_2627);
and U3406 (N_3406,N_2692,N_2301);
xnor U3407 (N_3407,N_2341,N_2546);
nor U3408 (N_3408,N_2617,N_2149);
nand U3409 (N_3409,N_2740,N_2735);
nand U3410 (N_3410,N_2684,N_2726);
nor U3411 (N_3411,N_2018,N_2910);
nor U3412 (N_3412,N_2807,N_2652);
or U3413 (N_3413,N_2572,N_2114);
or U3414 (N_3414,N_2498,N_2067);
xor U3415 (N_3415,N_2406,N_2202);
nand U3416 (N_3416,N_2024,N_2439);
or U3417 (N_3417,N_2947,N_2253);
xnor U3418 (N_3418,N_2147,N_2502);
xnor U3419 (N_3419,N_2450,N_2159);
xnor U3420 (N_3420,N_2446,N_2434);
and U3421 (N_3421,N_2289,N_2022);
and U3422 (N_3422,N_2859,N_2330);
xnor U3423 (N_3423,N_2088,N_2805);
xnor U3424 (N_3424,N_2079,N_2932);
xor U3425 (N_3425,N_2901,N_2029);
or U3426 (N_3426,N_2006,N_2248);
nor U3427 (N_3427,N_2125,N_2562);
nor U3428 (N_3428,N_2468,N_2478);
or U3429 (N_3429,N_2233,N_2440);
nor U3430 (N_3430,N_2691,N_2190);
and U3431 (N_3431,N_2137,N_2062);
xnor U3432 (N_3432,N_2797,N_2462);
or U3433 (N_3433,N_2971,N_2408);
nand U3434 (N_3434,N_2775,N_2407);
nor U3435 (N_3435,N_2020,N_2660);
xnor U3436 (N_3436,N_2504,N_2778);
nand U3437 (N_3437,N_2433,N_2247);
nand U3438 (N_3438,N_2650,N_2210);
xor U3439 (N_3439,N_2093,N_2558);
xnor U3440 (N_3440,N_2574,N_2827);
or U3441 (N_3441,N_2945,N_2308);
and U3442 (N_3442,N_2611,N_2940);
nand U3443 (N_3443,N_2958,N_2103);
or U3444 (N_3444,N_2413,N_2484);
or U3445 (N_3445,N_2854,N_2048);
xor U3446 (N_3446,N_2065,N_2874);
nor U3447 (N_3447,N_2344,N_2453);
nor U3448 (N_3448,N_2016,N_2841);
nor U3449 (N_3449,N_2226,N_2242);
or U3450 (N_3450,N_2833,N_2118);
xnor U3451 (N_3451,N_2926,N_2984);
nor U3452 (N_3452,N_2348,N_2292);
nand U3453 (N_3453,N_2747,N_2819);
xnor U3454 (N_3454,N_2059,N_2830);
or U3455 (N_3455,N_2417,N_2973);
nor U3456 (N_3456,N_2763,N_2986);
xnor U3457 (N_3457,N_2236,N_2565);
or U3458 (N_3458,N_2381,N_2489);
nor U3459 (N_3459,N_2077,N_2848);
or U3460 (N_3460,N_2549,N_2849);
or U3461 (N_3461,N_2186,N_2561);
xor U3462 (N_3462,N_2612,N_2990);
and U3463 (N_3463,N_2152,N_2607);
nand U3464 (N_3464,N_2729,N_2651);
and U3465 (N_3465,N_2467,N_2234);
nand U3466 (N_3466,N_2425,N_2482);
xor U3467 (N_3467,N_2153,N_2537);
nor U3468 (N_3468,N_2580,N_2246);
or U3469 (N_3469,N_2818,N_2804);
nand U3470 (N_3470,N_2111,N_2191);
and U3471 (N_3471,N_2094,N_2774);
or U3472 (N_3472,N_2452,N_2371);
xor U3473 (N_3473,N_2055,N_2769);
nor U3474 (N_3474,N_2238,N_2222);
and U3475 (N_3475,N_2884,N_2871);
or U3476 (N_3476,N_2085,N_2491);
nand U3477 (N_3477,N_2593,N_2076);
or U3478 (N_3478,N_2741,N_2505);
and U3479 (N_3479,N_2340,N_2483);
nand U3480 (N_3480,N_2664,N_2310);
nor U3481 (N_3481,N_2228,N_2638);
xnor U3482 (N_3482,N_2070,N_2589);
and U3483 (N_3483,N_2983,N_2170);
xor U3484 (N_3484,N_2199,N_2457);
and U3485 (N_3485,N_2160,N_2464);
and U3486 (N_3486,N_2097,N_2058);
or U3487 (N_3487,N_2632,N_2172);
and U3488 (N_3488,N_2720,N_2966);
nor U3489 (N_3489,N_2715,N_2764);
xnor U3490 (N_3490,N_2410,N_2012);
xnor U3491 (N_3491,N_2444,N_2378);
xor U3492 (N_3492,N_2954,N_2432);
nand U3493 (N_3493,N_2257,N_2138);
nand U3494 (N_3494,N_2696,N_2367);
or U3495 (N_3495,N_2069,N_2409);
nor U3496 (N_3496,N_2564,N_2033);
or U3497 (N_3497,N_2563,N_2394);
xor U3498 (N_3498,N_2358,N_2364);
or U3499 (N_3499,N_2745,N_2913);
nor U3500 (N_3500,N_2500,N_2738);
nor U3501 (N_3501,N_2132,N_2022);
nand U3502 (N_3502,N_2333,N_2640);
or U3503 (N_3503,N_2674,N_2227);
xnor U3504 (N_3504,N_2581,N_2433);
and U3505 (N_3505,N_2960,N_2418);
or U3506 (N_3506,N_2087,N_2147);
or U3507 (N_3507,N_2237,N_2842);
nand U3508 (N_3508,N_2688,N_2627);
or U3509 (N_3509,N_2814,N_2420);
and U3510 (N_3510,N_2412,N_2080);
nor U3511 (N_3511,N_2983,N_2639);
or U3512 (N_3512,N_2418,N_2557);
xnor U3513 (N_3513,N_2729,N_2898);
or U3514 (N_3514,N_2291,N_2990);
or U3515 (N_3515,N_2780,N_2678);
nor U3516 (N_3516,N_2267,N_2084);
nor U3517 (N_3517,N_2856,N_2027);
and U3518 (N_3518,N_2908,N_2328);
nor U3519 (N_3519,N_2101,N_2534);
xor U3520 (N_3520,N_2837,N_2051);
nand U3521 (N_3521,N_2726,N_2151);
nand U3522 (N_3522,N_2637,N_2651);
xor U3523 (N_3523,N_2214,N_2404);
nor U3524 (N_3524,N_2013,N_2971);
or U3525 (N_3525,N_2676,N_2494);
nor U3526 (N_3526,N_2051,N_2778);
xnor U3527 (N_3527,N_2638,N_2013);
or U3528 (N_3528,N_2351,N_2574);
xnor U3529 (N_3529,N_2937,N_2270);
or U3530 (N_3530,N_2677,N_2938);
nor U3531 (N_3531,N_2421,N_2418);
or U3532 (N_3532,N_2147,N_2309);
nand U3533 (N_3533,N_2428,N_2374);
xor U3534 (N_3534,N_2460,N_2767);
and U3535 (N_3535,N_2202,N_2253);
nand U3536 (N_3536,N_2197,N_2023);
xnor U3537 (N_3537,N_2698,N_2716);
or U3538 (N_3538,N_2460,N_2750);
nand U3539 (N_3539,N_2496,N_2388);
nor U3540 (N_3540,N_2140,N_2194);
or U3541 (N_3541,N_2373,N_2475);
nand U3542 (N_3542,N_2009,N_2290);
and U3543 (N_3543,N_2543,N_2082);
or U3544 (N_3544,N_2573,N_2043);
or U3545 (N_3545,N_2268,N_2694);
nor U3546 (N_3546,N_2370,N_2628);
nand U3547 (N_3547,N_2517,N_2691);
nand U3548 (N_3548,N_2088,N_2567);
nor U3549 (N_3549,N_2447,N_2425);
and U3550 (N_3550,N_2267,N_2123);
or U3551 (N_3551,N_2700,N_2327);
or U3552 (N_3552,N_2594,N_2311);
nor U3553 (N_3553,N_2638,N_2127);
and U3554 (N_3554,N_2516,N_2050);
xnor U3555 (N_3555,N_2817,N_2250);
or U3556 (N_3556,N_2715,N_2298);
nand U3557 (N_3557,N_2110,N_2058);
xor U3558 (N_3558,N_2641,N_2974);
and U3559 (N_3559,N_2257,N_2399);
nand U3560 (N_3560,N_2378,N_2765);
and U3561 (N_3561,N_2263,N_2483);
and U3562 (N_3562,N_2594,N_2000);
or U3563 (N_3563,N_2280,N_2406);
and U3564 (N_3564,N_2100,N_2368);
and U3565 (N_3565,N_2132,N_2224);
nor U3566 (N_3566,N_2975,N_2940);
nand U3567 (N_3567,N_2786,N_2569);
xnor U3568 (N_3568,N_2439,N_2244);
and U3569 (N_3569,N_2655,N_2870);
xor U3570 (N_3570,N_2559,N_2876);
nor U3571 (N_3571,N_2650,N_2054);
or U3572 (N_3572,N_2528,N_2075);
or U3573 (N_3573,N_2215,N_2514);
nor U3574 (N_3574,N_2511,N_2467);
nor U3575 (N_3575,N_2682,N_2775);
nor U3576 (N_3576,N_2307,N_2984);
or U3577 (N_3577,N_2953,N_2626);
or U3578 (N_3578,N_2573,N_2867);
or U3579 (N_3579,N_2656,N_2922);
xor U3580 (N_3580,N_2679,N_2303);
xor U3581 (N_3581,N_2304,N_2193);
or U3582 (N_3582,N_2952,N_2488);
nor U3583 (N_3583,N_2334,N_2930);
or U3584 (N_3584,N_2470,N_2110);
nor U3585 (N_3585,N_2857,N_2881);
nand U3586 (N_3586,N_2970,N_2865);
nor U3587 (N_3587,N_2898,N_2613);
nand U3588 (N_3588,N_2173,N_2270);
nand U3589 (N_3589,N_2868,N_2845);
or U3590 (N_3590,N_2626,N_2235);
xnor U3591 (N_3591,N_2674,N_2873);
and U3592 (N_3592,N_2238,N_2350);
xnor U3593 (N_3593,N_2839,N_2486);
nor U3594 (N_3594,N_2805,N_2375);
nor U3595 (N_3595,N_2831,N_2126);
or U3596 (N_3596,N_2012,N_2354);
and U3597 (N_3597,N_2945,N_2958);
nand U3598 (N_3598,N_2039,N_2243);
xnor U3599 (N_3599,N_2161,N_2800);
xnor U3600 (N_3600,N_2215,N_2576);
nor U3601 (N_3601,N_2295,N_2026);
or U3602 (N_3602,N_2272,N_2056);
xnor U3603 (N_3603,N_2408,N_2606);
nand U3604 (N_3604,N_2679,N_2557);
xnor U3605 (N_3605,N_2574,N_2433);
nand U3606 (N_3606,N_2734,N_2710);
nor U3607 (N_3607,N_2376,N_2511);
nor U3608 (N_3608,N_2546,N_2687);
nand U3609 (N_3609,N_2865,N_2198);
xor U3610 (N_3610,N_2722,N_2641);
nand U3611 (N_3611,N_2902,N_2491);
or U3612 (N_3612,N_2053,N_2162);
or U3613 (N_3613,N_2313,N_2824);
or U3614 (N_3614,N_2770,N_2657);
and U3615 (N_3615,N_2828,N_2159);
nor U3616 (N_3616,N_2053,N_2456);
nor U3617 (N_3617,N_2709,N_2585);
nor U3618 (N_3618,N_2063,N_2908);
and U3619 (N_3619,N_2453,N_2319);
nand U3620 (N_3620,N_2140,N_2630);
nand U3621 (N_3621,N_2199,N_2426);
or U3622 (N_3622,N_2897,N_2170);
and U3623 (N_3623,N_2364,N_2906);
nand U3624 (N_3624,N_2688,N_2335);
or U3625 (N_3625,N_2291,N_2544);
xor U3626 (N_3626,N_2695,N_2304);
nand U3627 (N_3627,N_2342,N_2652);
and U3628 (N_3628,N_2684,N_2663);
or U3629 (N_3629,N_2610,N_2488);
and U3630 (N_3630,N_2148,N_2864);
or U3631 (N_3631,N_2856,N_2010);
nand U3632 (N_3632,N_2734,N_2701);
nor U3633 (N_3633,N_2554,N_2608);
nor U3634 (N_3634,N_2555,N_2965);
xnor U3635 (N_3635,N_2683,N_2614);
nor U3636 (N_3636,N_2816,N_2796);
xnor U3637 (N_3637,N_2289,N_2787);
and U3638 (N_3638,N_2836,N_2649);
or U3639 (N_3639,N_2936,N_2661);
xor U3640 (N_3640,N_2132,N_2878);
nand U3641 (N_3641,N_2710,N_2383);
xnor U3642 (N_3642,N_2420,N_2790);
and U3643 (N_3643,N_2185,N_2111);
xor U3644 (N_3644,N_2838,N_2942);
xnor U3645 (N_3645,N_2282,N_2663);
nor U3646 (N_3646,N_2086,N_2099);
and U3647 (N_3647,N_2526,N_2409);
nand U3648 (N_3648,N_2153,N_2611);
nor U3649 (N_3649,N_2088,N_2419);
xnor U3650 (N_3650,N_2512,N_2933);
or U3651 (N_3651,N_2646,N_2956);
nor U3652 (N_3652,N_2356,N_2422);
xor U3653 (N_3653,N_2304,N_2576);
and U3654 (N_3654,N_2351,N_2233);
xor U3655 (N_3655,N_2319,N_2154);
nand U3656 (N_3656,N_2852,N_2201);
nand U3657 (N_3657,N_2521,N_2005);
xnor U3658 (N_3658,N_2900,N_2634);
xor U3659 (N_3659,N_2344,N_2970);
nand U3660 (N_3660,N_2868,N_2174);
or U3661 (N_3661,N_2997,N_2954);
and U3662 (N_3662,N_2057,N_2913);
nand U3663 (N_3663,N_2926,N_2318);
and U3664 (N_3664,N_2458,N_2461);
or U3665 (N_3665,N_2663,N_2105);
or U3666 (N_3666,N_2454,N_2416);
nor U3667 (N_3667,N_2984,N_2656);
nor U3668 (N_3668,N_2314,N_2822);
or U3669 (N_3669,N_2076,N_2357);
or U3670 (N_3670,N_2861,N_2298);
or U3671 (N_3671,N_2015,N_2405);
or U3672 (N_3672,N_2821,N_2731);
nor U3673 (N_3673,N_2134,N_2911);
nand U3674 (N_3674,N_2407,N_2955);
xnor U3675 (N_3675,N_2539,N_2843);
or U3676 (N_3676,N_2248,N_2157);
nand U3677 (N_3677,N_2316,N_2445);
nand U3678 (N_3678,N_2971,N_2990);
xnor U3679 (N_3679,N_2535,N_2396);
and U3680 (N_3680,N_2619,N_2084);
nand U3681 (N_3681,N_2131,N_2858);
and U3682 (N_3682,N_2312,N_2386);
or U3683 (N_3683,N_2305,N_2063);
xor U3684 (N_3684,N_2894,N_2416);
and U3685 (N_3685,N_2267,N_2268);
or U3686 (N_3686,N_2691,N_2003);
and U3687 (N_3687,N_2269,N_2230);
xor U3688 (N_3688,N_2727,N_2484);
or U3689 (N_3689,N_2900,N_2249);
nand U3690 (N_3690,N_2763,N_2645);
and U3691 (N_3691,N_2182,N_2948);
or U3692 (N_3692,N_2549,N_2206);
nor U3693 (N_3693,N_2527,N_2776);
nand U3694 (N_3694,N_2633,N_2732);
or U3695 (N_3695,N_2468,N_2072);
or U3696 (N_3696,N_2050,N_2311);
or U3697 (N_3697,N_2033,N_2693);
and U3698 (N_3698,N_2904,N_2648);
xor U3699 (N_3699,N_2213,N_2999);
and U3700 (N_3700,N_2276,N_2510);
or U3701 (N_3701,N_2425,N_2904);
and U3702 (N_3702,N_2440,N_2739);
nor U3703 (N_3703,N_2128,N_2498);
nor U3704 (N_3704,N_2877,N_2222);
nor U3705 (N_3705,N_2421,N_2502);
and U3706 (N_3706,N_2879,N_2070);
or U3707 (N_3707,N_2094,N_2863);
nand U3708 (N_3708,N_2370,N_2509);
and U3709 (N_3709,N_2100,N_2261);
or U3710 (N_3710,N_2618,N_2626);
nor U3711 (N_3711,N_2982,N_2094);
nor U3712 (N_3712,N_2044,N_2878);
nor U3713 (N_3713,N_2386,N_2742);
or U3714 (N_3714,N_2177,N_2338);
xor U3715 (N_3715,N_2349,N_2222);
and U3716 (N_3716,N_2662,N_2203);
nand U3717 (N_3717,N_2270,N_2517);
nand U3718 (N_3718,N_2446,N_2535);
nor U3719 (N_3719,N_2407,N_2405);
or U3720 (N_3720,N_2883,N_2093);
xor U3721 (N_3721,N_2887,N_2201);
or U3722 (N_3722,N_2134,N_2682);
or U3723 (N_3723,N_2402,N_2015);
nor U3724 (N_3724,N_2176,N_2034);
xor U3725 (N_3725,N_2972,N_2814);
xnor U3726 (N_3726,N_2644,N_2404);
nand U3727 (N_3727,N_2928,N_2675);
or U3728 (N_3728,N_2264,N_2828);
or U3729 (N_3729,N_2744,N_2048);
xor U3730 (N_3730,N_2786,N_2882);
xnor U3731 (N_3731,N_2439,N_2503);
nand U3732 (N_3732,N_2478,N_2580);
xor U3733 (N_3733,N_2339,N_2664);
xnor U3734 (N_3734,N_2460,N_2539);
or U3735 (N_3735,N_2955,N_2272);
nor U3736 (N_3736,N_2640,N_2181);
or U3737 (N_3737,N_2208,N_2082);
or U3738 (N_3738,N_2977,N_2971);
xnor U3739 (N_3739,N_2759,N_2436);
or U3740 (N_3740,N_2399,N_2611);
and U3741 (N_3741,N_2862,N_2875);
or U3742 (N_3742,N_2326,N_2750);
xnor U3743 (N_3743,N_2398,N_2873);
and U3744 (N_3744,N_2658,N_2438);
or U3745 (N_3745,N_2849,N_2290);
or U3746 (N_3746,N_2288,N_2557);
xnor U3747 (N_3747,N_2007,N_2187);
nor U3748 (N_3748,N_2626,N_2001);
nand U3749 (N_3749,N_2884,N_2792);
nor U3750 (N_3750,N_2627,N_2117);
nand U3751 (N_3751,N_2573,N_2822);
nor U3752 (N_3752,N_2706,N_2723);
and U3753 (N_3753,N_2762,N_2758);
nor U3754 (N_3754,N_2394,N_2847);
and U3755 (N_3755,N_2054,N_2861);
nor U3756 (N_3756,N_2116,N_2722);
or U3757 (N_3757,N_2815,N_2523);
xnor U3758 (N_3758,N_2223,N_2268);
nand U3759 (N_3759,N_2402,N_2796);
or U3760 (N_3760,N_2989,N_2389);
xor U3761 (N_3761,N_2266,N_2700);
or U3762 (N_3762,N_2796,N_2653);
nor U3763 (N_3763,N_2344,N_2503);
nand U3764 (N_3764,N_2663,N_2323);
xnor U3765 (N_3765,N_2612,N_2846);
nor U3766 (N_3766,N_2931,N_2238);
or U3767 (N_3767,N_2391,N_2196);
xor U3768 (N_3768,N_2424,N_2471);
or U3769 (N_3769,N_2694,N_2781);
xor U3770 (N_3770,N_2519,N_2804);
nor U3771 (N_3771,N_2123,N_2795);
nand U3772 (N_3772,N_2377,N_2875);
or U3773 (N_3773,N_2146,N_2802);
nand U3774 (N_3774,N_2338,N_2248);
xor U3775 (N_3775,N_2601,N_2370);
nand U3776 (N_3776,N_2874,N_2272);
and U3777 (N_3777,N_2003,N_2512);
or U3778 (N_3778,N_2891,N_2791);
nor U3779 (N_3779,N_2350,N_2508);
nand U3780 (N_3780,N_2875,N_2743);
nor U3781 (N_3781,N_2466,N_2099);
nand U3782 (N_3782,N_2451,N_2341);
and U3783 (N_3783,N_2965,N_2425);
xor U3784 (N_3784,N_2152,N_2970);
nor U3785 (N_3785,N_2870,N_2480);
nand U3786 (N_3786,N_2087,N_2786);
and U3787 (N_3787,N_2531,N_2522);
xor U3788 (N_3788,N_2528,N_2920);
xor U3789 (N_3789,N_2476,N_2502);
xnor U3790 (N_3790,N_2568,N_2926);
xnor U3791 (N_3791,N_2962,N_2910);
nor U3792 (N_3792,N_2718,N_2668);
xnor U3793 (N_3793,N_2693,N_2400);
xor U3794 (N_3794,N_2075,N_2725);
or U3795 (N_3795,N_2640,N_2454);
nand U3796 (N_3796,N_2322,N_2434);
nor U3797 (N_3797,N_2236,N_2957);
and U3798 (N_3798,N_2766,N_2027);
and U3799 (N_3799,N_2406,N_2878);
nand U3800 (N_3800,N_2633,N_2690);
nor U3801 (N_3801,N_2493,N_2672);
and U3802 (N_3802,N_2531,N_2962);
or U3803 (N_3803,N_2860,N_2240);
xor U3804 (N_3804,N_2875,N_2272);
nor U3805 (N_3805,N_2303,N_2341);
or U3806 (N_3806,N_2610,N_2591);
nor U3807 (N_3807,N_2584,N_2249);
and U3808 (N_3808,N_2415,N_2414);
nand U3809 (N_3809,N_2081,N_2594);
xnor U3810 (N_3810,N_2344,N_2856);
or U3811 (N_3811,N_2987,N_2518);
or U3812 (N_3812,N_2372,N_2913);
nand U3813 (N_3813,N_2422,N_2953);
xnor U3814 (N_3814,N_2838,N_2334);
nand U3815 (N_3815,N_2996,N_2376);
nor U3816 (N_3816,N_2517,N_2449);
or U3817 (N_3817,N_2755,N_2323);
xnor U3818 (N_3818,N_2851,N_2948);
nand U3819 (N_3819,N_2104,N_2649);
or U3820 (N_3820,N_2475,N_2366);
and U3821 (N_3821,N_2481,N_2435);
nor U3822 (N_3822,N_2930,N_2418);
nand U3823 (N_3823,N_2294,N_2496);
or U3824 (N_3824,N_2873,N_2621);
nor U3825 (N_3825,N_2212,N_2935);
nor U3826 (N_3826,N_2607,N_2217);
xnor U3827 (N_3827,N_2061,N_2341);
xnor U3828 (N_3828,N_2723,N_2830);
xnor U3829 (N_3829,N_2886,N_2169);
xor U3830 (N_3830,N_2120,N_2444);
nor U3831 (N_3831,N_2623,N_2947);
and U3832 (N_3832,N_2071,N_2068);
nand U3833 (N_3833,N_2119,N_2538);
nor U3834 (N_3834,N_2634,N_2867);
nand U3835 (N_3835,N_2426,N_2304);
and U3836 (N_3836,N_2208,N_2624);
nand U3837 (N_3837,N_2604,N_2569);
and U3838 (N_3838,N_2640,N_2380);
or U3839 (N_3839,N_2748,N_2893);
nand U3840 (N_3840,N_2158,N_2008);
or U3841 (N_3841,N_2540,N_2168);
nand U3842 (N_3842,N_2179,N_2483);
xor U3843 (N_3843,N_2881,N_2154);
nor U3844 (N_3844,N_2941,N_2601);
nor U3845 (N_3845,N_2573,N_2241);
or U3846 (N_3846,N_2196,N_2057);
xor U3847 (N_3847,N_2820,N_2231);
nor U3848 (N_3848,N_2980,N_2519);
nand U3849 (N_3849,N_2581,N_2549);
xor U3850 (N_3850,N_2781,N_2501);
xor U3851 (N_3851,N_2534,N_2682);
and U3852 (N_3852,N_2825,N_2278);
nand U3853 (N_3853,N_2944,N_2095);
nand U3854 (N_3854,N_2119,N_2392);
nor U3855 (N_3855,N_2499,N_2767);
nand U3856 (N_3856,N_2320,N_2743);
nand U3857 (N_3857,N_2909,N_2457);
nand U3858 (N_3858,N_2688,N_2234);
or U3859 (N_3859,N_2143,N_2788);
nor U3860 (N_3860,N_2667,N_2115);
nor U3861 (N_3861,N_2576,N_2850);
xnor U3862 (N_3862,N_2156,N_2256);
or U3863 (N_3863,N_2659,N_2039);
xor U3864 (N_3864,N_2473,N_2930);
and U3865 (N_3865,N_2273,N_2433);
and U3866 (N_3866,N_2428,N_2040);
xnor U3867 (N_3867,N_2514,N_2300);
or U3868 (N_3868,N_2516,N_2022);
nand U3869 (N_3869,N_2436,N_2221);
nand U3870 (N_3870,N_2848,N_2678);
and U3871 (N_3871,N_2014,N_2725);
xnor U3872 (N_3872,N_2355,N_2703);
or U3873 (N_3873,N_2781,N_2159);
xor U3874 (N_3874,N_2200,N_2363);
nor U3875 (N_3875,N_2129,N_2258);
nand U3876 (N_3876,N_2045,N_2282);
and U3877 (N_3877,N_2285,N_2973);
and U3878 (N_3878,N_2605,N_2488);
xnor U3879 (N_3879,N_2691,N_2904);
nor U3880 (N_3880,N_2946,N_2717);
or U3881 (N_3881,N_2519,N_2329);
and U3882 (N_3882,N_2628,N_2938);
or U3883 (N_3883,N_2047,N_2491);
and U3884 (N_3884,N_2834,N_2341);
xnor U3885 (N_3885,N_2513,N_2844);
or U3886 (N_3886,N_2210,N_2036);
nand U3887 (N_3887,N_2216,N_2128);
or U3888 (N_3888,N_2625,N_2298);
nor U3889 (N_3889,N_2217,N_2689);
and U3890 (N_3890,N_2831,N_2512);
or U3891 (N_3891,N_2022,N_2050);
xnor U3892 (N_3892,N_2757,N_2735);
xor U3893 (N_3893,N_2511,N_2150);
and U3894 (N_3894,N_2687,N_2772);
and U3895 (N_3895,N_2355,N_2487);
nor U3896 (N_3896,N_2034,N_2821);
nor U3897 (N_3897,N_2712,N_2608);
and U3898 (N_3898,N_2545,N_2754);
or U3899 (N_3899,N_2095,N_2006);
nand U3900 (N_3900,N_2237,N_2988);
nor U3901 (N_3901,N_2089,N_2297);
nor U3902 (N_3902,N_2133,N_2237);
or U3903 (N_3903,N_2180,N_2306);
nor U3904 (N_3904,N_2798,N_2478);
and U3905 (N_3905,N_2417,N_2845);
and U3906 (N_3906,N_2244,N_2111);
nor U3907 (N_3907,N_2865,N_2849);
nand U3908 (N_3908,N_2860,N_2357);
nor U3909 (N_3909,N_2461,N_2205);
nand U3910 (N_3910,N_2200,N_2805);
or U3911 (N_3911,N_2472,N_2963);
nand U3912 (N_3912,N_2455,N_2468);
and U3913 (N_3913,N_2790,N_2294);
nand U3914 (N_3914,N_2700,N_2766);
nand U3915 (N_3915,N_2100,N_2332);
nand U3916 (N_3916,N_2836,N_2609);
nand U3917 (N_3917,N_2028,N_2860);
nor U3918 (N_3918,N_2891,N_2916);
or U3919 (N_3919,N_2650,N_2939);
nand U3920 (N_3920,N_2705,N_2172);
nand U3921 (N_3921,N_2040,N_2579);
nand U3922 (N_3922,N_2281,N_2444);
and U3923 (N_3923,N_2803,N_2341);
nor U3924 (N_3924,N_2143,N_2833);
and U3925 (N_3925,N_2985,N_2989);
xnor U3926 (N_3926,N_2976,N_2130);
xor U3927 (N_3927,N_2536,N_2907);
and U3928 (N_3928,N_2948,N_2320);
or U3929 (N_3929,N_2587,N_2835);
xor U3930 (N_3930,N_2904,N_2736);
nor U3931 (N_3931,N_2132,N_2832);
or U3932 (N_3932,N_2095,N_2715);
nand U3933 (N_3933,N_2610,N_2287);
xnor U3934 (N_3934,N_2784,N_2894);
xor U3935 (N_3935,N_2584,N_2972);
or U3936 (N_3936,N_2842,N_2642);
xnor U3937 (N_3937,N_2230,N_2361);
nor U3938 (N_3938,N_2721,N_2895);
and U3939 (N_3939,N_2689,N_2426);
nand U3940 (N_3940,N_2399,N_2245);
xnor U3941 (N_3941,N_2530,N_2650);
or U3942 (N_3942,N_2393,N_2930);
and U3943 (N_3943,N_2928,N_2771);
and U3944 (N_3944,N_2482,N_2463);
nand U3945 (N_3945,N_2141,N_2737);
xnor U3946 (N_3946,N_2312,N_2303);
or U3947 (N_3947,N_2924,N_2494);
or U3948 (N_3948,N_2048,N_2709);
xor U3949 (N_3949,N_2486,N_2069);
nand U3950 (N_3950,N_2913,N_2016);
xnor U3951 (N_3951,N_2679,N_2485);
xor U3952 (N_3952,N_2083,N_2377);
nor U3953 (N_3953,N_2733,N_2679);
nand U3954 (N_3954,N_2404,N_2411);
xnor U3955 (N_3955,N_2166,N_2629);
xor U3956 (N_3956,N_2688,N_2108);
nand U3957 (N_3957,N_2820,N_2361);
and U3958 (N_3958,N_2098,N_2606);
xnor U3959 (N_3959,N_2524,N_2049);
or U3960 (N_3960,N_2817,N_2643);
or U3961 (N_3961,N_2782,N_2017);
xnor U3962 (N_3962,N_2934,N_2463);
xor U3963 (N_3963,N_2105,N_2700);
nor U3964 (N_3964,N_2492,N_2355);
or U3965 (N_3965,N_2447,N_2615);
or U3966 (N_3966,N_2081,N_2778);
nor U3967 (N_3967,N_2798,N_2891);
nand U3968 (N_3968,N_2717,N_2172);
or U3969 (N_3969,N_2191,N_2198);
xnor U3970 (N_3970,N_2481,N_2866);
nand U3971 (N_3971,N_2529,N_2637);
xnor U3972 (N_3972,N_2028,N_2867);
or U3973 (N_3973,N_2871,N_2693);
xnor U3974 (N_3974,N_2866,N_2881);
and U3975 (N_3975,N_2317,N_2476);
xnor U3976 (N_3976,N_2304,N_2707);
or U3977 (N_3977,N_2333,N_2020);
nor U3978 (N_3978,N_2711,N_2646);
or U3979 (N_3979,N_2100,N_2643);
nand U3980 (N_3980,N_2810,N_2498);
and U3981 (N_3981,N_2622,N_2168);
nor U3982 (N_3982,N_2938,N_2896);
nand U3983 (N_3983,N_2642,N_2228);
or U3984 (N_3984,N_2427,N_2596);
xor U3985 (N_3985,N_2798,N_2405);
nor U3986 (N_3986,N_2069,N_2317);
xor U3987 (N_3987,N_2778,N_2367);
nor U3988 (N_3988,N_2263,N_2508);
and U3989 (N_3989,N_2290,N_2675);
xor U3990 (N_3990,N_2907,N_2353);
nor U3991 (N_3991,N_2293,N_2143);
nand U3992 (N_3992,N_2738,N_2674);
or U3993 (N_3993,N_2803,N_2113);
and U3994 (N_3994,N_2231,N_2833);
or U3995 (N_3995,N_2541,N_2628);
and U3996 (N_3996,N_2797,N_2285);
and U3997 (N_3997,N_2192,N_2028);
nand U3998 (N_3998,N_2591,N_2942);
and U3999 (N_3999,N_2872,N_2052);
nor U4000 (N_4000,N_3497,N_3671);
and U4001 (N_4001,N_3188,N_3776);
nor U4002 (N_4002,N_3589,N_3768);
or U4003 (N_4003,N_3753,N_3332);
or U4004 (N_4004,N_3216,N_3068);
nor U4005 (N_4005,N_3949,N_3160);
and U4006 (N_4006,N_3979,N_3205);
nor U4007 (N_4007,N_3839,N_3481);
xor U4008 (N_4008,N_3941,N_3348);
nand U4009 (N_4009,N_3178,N_3569);
nor U4010 (N_4010,N_3455,N_3451);
nand U4011 (N_4011,N_3807,N_3651);
xnor U4012 (N_4012,N_3211,N_3145);
or U4013 (N_4013,N_3608,N_3822);
nand U4014 (N_4014,N_3241,N_3648);
xor U4015 (N_4015,N_3152,N_3040);
nand U4016 (N_4016,N_3620,N_3889);
and U4017 (N_4017,N_3149,N_3028);
nor U4018 (N_4018,N_3502,N_3645);
nand U4019 (N_4019,N_3765,N_3408);
nand U4020 (N_4020,N_3952,N_3225);
and U4021 (N_4021,N_3245,N_3985);
nand U4022 (N_4022,N_3132,N_3126);
nand U4023 (N_4023,N_3975,N_3785);
nand U4024 (N_4024,N_3486,N_3454);
nor U4025 (N_4025,N_3082,N_3505);
xor U4026 (N_4026,N_3668,N_3107);
xor U4027 (N_4027,N_3311,N_3067);
or U4028 (N_4028,N_3223,N_3854);
nand U4029 (N_4029,N_3744,N_3898);
xor U4030 (N_4030,N_3037,N_3795);
nand U4031 (N_4031,N_3432,N_3324);
and U4032 (N_4032,N_3006,N_3970);
nand U4033 (N_4033,N_3009,N_3075);
or U4034 (N_4034,N_3129,N_3182);
nor U4035 (N_4035,N_3409,N_3704);
nand U4036 (N_4036,N_3196,N_3088);
nor U4037 (N_4037,N_3260,N_3147);
xnor U4038 (N_4038,N_3515,N_3279);
or U4039 (N_4039,N_3108,N_3294);
xor U4040 (N_4040,N_3352,N_3389);
or U4041 (N_4041,N_3093,N_3708);
nor U4042 (N_4042,N_3681,N_3884);
and U4043 (N_4043,N_3299,N_3042);
nand U4044 (N_4044,N_3215,N_3456);
nor U4045 (N_4045,N_3619,N_3894);
or U4046 (N_4046,N_3287,N_3934);
xor U4047 (N_4047,N_3853,N_3448);
xor U4048 (N_4048,N_3010,N_3468);
nand U4049 (N_4049,N_3832,N_3046);
nor U4050 (N_4050,N_3122,N_3403);
and U4051 (N_4051,N_3254,N_3269);
nor U4052 (N_4052,N_3405,N_3531);
nand U4053 (N_4053,N_3388,N_3435);
nor U4054 (N_4054,N_3943,N_3399);
and U4055 (N_4055,N_3396,N_3304);
or U4056 (N_4056,N_3752,N_3238);
xor U4057 (N_4057,N_3746,N_3772);
nand U4058 (N_4058,N_3715,N_3001);
and U4059 (N_4059,N_3394,N_3367);
nand U4060 (N_4060,N_3778,N_3242);
nor U4061 (N_4061,N_3354,N_3818);
and U4062 (N_4062,N_3197,N_3100);
nand U4063 (N_4063,N_3901,N_3802);
or U4064 (N_4064,N_3548,N_3165);
nand U4065 (N_4065,N_3053,N_3076);
nor U4066 (N_4066,N_3113,N_3727);
xor U4067 (N_4067,N_3098,N_3106);
nor U4068 (N_4068,N_3919,N_3218);
xnor U4069 (N_4069,N_3317,N_3912);
nor U4070 (N_4070,N_3891,N_3118);
xnor U4071 (N_4071,N_3123,N_3071);
or U4072 (N_4072,N_3929,N_3667);
nor U4073 (N_4073,N_3699,N_3716);
nand U4074 (N_4074,N_3390,N_3618);
nor U4075 (N_4075,N_3236,N_3757);
xor U4076 (N_4076,N_3641,N_3433);
xor U4077 (N_4077,N_3494,N_3957);
nand U4078 (N_4078,N_3411,N_3457);
nor U4079 (N_4079,N_3315,N_3379);
nand U4080 (N_4080,N_3984,N_3686);
nand U4081 (N_4081,N_3282,N_3909);
nor U4082 (N_4082,N_3942,N_3692);
or U4083 (N_4083,N_3110,N_3518);
or U4084 (N_4084,N_3714,N_3597);
or U4085 (N_4085,N_3265,N_3339);
nor U4086 (N_4086,N_3888,N_3077);
nor U4087 (N_4087,N_3228,N_3740);
nand U4088 (N_4088,N_3356,N_3639);
nor U4089 (N_4089,N_3091,N_3138);
or U4090 (N_4090,N_3207,N_3580);
and U4091 (N_4091,N_3950,N_3120);
or U4092 (N_4092,N_3463,N_3925);
xnor U4093 (N_4093,N_3532,N_3217);
nand U4094 (N_4094,N_3858,N_3425);
nor U4095 (N_4095,N_3192,N_3868);
nand U4096 (N_4096,N_3094,N_3991);
or U4097 (N_4097,N_3964,N_3939);
and U4098 (N_4098,N_3141,N_3176);
xnor U4099 (N_4099,N_3109,N_3840);
and U4100 (N_4100,N_3755,N_3285);
and U4101 (N_4101,N_3137,N_3688);
xor U4102 (N_4102,N_3475,N_3173);
or U4103 (N_4103,N_3292,N_3836);
nor U4104 (N_4104,N_3660,N_3200);
nand U4105 (N_4105,N_3927,N_3575);
xnor U4106 (N_4106,N_3658,N_3695);
and U4107 (N_4107,N_3250,N_3751);
nand U4108 (N_4108,N_3310,N_3599);
and U4109 (N_4109,N_3896,N_3848);
or U4110 (N_4110,N_3972,N_3421);
nor U4111 (N_4111,N_3366,N_3144);
nand U4112 (N_4112,N_3773,N_3321);
nor U4113 (N_4113,N_3874,N_3043);
nand U4114 (N_4114,N_3125,N_3789);
nand U4115 (N_4115,N_3978,N_3210);
and U4116 (N_4116,N_3442,N_3737);
or U4117 (N_4117,N_3032,N_3541);
and U4118 (N_4118,N_3903,N_3081);
nand U4119 (N_4119,N_3437,N_3257);
or U4120 (N_4120,N_3290,N_3627);
nand U4121 (N_4121,N_3872,N_3607);
or U4122 (N_4122,N_3582,N_3664);
and U4123 (N_4123,N_3466,N_3823);
xnor U4124 (N_4124,N_3092,N_3229);
nor U4125 (N_4125,N_3097,N_3027);
or U4126 (N_4126,N_3361,N_3696);
nand U4127 (N_4127,N_3380,N_3048);
xor U4128 (N_4128,N_3499,N_3246);
or U4129 (N_4129,N_3343,N_3169);
nor U4130 (N_4130,N_3382,N_3997);
nand U4131 (N_4131,N_3490,N_3560);
nor U4132 (N_4132,N_3272,N_3512);
xor U4133 (N_4133,N_3924,N_3819);
or U4134 (N_4134,N_3312,N_3146);
or U4135 (N_4135,N_3498,N_3710);
nand U4136 (N_4136,N_3665,N_3923);
and U4137 (N_4137,N_3522,N_3351);
or U4138 (N_4138,N_3980,N_3690);
nor U4139 (N_4139,N_3221,N_3488);
nor U4140 (N_4140,N_3801,N_3038);
nor U4141 (N_4141,N_3025,N_3018);
nor U4142 (N_4142,N_3732,N_3669);
or U4143 (N_4143,N_3763,N_3267);
xor U4144 (N_4144,N_3637,N_3111);
nor U4145 (N_4145,N_3759,N_3820);
nor U4146 (N_4146,N_3434,N_3600);
nor U4147 (N_4147,N_3673,N_3349);
nor U4148 (N_4148,N_3771,N_3917);
nor U4149 (N_4149,N_3328,N_3535);
nor U4150 (N_4150,N_3712,N_3206);
xnor U4151 (N_4151,N_3322,N_3213);
and U4152 (N_4152,N_3609,N_3309);
nand U4153 (N_4153,N_3058,N_3799);
and U4154 (N_4154,N_3817,N_3266);
nand U4155 (N_4155,N_3882,N_3844);
nand U4156 (N_4156,N_3195,N_3446);
and U4157 (N_4157,N_3632,N_3362);
and U4158 (N_4158,N_3656,N_3533);
and U4159 (N_4159,N_3417,N_3056);
xor U4160 (N_4160,N_3798,N_3705);
nor U4161 (N_4161,N_3181,N_3766);
xnor U4162 (N_4162,N_3459,N_3041);
nand U4163 (N_4163,N_3509,N_3302);
nand U4164 (N_4164,N_3143,N_3371);
nand U4165 (N_4165,N_3430,N_3833);
or U4166 (N_4166,N_3275,N_3030);
nor U4167 (N_4167,N_3150,N_3930);
or U4168 (N_4168,N_3625,N_3724);
xor U4169 (N_4169,N_3177,N_3954);
xor U4170 (N_4170,N_3372,N_3480);
xor U4171 (N_4171,N_3958,N_3020);
nor U4172 (N_4172,N_3662,N_3513);
nand U4173 (N_4173,N_3762,N_3545);
nor U4174 (N_4174,N_3635,N_3406);
and U4175 (N_4175,N_3326,N_3174);
nand U4176 (N_4176,N_3615,N_3014);
and U4177 (N_4177,N_3557,N_3186);
or U4178 (N_4178,N_3460,N_3825);
xnor U4179 (N_4179,N_3171,N_3105);
nand U4180 (N_4180,N_3815,N_3910);
nor U4181 (N_4181,N_3377,N_3418);
xor U4182 (N_4182,N_3095,N_3445);
xnor U4183 (N_4183,N_3654,N_3947);
nor U4184 (N_4184,N_3689,N_3555);
xnor U4185 (N_4185,N_3059,N_3065);
xor U4186 (N_4186,N_3846,N_3087);
and U4187 (N_4187,N_3374,N_3342);
xnor U4188 (N_4188,N_3938,N_3567);
nor U4189 (N_4189,N_3426,N_3702);
nand U4190 (N_4190,N_3598,N_3892);
nor U4191 (N_4191,N_3542,N_3646);
and U4192 (N_4192,N_3274,N_3543);
nor U4193 (N_4193,N_3537,N_3993);
xor U4194 (N_4194,N_3167,N_3251);
xor U4195 (N_4195,N_3538,N_3381);
or U4196 (N_4196,N_3162,N_3968);
nand U4197 (N_4197,N_3774,N_3792);
xnor U4198 (N_4198,N_3517,N_3860);
nand U4199 (N_4199,N_3099,N_3491);
and U4200 (N_4200,N_3239,N_3590);
and U4201 (N_4201,N_3298,N_3603);
nand U4202 (N_4202,N_3526,N_3775);
nand U4203 (N_4203,N_3592,N_3742);
and U4204 (N_4204,N_3002,N_3011);
and U4205 (N_4205,N_3295,N_3866);
nand U4206 (N_4206,N_3156,N_3423);
or U4207 (N_4207,N_3300,N_3139);
nand U4208 (N_4208,N_3837,N_3035);
nand U4209 (N_4209,N_3482,N_3358);
or U4210 (N_4210,N_3754,N_3350);
nor U4211 (N_4211,N_3029,N_3741);
nor U4212 (N_4212,N_3489,N_3333);
or U4213 (N_4213,N_3931,N_3700);
or U4214 (N_4214,N_3697,N_3331);
or U4215 (N_4215,N_3487,N_3520);
and U4216 (N_4216,N_3222,N_3805);
and U4217 (N_4217,N_3201,N_3220);
nor U4218 (N_4218,N_3624,N_3248);
and U4219 (N_4219,N_3391,N_3899);
nor U4220 (N_4220,N_3325,N_3826);
nor U4221 (N_4221,N_3202,N_3887);
nor U4222 (N_4222,N_3360,N_3895);
or U4223 (N_4223,N_3297,N_3440);
nor U4224 (N_4224,N_3786,N_3303);
and U4225 (N_4225,N_3187,N_3640);
nor U4226 (N_4226,N_3429,N_3679);
and U4227 (N_4227,N_3231,N_3190);
nor U4228 (N_4228,N_3676,N_3469);
and U4229 (N_4229,N_3074,N_3008);
xnor U4230 (N_4230,N_3255,N_3227);
xnor U4231 (N_4231,N_3530,N_3722);
nand U4232 (N_4232,N_3133,N_3472);
and U4233 (N_4233,N_3605,N_3036);
nand U4234 (N_4234,N_3990,N_3155);
and U4235 (N_4235,N_3470,N_3511);
or U4236 (N_4236,N_3316,N_3586);
nor U4237 (N_4237,N_3687,N_3516);
nor U4238 (N_4238,N_3612,N_3063);
nor U4239 (N_4239,N_3674,N_3631);
nand U4240 (N_4240,N_3698,N_3412);
and U4241 (N_4241,N_3988,N_3571);
or U4242 (N_4242,N_3277,N_3034);
nand U4243 (N_4243,N_3420,N_3359);
and U4244 (N_4244,N_3334,N_3747);
nand U4245 (N_4245,N_3050,N_3284);
nand U4246 (N_4246,N_3636,N_3527);
xnor U4247 (N_4247,N_3718,N_3345);
nand U4248 (N_4248,N_3999,N_3525);
and U4249 (N_4249,N_3682,N_3208);
nand U4250 (N_4250,N_3004,N_3280);
and U4251 (N_4251,N_3613,N_3314);
nor U4252 (N_4252,N_3344,N_3655);
nor U4253 (N_4253,N_3606,N_3449);
xnor U4254 (N_4254,N_3249,N_3552);
or U4255 (N_4255,N_3928,N_3305);
or U4256 (N_4256,N_3383,N_3989);
nand U4257 (N_4257,N_3761,N_3869);
xor U4258 (N_4258,N_3581,N_3738);
or U4259 (N_4259,N_3735,N_3831);
or U4260 (N_4260,N_3871,N_3961);
or U4261 (N_4261,N_3769,N_3337);
xnor U4262 (N_4262,N_3528,N_3852);
nor U4263 (N_4263,N_3570,N_3378);
or U4264 (N_4264,N_3666,N_3749);
nand U4265 (N_4265,N_3493,N_3393);
nor U4266 (N_4266,N_3680,N_3812);
xor U4267 (N_4267,N_3725,N_3386);
and U4268 (N_4268,N_3783,N_3397);
xor U4269 (N_4269,N_3524,N_3628);
nor U4270 (N_4270,N_3047,N_3083);
nand U4271 (N_4271,N_3998,N_3838);
nor U4272 (N_4272,N_3370,N_3264);
or U4273 (N_4273,N_3614,N_3610);
nand U4274 (N_4274,N_3638,N_3758);
nor U4275 (N_4275,N_3547,N_3562);
or U4276 (N_4276,N_3085,N_3153);
nand U4277 (N_4277,N_3551,N_3353);
nand U4278 (N_4278,N_3230,N_3368);
and U4279 (N_4279,N_3994,N_3670);
nor U4280 (N_4280,N_3583,N_3920);
or U4281 (N_4281,N_3711,N_3478);
or U4282 (N_4282,N_3946,N_3070);
or U4283 (N_4283,N_3276,N_3566);
and U4284 (N_4284,N_3116,N_3955);
or U4285 (N_4285,N_3723,N_3849);
or U4286 (N_4286,N_3626,N_3452);
xnor U4287 (N_4287,N_3835,N_3616);
nand U4288 (N_4288,N_3387,N_3080);
and U4289 (N_4289,N_3507,N_3465);
or U4290 (N_4290,N_3788,N_3154);
nand U4291 (N_4291,N_3338,N_3963);
nand U4292 (N_4292,N_3734,N_3701);
xor U4293 (N_4293,N_3096,N_3444);
nor U4294 (N_4294,N_3707,N_3184);
or U4295 (N_4295,N_3536,N_3506);
nor U4296 (N_4296,N_3007,N_3045);
xor U4297 (N_4297,N_3862,N_3293);
or U4298 (N_4298,N_3436,N_3890);
nand U4299 (N_4299,N_3384,N_3717);
or U4300 (N_4300,N_3851,N_3720);
nor U4301 (N_4301,N_3336,N_3739);
nor U4302 (N_4302,N_3289,N_3424);
and U4303 (N_4303,N_3703,N_3128);
xor U4304 (N_4304,N_3464,N_3878);
nor U4305 (N_4305,N_3604,N_3811);
or U4306 (N_4306,N_3797,N_3024);
nor U4307 (N_4307,N_3209,N_3573);
or U4308 (N_4308,N_3031,N_3049);
and U4309 (N_4309,N_3810,N_3951);
or U4310 (N_4310,N_3484,N_3185);
or U4311 (N_4311,N_3678,N_3905);
and U4312 (N_4312,N_3226,N_3079);
nand U4313 (N_4313,N_3164,N_3170);
xor U4314 (N_4314,N_3234,N_3623);
xnor U4315 (N_4315,N_3373,N_3501);
or U4316 (N_4316,N_3427,N_3115);
xor U4317 (N_4317,N_3659,N_3602);
or U4318 (N_4318,N_3830,N_3175);
nand U4319 (N_4319,N_3796,N_3503);
or U4320 (N_4320,N_3987,N_3861);
xnor U4321 (N_4321,N_3915,N_3911);
nor U4322 (N_4322,N_3719,N_3307);
or U4323 (N_4323,N_3415,N_3845);
xnor U4324 (N_4324,N_3219,N_3346);
or U4325 (N_4325,N_3885,N_3240);
nand U4326 (N_4326,N_3780,N_3431);
or U4327 (N_4327,N_3847,N_3458);
xnor U4328 (N_4328,N_3060,N_3453);
xor U4329 (N_4329,N_3233,N_3232);
or U4330 (N_4330,N_3398,N_3114);
and U4331 (N_4331,N_3330,N_3450);
and U4332 (N_4332,N_3086,N_3496);
or U4333 (N_4333,N_3318,N_3395);
xor U4334 (N_4334,N_3824,N_3023);
and U4335 (N_4335,N_3301,N_3565);
nand U4336 (N_4336,N_3743,N_3568);
xnor U4337 (N_4337,N_3881,N_3617);
and U4338 (N_4338,N_3561,N_3601);
xnor U4339 (N_4339,N_3514,N_3995);
nand U4340 (N_4340,N_3012,N_3474);
and U4341 (N_4341,N_3564,N_3584);
nor U4342 (N_4342,N_3808,N_3119);
nor U4343 (N_4343,N_3033,N_3856);
nor U4344 (N_4344,N_3966,N_3981);
xnor U4345 (N_4345,N_3706,N_3691);
nand U4346 (N_4346,N_3694,N_3183);
nor U4347 (N_4347,N_3558,N_3323);
nor U4348 (N_4348,N_3319,N_3404);
nor U4349 (N_4349,N_3244,N_3504);
and U4350 (N_4350,N_3843,N_3713);
xor U4351 (N_4351,N_3278,N_3880);
nor U4352 (N_4352,N_3320,N_3883);
or U4353 (N_4353,N_3015,N_3829);
nor U4354 (N_4354,N_3363,N_3685);
or U4355 (N_4355,N_3959,N_3926);
and U4356 (N_4356,N_3574,N_3657);
nand U4357 (N_4357,N_3933,N_3945);
and U4358 (N_4358,N_3893,N_3629);
nor U4359 (N_4359,N_3967,N_3179);
xor U4360 (N_4360,N_3414,N_3992);
nor U4361 (N_4361,N_3976,N_3633);
xor U4362 (N_4362,N_3977,N_3039);
and U4363 (N_4363,N_3485,N_3443);
or U4364 (N_4364,N_3313,N_3864);
xnor U4365 (N_4365,N_3365,N_3283);
xor U4366 (N_4366,N_3983,N_3168);
xor U4367 (N_4367,N_3510,N_3103);
or U4368 (N_4368,N_3212,N_3180);
and U4369 (N_4369,N_3587,N_3407);
or U4370 (N_4370,N_3112,N_3729);
nand U4371 (N_4371,N_3529,N_3794);
and U4372 (N_4372,N_3828,N_3935);
nor U4373 (N_4373,N_3906,N_3044);
or U4374 (N_4374,N_3090,N_3982);
xor U4375 (N_4375,N_3288,N_3948);
xor U4376 (N_4376,N_3495,N_3721);
or U4377 (N_4377,N_3973,N_3483);
or U4378 (N_4378,N_3447,N_3733);
nand U4379 (N_4379,N_3770,N_3335);
or U4380 (N_4380,N_3140,N_3588);
nor U4381 (N_4381,N_3369,N_3726);
xnor U4382 (N_4382,N_3261,N_3523);
nor U4383 (N_4383,N_3579,N_3142);
nor U4384 (N_4384,N_3539,N_3055);
xnor U4385 (N_4385,N_3492,N_3413);
nand U4386 (N_4386,N_3062,N_3821);
xor U4387 (N_4387,N_3634,N_3017);
and U4388 (N_4388,N_3867,N_3953);
or U4389 (N_4389,N_3003,N_3902);
or U4390 (N_4390,N_3401,N_3827);
nand U4391 (N_4391,N_3736,N_3791);
or U4392 (N_4392,N_3462,N_3556);
nand U4393 (N_4393,N_3476,N_3730);
and U4394 (N_4394,N_3341,N_3376);
and U4395 (N_4395,N_3422,N_3760);
and U4396 (N_4396,N_3130,N_3932);
or U4397 (N_4397,N_3577,N_3019);
and U4398 (N_4398,N_3675,N_3653);
and U4399 (N_4399,N_3649,N_3784);
and U4400 (N_4400,N_3937,N_3131);
xor U4401 (N_4401,N_3611,N_3875);
and U4402 (N_4402,N_3803,N_3806);
and U4403 (N_4403,N_3163,N_3916);
xor U4404 (N_4404,N_3273,N_3064);
xnor U4405 (N_4405,N_3809,N_3642);
nand U4406 (N_4406,N_3364,N_3270);
nor U4407 (N_4407,N_3259,N_3559);
nand U4408 (N_4408,N_3750,N_3135);
nor U4409 (N_4409,N_3340,N_3199);
nor U4410 (N_4410,N_3473,N_3268);
xnor U4411 (N_4411,N_3622,N_3439);
nand U4412 (N_4412,N_3385,N_3936);
or U4413 (N_4413,N_3907,N_3479);
xor U4414 (N_4414,N_3237,N_3777);
nor U4415 (N_4415,N_3329,N_3879);
and U4416 (N_4416,N_3419,N_3519);
nor U4417 (N_4417,N_3652,N_3804);
or U4418 (N_4418,N_3089,N_3918);
or U4419 (N_4419,N_3005,N_3148);
nor U4420 (N_4420,N_3521,N_3863);
and U4421 (N_4421,N_3572,N_3247);
xnor U4422 (N_4422,N_3101,N_3072);
nand U4423 (N_4423,N_3235,N_3800);
xor U4424 (N_4424,N_3986,N_3327);
or U4425 (N_4425,N_3286,N_3576);
or U4426 (N_4426,N_3940,N_3243);
xnor U4427 (N_4427,N_3962,N_3084);
and U4428 (N_4428,N_3203,N_3016);
or U4429 (N_4429,N_3728,N_3855);
nor U4430 (N_4430,N_3540,N_3136);
nand U4431 (N_4431,N_3224,N_3793);
nand U4432 (N_4432,N_3416,N_3172);
nand U4433 (N_4433,N_3271,N_3544);
xnor U4434 (N_4434,N_3886,N_3392);
nand U4435 (N_4435,N_3355,N_3159);
xnor U4436 (N_4436,N_3870,N_3709);
nand U4437 (N_4437,N_3308,N_3585);
nor U4438 (N_4438,N_3263,N_3441);
or U4439 (N_4439,N_3960,N_3508);
and U4440 (N_4440,N_3438,N_3000);
or U4441 (N_4441,N_3914,N_3121);
nor U4442 (N_4442,N_3252,N_3296);
nor U4443 (N_4443,N_3974,N_3921);
or U4444 (N_4444,N_3781,N_3051);
nor U4445 (N_4445,N_3683,N_3198);
xor U4446 (N_4446,N_3134,N_3281);
xor U4447 (N_4447,N_3873,N_3661);
nor U4448 (N_4448,N_3104,N_3814);
nor U4449 (N_4449,N_3073,N_3779);
nor U4450 (N_4450,N_3102,N_3850);
or U4451 (N_4451,N_3054,N_3865);
xnor U4452 (N_4452,N_3262,N_3677);
nand U4453 (N_4453,N_3347,N_3022);
xor U4454 (N_4454,N_3402,N_3593);
xor U4455 (N_4455,N_3428,N_3834);
nor U4456 (N_4456,N_3859,N_3256);
xnor U4457 (N_4457,N_3790,N_3066);
or U4458 (N_4458,N_3553,N_3944);
and U4459 (N_4459,N_3117,N_3647);
nor U4460 (N_4460,N_3971,N_3375);
nor U4461 (N_4461,N_3069,N_3877);
xor U4462 (N_4462,N_3596,N_3052);
nor U4463 (N_4463,N_3400,N_3630);
xor U4464 (N_4464,N_3550,N_3969);
or U4465 (N_4465,N_3897,N_3693);
nor U4466 (N_4466,N_3061,N_3594);
nor U4467 (N_4467,N_3908,N_3214);
nor U4468 (N_4468,N_3684,N_3258);
xor U4469 (N_4469,N_3021,N_3151);
or U4470 (N_4470,N_3291,N_3549);
or U4471 (N_4471,N_3756,N_3078);
and U4472 (N_4472,N_3857,N_3672);
and U4473 (N_4473,N_3467,N_3748);
or U4474 (N_4474,N_3026,N_3913);
and U4475 (N_4475,N_3745,N_3767);
nand U4476 (N_4476,N_3194,N_3876);
nand U4477 (N_4477,N_3965,N_3357);
or U4478 (N_4478,N_3546,N_3731);
or U4479 (N_4479,N_3127,N_3904);
xor U4480 (N_4480,N_3841,N_3534);
xnor U4481 (N_4481,N_3410,N_3204);
xnor U4482 (N_4482,N_3500,N_3644);
xnor U4483 (N_4483,N_3471,N_3787);
nand U4484 (N_4484,N_3764,N_3663);
or U4485 (N_4485,N_3193,N_3306);
and U4486 (N_4486,N_3922,N_3621);
or U4487 (N_4487,N_3124,N_3013);
nor U4488 (N_4488,N_3253,N_3842);
xor U4489 (N_4489,N_3158,N_3189);
and U4490 (N_4490,N_3057,N_3554);
nor U4491 (N_4491,N_3900,N_3650);
nand U4492 (N_4492,N_3578,N_3166);
or U4493 (N_4493,N_3643,N_3813);
nand U4494 (N_4494,N_3161,N_3595);
nand U4495 (N_4495,N_3563,N_3956);
nor U4496 (N_4496,N_3816,N_3157);
nand U4497 (N_4497,N_3191,N_3477);
and U4498 (N_4498,N_3461,N_3996);
and U4499 (N_4499,N_3782,N_3591);
nor U4500 (N_4500,N_3076,N_3665);
nor U4501 (N_4501,N_3820,N_3591);
nor U4502 (N_4502,N_3922,N_3904);
or U4503 (N_4503,N_3466,N_3570);
and U4504 (N_4504,N_3836,N_3540);
or U4505 (N_4505,N_3810,N_3610);
xor U4506 (N_4506,N_3495,N_3586);
nand U4507 (N_4507,N_3968,N_3123);
nand U4508 (N_4508,N_3063,N_3680);
or U4509 (N_4509,N_3903,N_3189);
nor U4510 (N_4510,N_3132,N_3138);
and U4511 (N_4511,N_3160,N_3101);
or U4512 (N_4512,N_3080,N_3170);
nor U4513 (N_4513,N_3137,N_3413);
xnor U4514 (N_4514,N_3553,N_3285);
and U4515 (N_4515,N_3208,N_3578);
or U4516 (N_4516,N_3130,N_3731);
nand U4517 (N_4517,N_3023,N_3889);
nand U4518 (N_4518,N_3386,N_3157);
or U4519 (N_4519,N_3364,N_3410);
nand U4520 (N_4520,N_3445,N_3099);
nand U4521 (N_4521,N_3674,N_3700);
xor U4522 (N_4522,N_3391,N_3057);
nand U4523 (N_4523,N_3365,N_3228);
and U4524 (N_4524,N_3667,N_3836);
xor U4525 (N_4525,N_3300,N_3903);
nand U4526 (N_4526,N_3782,N_3164);
xor U4527 (N_4527,N_3781,N_3570);
nand U4528 (N_4528,N_3974,N_3911);
nand U4529 (N_4529,N_3774,N_3450);
nand U4530 (N_4530,N_3436,N_3037);
or U4531 (N_4531,N_3756,N_3582);
and U4532 (N_4532,N_3216,N_3064);
or U4533 (N_4533,N_3501,N_3508);
nor U4534 (N_4534,N_3287,N_3776);
nor U4535 (N_4535,N_3031,N_3499);
or U4536 (N_4536,N_3174,N_3199);
and U4537 (N_4537,N_3331,N_3338);
and U4538 (N_4538,N_3103,N_3701);
and U4539 (N_4539,N_3497,N_3905);
nor U4540 (N_4540,N_3506,N_3356);
xor U4541 (N_4541,N_3497,N_3359);
or U4542 (N_4542,N_3902,N_3222);
nand U4543 (N_4543,N_3560,N_3275);
xor U4544 (N_4544,N_3078,N_3638);
and U4545 (N_4545,N_3716,N_3634);
and U4546 (N_4546,N_3286,N_3392);
nand U4547 (N_4547,N_3958,N_3437);
or U4548 (N_4548,N_3684,N_3325);
and U4549 (N_4549,N_3938,N_3165);
and U4550 (N_4550,N_3261,N_3870);
and U4551 (N_4551,N_3962,N_3064);
or U4552 (N_4552,N_3300,N_3334);
and U4553 (N_4553,N_3758,N_3415);
nor U4554 (N_4554,N_3844,N_3903);
or U4555 (N_4555,N_3098,N_3005);
nand U4556 (N_4556,N_3824,N_3301);
xnor U4557 (N_4557,N_3688,N_3917);
or U4558 (N_4558,N_3286,N_3506);
nor U4559 (N_4559,N_3680,N_3321);
or U4560 (N_4560,N_3583,N_3154);
nand U4561 (N_4561,N_3212,N_3963);
nor U4562 (N_4562,N_3899,N_3002);
nor U4563 (N_4563,N_3166,N_3328);
and U4564 (N_4564,N_3802,N_3495);
and U4565 (N_4565,N_3024,N_3132);
nand U4566 (N_4566,N_3070,N_3321);
nand U4567 (N_4567,N_3233,N_3865);
and U4568 (N_4568,N_3565,N_3886);
or U4569 (N_4569,N_3571,N_3749);
xor U4570 (N_4570,N_3367,N_3760);
or U4571 (N_4571,N_3324,N_3403);
xnor U4572 (N_4572,N_3363,N_3128);
nor U4573 (N_4573,N_3890,N_3444);
and U4574 (N_4574,N_3901,N_3940);
nand U4575 (N_4575,N_3272,N_3384);
nand U4576 (N_4576,N_3343,N_3374);
nand U4577 (N_4577,N_3339,N_3904);
nand U4578 (N_4578,N_3284,N_3642);
nor U4579 (N_4579,N_3925,N_3227);
nor U4580 (N_4580,N_3360,N_3620);
nand U4581 (N_4581,N_3542,N_3236);
and U4582 (N_4582,N_3955,N_3853);
nand U4583 (N_4583,N_3996,N_3808);
and U4584 (N_4584,N_3660,N_3195);
xnor U4585 (N_4585,N_3800,N_3394);
nor U4586 (N_4586,N_3689,N_3300);
or U4587 (N_4587,N_3399,N_3717);
xor U4588 (N_4588,N_3108,N_3550);
nand U4589 (N_4589,N_3458,N_3759);
nor U4590 (N_4590,N_3667,N_3383);
nand U4591 (N_4591,N_3019,N_3413);
nand U4592 (N_4592,N_3526,N_3896);
nand U4593 (N_4593,N_3758,N_3497);
nand U4594 (N_4594,N_3315,N_3702);
or U4595 (N_4595,N_3323,N_3636);
nor U4596 (N_4596,N_3934,N_3507);
nor U4597 (N_4597,N_3312,N_3974);
or U4598 (N_4598,N_3505,N_3721);
or U4599 (N_4599,N_3744,N_3781);
nand U4600 (N_4600,N_3971,N_3735);
xor U4601 (N_4601,N_3602,N_3019);
nand U4602 (N_4602,N_3994,N_3091);
nand U4603 (N_4603,N_3507,N_3685);
nand U4604 (N_4604,N_3586,N_3075);
nor U4605 (N_4605,N_3919,N_3166);
nand U4606 (N_4606,N_3293,N_3868);
and U4607 (N_4607,N_3177,N_3447);
and U4608 (N_4608,N_3769,N_3404);
or U4609 (N_4609,N_3134,N_3698);
xnor U4610 (N_4610,N_3024,N_3984);
nand U4611 (N_4611,N_3012,N_3303);
nor U4612 (N_4612,N_3738,N_3521);
nor U4613 (N_4613,N_3087,N_3375);
xnor U4614 (N_4614,N_3766,N_3268);
or U4615 (N_4615,N_3716,N_3601);
nor U4616 (N_4616,N_3569,N_3262);
xnor U4617 (N_4617,N_3018,N_3474);
and U4618 (N_4618,N_3121,N_3108);
and U4619 (N_4619,N_3202,N_3914);
or U4620 (N_4620,N_3723,N_3857);
or U4621 (N_4621,N_3579,N_3494);
or U4622 (N_4622,N_3787,N_3365);
nand U4623 (N_4623,N_3608,N_3714);
nand U4624 (N_4624,N_3637,N_3740);
and U4625 (N_4625,N_3257,N_3181);
or U4626 (N_4626,N_3268,N_3988);
xor U4627 (N_4627,N_3948,N_3906);
xor U4628 (N_4628,N_3343,N_3845);
nand U4629 (N_4629,N_3124,N_3096);
nand U4630 (N_4630,N_3956,N_3897);
and U4631 (N_4631,N_3257,N_3528);
or U4632 (N_4632,N_3971,N_3802);
or U4633 (N_4633,N_3336,N_3522);
xor U4634 (N_4634,N_3079,N_3600);
and U4635 (N_4635,N_3580,N_3038);
xnor U4636 (N_4636,N_3819,N_3919);
or U4637 (N_4637,N_3580,N_3405);
or U4638 (N_4638,N_3050,N_3420);
and U4639 (N_4639,N_3278,N_3223);
and U4640 (N_4640,N_3673,N_3337);
nand U4641 (N_4641,N_3389,N_3685);
nor U4642 (N_4642,N_3059,N_3227);
nand U4643 (N_4643,N_3684,N_3510);
nor U4644 (N_4644,N_3221,N_3381);
nor U4645 (N_4645,N_3833,N_3039);
nor U4646 (N_4646,N_3719,N_3636);
xnor U4647 (N_4647,N_3413,N_3143);
and U4648 (N_4648,N_3866,N_3055);
or U4649 (N_4649,N_3886,N_3805);
and U4650 (N_4650,N_3341,N_3968);
or U4651 (N_4651,N_3245,N_3279);
nand U4652 (N_4652,N_3154,N_3498);
nand U4653 (N_4653,N_3617,N_3687);
and U4654 (N_4654,N_3026,N_3007);
nand U4655 (N_4655,N_3843,N_3381);
xor U4656 (N_4656,N_3048,N_3014);
nor U4657 (N_4657,N_3237,N_3820);
nor U4658 (N_4658,N_3687,N_3180);
nor U4659 (N_4659,N_3340,N_3908);
xor U4660 (N_4660,N_3494,N_3265);
or U4661 (N_4661,N_3282,N_3501);
xor U4662 (N_4662,N_3932,N_3296);
nand U4663 (N_4663,N_3319,N_3971);
xor U4664 (N_4664,N_3451,N_3719);
xor U4665 (N_4665,N_3096,N_3475);
and U4666 (N_4666,N_3299,N_3217);
nor U4667 (N_4667,N_3195,N_3594);
and U4668 (N_4668,N_3855,N_3176);
nand U4669 (N_4669,N_3692,N_3796);
nor U4670 (N_4670,N_3249,N_3000);
and U4671 (N_4671,N_3316,N_3702);
and U4672 (N_4672,N_3810,N_3950);
nand U4673 (N_4673,N_3319,N_3020);
or U4674 (N_4674,N_3048,N_3806);
xor U4675 (N_4675,N_3098,N_3998);
nor U4676 (N_4676,N_3879,N_3043);
nor U4677 (N_4677,N_3362,N_3481);
nor U4678 (N_4678,N_3594,N_3123);
and U4679 (N_4679,N_3714,N_3856);
and U4680 (N_4680,N_3910,N_3147);
nor U4681 (N_4681,N_3992,N_3869);
nand U4682 (N_4682,N_3724,N_3617);
or U4683 (N_4683,N_3685,N_3900);
or U4684 (N_4684,N_3484,N_3302);
xor U4685 (N_4685,N_3586,N_3147);
and U4686 (N_4686,N_3072,N_3015);
xor U4687 (N_4687,N_3453,N_3429);
nand U4688 (N_4688,N_3200,N_3672);
and U4689 (N_4689,N_3713,N_3012);
or U4690 (N_4690,N_3997,N_3555);
nand U4691 (N_4691,N_3017,N_3360);
or U4692 (N_4692,N_3415,N_3789);
and U4693 (N_4693,N_3043,N_3192);
xnor U4694 (N_4694,N_3192,N_3827);
nor U4695 (N_4695,N_3472,N_3132);
or U4696 (N_4696,N_3756,N_3816);
xor U4697 (N_4697,N_3461,N_3786);
xor U4698 (N_4698,N_3192,N_3527);
xnor U4699 (N_4699,N_3435,N_3840);
xnor U4700 (N_4700,N_3064,N_3797);
xnor U4701 (N_4701,N_3554,N_3387);
nor U4702 (N_4702,N_3013,N_3511);
xnor U4703 (N_4703,N_3489,N_3492);
nand U4704 (N_4704,N_3750,N_3756);
and U4705 (N_4705,N_3215,N_3430);
nand U4706 (N_4706,N_3699,N_3471);
nand U4707 (N_4707,N_3036,N_3055);
and U4708 (N_4708,N_3223,N_3233);
nor U4709 (N_4709,N_3522,N_3490);
xnor U4710 (N_4710,N_3892,N_3757);
xnor U4711 (N_4711,N_3888,N_3323);
xor U4712 (N_4712,N_3769,N_3427);
or U4713 (N_4713,N_3657,N_3388);
or U4714 (N_4714,N_3729,N_3129);
xor U4715 (N_4715,N_3007,N_3392);
or U4716 (N_4716,N_3762,N_3140);
and U4717 (N_4717,N_3945,N_3401);
and U4718 (N_4718,N_3269,N_3052);
or U4719 (N_4719,N_3253,N_3835);
or U4720 (N_4720,N_3860,N_3426);
xnor U4721 (N_4721,N_3731,N_3238);
nand U4722 (N_4722,N_3647,N_3100);
or U4723 (N_4723,N_3042,N_3722);
nand U4724 (N_4724,N_3371,N_3319);
xnor U4725 (N_4725,N_3690,N_3226);
nand U4726 (N_4726,N_3185,N_3573);
nand U4727 (N_4727,N_3683,N_3363);
nor U4728 (N_4728,N_3138,N_3360);
nor U4729 (N_4729,N_3494,N_3935);
nor U4730 (N_4730,N_3278,N_3248);
and U4731 (N_4731,N_3774,N_3972);
nor U4732 (N_4732,N_3989,N_3753);
nor U4733 (N_4733,N_3800,N_3554);
and U4734 (N_4734,N_3058,N_3966);
nand U4735 (N_4735,N_3688,N_3732);
and U4736 (N_4736,N_3208,N_3193);
nand U4737 (N_4737,N_3034,N_3665);
or U4738 (N_4738,N_3392,N_3020);
nand U4739 (N_4739,N_3704,N_3444);
and U4740 (N_4740,N_3431,N_3734);
and U4741 (N_4741,N_3930,N_3698);
or U4742 (N_4742,N_3608,N_3331);
nor U4743 (N_4743,N_3749,N_3661);
and U4744 (N_4744,N_3455,N_3857);
nand U4745 (N_4745,N_3323,N_3236);
or U4746 (N_4746,N_3641,N_3244);
and U4747 (N_4747,N_3476,N_3824);
nor U4748 (N_4748,N_3413,N_3389);
or U4749 (N_4749,N_3580,N_3019);
and U4750 (N_4750,N_3074,N_3807);
nor U4751 (N_4751,N_3167,N_3415);
or U4752 (N_4752,N_3567,N_3515);
xnor U4753 (N_4753,N_3104,N_3781);
xnor U4754 (N_4754,N_3123,N_3747);
nand U4755 (N_4755,N_3021,N_3381);
and U4756 (N_4756,N_3625,N_3044);
nor U4757 (N_4757,N_3878,N_3990);
nand U4758 (N_4758,N_3894,N_3987);
nand U4759 (N_4759,N_3819,N_3002);
xnor U4760 (N_4760,N_3036,N_3428);
and U4761 (N_4761,N_3656,N_3697);
and U4762 (N_4762,N_3254,N_3345);
nand U4763 (N_4763,N_3637,N_3678);
or U4764 (N_4764,N_3695,N_3403);
or U4765 (N_4765,N_3106,N_3587);
or U4766 (N_4766,N_3634,N_3438);
or U4767 (N_4767,N_3983,N_3128);
and U4768 (N_4768,N_3627,N_3767);
nor U4769 (N_4769,N_3637,N_3203);
xnor U4770 (N_4770,N_3383,N_3061);
xor U4771 (N_4771,N_3111,N_3438);
xor U4772 (N_4772,N_3143,N_3474);
and U4773 (N_4773,N_3857,N_3527);
or U4774 (N_4774,N_3839,N_3288);
xor U4775 (N_4775,N_3745,N_3631);
or U4776 (N_4776,N_3624,N_3801);
or U4777 (N_4777,N_3317,N_3517);
nor U4778 (N_4778,N_3226,N_3854);
nor U4779 (N_4779,N_3125,N_3663);
xor U4780 (N_4780,N_3383,N_3088);
xor U4781 (N_4781,N_3081,N_3479);
and U4782 (N_4782,N_3484,N_3864);
or U4783 (N_4783,N_3918,N_3791);
nand U4784 (N_4784,N_3144,N_3632);
nor U4785 (N_4785,N_3106,N_3292);
nor U4786 (N_4786,N_3360,N_3757);
nand U4787 (N_4787,N_3628,N_3254);
xnor U4788 (N_4788,N_3573,N_3646);
and U4789 (N_4789,N_3027,N_3031);
and U4790 (N_4790,N_3010,N_3413);
xnor U4791 (N_4791,N_3249,N_3841);
and U4792 (N_4792,N_3277,N_3953);
or U4793 (N_4793,N_3481,N_3910);
nor U4794 (N_4794,N_3845,N_3130);
or U4795 (N_4795,N_3095,N_3150);
or U4796 (N_4796,N_3660,N_3190);
nand U4797 (N_4797,N_3000,N_3724);
xor U4798 (N_4798,N_3616,N_3018);
nor U4799 (N_4799,N_3684,N_3733);
and U4800 (N_4800,N_3168,N_3461);
and U4801 (N_4801,N_3103,N_3353);
and U4802 (N_4802,N_3114,N_3516);
nor U4803 (N_4803,N_3165,N_3890);
nand U4804 (N_4804,N_3439,N_3459);
nor U4805 (N_4805,N_3919,N_3501);
nand U4806 (N_4806,N_3522,N_3446);
xnor U4807 (N_4807,N_3552,N_3044);
or U4808 (N_4808,N_3732,N_3711);
nor U4809 (N_4809,N_3152,N_3256);
xor U4810 (N_4810,N_3710,N_3772);
xor U4811 (N_4811,N_3433,N_3470);
nor U4812 (N_4812,N_3990,N_3689);
or U4813 (N_4813,N_3193,N_3018);
nand U4814 (N_4814,N_3760,N_3016);
or U4815 (N_4815,N_3054,N_3400);
nor U4816 (N_4816,N_3499,N_3336);
xnor U4817 (N_4817,N_3276,N_3636);
or U4818 (N_4818,N_3807,N_3888);
xnor U4819 (N_4819,N_3718,N_3010);
or U4820 (N_4820,N_3933,N_3824);
nor U4821 (N_4821,N_3913,N_3893);
nand U4822 (N_4822,N_3099,N_3279);
xnor U4823 (N_4823,N_3730,N_3464);
or U4824 (N_4824,N_3548,N_3927);
xor U4825 (N_4825,N_3558,N_3629);
and U4826 (N_4826,N_3471,N_3242);
and U4827 (N_4827,N_3131,N_3533);
nand U4828 (N_4828,N_3356,N_3952);
or U4829 (N_4829,N_3137,N_3125);
or U4830 (N_4830,N_3732,N_3259);
and U4831 (N_4831,N_3229,N_3464);
and U4832 (N_4832,N_3295,N_3906);
or U4833 (N_4833,N_3314,N_3471);
xor U4834 (N_4834,N_3887,N_3267);
or U4835 (N_4835,N_3765,N_3757);
nor U4836 (N_4836,N_3381,N_3806);
nor U4837 (N_4837,N_3238,N_3569);
and U4838 (N_4838,N_3244,N_3827);
or U4839 (N_4839,N_3870,N_3323);
nand U4840 (N_4840,N_3035,N_3199);
and U4841 (N_4841,N_3245,N_3033);
or U4842 (N_4842,N_3477,N_3171);
xnor U4843 (N_4843,N_3079,N_3933);
or U4844 (N_4844,N_3859,N_3774);
xor U4845 (N_4845,N_3270,N_3182);
nor U4846 (N_4846,N_3270,N_3504);
nand U4847 (N_4847,N_3478,N_3969);
and U4848 (N_4848,N_3804,N_3501);
xnor U4849 (N_4849,N_3230,N_3510);
nand U4850 (N_4850,N_3492,N_3208);
or U4851 (N_4851,N_3387,N_3206);
nand U4852 (N_4852,N_3293,N_3206);
xor U4853 (N_4853,N_3717,N_3996);
or U4854 (N_4854,N_3096,N_3546);
nand U4855 (N_4855,N_3255,N_3015);
xnor U4856 (N_4856,N_3670,N_3931);
nor U4857 (N_4857,N_3351,N_3375);
or U4858 (N_4858,N_3268,N_3479);
and U4859 (N_4859,N_3564,N_3808);
xnor U4860 (N_4860,N_3006,N_3751);
nor U4861 (N_4861,N_3067,N_3894);
nor U4862 (N_4862,N_3269,N_3105);
nand U4863 (N_4863,N_3172,N_3379);
xor U4864 (N_4864,N_3858,N_3419);
and U4865 (N_4865,N_3210,N_3625);
xnor U4866 (N_4866,N_3346,N_3521);
xor U4867 (N_4867,N_3656,N_3551);
xnor U4868 (N_4868,N_3206,N_3475);
nor U4869 (N_4869,N_3807,N_3041);
and U4870 (N_4870,N_3971,N_3330);
nor U4871 (N_4871,N_3161,N_3652);
xnor U4872 (N_4872,N_3824,N_3595);
or U4873 (N_4873,N_3836,N_3234);
nand U4874 (N_4874,N_3186,N_3372);
nand U4875 (N_4875,N_3706,N_3757);
or U4876 (N_4876,N_3128,N_3074);
xor U4877 (N_4877,N_3311,N_3094);
and U4878 (N_4878,N_3740,N_3079);
xor U4879 (N_4879,N_3743,N_3768);
nand U4880 (N_4880,N_3213,N_3255);
and U4881 (N_4881,N_3983,N_3541);
xor U4882 (N_4882,N_3676,N_3679);
nand U4883 (N_4883,N_3341,N_3946);
nor U4884 (N_4884,N_3251,N_3849);
and U4885 (N_4885,N_3831,N_3860);
or U4886 (N_4886,N_3280,N_3982);
or U4887 (N_4887,N_3376,N_3580);
xor U4888 (N_4888,N_3272,N_3778);
nor U4889 (N_4889,N_3451,N_3288);
nor U4890 (N_4890,N_3047,N_3187);
nor U4891 (N_4891,N_3303,N_3398);
xor U4892 (N_4892,N_3692,N_3515);
nand U4893 (N_4893,N_3061,N_3554);
nand U4894 (N_4894,N_3812,N_3376);
or U4895 (N_4895,N_3962,N_3534);
nand U4896 (N_4896,N_3106,N_3504);
or U4897 (N_4897,N_3811,N_3127);
nor U4898 (N_4898,N_3598,N_3691);
nor U4899 (N_4899,N_3593,N_3559);
nor U4900 (N_4900,N_3389,N_3968);
or U4901 (N_4901,N_3176,N_3942);
nand U4902 (N_4902,N_3666,N_3139);
nand U4903 (N_4903,N_3383,N_3007);
and U4904 (N_4904,N_3523,N_3550);
and U4905 (N_4905,N_3898,N_3237);
nor U4906 (N_4906,N_3801,N_3327);
or U4907 (N_4907,N_3182,N_3436);
nand U4908 (N_4908,N_3901,N_3862);
nand U4909 (N_4909,N_3570,N_3279);
nor U4910 (N_4910,N_3794,N_3337);
nor U4911 (N_4911,N_3762,N_3073);
or U4912 (N_4912,N_3453,N_3180);
xor U4913 (N_4913,N_3365,N_3595);
nor U4914 (N_4914,N_3777,N_3904);
nor U4915 (N_4915,N_3883,N_3926);
xnor U4916 (N_4916,N_3101,N_3065);
or U4917 (N_4917,N_3384,N_3660);
or U4918 (N_4918,N_3469,N_3617);
xnor U4919 (N_4919,N_3572,N_3082);
or U4920 (N_4920,N_3689,N_3131);
xnor U4921 (N_4921,N_3345,N_3550);
and U4922 (N_4922,N_3745,N_3289);
nand U4923 (N_4923,N_3998,N_3212);
nor U4924 (N_4924,N_3091,N_3481);
or U4925 (N_4925,N_3793,N_3000);
and U4926 (N_4926,N_3557,N_3566);
nand U4927 (N_4927,N_3428,N_3388);
nand U4928 (N_4928,N_3119,N_3795);
nor U4929 (N_4929,N_3147,N_3738);
and U4930 (N_4930,N_3828,N_3892);
nor U4931 (N_4931,N_3041,N_3861);
and U4932 (N_4932,N_3286,N_3580);
and U4933 (N_4933,N_3930,N_3846);
or U4934 (N_4934,N_3514,N_3314);
nor U4935 (N_4935,N_3760,N_3914);
xor U4936 (N_4936,N_3840,N_3789);
or U4937 (N_4937,N_3322,N_3742);
or U4938 (N_4938,N_3088,N_3061);
xor U4939 (N_4939,N_3748,N_3020);
or U4940 (N_4940,N_3545,N_3748);
nor U4941 (N_4941,N_3837,N_3349);
nand U4942 (N_4942,N_3514,N_3190);
or U4943 (N_4943,N_3985,N_3558);
nand U4944 (N_4944,N_3075,N_3785);
nor U4945 (N_4945,N_3071,N_3555);
nand U4946 (N_4946,N_3767,N_3219);
xor U4947 (N_4947,N_3860,N_3429);
nand U4948 (N_4948,N_3866,N_3017);
xnor U4949 (N_4949,N_3793,N_3979);
nand U4950 (N_4950,N_3518,N_3285);
and U4951 (N_4951,N_3007,N_3128);
and U4952 (N_4952,N_3249,N_3876);
and U4953 (N_4953,N_3876,N_3633);
and U4954 (N_4954,N_3506,N_3135);
xnor U4955 (N_4955,N_3765,N_3854);
xor U4956 (N_4956,N_3073,N_3166);
or U4957 (N_4957,N_3558,N_3702);
nor U4958 (N_4958,N_3517,N_3472);
and U4959 (N_4959,N_3092,N_3423);
nor U4960 (N_4960,N_3927,N_3684);
xor U4961 (N_4961,N_3207,N_3493);
and U4962 (N_4962,N_3451,N_3407);
nand U4963 (N_4963,N_3977,N_3666);
or U4964 (N_4964,N_3159,N_3748);
nor U4965 (N_4965,N_3687,N_3902);
and U4966 (N_4966,N_3274,N_3938);
nor U4967 (N_4967,N_3735,N_3117);
xnor U4968 (N_4968,N_3928,N_3395);
xnor U4969 (N_4969,N_3088,N_3908);
xor U4970 (N_4970,N_3846,N_3305);
xor U4971 (N_4971,N_3269,N_3752);
and U4972 (N_4972,N_3440,N_3832);
nand U4973 (N_4973,N_3845,N_3335);
or U4974 (N_4974,N_3856,N_3124);
or U4975 (N_4975,N_3669,N_3647);
nor U4976 (N_4976,N_3545,N_3632);
nand U4977 (N_4977,N_3924,N_3899);
nand U4978 (N_4978,N_3956,N_3731);
nor U4979 (N_4979,N_3951,N_3083);
and U4980 (N_4980,N_3964,N_3322);
xor U4981 (N_4981,N_3225,N_3117);
xor U4982 (N_4982,N_3615,N_3870);
nor U4983 (N_4983,N_3828,N_3498);
xnor U4984 (N_4984,N_3502,N_3878);
or U4985 (N_4985,N_3429,N_3812);
and U4986 (N_4986,N_3977,N_3676);
nor U4987 (N_4987,N_3645,N_3082);
nor U4988 (N_4988,N_3394,N_3468);
and U4989 (N_4989,N_3149,N_3940);
or U4990 (N_4990,N_3218,N_3077);
nor U4991 (N_4991,N_3555,N_3098);
and U4992 (N_4992,N_3391,N_3382);
or U4993 (N_4993,N_3218,N_3486);
xor U4994 (N_4994,N_3890,N_3616);
xnor U4995 (N_4995,N_3028,N_3286);
nor U4996 (N_4996,N_3288,N_3042);
and U4997 (N_4997,N_3808,N_3460);
or U4998 (N_4998,N_3905,N_3713);
xor U4999 (N_4999,N_3239,N_3561);
nor U5000 (N_5000,N_4423,N_4391);
or U5001 (N_5001,N_4239,N_4351);
and U5002 (N_5002,N_4542,N_4537);
nand U5003 (N_5003,N_4762,N_4763);
nor U5004 (N_5004,N_4125,N_4343);
nand U5005 (N_5005,N_4493,N_4964);
nor U5006 (N_5006,N_4393,N_4828);
and U5007 (N_5007,N_4637,N_4352);
nand U5008 (N_5008,N_4517,N_4134);
and U5009 (N_5009,N_4363,N_4106);
or U5010 (N_5010,N_4751,N_4174);
nand U5011 (N_5011,N_4266,N_4460);
nor U5012 (N_5012,N_4663,N_4236);
xnor U5013 (N_5013,N_4317,N_4742);
xor U5014 (N_5014,N_4670,N_4107);
and U5015 (N_5015,N_4313,N_4576);
or U5016 (N_5016,N_4212,N_4782);
and U5017 (N_5017,N_4092,N_4028);
xor U5018 (N_5018,N_4556,N_4540);
nand U5019 (N_5019,N_4585,N_4318);
and U5020 (N_5020,N_4648,N_4740);
xor U5021 (N_5021,N_4781,N_4987);
and U5022 (N_5022,N_4717,N_4533);
xor U5023 (N_5023,N_4187,N_4366);
nand U5024 (N_5024,N_4922,N_4095);
nand U5025 (N_5025,N_4864,N_4120);
nor U5026 (N_5026,N_4735,N_4579);
xor U5027 (N_5027,N_4729,N_4350);
and U5028 (N_5028,N_4721,N_4892);
or U5029 (N_5029,N_4226,N_4872);
nor U5030 (N_5030,N_4386,N_4645);
nor U5031 (N_5031,N_4432,N_4845);
nor U5032 (N_5032,N_4060,N_4815);
nor U5033 (N_5033,N_4247,N_4611);
nand U5034 (N_5034,N_4688,N_4691);
nor U5035 (N_5035,N_4957,N_4859);
nor U5036 (N_5036,N_4652,N_4941);
or U5037 (N_5037,N_4230,N_4622);
xnor U5038 (N_5038,N_4179,N_4029);
xor U5039 (N_5039,N_4019,N_4241);
and U5040 (N_5040,N_4405,N_4961);
or U5041 (N_5041,N_4246,N_4639);
nor U5042 (N_5042,N_4039,N_4056);
and U5043 (N_5043,N_4695,N_4726);
nand U5044 (N_5044,N_4501,N_4018);
nor U5045 (N_5045,N_4249,N_4122);
nand U5046 (N_5046,N_4903,N_4888);
and U5047 (N_5047,N_4114,N_4720);
and U5048 (N_5048,N_4080,N_4368);
and U5049 (N_5049,N_4306,N_4188);
nand U5050 (N_5050,N_4597,N_4111);
or U5051 (N_5051,N_4527,N_4243);
nand U5052 (N_5052,N_4298,N_4562);
or U5053 (N_5053,N_4422,N_4974);
and U5054 (N_5054,N_4671,N_4984);
xnor U5055 (N_5055,N_4618,N_4287);
nor U5056 (N_5056,N_4673,N_4176);
and U5057 (N_5057,N_4248,N_4148);
xor U5058 (N_5058,N_4965,N_4098);
nor U5059 (N_5059,N_4950,N_4299);
or U5060 (N_5060,N_4127,N_4307);
xor U5061 (N_5061,N_4335,N_4788);
xnor U5062 (N_5062,N_4659,N_4012);
nand U5063 (N_5063,N_4764,N_4606);
or U5064 (N_5064,N_4678,N_4996);
and U5065 (N_5065,N_4117,N_4336);
or U5066 (N_5066,N_4676,N_4147);
or U5067 (N_5067,N_4087,N_4449);
nand U5068 (N_5068,N_4103,N_4768);
nand U5069 (N_5069,N_4817,N_4858);
and U5070 (N_5070,N_4599,N_4654);
and U5071 (N_5071,N_4909,N_4936);
or U5072 (N_5072,N_4172,N_4031);
or U5073 (N_5073,N_4733,N_4427);
nand U5074 (N_5074,N_4059,N_4337);
xnor U5075 (N_5075,N_4235,N_4870);
xnor U5076 (N_5076,N_4710,N_4975);
xor U5077 (N_5077,N_4590,N_4371);
nor U5078 (N_5078,N_4837,N_4008);
and U5079 (N_5079,N_4309,N_4348);
nand U5080 (N_5080,N_4388,N_4444);
nand U5081 (N_5081,N_4392,N_4536);
xor U5082 (N_5082,N_4508,N_4617);
or U5083 (N_5083,N_4704,N_4398);
nand U5084 (N_5084,N_4474,N_4412);
and U5085 (N_5085,N_4473,N_4948);
xnor U5086 (N_5086,N_4582,N_4951);
or U5087 (N_5087,N_4602,N_4158);
nand U5088 (N_5088,N_4373,N_4455);
xnor U5089 (N_5089,N_4206,N_4598);
or U5090 (N_5090,N_4030,N_4826);
xor U5091 (N_5091,N_4549,N_4133);
nand U5092 (N_5092,N_4963,N_4138);
xor U5093 (N_5093,N_4390,N_4960);
or U5094 (N_5094,N_4901,N_4032);
xor U5095 (N_5095,N_4580,N_4048);
and U5096 (N_5096,N_4842,N_4015);
nand U5097 (N_5097,N_4310,N_4271);
nand U5098 (N_5098,N_4101,N_4384);
or U5099 (N_5099,N_4433,N_4958);
nor U5100 (N_5100,N_4989,N_4969);
or U5101 (N_5101,N_4642,N_4701);
nand U5102 (N_5102,N_4970,N_4777);
xor U5103 (N_5103,N_4478,N_4042);
nand U5104 (N_5104,N_4943,N_4441);
nand U5105 (N_5105,N_4340,N_4785);
nor U5106 (N_5106,N_4213,N_4467);
and U5107 (N_5107,N_4126,N_4001);
xnor U5108 (N_5108,N_4291,N_4732);
nand U5109 (N_5109,N_4083,N_4369);
nand U5110 (N_5110,N_4380,N_4112);
nand U5111 (N_5111,N_4516,N_4857);
or U5112 (N_5112,N_4578,N_4166);
nor U5113 (N_5113,N_4833,N_4897);
xnor U5114 (N_5114,N_4865,N_4813);
xor U5115 (N_5115,N_4069,N_4035);
nor U5116 (N_5116,N_4899,N_4486);
and U5117 (N_5117,N_4853,N_4852);
and U5118 (N_5118,N_4711,N_4672);
xnor U5119 (N_5119,N_4719,N_4534);
and U5120 (N_5120,N_4295,N_4435);
xor U5121 (N_5121,N_4472,N_4468);
xnor U5122 (N_5122,N_4128,N_4041);
nor U5123 (N_5123,N_4811,N_4500);
nand U5124 (N_5124,N_4697,N_4314);
or U5125 (N_5125,N_4685,N_4605);
nand U5126 (N_5126,N_4417,N_4219);
nor U5127 (N_5127,N_4144,N_4354);
and U5128 (N_5128,N_4929,N_4448);
nor U5129 (N_5129,N_4322,N_4196);
or U5130 (N_5130,N_4090,N_4862);
nor U5131 (N_5131,N_4358,N_4481);
nand U5132 (N_5132,N_4553,N_4917);
xnor U5133 (N_5133,N_4497,N_4947);
or U5134 (N_5134,N_4382,N_4331);
nand U5135 (N_5135,N_4274,N_4918);
nor U5136 (N_5136,N_4666,N_4806);
and U5137 (N_5137,N_4829,N_4883);
xor U5138 (N_5138,N_4752,N_4223);
xnor U5139 (N_5139,N_4278,N_4082);
nand U5140 (N_5140,N_4362,N_4292);
nand U5141 (N_5141,N_4904,N_4430);
nor U5142 (N_5142,N_4300,N_4779);
and U5143 (N_5143,N_4660,N_4926);
or U5144 (N_5144,N_4007,N_4634);
and U5145 (N_5145,N_4066,N_4203);
and U5146 (N_5146,N_4630,N_4277);
and U5147 (N_5147,N_4739,N_4476);
or U5148 (N_5148,N_4400,N_4966);
and U5149 (N_5149,N_4184,N_4669);
and U5150 (N_5150,N_4071,N_4237);
or U5151 (N_5151,N_4968,N_4413);
nor U5152 (N_5152,N_4381,N_4320);
and U5153 (N_5153,N_4577,N_4426);
or U5154 (N_5154,N_4442,N_4357);
or U5155 (N_5155,N_4905,N_4631);
xnor U5156 (N_5156,N_4689,N_4131);
or U5157 (N_5157,N_4329,N_4210);
xor U5158 (N_5158,N_4410,N_4286);
and U5159 (N_5159,N_4022,N_4934);
nand U5160 (N_5160,N_4139,N_4208);
and U5161 (N_5161,N_4195,N_4548);
nand U5162 (N_5162,N_4667,N_4175);
nand U5163 (N_5163,N_4067,N_4755);
nor U5164 (N_5164,N_4263,N_4070);
xnor U5165 (N_5165,N_4635,N_4462);
or U5166 (N_5166,N_4531,N_4167);
nor U5167 (N_5167,N_4954,N_4461);
and U5168 (N_5168,N_4170,N_4510);
xnor U5169 (N_5169,N_4457,N_4894);
xor U5170 (N_5170,N_4428,N_4898);
or U5171 (N_5171,N_4055,N_4332);
xor U5172 (N_5172,N_4529,N_4896);
xor U5173 (N_5173,N_4159,N_4973);
or U5174 (N_5174,N_4803,N_4315);
nor U5175 (N_5175,N_4955,N_4094);
or U5176 (N_5176,N_4925,N_4293);
or U5177 (N_5177,N_4401,N_4915);
and U5178 (N_5178,N_4923,N_4992);
nor U5179 (N_5179,N_4265,N_4372);
nand U5180 (N_5180,N_4222,N_4566);
or U5181 (N_5181,N_4728,N_4783);
nand U5182 (N_5182,N_4543,N_4044);
and U5183 (N_5183,N_4620,N_4054);
nor U5184 (N_5184,N_4123,N_4919);
xor U5185 (N_5185,N_4770,N_4805);
nand U5186 (N_5186,N_4604,N_4308);
and U5187 (N_5187,N_4301,N_4712);
and U5188 (N_5188,N_4831,N_4339);
or U5189 (N_5189,N_4270,N_4503);
nor U5190 (N_5190,N_4253,N_4003);
xnor U5191 (N_5191,N_4181,N_4465);
nand U5192 (N_5192,N_4713,N_4827);
or U5193 (N_5193,N_4623,N_4743);
nor U5194 (N_5194,N_4985,N_4312);
or U5195 (N_5195,N_4484,N_4229);
or U5196 (N_5196,N_4932,N_4355);
and U5197 (N_5197,N_4698,N_4102);
xnor U5198 (N_5198,N_4784,N_4953);
and U5199 (N_5199,N_4871,N_4215);
xor U5200 (N_5200,N_4220,N_4438);
nand U5201 (N_5201,N_4737,N_4108);
and U5202 (N_5202,N_4482,N_4569);
nand U5203 (N_5203,N_4769,N_4397);
xor U5204 (N_5204,N_4451,N_4010);
nor U5205 (N_5205,N_4256,N_4884);
or U5206 (N_5206,N_4940,N_4024);
nor U5207 (N_5207,N_4443,N_4479);
xnor U5208 (N_5208,N_4745,N_4047);
xnor U5209 (N_5209,N_4696,N_4808);
xor U5210 (N_5210,N_4110,N_4924);
xnor U5211 (N_5211,N_4023,N_4233);
and U5212 (N_5212,N_4570,N_4601);
nand U5213 (N_5213,N_4281,N_4004);
or U5214 (N_5214,N_4771,N_4496);
and U5215 (N_5215,N_4703,N_4708);
nor U5216 (N_5216,N_4025,N_4981);
xor U5217 (N_5217,N_4690,N_4945);
nand U5218 (N_5218,N_4586,N_4261);
nand U5219 (N_5219,N_4628,N_4135);
xnor U5220 (N_5220,N_4855,N_4458);
or U5221 (N_5221,N_4952,N_4538);
or U5222 (N_5222,N_4773,N_4545);
nor U5223 (N_5223,N_4000,N_4072);
or U5224 (N_5224,N_4641,N_4843);
nand U5225 (N_5225,N_4902,N_4880);
and U5226 (N_5226,N_4259,N_4600);
xnor U5227 (N_5227,N_4150,N_4559);
and U5228 (N_5228,N_4323,N_4319);
nand U5229 (N_5229,N_4061,N_4456);
nor U5230 (N_5230,N_4376,N_4284);
xnor U5231 (N_5231,N_4668,N_4205);
or U5232 (N_5232,N_4789,N_4891);
nand U5233 (N_5233,N_4440,N_4504);
nand U5234 (N_5234,N_4296,N_4420);
or U5235 (N_5235,N_4825,N_4279);
or U5236 (N_5236,N_4571,N_4608);
or U5237 (N_5237,N_4214,N_4183);
nor U5238 (N_5238,N_4252,N_4959);
nand U5239 (N_5239,N_4353,N_4492);
xnor U5240 (N_5240,N_4136,N_4804);
nor U5241 (N_5241,N_4991,N_4521);
and U5242 (N_5242,N_4040,N_4129);
xnor U5243 (N_5243,N_4861,N_4491);
or U5244 (N_5244,N_4034,N_4629);
xor U5245 (N_5245,N_4514,N_4077);
and U5246 (N_5246,N_4658,N_4574);
and U5247 (N_5247,N_4887,N_4119);
nand U5248 (N_5248,N_4885,N_4850);
or U5249 (N_5249,N_4304,N_4038);
nor U5250 (N_5250,N_4723,N_4665);
and U5251 (N_5251,N_4342,N_4242);
nor U5252 (N_5252,N_4824,N_4627);
xor U5253 (N_5253,N_4589,N_4979);
or U5254 (N_5254,N_4847,N_4509);
or U5255 (N_5255,N_4624,N_4447);
and U5256 (N_5256,N_4844,N_4065);
or U5257 (N_5257,N_4583,N_4809);
and U5258 (N_5258,N_4749,N_4778);
or U5259 (N_5259,N_4794,N_4552);
nand U5260 (N_5260,N_4873,N_4882);
nor U5261 (N_5261,N_4976,N_4879);
or U5262 (N_5262,N_4716,N_4480);
or U5263 (N_5263,N_4063,N_4999);
xnor U5264 (N_5264,N_4483,N_4581);
nor U5265 (N_5265,N_4801,N_4105);
xor U5266 (N_5266,N_4334,N_4986);
nand U5267 (N_5267,N_4238,N_4408);
nor U5268 (N_5268,N_4240,N_4646);
and U5269 (N_5269,N_4192,N_4734);
nand U5270 (N_5270,N_4209,N_4211);
nand U5271 (N_5271,N_4560,N_4787);
nor U5272 (N_5272,N_4093,N_4568);
or U5273 (N_5273,N_4164,N_4452);
nor U5274 (N_5274,N_4191,N_4725);
xor U5275 (N_5275,N_4962,N_4889);
or U5276 (N_5276,N_4201,N_4983);
or U5277 (N_5277,N_4526,N_4445);
or U5278 (N_5278,N_4816,N_4874);
or U5279 (N_5279,N_4881,N_4555);
and U5280 (N_5280,N_4200,N_4463);
and U5281 (N_5281,N_4109,N_4632);
xnor U5282 (N_5282,N_4361,N_4650);
or U5283 (N_5283,N_4613,N_4683);
and U5284 (N_5284,N_4027,N_4610);
xor U5285 (N_5285,N_4377,N_4994);
nor U5286 (N_5286,N_4193,N_4793);
nor U5287 (N_5287,N_4615,N_4835);
or U5288 (N_5288,N_4705,N_4868);
xnor U5289 (N_5289,N_4100,N_4772);
xor U5290 (N_5290,N_4050,N_4524);
and U5291 (N_5291,N_4268,N_4561);
xnor U5292 (N_5292,N_4169,N_4655);
and U5293 (N_5293,N_4792,N_4812);
xor U5294 (N_5294,N_4906,N_4282);
xor U5295 (N_5295,N_4832,N_4890);
xnor U5296 (N_5296,N_4978,N_4541);
nand U5297 (N_5297,N_4411,N_4033);
xor U5298 (N_5298,N_4823,N_4692);
nand U5299 (N_5299,N_4190,N_4402);
nor U5300 (N_5300,N_4152,N_4928);
and U5301 (N_5301,N_4914,N_4140);
nor U5302 (N_5302,N_4851,N_4619);
nand U5303 (N_5303,N_4429,N_4385);
nor U5304 (N_5304,N_4026,N_4621);
xor U5305 (N_5305,N_4475,N_4765);
or U5306 (N_5306,N_4394,N_4488);
xnor U5307 (N_5307,N_4796,N_4021);
nor U5308 (N_5308,N_4244,N_4748);
or U5309 (N_5309,N_4194,N_4609);
xnor U5310 (N_5310,N_4389,N_4840);
xnor U5311 (N_5311,N_4178,N_4849);
and U5312 (N_5312,N_4730,N_4416);
nor U5313 (N_5313,N_4694,N_4005);
and U5314 (N_5314,N_4116,N_4780);
or U5315 (N_5315,N_4346,N_4997);
and U5316 (N_5316,N_4378,N_4834);
nor U5317 (N_5317,N_4137,N_4995);
xnor U5318 (N_5318,N_4546,N_4738);
or U5319 (N_5319,N_4328,N_4349);
xnor U5320 (N_5320,N_4113,N_4636);
nand U5321 (N_5321,N_4535,N_4370);
nor U5322 (N_5322,N_4155,N_4550);
and U5323 (N_5323,N_4217,N_4283);
and U5324 (N_5324,N_4724,N_4564);
xor U5325 (N_5325,N_4406,N_4900);
xnor U5326 (N_5326,N_4747,N_4907);
xnor U5327 (N_5327,N_4437,N_4614);
nand U5328 (N_5328,N_4797,N_4640);
xnor U5329 (N_5329,N_4439,N_4911);
nand U5330 (N_5330,N_4020,N_4551);
and U5331 (N_5331,N_4511,N_4130);
or U5332 (N_5332,N_4626,N_4643);
xor U5333 (N_5333,N_4707,N_4625);
nor U5334 (N_5334,N_4939,N_4799);
and U5335 (N_5335,N_4185,N_4036);
xnor U5336 (N_5336,N_4664,N_4846);
or U5337 (N_5337,N_4592,N_4702);
nor U5338 (N_5338,N_4588,N_4518);
nand U5339 (N_5339,N_4736,N_4324);
nor U5340 (N_5340,N_4199,N_4333);
or U5341 (N_5341,N_4767,N_4260);
nand U5342 (N_5342,N_4180,N_4177);
nand U5343 (N_5343,N_4168,N_4878);
nor U5344 (N_5344,N_4424,N_4446);
nor U5345 (N_5345,N_4856,N_4819);
xnor U5346 (N_5346,N_4251,N_4595);
xor U5347 (N_5347,N_4303,N_4189);
and U5348 (N_5348,N_4163,N_4949);
nand U5349 (N_5349,N_4754,N_4662);
nand U5350 (N_5350,N_4656,N_4046);
xnor U5351 (N_5351,N_4280,N_4638);
xor U5352 (N_5352,N_4151,N_4972);
xor U5353 (N_5353,N_4273,N_4225);
or U5354 (N_5354,N_4075,N_4866);
nor U5355 (N_5355,N_4913,N_4741);
nand U5356 (N_5356,N_4775,N_4776);
xor U5357 (N_5357,N_4450,N_4593);
nor U5358 (N_5358,N_4267,N_4786);
nand U5359 (N_5359,N_4414,N_4587);
or U5360 (N_5360,N_4058,N_4316);
and U5361 (N_5361,N_4507,N_4407);
or U5362 (N_5362,N_4675,N_4869);
xor U5363 (N_5363,N_4718,N_4289);
nand U5364 (N_5364,N_4532,N_4436);
and U5365 (N_5365,N_4375,N_4774);
xor U5366 (N_5366,N_4761,N_4146);
nor U5367 (N_5367,N_4104,N_4074);
or U5368 (N_5368,N_4810,N_4231);
nand U5369 (N_5369,N_4379,N_4097);
or U5370 (N_5370,N_4927,N_4272);
nand U5371 (N_5371,N_4197,N_4469);
or U5372 (N_5372,N_4453,N_4512);
or U5373 (N_5373,N_4224,N_4431);
or U5374 (N_5374,N_4766,N_4182);
nor U5375 (N_5375,N_4791,N_4750);
nand U5376 (N_5376,N_4993,N_4173);
xor U5377 (N_5377,N_4285,N_4078);
or U5378 (N_5378,N_4043,N_4714);
or U5379 (N_5379,N_4679,N_4245);
or U5380 (N_5380,N_4933,N_4800);
or U5381 (N_5381,N_4297,N_4115);
xor U5382 (N_5382,N_4326,N_4434);
nor U5383 (N_5383,N_4502,N_4607);
nand U5384 (N_5384,N_4171,N_4344);
or U5385 (N_5385,N_4544,N_4325);
nand U5386 (N_5386,N_4674,N_4202);
nand U5387 (N_5387,N_4495,N_4228);
or U5388 (N_5388,N_4760,N_4143);
nand U5389 (N_5389,N_4099,N_4421);
xnor U5390 (N_5390,N_4498,N_4715);
and U5391 (N_5391,N_4523,N_4360);
nor U5392 (N_5392,N_4633,N_4269);
nand U5393 (N_5393,N_4338,N_4980);
or U5394 (N_5394,N_4255,N_4876);
and U5395 (N_5395,N_4687,N_4931);
xnor U5396 (N_5396,N_4795,N_4506);
and U5397 (N_5397,N_4470,N_4731);
nand U5398 (N_5398,N_4649,N_4367);
nand U5399 (N_5399,N_4403,N_4937);
or U5400 (N_5400,N_4085,N_4294);
xnor U5401 (N_5401,N_4330,N_4557);
nor U5402 (N_5402,N_4596,N_4364);
or U5403 (N_5403,N_4700,N_4684);
or U5404 (N_5404,N_4161,N_4982);
nor U5405 (N_5405,N_4490,N_4830);
nand U5406 (N_5406,N_4820,N_4198);
and U5407 (N_5407,N_4204,N_4584);
nand U5408 (N_5408,N_4073,N_4612);
xor U5409 (N_5409,N_4227,N_4935);
xnor U5410 (N_5410,N_4053,N_4356);
or U5411 (N_5411,N_4057,N_4591);
nor U5412 (N_5412,N_4002,N_4345);
or U5413 (N_5413,N_4867,N_4374);
nor U5414 (N_5414,N_4311,N_4758);
and U5415 (N_5415,N_4554,N_4839);
nand U5416 (N_5416,N_4154,N_4016);
nor U5417 (N_5417,N_4014,N_4942);
nor U5418 (N_5418,N_4258,N_4096);
and U5419 (N_5419,N_4207,N_4276);
and U5420 (N_5420,N_4647,N_4798);
nand U5421 (N_5421,N_4347,N_4464);
or U5422 (N_5422,N_4807,N_4409);
and U5423 (N_5423,N_4946,N_4162);
nor U5424 (N_5424,N_4013,N_4938);
nor U5425 (N_5425,N_4232,N_4988);
or U5426 (N_5426,N_4321,N_4860);
nor U5427 (N_5427,N_4466,N_4528);
or U5428 (N_5428,N_4722,N_4499);
xor U5429 (N_5429,N_4037,N_4744);
nor U5430 (N_5430,N_4489,N_4603);
xor U5431 (N_5431,N_4153,N_4753);
and U5432 (N_5432,N_4365,N_4288);
nand U5433 (N_5433,N_4539,N_4944);
nand U5434 (N_5434,N_4573,N_4863);
nor U5435 (N_5435,N_4383,N_4088);
and U5436 (N_5436,N_4477,N_4686);
nor U5437 (N_5437,N_4485,N_4575);
and U5438 (N_5438,N_4305,N_4912);
and U5439 (N_5439,N_4836,N_4399);
and U5440 (N_5440,N_4567,N_4257);
and U5441 (N_5441,N_4049,N_4149);
nand U5442 (N_5442,N_4089,N_4790);
xor U5443 (N_5443,N_4920,N_4009);
and U5444 (N_5444,N_4756,N_4875);
and U5445 (N_5445,N_4814,N_4657);
or U5446 (N_5446,N_4977,N_4572);
or U5447 (N_5447,N_4644,N_4616);
or U5448 (N_5448,N_4145,N_4459);
nand U5449 (N_5449,N_4045,N_4519);
or U5450 (N_5450,N_4395,N_4221);
nand U5451 (N_5451,N_4746,N_4404);
nor U5452 (N_5452,N_4956,N_4142);
nor U5453 (N_5453,N_4156,N_4419);
and U5454 (N_5454,N_4359,N_4017);
nand U5455 (N_5455,N_4079,N_4522);
xnor U5456 (N_5456,N_4921,N_4091);
nor U5457 (N_5457,N_4505,N_4425);
nand U5458 (N_5458,N_4157,N_4121);
xnor U5459 (N_5459,N_4530,N_4699);
and U5460 (N_5460,N_4525,N_4132);
or U5461 (N_5461,N_4759,N_4186);
nor U5462 (N_5462,N_4341,N_4594);
nor U5463 (N_5463,N_4854,N_4680);
xor U5464 (N_5464,N_4415,N_4681);
nor U5465 (N_5465,N_4302,N_4471);
xor U5466 (N_5466,N_4706,N_4677);
or U5467 (N_5467,N_4254,N_4990);
or U5468 (N_5468,N_4910,N_4141);
and U5469 (N_5469,N_4709,N_4262);
nand U5470 (N_5470,N_4081,N_4821);
and U5471 (N_5471,N_4886,N_4893);
nor U5472 (N_5472,N_4494,N_4124);
nand U5473 (N_5473,N_4250,N_4757);
or U5474 (N_5474,N_4418,N_4727);
nand U5475 (N_5475,N_4565,N_4877);
xor U5476 (N_5476,N_4076,N_4682);
or U5477 (N_5477,N_4651,N_4895);
nor U5478 (N_5478,N_4848,N_4290);
xor U5479 (N_5479,N_4216,N_4693);
and U5480 (N_5480,N_4822,N_4062);
nor U5481 (N_5481,N_4520,N_4661);
and U5482 (N_5482,N_4387,N_4011);
nor U5483 (N_5483,N_4841,N_4971);
and U5484 (N_5484,N_4006,N_4653);
nand U5485 (N_5485,N_4327,N_4118);
nand U5486 (N_5486,N_4275,N_4547);
xor U5487 (N_5487,N_4838,N_4563);
xor U5488 (N_5488,N_4802,N_4487);
and U5489 (N_5489,N_4930,N_4916);
and U5490 (N_5490,N_4084,N_4967);
nand U5491 (N_5491,N_4513,N_4234);
nor U5492 (N_5492,N_4165,N_4160);
or U5493 (N_5493,N_4068,N_4264);
nor U5494 (N_5494,N_4396,N_4086);
and U5495 (N_5495,N_4515,N_4454);
xnor U5496 (N_5496,N_4558,N_4051);
nor U5497 (N_5497,N_4064,N_4052);
and U5498 (N_5498,N_4218,N_4818);
or U5499 (N_5499,N_4998,N_4908);
nand U5500 (N_5500,N_4087,N_4113);
nor U5501 (N_5501,N_4836,N_4427);
and U5502 (N_5502,N_4042,N_4832);
nor U5503 (N_5503,N_4919,N_4412);
xnor U5504 (N_5504,N_4711,N_4259);
nor U5505 (N_5505,N_4149,N_4984);
and U5506 (N_5506,N_4475,N_4719);
xor U5507 (N_5507,N_4992,N_4028);
nand U5508 (N_5508,N_4599,N_4574);
nor U5509 (N_5509,N_4184,N_4651);
nand U5510 (N_5510,N_4423,N_4730);
and U5511 (N_5511,N_4896,N_4172);
nand U5512 (N_5512,N_4382,N_4098);
nand U5513 (N_5513,N_4298,N_4631);
nor U5514 (N_5514,N_4033,N_4115);
nand U5515 (N_5515,N_4681,N_4523);
nand U5516 (N_5516,N_4582,N_4930);
or U5517 (N_5517,N_4978,N_4746);
and U5518 (N_5518,N_4026,N_4346);
xnor U5519 (N_5519,N_4162,N_4988);
and U5520 (N_5520,N_4887,N_4600);
or U5521 (N_5521,N_4925,N_4090);
or U5522 (N_5522,N_4832,N_4605);
nor U5523 (N_5523,N_4763,N_4289);
nand U5524 (N_5524,N_4660,N_4121);
nand U5525 (N_5525,N_4309,N_4914);
nand U5526 (N_5526,N_4260,N_4135);
nor U5527 (N_5527,N_4035,N_4212);
and U5528 (N_5528,N_4636,N_4536);
nor U5529 (N_5529,N_4620,N_4541);
nor U5530 (N_5530,N_4497,N_4802);
and U5531 (N_5531,N_4625,N_4080);
or U5532 (N_5532,N_4263,N_4180);
and U5533 (N_5533,N_4188,N_4662);
and U5534 (N_5534,N_4559,N_4091);
and U5535 (N_5535,N_4314,N_4372);
nand U5536 (N_5536,N_4481,N_4598);
and U5537 (N_5537,N_4142,N_4831);
nand U5538 (N_5538,N_4292,N_4484);
xnor U5539 (N_5539,N_4290,N_4160);
nor U5540 (N_5540,N_4745,N_4548);
or U5541 (N_5541,N_4172,N_4632);
nand U5542 (N_5542,N_4266,N_4295);
xor U5543 (N_5543,N_4394,N_4246);
nor U5544 (N_5544,N_4745,N_4840);
and U5545 (N_5545,N_4110,N_4322);
nor U5546 (N_5546,N_4341,N_4299);
nand U5547 (N_5547,N_4856,N_4347);
nand U5548 (N_5548,N_4340,N_4983);
xnor U5549 (N_5549,N_4808,N_4123);
and U5550 (N_5550,N_4122,N_4502);
xnor U5551 (N_5551,N_4308,N_4922);
xor U5552 (N_5552,N_4150,N_4925);
xnor U5553 (N_5553,N_4379,N_4333);
and U5554 (N_5554,N_4349,N_4507);
or U5555 (N_5555,N_4470,N_4426);
or U5556 (N_5556,N_4579,N_4793);
nand U5557 (N_5557,N_4471,N_4539);
xor U5558 (N_5558,N_4971,N_4834);
or U5559 (N_5559,N_4784,N_4772);
and U5560 (N_5560,N_4731,N_4754);
xnor U5561 (N_5561,N_4100,N_4445);
xnor U5562 (N_5562,N_4857,N_4800);
nor U5563 (N_5563,N_4251,N_4774);
nor U5564 (N_5564,N_4330,N_4771);
nand U5565 (N_5565,N_4381,N_4836);
xor U5566 (N_5566,N_4449,N_4608);
and U5567 (N_5567,N_4592,N_4972);
nand U5568 (N_5568,N_4200,N_4603);
nand U5569 (N_5569,N_4631,N_4397);
or U5570 (N_5570,N_4420,N_4773);
nor U5571 (N_5571,N_4951,N_4223);
xor U5572 (N_5572,N_4139,N_4594);
xor U5573 (N_5573,N_4524,N_4360);
nand U5574 (N_5574,N_4948,N_4038);
and U5575 (N_5575,N_4683,N_4655);
xor U5576 (N_5576,N_4074,N_4352);
or U5577 (N_5577,N_4198,N_4805);
xnor U5578 (N_5578,N_4878,N_4472);
nand U5579 (N_5579,N_4597,N_4838);
xnor U5580 (N_5580,N_4120,N_4874);
and U5581 (N_5581,N_4504,N_4589);
nor U5582 (N_5582,N_4889,N_4340);
nand U5583 (N_5583,N_4036,N_4275);
nand U5584 (N_5584,N_4454,N_4188);
nand U5585 (N_5585,N_4452,N_4849);
or U5586 (N_5586,N_4898,N_4176);
nand U5587 (N_5587,N_4996,N_4561);
nor U5588 (N_5588,N_4433,N_4290);
and U5589 (N_5589,N_4674,N_4730);
xnor U5590 (N_5590,N_4106,N_4506);
and U5591 (N_5591,N_4997,N_4694);
or U5592 (N_5592,N_4017,N_4127);
and U5593 (N_5593,N_4173,N_4523);
nand U5594 (N_5594,N_4087,N_4751);
or U5595 (N_5595,N_4595,N_4748);
xnor U5596 (N_5596,N_4271,N_4598);
nor U5597 (N_5597,N_4608,N_4857);
nor U5598 (N_5598,N_4802,N_4270);
and U5599 (N_5599,N_4496,N_4906);
or U5600 (N_5600,N_4280,N_4695);
and U5601 (N_5601,N_4815,N_4148);
and U5602 (N_5602,N_4453,N_4798);
xnor U5603 (N_5603,N_4103,N_4628);
nand U5604 (N_5604,N_4576,N_4737);
nor U5605 (N_5605,N_4769,N_4490);
or U5606 (N_5606,N_4120,N_4602);
xnor U5607 (N_5607,N_4624,N_4814);
nand U5608 (N_5608,N_4591,N_4074);
or U5609 (N_5609,N_4966,N_4518);
or U5610 (N_5610,N_4932,N_4338);
or U5611 (N_5611,N_4867,N_4987);
or U5612 (N_5612,N_4878,N_4710);
nor U5613 (N_5613,N_4523,N_4203);
nand U5614 (N_5614,N_4133,N_4816);
xor U5615 (N_5615,N_4252,N_4351);
or U5616 (N_5616,N_4560,N_4264);
and U5617 (N_5617,N_4924,N_4388);
xnor U5618 (N_5618,N_4471,N_4889);
nand U5619 (N_5619,N_4192,N_4658);
nor U5620 (N_5620,N_4396,N_4261);
nor U5621 (N_5621,N_4915,N_4757);
nand U5622 (N_5622,N_4816,N_4399);
xnor U5623 (N_5623,N_4311,N_4505);
nand U5624 (N_5624,N_4260,N_4375);
xor U5625 (N_5625,N_4204,N_4916);
and U5626 (N_5626,N_4312,N_4884);
nor U5627 (N_5627,N_4868,N_4768);
nor U5628 (N_5628,N_4913,N_4108);
nor U5629 (N_5629,N_4030,N_4428);
xnor U5630 (N_5630,N_4209,N_4497);
or U5631 (N_5631,N_4012,N_4535);
nor U5632 (N_5632,N_4095,N_4710);
nand U5633 (N_5633,N_4972,N_4028);
and U5634 (N_5634,N_4427,N_4779);
and U5635 (N_5635,N_4945,N_4014);
and U5636 (N_5636,N_4138,N_4371);
or U5637 (N_5637,N_4361,N_4088);
nor U5638 (N_5638,N_4672,N_4277);
xnor U5639 (N_5639,N_4296,N_4147);
xor U5640 (N_5640,N_4007,N_4396);
xor U5641 (N_5641,N_4649,N_4267);
and U5642 (N_5642,N_4789,N_4593);
nand U5643 (N_5643,N_4080,N_4045);
and U5644 (N_5644,N_4692,N_4146);
or U5645 (N_5645,N_4312,N_4367);
and U5646 (N_5646,N_4756,N_4370);
nand U5647 (N_5647,N_4443,N_4534);
nor U5648 (N_5648,N_4264,N_4147);
nand U5649 (N_5649,N_4432,N_4005);
or U5650 (N_5650,N_4150,N_4786);
nand U5651 (N_5651,N_4348,N_4703);
and U5652 (N_5652,N_4693,N_4304);
nand U5653 (N_5653,N_4240,N_4265);
nand U5654 (N_5654,N_4781,N_4001);
or U5655 (N_5655,N_4774,N_4966);
nand U5656 (N_5656,N_4048,N_4503);
and U5657 (N_5657,N_4460,N_4177);
and U5658 (N_5658,N_4877,N_4334);
xor U5659 (N_5659,N_4779,N_4166);
xnor U5660 (N_5660,N_4765,N_4144);
or U5661 (N_5661,N_4629,N_4159);
xnor U5662 (N_5662,N_4344,N_4388);
or U5663 (N_5663,N_4288,N_4623);
or U5664 (N_5664,N_4762,N_4631);
and U5665 (N_5665,N_4041,N_4985);
xor U5666 (N_5666,N_4422,N_4754);
nor U5667 (N_5667,N_4521,N_4952);
nand U5668 (N_5668,N_4685,N_4361);
nand U5669 (N_5669,N_4391,N_4569);
nand U5670 (N_5670,N_4282,N_4206);
or U5671 (N_5671,N_4482,N_4619);
nand U5672 (N_5672,N_4266,N_4599);
and U5673 (N_5673,N_4269,N_4903);
xor U5674 (N_5674,N_4287,N_4379);
xor U5675 (N_5675,N_4959,N_4551);
nand U5676 (N_5676,N_4009,N_4474);
xnor U5677 (N_5677,N_4741,N_4154);
nand U5678 (N_5678,N_4604,N_4381);
nand U5679 (N_5679,N_4208,N_4123);
nor U5680 (N_5680,N_4840,N_4732);
nand U5681 (N_5681,N_4575,N_4030);
nand U5682 (N_5682,N_4441,N_4348);
xnor U5683 (N_5683,N_4246,N_4069);
and U5684 (N_5684,N_4993,N_4302);
nor U5685 (N_5685,N_4601,N_4374);
or U5686 (N_5686,N_4649,N_4671);
and U5687 (N_5687,N_4249,N_4671);
nand U5688 (N_5688,N_4927,N_4566);
nand U5689 (N_5689,N_4913,N_4955);
or U5690 (N_5690,N_4813,N_4902);
and U5691 (N_5691,N_4389,N_4205);
and U5692 (N_5692,N_4550,N_4663);
xor U5693 (N_5693,N_4314,N_4596);
or U5694 (N_5694,N_4516,N_4791);
and U5695 (N_5695,N_4942,N_4915);
nand U5696 (N_5696,N_4955,N_4533);
xnor U5697 (N_5697,N_4438,N_4965);
xnor U5698 (N_5698,N_4454,N_4323);
nor U5699 (N_5699,N_4767,N_4793);
xor U5700 (N_5700,N_4478,N_4948);
or U5701 (N_5701,N_4725,N_4781);
or U5702 (N_5702,N_4357,N_4129);
nand U5703 (N_5703,N_4241,N_4843);
or U5704 (N_5704,N_4836,N_4759);
and U5705 (N_5705,N_4309,N_4891);
or U5706 (N_5706,N_4545,N_4200);
nor U5707 (N_5707,N_4219,N_4507);
and U5708 (N_5708,N_4559,N_4060);
or U5709 (N_5709,N_4682,N_4403);
nor U5710 (N_5710,N_4246,N_4354);
and U5711 (N_5711,N_4786,N_4565);
xnor U5712 (N_5712,N_4778,N_4051);
xor U5713 (N_5713,N_4277,N_4273);
nor U5714 (N_5714,N_4866,N_4229);
nand U5715 (N_5715,N_4678,N_4623);
xor U5716 (N_5716,N_4870,N_4928);
nand U5717 (N_5717,N_4793,N_4504);
nand U5718 (N_5718,N_4606,N_4753);
nor U5719 (N_5719,N_4509,N_4313);
nor U5720 (N_5720,N_4994,N_4597);
and U5721 (N_5721,N_4137,N_4721);
or U5722 (N_5722,N_4918,N_4239);
and U5723 (N_5723,N_4730,N_4846);
nand U5724 (N_5724,N_4693,N_4013);
and U5725 (N_5725,N_4369,N_4759);
xor U5726 (N_5726,N_4997,N_4440);
nand U5727 (N_5727,N_4702,N_4500);
nand U5728 (N_5728,N_4749,N_4159);
nand U5729 (N_5729,N_4702,N_4988);
xor U5730 (N_5730,N_4822,N_4322);
and U5731 (N_5731,N_4754,N_4069);
nand U5732 (N_5732,N_4090,N_4251);
and U5733 (N_5733,N_4644,N_4718);
nand U5734 (N_5734,N_4056,N_4404);
or U5735 (N_5735,N_4094,N_4098);
and U5736 (N_5736,N_4444,N_4749);
or U5737 (N_5737,N_4280,N_4386);
nor U5738 (N_5738,N_4494,N_4021);
xor U5739 (N_5739,N_4208,N_4847);
and U5740 (N_5740,N_4197,N_4772);
or U5741 (N_5741,N_4418,N_4079);
nor U5742 (N_5742,N_4270,N_4642);
and U5743 (N_5743,N_4175,N_4690);
nand U5744 (N_5744,N_4285,N_4893);
and U5745 (N_5745,N_4363,N_4684);
and U5746 (N_5746,N_4690,N_4176);
nand U5747 (N_5747,N_4843,N_4694);
xnor U5748 (N_5748,N_4198,N_4899);
or U5749 (N_5749,N_4629,N_4013);
and U5750 (N_5750,N_4187,N_4602);
and U5751 (N_5751,N_4980,N_4252);
nor U5752 (N_5752,N_4430,N_4643);
nand U5753 (N_5753,N_4462,N_4527);
nand U5754 (N_5754,N_4526,N_4093);
and U5755 (N_5755,N_4167,N_4346);
xor U5756 (N_5756,N_4304,N_4501);
nand U5757 (N_5757,N_4930,N_4667);
nand U5758 (N_5758,N_4540,N_4847);
nand U5759 (N_5759,N_4402,N_4860);
nor U5760 (N_5760,N_4615,N_4867);
nor U5761 (N_5761,N_4548,N_4198);
nor U5762 (N_5762,N_4974,N_4464);
and U5763 (N_5763,N_4958,N_4125);
xor U5764 (N_5764,N_4695,N_4227);
xnor U5765 (N_5765,N_4891,N_4354);
nand U5766 (N_5766,N_4020,N_4566);
nor U5767 (N_5767,N_4627,N_4328);
or U5768 (N_5768,N_4699,N_4729);
and U5769 (N_5769,N_4356,N_4740);
nor U5770 (N_5770,N_4202,N_4019);
nand U5771 (N_5771,N_4077,N_4416);
and U5772 (N_5772,N_4281,N_4297);
nor U5773 (N_5773,N_4588,N_4169);
nand U5774 (N_5774,N_4250,N_4376);
nor U5775 (N_5775,N_4210,N_4616);
or U5776 (N_5776,N_4168,N_4651);
nor U5777 (N_5777,N_4134,N_4824);
nor U5778 (N_5778,N_4979,N_4395);
and U5779 (N_5779,N_4627,N_4378);
or U5780 (N_5780,N_4483,N_4567);
xnor U5781 (N_5781,N_4859,N_4707);
xnor U5782 (N_5782,N_4127,N_4648);
and U5783 (N_5783,N_4494,N_4526);
nand U5784 (N_5784,N_4615,N_4750);
or U5785 (N_5785,N_4336,N_4023);
or U5786 (N_5786,N_4024,N_4522);
and U5787 (N_5787,N_4136,N_4454);
nor U5788 (N_5788,N_4692,N_4999);
nand U5789 (N_5789,N_4692,N_4629);
nor U5790 (N_5790,N_4166,N_4905);
nor U5791 (N_5791,N_4149,N_4320);
nand U5792 (N_5792,N_4009,N_4566);
or U5793 (N_5793,N_4893,N_4875);
nor U5794 (N_5794,N_4896,N_4195);
xnor U5795 (N_5795,N_4142,N_4940);
and U5796 (N_5796,N_4939,N_4774);
nor U5797 (N_5797,N_4423,N_4644);
xnor U5798 (N_5798,N_4202,N_4523);
or U5799 (N_5799,N_4069,N_4920);
nor U5800 (N_5800,N_4812,N_4158);
xnor U5801 (N_5801,N_4552,N_4857);
nor U5802 (N_5802,N_4392,N_4817);
xor U5803 (N_5803,N_4333,N_4570);
xnor U5804 (N_5804,N_4767,N_4774);
or U5805 (N_5805,N_4736,N_4146);
nor U5806 (N_5806,N_4410,N_4220);
and U5807 (N_5807,N_4324,N_4727);
nor U5808 (N_5808,N_4615,N_4226);
nor U5809 (N_5809,N_4166,N_4702);
or U5810 (N_5810,N_4876,N_4804);
nor U5811 (N_5811,N_4460,N_4871);
or U5812 (N_5812,N_4791,N_4563);
and U5813 (N_5813,N_4548,N_4370);
nand U5814 (N_5814,N_4464,N_4243);
xnor U5815 (N_5815,N_4177,N_4067);
or U5816 (N_5816,N_4958,N_4091);
or U5817 (N_5817,N_4975,N_4885);
nor U5818 (N_5818,N_4371,N_4408);
or U5819 (N_5819,N_4279,N_4455);
nand U5820 (N_5820,N_4336,N_4140);
and U5821 (N_5821,N_4171,N_4433);
xor U5822 (N_5822,N_4601,N_4456);
xor U5823 (N_5823,N_4303,N_4103);
or U5824 (N_5824,N_4669,N_4780);
nand U5825 (N_5825,N_4389,N_4479);
nand U5826 (N_5826,N_4540,N_4503);
or U5827 (N_5827,N_4395,N_4113);
and U5828 (N_5828,N_4160,N_4443);
or U5829 (N_5829,N_4474,N_4510);
nor U5830 (N_5830,N_4426,N_4643);
xnor U5831 (N_5831,N_4950,N_4154);
nand U5832 (N_5832,N_4767,N_4732);
xnor U5833 (N_5833,N_4751,N_4512);
xor U5834 (N_5834,N_4968,N_4233);
or U5835 (N_5835,N_4959,N_4331);
and U5836 (N_5836,N_4079,N_4177);
nand U5837 (N_5837,N_4747,N_4916);
and U5838 (N_5838,N_4704,N_4016);
and U5839 (N_5839,N_4290,N_4929);
nor U5840 (N_5840,N_4657,N_4222);
and U5841 (N_5841,N_4840,N_4683);
nand U5842 (N_5842,N_4561,N_4880);
xnor U5843 (N_5843,N_4953,N_4974);
or U5844 (N_5844,N_4605,N_4030);
xor U5845 (N_5845,N_4088,N_4576);
and U5846 (N_5846,N_4601,N_4449);
xnor U5847 (N_5847,N_4295,N_4140);
xnor U5848 (N_5848,N_4812,N_4848);
or U5849 (N_5849,N_4614,N_4648);
nor U5850 (N_5850,N_4913,N_4530);
nor U5851 (N_5851,N_4668,N_4990);
xor U5852 (N_5852,N_4029,N_4866);
xnor U5853 (N_5853,N_4636,N_4187);
or U5854 (N_5854,N_4818,N_4518);
nor U5855 (N_5855,N_4561,N_4584);
or U5856 (N_5856,N_4820,N_4203);
and U5857 (N_5857,N_4872,N_4363);
nor U5858 (N_5858,N_4722,N_4262);
nand U5859 (N_5859,N_4746,N_4595);
xor U5860 (N_5860,N_4564,N_4304);
xnor U5861 (N_5861,N_4307,N_4525);
nand U5862 (N_5862,N_4826,N_4362);
and U5863 (N_5863,N_4519,N_4812);
nor U5864 (N_5864,N_4180,N_4700);
or U5865 (N_5865,N_4057,N_4341);
xnor U5866 (N_5866,N_4436,N_4031);
and U5867 (N_5867,N_4130,N_4265);
xor U5868 (N_5868,N_4790,N_4956);
and U5869 (N_5869,N_4262,N_4994);
xnor U5870 (N_5870,N_4368,N_4389);
xor U5871 (N_5871,N_4188,N_4239);
or U5872 (N_5872,N_4385,N_4321);
or U5873 (N_5873,N_4698,N_4740);
nand U5874 (N_5874,N_4010,N_4071);
nor U5875 (N_5875,N_4688,N_4575);
xor U5876 (N_5876,N_4762,N_4230);
xnor U5877 (N_5877,N_4089,N_4311);
and U5878 (N_5878,N_4799,N_4065);
and U5879 (N_5879,N_4036,N_4796);
or U5880 (N_5880,N_4191,N_4414);
nor U5881 (N_5881,N_4823,N_4722);
xor U5882 (N_5882,N_4200,N_4094);
xnor U5883 (N_5883,N_4823,N_4941);
nand U5884 (N_5884,N_4535,N_4247);
or U5885 (N_5885,N_4303,N_4678);
nor U5886 (N_5886,N_4579,N_4947);
xor U5887 (N_5887,N_4518,N_4808);
or U5888 (N_5888,N_4188,N_4358);
or U5889 (N_5889,N_4119,N_4990);
and U5890 (N_5890,N_4827,N_4282);
or U5891 (N_5891,N_4910,N_4248);
xor U5892 (N_5892,N_4955,N_4334);
nor U5893 (N_5893,N_4362,N_4698);
or U5894 (N_5894,N_4893,N_4538);
and U5895 (N_5895,N_4502,N_4660);
and U5896 (N_5896,N_4822,N_4925);
or U5897 (N_5897,N_4069,N_4097);
xor U5898 (N_5898,N_4146,N_4536);
or U5899 (N_5899,N_4442,N_4726);
nor U5900 (N_5900,N_4853,N_4357);
and U5901 (N_5901,N_4773,N_4097);
xor U5902 (N_5902,N_4193,N_4076);
nand U5903 (N_5903,N_4024,N_4027);
or U5904 (N_5904,N_4393,N_4783);
xnor U5905 (N_5905,N_4222,N_4251);
and U5906 (N_5906,N_4416,N_4070);
nand U5907 (N_5907,N_4155,N_4175);
or U5908 (N_5908,N_4877,N_4243);
nand U5909 (N_5909,N_4804,N_4765);
nor U5910 (N_5910,N_4987,N_4961);
and U5911 (N_5911,N_4936,N_4379);
and U5912 (N_5912,N_4459,N_4200);
xnor U5913 (N_5913,N_4252,N_4132);
or U5914 (N_5914,N_4819,N_4704);
nand U5915 (N_5915,N_4600,N_4661);
xnor U5916 (N_5916,N_4208,N_4555);
xor U5917 (N_5917,N_4268,N_4622);
nand U5918 (N_5918,N_4071,N_4847);
nor U5919 (N_5919,N_4407,N_4066);
nand U5920 (N_5920,N_4360,N_4519);
nor U5921 (N_5921,N_4496,N_4533);
or U5922 (N_5922,N_4353,N_4319);
xnor U5923 (N_5923,N_4551,N_4371);
nand U5924 (N_5924,N_4648,N_4171);
or U5925 (N_5925,N_4663,N_4116);
or U5926 (N_5926,N_4296,N_4864);
or U5927 (N_5927,N_4828,N_4815);
nor U5928 (N_5928,N_4366,N_4602);
and U5929 (N_5929,N_4296,N_4268);
nor U5930 (N_5930,N_4372,N_4298);
nor U5931 (N_5931,N_4086,N_4407);
nor U5932 (N_5932,N_4454,N_4166);
nor U5933 (N_5933,N_4727,N_4500);
nor U5934 (N_5934,N_4176,N_4993);
nor U5935 (N_5935,N_4425,N_4363);
nor U5936 (N_5936,N_4895,N_4320);
nand U5937 (N_5937,N_4887,N_4615);
nor U5938 (N_5938,N_4244,N_4497);
or U5939 (N_5939,N_4241,N_4068);
or U5940 (N_5940,N_4042,N_4407);
xor U5941 (N_5941,N_4239,N_4270);
nand U5942 (N_5942,N_4661,N_4611);
nor U5943 (N_5943,N_4197,N_4405);
nor U5944 (N_5944,N_4725,N_4157);
and U5945 (N_5945,N_4240,N_4979);
xnor U5946 (N_5946,N_4570,N_4409);
nor U5947 (N_5947,N_4875,N_4864);
nand U5948 (N_5948,N_4225,N_4196);
and U5949 (N_5949,N_4699,N_4804);
nand U5950 (N_5950,N_4372,N_4801);
nand U5951 (N_5951,N_4212,N_4367);
nand U5952 (N_5952,N_4112,N_4944);
nor U5953 (N_5953,N_4126,N_4045);
and U5954 (N_5954,N_4057,N_4869);
or U5955 (N_5955,N_4355,N_4874);
or U5956 (N_5956,N_4168,N_4296);
and U5957 (N_5957,N_4546,N_4899);
and U5958 (N_5958,N_4447,N_4534);
nor U5959 (N_5959,N_4204,N_4228);
nand U5960 (N_5960,N_4956,N_4119);
and U5961 (N_5961,N_4231,N_4130);
or U5962 (N_5962,N_4376,N_4933);
and U5963 (N_5963,N_4547,N_4364);
nand U5964 (N_5964,N_4606,N_4338);
xnor U5965 (N_5965,N_4460,N_4230);
nand U5966 (N_5966,N_4239,N_4121);
or U5967 (N_5967,N_4116,N_4135);
nor U5968 (N_5968,N_4953,N_4635);
and U5969 (N_5969,N_4799,N_4594);
xor U5970 (N_5970,N_4351,N_4912);
nor U5971 (N_5971,N_4300,N_4658);
xnor U5972 (N_5972,N_4634,N_4662);
nand U5973 (N_5973,N_4129,N_4054);
and U5974 (N_5974,N_4927,N_4614);
and U5975 (N_5975,N_4963,N_4865);
nand U5976 (N_5976,N_4654,N_4081);
nand U5977 (N_5977,N_4269,N_4165);
xnor U5978 (N_5978,N_4433,N_4231);
or U5979 (N_5979,N_4299,N_4720);
xnor U5980 (N_5980,N_4149,N_4625);
or U5981 (N_5981,N_4097,N_4659);
and U5982 (N_5982,N_4328,N_4299);
and U5983 (N_5983,N_4268,N_4942);
and U5984 (N_5984,N_4829,N_4249);
nand U5985 (N_5985,N_4158,N_4234);
nand U5986 (N_5986,N_4672,N_4430);
xnor U5987 (N_5987,N_4739,N_4466);
xnor U5988 (N_5988,N_4657,N_4957);
xnor U5989 (N_5989,N_4693,N_4425);
xnor U5990 (N_5990,N_4442,N_4186);
or U5991 (N_5991,N_4112,N_4194);
or U5992 (N_5992,N_4454,N_4312);
nor U5993 (N_5993,N_4998,N_4558);
and U5994 (N_5994,N_4805,N_4609);
nand U5995 (N_5995,N_4276,N_4089);
and U5996 (N_5996,N_4685,N_4641);
or U5997 (N_5997,N_4369,N_4738);
nand U5998 (N_5998,N_4085,N_4000);
nand U5999 (N_5999,N_4492,N_4369);
xor U6000 (N_6000,N_5591,N_5063);
or U6001 (N_6001,N_5315,N_5562);
or U6002 (N_6002,N_5766,N_5191);
or U6003 (N_6003,N_5006,N_5004);
nand U6004 (N_6004,N_5199,N_5623);
or U6005 (N_6005,N_5327,N_5780);
or U6006 (N_6006,N_5078,N_5155);
and U6007 (N_6007,N_5894,N_5776);
nor U6008 (N_6008,N_5292,N_5380);
and U6009 (N_6009,N_5201,N_5885);
nor U6010 (N_6010,N_5851,N_5092);
or U6011 (N_6011,N_5332,N_5625);
nand U6012 (N_6012,N_5844,N_5284);
or U6013 (N_6013,N_5480,N_5349);
or U6014 (N_6014,N_5121,N_5320);
nor U6015 (N_6015,N_5639,N_5627);
and U6016 (N_6016,N_5041,N_5048);
nand U6017 (N_6017,N_5364,N_5813);
nand U6018 (N_6018,N_5996,N_5599);
xnor U6019 (N_6019,N_5356,N_5317);
nand U6020 (N_6020,N_5210,N_5278);
or U6021 (N_6021,N_5283,N_5664);
nand U6022 (N_6022,N_5207,N_5868);
nor U6023 (N_6023,N_5496,N_5059);
and U6024 (N_6024,N_5802,N_5412);
or U6025 (N_6025,N_5864,N_5857);
or U6026 (N_6026,N_5072,N_5878);
nand U6027 (N_6027,N_5093,N_5335);
nor U6028 (N_6028,N_5822,N_5202);
xnor U6029 (N_6029,N_5212,N_5451);
xnor U6030 (N_6030,N_5019,N_5989);
nand U6031 (N_6031,N_5637,N_5262);
or U6032 (N_6032,N_5365,N_5785);
nand U6033 (N_6033,N_5512,N_5217);
nor U6034 (N_6034,N_5460,N_5643);
xnor U6035 (N_6035,N_5389,N_5406);
or U6036 (N_6036,N_5969,N_5914);
nand U6037 (N_6037,N_5694,N_5267);
xor U6038 (N_6038,N_5732,N_5114);
nor U6039 (N_6039,N_5000,N_5951);
xnor U6040 (N_6040,N_5721,N_5127);
and U6041 (N_6041,N_5630,N_5848);
and U6042 (N_6042,N_5130,N_5696);
or U6043 (N_6043,N_5569,N_5456);
xor U6044 (N_6044,N_5531,N_5386);
nand U6045 (N_6045,N_5464,N_5892);
and U6046 (N_6046,N_5146,N_5449);
or U6047 (N_6047,N_5368,N_5974);
xor U6048 (N_6048,N_5045,N_5959);
nand U6049 (N_6049,N_5757,N_5036);
nand U6050 (N_6050,N_5624,N_5076);
or U6051 (N_6051,N_5177,N_5738);
or U6052 (N_6052,N_5617,N_5887);
and U6053 (N_6053,N_5580,N_5972);
and U6054 (N_6054,N_5872,N_5180);
or U6055 (N_6055,N_5106,N_5331);
nor U6056 (N_6056,N_5519,N_5919);
or U6057 (N_6057,N_5251,N_5051);
or U6058 (N_6058,N_5920,N_5502);
or U6059 (N_6059,N_5622,N_5925);
xor U6060 (N_6060,N_5265,N_5174);
and U6061 (N_6061,N_5084,N_5835);
xor U6062 (N_6062,N_5582,N_5376);
nor U6063 (N_6063,N_5646,N_5960);
nor U6064 (N_6064,N_5438,N_5043);
or U6065 (N_6065,N_5908,N_5884);
nand U6066 (N_6066,N_5156,N_5903);
nand U6067 (N_6067,N_5240,N_5410);
xnor U6068 (N_6068,N_5746,N_5466);
and U6069 (N_6069,N_5706,N_5444);
nand U6070 (N_6070,N_5508,N_5940);
nand U6071 (N_6071,N_5577,N_5606);
nor U6072 (N_6072,N_5518,N_5465);
nor U6073 (N_6073,N_5831,N_5269);
or U6074 (N_6074,N_5398,N_5268);
nor U6075 (N_6075,N_5392,N_5521);
or U6076 (N_6076,N_5533,N_5091);
nand U6077 (N_6077,N_5977,N_5472);
nor U6078 (N_6078,N_5129,N_5160);
and U6079 (N_6079,N_5642,N_5904);
or U6080 (N_6080,N_5939,N_5397);
nand U6081 (N_6081,N_5856,N_5353);
or U6082 (N_6082,N_5401,N_5657);
and U6083 (N_6083,N_5101,N_5017);
or U6084 (N_6084,N_5455,N_5289);
xnor U6085 (N_6085,N_5681,N_5205);
and U6086 (N_6086,N_5970,N_5243);
xor U6087 (N_6087,N_5812,N_5470);
and U6088 (N_6088,N_5462,N_5105);
and U6089 (N_6089,N_5228,N_5366);
or U6090 (N_6090,N_5545,N_5404);
nor U6091 (N_6091,N_5286,N_5382);
nand U6092 (N_6092,N_5170,N_5786);
nor U6093 (N_6093,N_5165,N_5816);
or U6094 (N_6094,N_5823,N_5836);
nand U6095 (N_6095,N_5291,N_5762);
nand U6096 (N_6096,N_5002,N_5066);
nor U6097 (N_6097,N_5138,N_5527);
and U6098 (N_6098,N_5244,N_5275);
or U6099 (N_6099,N_5215,N_5337);
xor U6100 (N_6100,N_5407,N_5071);
or U6101 (N_6101,N_5081,N_5481);
nand U6102 (N_6102,N_5737,N_5733);
or U6103 (N_6103,N_5687,N_5719);
xnor U6104 (N_6104,N_5307,N_5390);
nand U6105 (N_6105,N_5369,N_5585);
nand U6106 (N_6106,N_5587,N_5383);
nand U6107 (N_6107,N_5126,N_5184);
and U6108 (N_6108,N_5538,N_5852);
xor U6109 (N_6109,N_5446,N_5628);
xor U6110 (N_6110,N_5858,N_5109);
or U6111 (N_6111,N_5497,N_5433);
nand U6112 (N_6112,N_5420,N_5697);
xor U6113 (N_6113,N_5375,N_5342);
nor U6114 (N_6114,N_5699,N_5689);
nand U6115 (N_6115,N_5612,N_5225);
or U6116 (N_6116,N_5610,N_5739);
nand U6117 (N_6117,N_5423,N_5552);
or U6118 (N_6118,N_5299,N_5988);
or U6119 (N_6119,N_5711,N_5361);
and U6120 (N_6120,N_5498,N_5992);
nor U6121 (N_6121,N_5902,N_5163);
nand U6122 (N_6122,N_5312,N_5718);
nand U6123 (N_6123,N_5613,N_5850);
xnor U6124 (N_6124,N_5351,N_5966);
nand U6125 (N_6125,N_5501,N_5341);
nand U6126 (N_6126,N_5149,N_5068);
xnor U6127 (N_6127,N_5221,N_5484);
or U6128 (N_6128,N_5104,N_5979);
nor U6129 (N_6129,N_5821,N_5842);
or U6130 (N_6130,N_5935,N_5021);
and U6131 (N_6131,N_5968,N_5633);
xor U6132 (N_6132,N_5115,N_5997);
or U6133 (N_6133,N_5564,N_5676);
and U6134 (N_6134,N_5791,N_5783);
or U6135 (N_6135,N_5226,N_5123);
xnor U6136 (N_6136,N_5488,N_5475);
nor U6137 (N_6137,N_5391,N_5428);
or U6138 (N_6138,N_5744,N_5300);
xnor U6139 (N_6139,N_5001,N_5861);
or U6140 (N_6140,N_5060,N_5551);
nand U6141 (N_6141,N_5980,N_5476);
and U6142 (N_6142,N_5399,N_5990);
nor U6143 (N_6143,N_5889,N_5425);
and U6144 (N_6144,N_5248,N_5660);
xor U6145 (N_6145,N_5937,N_5408);
or U6146 (N_6146,N_5578,N_5705);
xor U6147 (N_6147,N_5800,N_5264);
nand U6148 (N_6148,N_5259,N_5012);
xor U6149 (N_6149,N_5758,N_5461);
nor U6150 (N_6150,N_5529,N_5429);
xnor U6151 (N_6151,N_5011,N_5586);
xor U6152 (N_6152,N_5702,N_5302);
nor U6153 (N_6153,N_5930,N_5318);
nor U6154 (N_6154,N_5125,N_5880);
nand U6155 (N_6155,N_5232,N_5952);
nand U6156 (N_6156,N_5654,N_5672);
or U6157 (N_6157,N_5448,N_5009);
xor U6158 (N_6158,N_5220,N_5741);
and U6159 (N_6159,N_5808,N_5094);
nand U6160 (N_6160,N_5249,N_5874);
nor U6161 (N_6161,N_5953,N_5526);
xnor U6162 (N_6162,N_5479,N_5805);
xor U6163 (N_6163,N_5928,N_5982);
xor U6164 (N_6164,N_5118,N_5439);
nand U6165 (N_6165,N_5541,N_5082);
nand U6166 (N_6166,N_5941,N_5279);
and U6167 (N_6167,N_5188,N_5136);
nand U6168 (N_6168,N_5157,N_5107);
and U6169 (N_6169,N_5905,N_5046);
nand U6170 (N_6170,N_5932,N_5325);
or U6171 (N_6171,N_5247,N_5729);
and U6172 (N_6172,N_5614,N_5566);
or U6173 (N_6173,N_5020,N_5704);
xnor U6174 (N_6174,N_5113,N_5881);
or U6175 (N_6175,N_5962,N_5352);
xor U6176 (N_6176,N_5897,N_5948);
nand U6177 (N_6177,N_5445,N_5034);
nor U6178 (N_6178,N_5186,N_5134);
or U6179 (N_6179,N_5023,N_5241);
nor U6180 (N_6180,N_5301,N_5073);
nor U6181 (N_6181,N_5112,N_5025);
nand U6182 (N_6182,N_5161,N_5028);
and U6183 (N_6183,N_5579,N_5354);
nor U6184 (N_6184,N_5634,N_5057);
or U6185 (N_6185,N_5590,N_5485);
and U6186 (N_6186,N_5505,N_5806);
or U6187 (N_6187,N_5373,N_5549);
nand U6188 (N_6188,N_5430,N_5159);
xnor U6189 (N_6189,N_5454,N_5840);
nor U6190 (N_6190,N_5819,N_5338);
or U6191 (N_6191,N_5148,N_5471);
or U6192 (N_6192,N_5058,N_5747);
nor U6193 (N_6193,N_5346,N_5888);
nor U6194 (N_6194,N_5877,N_5945);
xnor U6195 (N_6195,N_5088,N_5061);
and U6196 (N_6196,N_5167,N_5635);
nand U6197 (N_6197,N_5145,N_5525);
and U6198 (N_6198,N_5477,N_5440);
or U6199 (N_6199,N_5506,N_5142);
xor U6200 (N_6200,N_5245,N_5467);
xnor U6201 (N_6201,N_5832,N_5916);
nand U6202 (N_6202,N_5603,N_5182);
xnor U6203 (N_6203,N_5363,N_5755);
and U6204 (N_6204,N_5804,N_5753);
or U6205 (N_6205,N_5434,N_5216);
and U6206 (N_6206,N_5764,N_5233);
xor U6207 (N_6207,N_5830,N_5333);
nor U6208 (N_6208,N_5108,N_5517);
nand U6209 (N_6209,N_5588,N_5098);
or U6210 (N_6210,N_5381,N_5649);
nand U6211 (N_6211,N_5743,N_5954);
nand U6212 (N_6212,N_5431,N_5814);
xnor U6213 (N_6213,N_5770,N_5867);
nor U6214 (N_6214,N_5978,N_5256);
or U6215 (N_6215,N_5695,N_5388);
or U6216 (N_6216,N_5597,N_5865);
nand U6217 (N_6217,N_5007,N_5871);
or U6218 (N_6218,N_5933,N_5782);
xnor U6219 (N_6219,N_5282,N_5504);
nand U6220 (N_6220,N_5294,N_5079);
nor U6221 (N_6221,N_5227,N_5097);
or U6222 (N_6222,N_5235,N_5074);
or U6223 (N_6223,N_5520,N_5487);
and U6224 (N_6224,N_5572,N_5385);
nand U6225 (N_6225,N_5372,N_5558);
nand U6226 (N_6226,N_5847,N_5324);
or U6227 (N_6227,N_5178,N_5260);
and U6228 (N_6228,N_5875,N_5542);
nor U6229 (N_6229,N_5211,N_5544);
and U6230 (N_6230,N_5133,N_5168);
or U6231 (N_6231,N_5665,N_5913);
nor U6232 (N_6232,N_5629,N_5298);
and U6233 (N_6233,N_5086,N_5956);
xor U6234 (N_6234,N_5272,N_5489);
or U6235 (N_6235,N_5795,N_5193);
nand U6236 (N_6236,N_5927,N_5931);
nand U6237 (N_6237,N_5749,N_5054);
xor U6238 (N_6238,N_5322,N_5285);
nand U6239 (N_6239,N_5055,N_5340);
and U6240 (N_6240,N_5547,N_5734);
and U6241 (N_6241,N_5550,N_5742);
nand U6242 (N_6242,N_5083,N_5828);
nand U6243 (N_6243,N_5026,N_5218);
nand U6244 (N_6244,N_5883,N_5185);
nor U6245 (N_6245,N_5616,N_5876);
or U6246 (N_6246,N_5474,N_5863);
nor U6247 (N_6247,N_5921,N_5700);
and U6248 (N_6248,N_5618,N_5064);
nand U6249 (N_6249,N_5117,N_5509);
nand U6250 (N_6250,N_5790,N_5608);
or U6251 (N_6251,N_5846,N_5468);
nor U6252 (N_6252,N_5172,N_5189);
and U6253 (N_6253,N_5581,N_5219);
nand U6254 (N_6254,N_5570,N_5656);
or U6255 (N_6255,N_5297,N_5473);
xor U6256 (N_6256,N_5103,N_5576);
xor U6257 (N_6257,N_5553,N_5457);
and U6258 (N_6258,N_5367,N_5419);
nor U6259 (N_6259,N_5815,N_5593);
nor U6260 (N_6260,N_5344,N_5378);
or U6261 (N_6261,N_5038,N_5250);
and U6262 (N_6262,N_5442,N_5246);
nor U6263 (N_6263,N_5253,N_5554);
nand U6264 (N_6264,N_5237,N_5273);
nand U6265 (N_6265,N_5709,N_5667);
nor U6266 (N_6266,N_5917,N_5416);
nor U6267 (N_6267,N_5065,N_5374);
or U6268 (N_6268,N_5037,N_5532);
or U6269 (N_6269,N_5132,N_5715);
nor U6270 (N_6270,N_5967,N_5140);
xnor U6271 (N_6271,N_5255,N_5958);
nand U6272 (N_6272,N_5304,N_5797);
or U6273 (N_6273,N_5432,N_5792);
xor U6274 (N_6274,N_5632,N_5619);
or U6275 (N_6275,N_5266,N_5756);
and U6276 (N_6276,N_5052,N_5173);
or U6277 (N_6277,N_5181,N_5929);
and U6278 (N_6278,N_5443,N_5886);
nor U6279 (N_6279,N_5834,N_5818);
xnor U6280 (N_6280,N_5609,N_5303);
nor U6281 (N_6281,N_5411,N_5100);
xor U6282 (N_6282,N_5405,N_5598);
xnor U6283 (N_6283,N_5224,N_5799);
nor U6284 (N_6284,N_5413,N_5056);
nor U6285 (N_6285,N_5309,N_5839);
xnor U6286 (N_6286,N_5452,N_5991);
or U6287 (N_6287,N_5280,N_5111);
or U6288 (N_6288,N_5415,N_5647);
nand U6289 (N_6289,N_5116,N_5370);
or U6290 (N_6290,N_5798,N_5018);
and U6291 (N_6291,N_5556,N_5854);
nor U6292 (N_6292,N_5447,N_5080);
xnor U6293 (N_6293,N_5720,N_5973);
xor U6294 (N_6294,N_5774,N_5321);
nor U6295 (N_6295,N_5949,N_5843);
or U6296 (N_6296,N_5120,N_5024);
and U6297 (N_6297,N_5663,N_5436);
nor U6298 (N_6298,N_5648,N_5825);
and U6299 (N_6299,N_5722,N_5214);
or U6300 (N_6300,N_5075,N_5143);
xor U6301 (N_6301,N_5393,N_5772);
and U6302 (N_6302,N_5675,N_5033);
nor U6303 (N_6303,N_5678,N_5651);
and U6304 (N_6304,N_5510,N_5491);
or U6305 (N_6305,N_5516,N_5032);
and U6306 (N_6306,N_5493,N_5557);
xor U6307 (N_6307,N_5677,N_5998);
and U6308 (N_6308,N_5010,N_5662);
nor U6309 (N_6309,N_5895,N_5230);
nor U6310 (N_6310,N_5592,N_5759);
nand U6311 (N_6311,N_5261,N_5723);
nand U6312 (N_6312,N_5934,N_5910);
nor U6313 (N_6313,N_5530,N_5882);
or U6314 (N_6314,N_5314,N_5652);
and U6315 (N_6315,N_5680,N_5206);
xnor U6316 (N_6316,N_5197,N_5964);
nor U6317 (N_6317,N_5195,N_5684);
xor U6318 (N_6318,N_5040,N_5169);
xor U6319 (N_6319,N_5987,N_5027);
or U6320 (N_6320,N_5070,N_5981);
nand U6321 (N_6321,N_5031,N_5767);
xnor U6322 (N_6322,N_5257,N_5152);
nor U6323 (N_6323,N_5306,N_5993);
nand U6324 (N_6324,N_5994,N_5740);
or U6325 (N_6325,N_5957,N_5922);
nor U6326 (N_6326,N_5906,N_5866);
nor U6327 (N_6327,N_5336,N_5131);
and U6328 (N_6328,N_5494,N_5511);
nor U6329 (N_6329,N_5555,N_5358);
or U6330 (N_6330,N_5644,N_5151);
and U6331 (N_6331,N_5085,N_5942);
or U6332 (N_6332,N_5898,N_5595);
or U6333 (N_6333,N_5809,N_5053);
or U6334 (N_6334,N_5548,N_5611);
and U6335 (N_6335,N_5424,N_5682);
xor U6336 (N_6336,N_5029,N_5621);
xor U6337 (N_6337,N_5596,N_5859);
nor U6338 (N_6338,N_5162,N_5089);
and U6339 (N_6339,N_5258,N_5926);
xor U6340 (N_6340,N_5175,N_5841);
or U6341 (N_6341,N_5890,N_5691);
or U6342 (N_6342,N_5763,N_5900);
nor U6343 (N_6343,N_5119,N_5698);
xnor U6344 (N_6344,N_5653,N_5985);
nor U6345 (N_6345,N_5685,N_5102);
nor U6346 (N_6346,N_5062,N_5158);
xnor U6347 (N_6347,N_5137,N_5674);
nand U6348 (N_6348,N_5963,N_5236);
or U6349 (N_6349,N_5513,N_5777);
nand U6350 (N_6350,N_5495,N_5845);
and U6351 (N_6351,N_5426,N_5343);
nor U6352 (N_6352,N_5971,N_5984);
and U6353 (N_6353,N_5500,N_5631);
nand U6354 (N_6354,N_5200,N_5400);
xnor U6355 (N_6355,N_5668,N_5329);
nor U6356 (N_6356,N_5748,N_5293);
or U6357 (N_6357,N_5717,N_5276);
xnor U6358 (N_6358,N_5670,N_5409);
or U6359 (N_6359,N_5042,N_5754);
nor U6360 (N_6360,N_5655,N_5150);
or U6361 (N_6361,N_5523,N_5166);
and U6362 (N_6362,N_5503,N_5090);
or U6363 (N_6363,N_5295,N_5077);
nor U6364 (N_6364,N_5290,N_5524);
xor U6365 (N_6365,N_5371,N_5463);
or U6366 (N_6366,N_5252,N_5752);
and U6367 (N_6367,N_5417,N_5396);
and U6368 (N_6368,N_5482,N_5190);
or U6369 (N_6369,N_5669,N_5707);
nand U6370 (N_6370,N_5620,N_5924);
nand U6371 (N_6371,N_5671,N_5801);
nor U6372 (N_6372,N_5661,N_5820);
nor U6373 (N_6373,N_5003,N_5710);
nor U6374 (N_6374,N_5833,N_5893);
or U6375 (N_6375,N_5849,N_5796);
nor U6376 (N_6376,N_5873,N_5005);
and U6377 (N_6377,N_5450,N_5514);
nor U6378 (N_6378,N_5016,N_5728);
and U6379 (N_6379,N_5522,N_5486);
and U6380 (N_6380,N_5422,N_5896);
nand U6381 (N_6381,N_5435,N_5794);
nor U6382 (N_6382,N_5658,N_5222);
or U6383 (N_6383,N_5688,N_5735);
or U6384 (N_6384,N_5458,N_5760);
or U6385 (N_6385,N_5965,N_5305);
xor U6386 (N_6386,N_5659,N_5147);
xor U6387 (N_6387,N_5316,N_5853);
nor U6388 (N_6388,N_5730,N_5239);
or U6389 (N_6389,N_5044,N_5975);
xnor U6390 (N_6390,N_5271,N_5141);
or U6391 (N_6391,N_5976,N_5793);
or U6392 (N_6392,N_5947,N_5673);
and U6393 (N_6393,N_5563,N_5571);
xnor U6394 (N_6394,N_5515,N_5022);
or U6395 (N_6395,N_5192,N_5014);
nor U6396 (N_6396,N_5441,N_5427);
nor U6397 (N_6397,N_5403,N_5826);
and U6398 (N_6398,N_5773,N_5499);
nor U6399 (N_6399,N_5650,N_5899);
nand U6400 (N_6400,N_5950,N_5751);
and U6401 (N_6401,N_5936,N_5153);
nor U6402 (N_6402,N_5418,N_5421);
xnor U6403 (N_6403,N_5645,N_5869);
xnor U6404 (N_6404,N_5263,N_5911);
or U6405 (N_6405,N_5918,N_5030);
xor U6406 (N_6406,N_5015,N_5779);
or U6407 (N_6407,N_5359,N_5231);
nor U6408 (N_6408,N_5537,N_5891);
nand U6409 (N_6409,N_5287,N_5810);
nand U6410 (N_6410,N_5198,N_5311);
nor U6411 (N_6411,N_5347,N_5961);
xor U6412 (N_6412,N_5328,N_5254);
xnor U6413 (N_6413,N_5855,N_5171);
nor U6414 (N_6414,N_5047,N_5714);
and U6415 (N_6415,N_5573,N_5229);
xor U6416 (N_6416,N_5242,N_5745);
nand U6417 (N_6417,N_5683,N_5223);
xor U6418 (N_6418,N_5769,N_5394);
nand U6419 (N_6419,N_5323,N_5870);
xnor U6420 (N_6420,N_5589,N_5686);
and U6421 (N_6421,N_5716,N_5277);
xor U6422 (N_6422,N_5384,N_5543);
nand U6423 (N_6423,N_5736,N_5128);
and U6424 (N_6424,N_5049,N_5679);
xnor U6425 (N_6425,N_5362,N_5050);
nor U6426 (N_6426,N_5559,N_5778);
nand U6427 (N_6427,N_5641,N_5803);
xnor U6428 (N_6428,N_5565,N_5536);
nor U6429 (N_6429,N_5360,N_5110);
xor U6430 (N_6430,N_5196,N_5605);
and U6431 (N_6431,N_5638,N_5690);
and U6432 (N_6432,N_5560,N_5395);
nor U6433 (N_6433,N_5807,N_5713);
xor U6434 (N_6434,N_5288,N_5459);
nor U6435 (N_6435,N_5490,N_5862);
or U6436 (N_6436,N_5194,N_5995);
or U6437 (N_6437,N_5453,N_5837);
nand U6438 (N_6438,N_5350,N_5203);
and U6439 (N_6439,N_5724,N_5901);
or U6440 (N_6440,N_5437,N_5528);
nor U6441 (N_6441,N_5095,N_5594);
nor U6442 (N_6442,N_5788,N_5731);
nand U6443 (N_6443,N_5765,N_5507);
nand U6444 (N_6444,N_5154,N_5583);
xor U6445 (N_6445,N_5838,N_5096);
or U6446 (N_6446,N_5983,N_5817);
and U6447 (N_6447,N_5124,N_5636);
or U6448 (N_6448,N_5334,N_5535);
or U6449 (N_6449,N_5909,N_5274);
or U6450 (N_6450,N_5584,N_5602);
or U6451 (N_6451,N_5829,N_5414);
nand U6452 (N_6452,N_5377,N_5946);
or U6453 (N_6453,N_5179,N_5923);
nand U6454 (N_6454,N_5238,N_5234);
or U6455 (N_6455,N_5008,N_5296);
and U6456 (N_6456,N_5860,N_5183);
and U6457 (N_6457,N_5703,N_5209);
or U6458 (N_6458,N_5750,N_5824);
nor U6459 (N_6459,N_5013,N_5539);
xnor U6460 (N_6460,N_5567,N_5640);
and U6461 (N_6461,N_5986,N_5345);
or U6462 (N_6462,N_5712,N_5478);
or U6463 (N_6463,N_5768,N_5781);
nand U6464 (N_6464,N_5319,N_5575);
nor U6465 (N_6465,N_5039,N_5213);
nand U6466 (N_6466,N_5492,N_5144);
or U6467 (N_6467,N_5604,N_5907);
xor U6468 (N_6468,N_5761,N_5540);
and U6469 (N_6469,N_5339,N_5727);
or U6470 (N_6470,N_5999,N_5912);
or U6471 (N_6471,N_5666,N_5164);
or U6472 (N_6472,N_5310,N_5469);
or U6473 (N_6473,N_5574,N_5938);
xor U6474 (N_6474,N_5708,N_5099);
and U6475 (N_6475,N_5811,N_5915);
xnor U6476 (N_6476,N_5546,N_5626);
nand U6477 (N_6477,N_5726,N_5944);
nor U6478 (N_6478,N_5122,N_5568);
nand U6479 (N_6479,N_5308,N_5330);
xor U6480 (N_6480,N_5534,N_5402);
or U6481 (N_6481,N_5601,N_5955);
nor U6482 (N_6482,N_5139,N_5379);
nor U6483 (N_6483,N_5879,N_5784);
or U6484 (N_6484,N_5725,N_5035);
nor U6485 (N_6485,N_5067,N_5607);
and U6486 (N_6486,N_5827,N_5600);
and U6487 (N_6487,N_5789,N_5135);
and U6488 (N_6488,N_5787,N_5348);
nand U6489 (N_6489,N_5693,N_5387);
or U6490 (N_6490,N_5270,N_5692);
and U6491 (N_6491,N_5313,N_5204);
nor U6492 (N_6492,N_5483,N_5069);
and U6493 (N_6493,N_5281,N_5208);
or U6494 (N_6494,N_5561,N_5775);
nand U6495 (N_6495,N_5355,N_5326);
and U6496 (N_6496,N_5943,N_5357);
nor U6497 (N_6497,N_5176,N_5087);
and U6498 (N_6498,N_5615,N_5701);
nand U6499 (N_6499,N_5187,N_5771);
xor U6500 (N_6500,N_5848,N_5514);
or U6501 (N_6501,N_5241,N_5049);
xnor U6502 (N_6502,N_5104,N_5301);
and U6503 (N_6503,N_5798,N_5963);
or U6504 (N_6504,N_5799,N_5123);
xor U6505 (N_6505,N_5770,N_5166);
and U6506 (N_6506,N_5814,N_5572);
xor U6507 (N_6507,N_5048,N_5680);
xnor U6508 (N_6508,N_5992,N_5877);
xnor U6509 (N_6509,N_5966,N_5701);
xor U6510 (N_6510,N_5332,N_5064);
nor U6511 (N_6511,N_5566,N_5616);
or U6512 (N_6512,N_5726,N_5443);
xor U6513 (N_6513,N_5551,N_5069);
and U6514 (N_6514,N_5560,N_5500);
or U6515 (N_6515,N_5408,N_5198);
and U6516 (N_6516,N_5864,N_5543);
nand U6517 (N_6517,N_5312,N_5684);
nor U6518 (N_6518,N_5973,N_5452);
nand U6519 (N_6519,N_5369,N_5539);
and U6520 (N_6520,N_5156,N_5016);
xor U6521 (N_6521,N_5252,N_5904);
nor U6522 (N_6522,N_5853,N_5539);
or U6523 (N_6523,N_5481,N_5795);
or U6524 (N_6524,N_5139,N_5771);
nand U6525 (N_6525,N_5073,N_5971);
nor U6526 (N_6526,N_5232,N_5972);
and U6527 (N_6527,N_5684,N_5052);
and U6528 (N_6528,N_5309,N_5217);
or U6529 (N_6529,N_5832,N_5532);
xor U6530 (N_6530,N_5035,N_5819);
xor U6531 (N_6531,N_5295,N_5192);
xor U6532 (N_6532,N_5604,N_5987);
nor U6533 (N_6533,N_5455,N_5208);
nand U6534 (N_6534,N_5024,N_5953);
and U6535 (N_6535,N_5328,N_5610);
nand U6536 (N_6536,N_5634,N_5463);
and U6537 (N_6537,N_5543,N_5002);
and U6538 (N_6538,N_5348,N_5130);
nand U6539 (N_6539,N_5156,N_5674);
xor U6540 (N_6540,N_5126,N_5548);
nor U6541 (N_6541,N_5769,N_5371);
nor U6542 (N_6542,N_5246,N_5981);
and U6543 (N_6543,N_5484,N_5005);
nor U6544 (N_6544,N_5654,N_5548);
or U6545 (N_6545,N_5638,N_5206);
or U6546 (N_6546,N_5019,N_5258);
nor U6547 (N_6547,N_5165,N_5804);
xnor U6548 (N_6548,N_5045,N_5740);
nand U6549 (N_6549,N_5125,N_5024);
xnor U6550 (N_6550,N_5992,N_5925);
or U6551 (N_6551,N_5943,N_5601);
and U6552 (N_6552,N_5227,N_5249);
nand U6553 (N_6553,N_5541,N_5670);
nor U6554 (N_6554,N_5689,N_5621);
nor U6555 (N_6555,N_5644,N_5871);
or U6556 (N_6556,N_5717,N_5713);
or U6557 (N_6557,N_5817,N_5953);
and U6558 (N_6558,N_5186,N_5503);
nand U6559 (N_6559,N_5362,N_5019);
xnor U6560 (N_6560,N_5788,N_5534);
xor U6561 (N_6561,N_5719,N_5049);
nor U6562 (N_6562,N_5047,N_5895);
and U6563 (N_6563,N_5300,N_5645);
nand U6564 (N_6564,N_5133,N_5050);
and U6565 (N_6565,N_5062,N_5584);
xnor U6566 (N_6566,N_5340,N_5605);
nand U6567 (N_6567,N_5414,N_5981);
and U6568 (N_6568,N_5016,N_5065);
nand U6569 (N_6569,N_5961,N_5149);
nor U6570 (N_6570,N_5077,N_5600);
nor U6571 (N_6571,N_5278,N_5387);
nand U6572 (N_6572,N_5033,N_5430);
or U6573 (N_6573,N_5147,N_5433);
or U6574 (N_6574,N_5714,N_5189);
nand U6575 (N_6575,N_5347,N_5281);
xnor U6576 (N_6576,N_5135,N_5519);
nor U6577 (N_6577,N_5781,N_5970);
xor U6578 (N_6578,N_5555,N_5759);
or U6579 (N_6579,N_5813,N_5598);
nor U6580 (N_6580,N_5773,N_5772);
xnor U6581 (N_6581,N_5534,N_5552);
xnor U6582 (N_6582,N_5043,N_5855);
or U6583 (N_6583,N_5605,N_5032);
nor U6584 (N_6584,N_5748,N_5544);
xnor U6585 (N_6585,N_5274,N_5141);
or U6586 (N_6586,N_5650,N_5747);
and U6587 (N_6587,N_5937,N_5952);
xor U6588 (N_6588,N_5469,N_5352);
nor U6589 (N_6589,N_5590,N_5497);
or U6590 (N_6590,N_5384,N_5839);
or U6591 (N_6591,N_5704,N_5460);
nand U6592 (N_6592,N_5111,N_5347);
or U6593 (N_6593,N_5211,N_5617);
and U6594 (N_6594,N_5078,N_5251);
nor U6595 (N_6595,N_5883,N_5972);
xnor U6596 (N_6596,N_5596,N_5537);
nor U6597 (N_6597,N_5233,N_5652);
nor U6598 (N_6598,N_5144,N_5414);
or U6599 (N_6599,N_5876,N_5859);
nand U6600 (N_6600,N_5416,N_5533);
nor U6601 (N_6601,N_5218,N_5443);
or U6602 (N_6602,N_5052,N_5993);
xor U6603 (N_6603,N_5247,N_5615);
nor U6604 (N_6604,N_5454,N_5615);
nor U6605 (N_6605,N_5199,N_5171);
xnor U6606 (N_6606,N_5353,N_5987);
nand U6607 (N_6607,N_5990,N_5531);
xnor U6608 (N_6608,N_5342,N_5577);
and U6609 (N_6609,N_5261,N_5547);
and U6610 (N_6610,N_5433,N_5157);
nor U6611 (N_6611,N_5347,N_5818);
and U6612 (N_6612,N_5637,N_5734);
and U6613 (N_6613,N_5568,N_5986);
and U6614 (N_6614,N_5129,N_5965);
xor U6615 (N_6615,N_5820,N_5044);
nor U6616 (N_6616,N_5793,N_5197);
or U6617 (N_6617,N_5924,N_5048);
nor U6618 (N_6618,N_5677,N_5834);
nand U6619 (N_6619,N_5613,N_5242);
nand U6620 (N_6620,N_5751,N_5147);
nand U6621 (N_6621,N_5814,N_5712);
and U6622 (N_6622,N_5392,N_5469);
or U6623 (N_6623,N_5886,N_5257);
nand U6624 (N_6624,N_5200,N_5837);
nand U6625 (N_6625,N_5405,N_5822);
nor U6626 (N_6626,N_5377,N_5703);
or U6627 (N_6627,N_5405,N_5916);
and U6628 (N_6628,N_5378,N_5616);
xnor U6629 (N_6629,N_5760,N_5987);
or U6630 (N_6630,N_5376,N_5176);
xor U6631 (N_6631,N_5528,N_5253);
nor U6632 (N_6632,N_5895,N_5522);
or U6633 (N_6633,N_5827,N_5326);
nand U6634 (N_6634,N_5235,N_5092);
or U6635 (N_6635,N_5854,N_5246);
and U6636 (N_6636,N_5760,N_5071);
and U6637 (N_6637,N_5510,N_5068);
nor U6638 (N_6638,N_5812,N_5461);
xnor U6639 (N_6639,N_5797,N_5849);
or U6640 (N_6640,N_5258,N_5975);
nand U6641 (N_6641,N_5424,N_5568);
nand U6642 (N_6642,N_5049,N_5309);
nand U6643 (N_6643,N_5461,N_5685);
nand U6644 (N_6644,N_5376,N_5786);
nand U6645 (N_6645,N_5709,N_5352);
and U6646 (N_6646,N_5829,N_5378);
nand U6647 (N_6647,N_5353,N_5798);
nand U6648 (N_6648,N_5984,N_5593);
and U6649 (N_6649,N_5206,N_5129);
and U6650 (N_6650,N_5204,N_5953);
nor U6651 (N_6651,N_5365,N_5115);
or U6652 (N_6652,N_5605,N_5125);
nor U6653 (N_6653,N_5275,N_5451);
and U6654 (N_6654,N_5547,N_5153);
or U6655 (N_6655,N_5461,N_5161);
or U6656 (N_6656,N_5874,N_5286);
and U6657 (N_6657,N_5237,N_5505);
nand U6658 (N_6658,N_5672,N_5721);
xnor U6659 (N_6659,N_5353,N_5546);
nor U6660 (N_6660,N_5103,N_5023);
nor U6661 (N_6661,N_5158,N_5990);
nand U6662 (N_6662,N_5235,N_5846);
nand U6663 (N_6663,N_5715,N_5363);
nand U6664 (N_6664,N_5608,N_5558);
and U6665 (N_6665,N_5233,N_5901);
nand U6666 (N_6666,N_5623,N_5922);
xnor U6667 (N_6667,N_5552,N_5266);
or U6668 (N_6668,N_5643,N_5739);
or U6669 (N_6669,N_5716,N_5016);
and U6670 (N_6670,N_5841,N_5814);
or U6671 (N_6671,N_5569,N_5816);
nor U6672 (N_6672,N_5489,N_5521);
or U6673 (N_6673,N_5163,N_5553);
nor U6674 (N_6674,N_5716,N_5824);
nand U6675 (N_6675,N_5007,N_5066);
or U6676 (N_6676,N_5342,N_5009);
nand U6677 (N_6677,N_5732,N_5744);
xor U6678 (N_6678,N_5600,N_5898);
and U6679 (N_6679,N_5366,N_5708);
or U6680 (N_6680,N_5472,N_5958);
xnor U6681 (N_6681,N_5518,N_5714);
or U6682 (N_6682,N_5732,N_5143);
or U6683 (N_6683,N_5731,N_5474);
or U6684 (N_6684,N_5007,N_5099);
nand U6685 (N_6685,N_5206,N_5900);
and U6686 (N_6686,N_5439,N_5302);
or U6687 (N_6687,N_5968,N_5626);
and U6688 (N_6688,N_5924,N_5215);
nor U6689 (N_6689,N_5782,N_5175);
xor U6690 (N_6690,N_5447,N_5546);
xor U6691 (N_6691,N_5476,N_5613);
nor U6692 (N_6692,N_5080,N_5514);
and U6693 (N_6693,N_5453,N_5118);
or U6694 (N_6694,N_5161,N_5926);
and U6695 (N_6695,N_5324,N_5370);
nand U6696 (N_6696,N_5898,N_5765);
xor U6697 (N_6697,N_5623,N_5297);
or U6698 (N_6698,N_5117,N_5883);
nand U6699 (N_6699,N_5364,N_5522);
nor U6700 (N_6700,N_5731,N_5004);
and U6701 (N_6701,N_5463,N_5402);
nand U6702 (N_6702,N_5700,N_5075);
nor U6703 (N_6703,N_5083,N_5989);
nor U6704 (N_6704,N_5038,N_5947);
nor U6705 (N_6705,N_5498,N_5020);
or U6706 (N_6706,N_5991,N_5269);
nand U6707 (N_6707,N_5635,N_5049);
nor U6708 (N_6708,N_5189,N_5681);
xnor U6709 (N_6709,N_5626,N_5741);
and U6710 (N_6710,N_5499,N_5981);
xnor U6711 (N_6711,N_5694,N_5518);
or U6712 (N_6712,N_5445,N_5759);
xor U6713 (N_6713,N_5081,N_5144);
and U6714 (N_6714,N_5299,N_5304);
xnor U6715 (N_6715,N_5080,N_5262);
xor U6716 (N_6716,N_5800,N_5771);
xor U6717 (N_6717,N_5038,N_5450);
nor U6718 (N_6718,N_5659,N_5629);
nor U6719 (N_6719,N_5293,N_5611);
and U6720 (N_6720,N_5589,N_5327);
nand U6721 (N_6721,N_5533,N_5858);
or U6722 (N_6722,N_5630,N_5148);
and U6723 (N_6723,N_5250,N_5579);
nor U6724 (N_6724,N_5520,N_5210);
and U6725 (N_6725,N_5516,N_5351);
nand U6726 (N_6726,N_5664,N_5776);
nand U6727 (N_6727,N_5035,N_5597);
nor U6728 (N_6728,N_5106,N_5749);
or U6729 (N_6729,N_5412,N_5462);
nand U6730 (N_6730,N_5205,N_5722);
nor U6731 (N_6731,N_5009,N_5901);
or U6732 (N_6732,N_5132,N_5284);
or U6733 (N_6733,N_5443,N_5795);
and U6734 (N_6734,N_5026,N_5735);
or U6735 (N_6735,N_5341,N_5832);
and U6736 (N_6736,N_5707,N_5818);
nand U6737 (N_6737,N_5983,N_5724);
nor U6738 (N_6738,N_5140,N_5556);
nand U6739 (N_6739,N_5988,N_5263);
xnor U6740 (N_6740,N_5573,N_5496);
nor U6741 (N_6741,N_5486,N_5343);
or U6742 (N_6742,N_5945,N_5169);
nand U6743 (N_6743,N_5476,N_5099);
or U6744 (N_6744,N_5347,N_5906);
or U6745 (N_6745,N_5880,N_5416);
nand U6746 (N_6746,N_5118,N_5242);
nand U6747 (N_6747,N_5535,N_5325);
or U6748 (N_6748,N_5378,N_5645);
nand U6749 (N_6749,N_5406,N_5303);
xor U6750 (N_6750,N_5182,N_5685);
or U6751 (N_6751,N_5694,N_5324);
or U6752 (N_6752,N_5079,N_5778);
or U6753 (N_6753,N_5319,N_5798);
nor U6754 (N_6754,N_5335,N_5569);
and U6755 (N_6755,N_5450,N_5139);
nor U6756 (N_6756,N_5757,N_5674);
nand U6757 (N_6757,N_5370,N_5847);
xor U6758 (N_6758,N_5697,N_5240);
nor U6759 (N_6759,N_5339,N_5981);
and U6760 (N_6760,N_5716,N_5340);
and U6761 (N_6761,N_5532,N_5398);
nor U6762 (N_6762,N_5739,N_5913);
xor U6763 (N_6763,N_5556,N_5067);
and U6764 (N_6764,N_5209,N_5113);
and U6765 (N_6765,N_5591,N_5588);
and U6766 (N_6766,N_5275,N_5249);
nor U6767 (N_6767,N_5313,N_5253);
or U6768 (N_6768,N_5216,N_5530);
nor U6769 (N_6769,N_5912,N_5082);
nand U6770 (N_6770,N_5832,N_5507);
and U6771 (N_6771,N_5293,N_5390);
xor U6772 (N_6772,N_5187,N_5448);
xnor U6773 (N_6773,N_5713,N_5950);
and U6774 (N_6774,N_5400,N_5774);
nor U6775 (N_6775,N_5013,N_5567);
nor U6776 (N_6776,N_5225,N_5920);
or U6777 (N_6777,N_5844,N_5108);
and U6778 (N_6778,N_5082,N_5067);
or U6779 (N_6779,N_5327,N_5041);
and U6780 (N_6780,N_5937,N_5130);
and U6781 (N_6781,N_5077,N_5401);
or U6782 (N_6782,N_5330,N_5125);
nand U6783 (N_6783,N_5341,N_5393);
or U6784 (N_6784,N_5291,N_5154);
nor U6785 (N_6785,N_5564,N_5215);
nand U6786 (N_6786,N_5235,N_5264);
or U6787 (N_6787,N_5361,N_5576);
or U6788 (N_6788,N_5751,N_5340);
xor U6789 (N_6789,N_5955,N_5213);
xnor U6790 (N_6790,N_5791,N_5563);
nand U6791 (N_6791,N_5116,N_5165);
nand U6792 (N_6792,N_5374,N_5912);
nor U6793 (N_6793,N_5984,N_5393);
or U6794 (N_6794,N_5381,N_5728);
and U6795 (N_6795,N_5251,N_5211);
nand U6796 (N_6796,N_5011,N_5024);
nor U6797 (N_6797,N_5110,N_5319);
nor U6798 (N_6798,N_5567,N_5156);
and U6799 (N_6799,N_5969,N_5345);
nand U6800 (N_6800,N_5017,N_5692);
nand U6801 (N_6801,N_5254,N_5778);
nor U6802 (N_6802,N_5645,N_5195);
xnor U6803 (N_6803,N_5368,N_5644);
nand U6804 (N_6804,N_5198,N_5716);
and U6805 (N_6805,N_5134,N_5399);
nor U6806 (N_6806,N_5869,N_5260);
or U6807 (N_6807,N_5353,N_5925);
xnor U6808 (N_6808,N_5013,N_5612);
or U6809 (N_6809,N_5804,N_5395);
xnor U6810 (N_6810,N_5986,N_5044);
xnor U6811 (N_6811,N_5359,N_5973);
and U6812 (N_6812,N_5665,N_5525);
nand U6813 (N_6813,N_5456,N_5514);
nor U6814 (N_6814,N_5117,N_5559);
or U6815 (N_6815,N_5590,N_5381);
nand U6816 (N_6816,N_5512,N_5013);
xor U6817 (N_6817,N_5585,N_5409);
or U6818 (N_6818,N_5805,N_5860);
or U6819 (N_6819,N_5308,N_5440);
nand U6820 (N_6820,N_5897,N_5879);
nor U6821 (N_6821,N_5645,N_5791);
xnor U6822 (N_6822,N_5830,N_5691);
or U6823 (N_6823,N_5430,N_5200);
nand U6824 (N_6824,N_5519,N_5173);
and U6825 (N_6825,N_5296,N_5787);
nor U6826 (N_6826,N_5780,N_5223);
or U6827 (N_6827,N_5631,N_5950);
and U6828 (N_6828,N_5336,N_5465);
or U6829 (N_6829,N_5104,N_5025);
and U6830 (N_6830,N_5449,N_5873);
or U6831 (N_6831,N_5988,N_5742);
and U6832 (N_6832,N_5146,N_5838);
nand U6833 (N_6833,N_5127,N_5761);
or U6834 (N_6834,N_5852,N_5054);
nor U6835 (N_6835,N_5482,N_5478);
and U6836 (N_6836,N_5050,N_5968);
and U6837 (N_6837,N_5820,N_5349);
xnor U6838 (N_6838,N_5779,N_5877);
and U6839 (N_6839,N_5701,N_5246);
xnor U6840 (N_6840,N_5712,N_5082);
nand U6841 (N_6841,N_5528,N_5148);
nor U6842 (N_6842,N_5266,N_5634);
nand U6843 (N_6843,N_5020,N_5481);
xor U6844 (N_6844,N_5431,N_5089);
xnor U6845 (N_6845,N_5615,N_5012);
nor U6846 (N_6846,N_5176,N_5130);
and U6847 (N_6847,N_5532,N_5693);
and U6848 (N_6848,N_5193,N_5944);
nand U6849 (N_6849,N_5086,N_5397);
nand U6850 (N_6850,N_5173,N_5909);
nor U6851 (N_6851,N_5409,N_5488);
or U6852 (N_6852,N_5367,N_5177);
xor U6853 (N_6853,N_5475,N_5743);
nand U6854 (N_6854,N_5722,N_5965);
or U6855 (N_6855,N_5746,N_5781);
nor U6856 (N_6856,N_5030,N_5380);
or U6857 (N_6857,N_5186,N_5489);
or U6858 (N_6858,N_5272,N_5876);
nor U6859 (N_6859,N_5150,N_5977);
or U6860 (N_6860,N_5302,N_5954);
nand U6861 (N_6861,N_5432,N_5355);
nand U6862 (N_6862,N_5526,N_5229);
nor U6863 (N_6863,N_5044,N_5252);
and U6864 (N_6864,N_5752,N_5765);
nor U6865 (N_6865,N_5249,N_5757);
nand U6866 (N_6866,N_5190,N_5241);
and U6867 (N_6867,N_5175,N_5402);
or U6868 (N_6868,N_5866,N_5137);
or U6869 (N_6869,N_5441,N_5615);
and U6870 (N_6870,N_5360,N_5926);
xnor U6871 (N_6871,N_5013,N_5399);
and U6872 (N_6872,N_5119,N_5328);
nor U6873 (N_6873,N_5953,N_5954);
nor U6874 (N_6874,N_5719,N_5894);
or U6875 (N_6875,N_5456,N_5043);
xor U6876 (N_6876,N_5641,N_5764);
nand U6877 (N_6877,N_5813,N_5728);
and U6878 (N_6878,N_5200,N_5533);
or U6879 (N_6879,N_5201,N_5635);
nand U6880 (N_6880,N_5974,N_5834);
nor U6881 (N_6881,N_5796,N_5222);
xnor U6882 (N_6882,N_5910,N_5573);
or U6883 (N_6883,N_5224,N_5991);
and U6884 (N_6884,N_5507,N_5857);
nor U6885 (N_6885,N_5546,N_5048);
and U6886 (N_6886,N_5230,N_5022);
nand U6887 (N_6887,N_5593,N_5591);
or U6888 (N_6888,N_5234,N_5541);
nand U6889 (N_6889,N_5058,N_5510);
nor U6890 (N_6890,N_5187,N_5806);
nand U6891 (N_6891,N_5567,N_5937);
xnor U6892 (N_6892,N_5740,N_5301);
nor U6893 (N_6893,N_5733,N_5924);
and U6894 (N_6894,N_5354,N_5441);
or U6895 (N_6895,N_5956,N_5217);
nand U6896 (N_6896,N_5403,N_5880);
nand U6897 (N_6897,N_5399,N_5855);
nor U6898 (N_6898,N_5587,N_5042);
nor U6899 (N_6899,N_5073,N_5386);
and U6900 (N_6900,N_5556,N_5252);
and U6901 (N_6901,N_5365,N_5755);
nor U6902 (N_6902,N_5526,N_5245);
xnor U6903 (N_6903,N_5637,N_5020);
and U6904 (N_6904,N_5897,N_5451);
xor U6905 (N_6905,N_5436,N_5871);
nor U6906 (N_6906,N_5134,N_5954);
nor U6907 (N_6907,N_5425,N_5435);
and U6908 (N_6908,N_5338,N_5600);
nand U6909 (N_6909,N_5953,N_5042);
or U6910 (N_6910,N_5319,N_5288);
and U6911 (N_6911,N_5340,N_5519);
nand U6912 (N_6912,N_5890,N_5028);
xnor U6913 (N_6913,N_5824,N_5585);
xor U6914 (N_6914,N_5301,N_5523);
or U6915 (N_6915,N_5570,N_5400);
nor U6916 (N_6916,N_5496,N_5786);
xor U6917 (N_6917,N_5198,N_5025);
nor U6918 (N_6918,N_5005,N_5229);
nand U6919 (N_6919,N_5905,N_5128);
nand U6920 (N_6920,N_5433,N_5102);
and U6921 (N_6921,N_5988,N_5866);
nand U6922 (N_6922,N_5253,N_5521);
xnor U6923 (N_6923,N_5922,N_5872);
nand U6924 (N_6924,N_5035,N_5745);
nor U6925 (N_6925,N_5458,N_5879);
nor U6926 (N_6926,N_5917,N_5421);
and U6927 (N_6927,N_5427,N_5822);
nor U6928 (N_6928,N_5596,N_5363);
and U6929 (N_6929,N_5943,N_5108);
xor U6930 (N_6930,N_5399,N_5773);
nor U6931 (N_6931,N_5774,N_5136);
and U6932 (N_6932,N_5887,N_5231);
nor U6933 (N_6933,N_5789,N_5838);
nor U6934 (N_6934,N_5566,N_5360);
and U6935 (N_6935,N_5978,N_5789);
nand U6936 (N_6936,N_5557,N_5201);
nor U6937 (N_6937,N_5097,N_5112);
and U6938 (N_6938,N_5485,N_5191);
nor U6939 (N_6939,N_5510,N_5668);
and U6940 (N_6940,N_5419,N_5910);
nor U6941 (N_6941,N_5881,N_5707);
or U6942 (N_6942,N_5186,N_5700);
and U6943 (N_6943,N_5182,N_5527);
xor U6944 (N_6944,N_5188,N_5249);
and U6945 (N_6945,N_5901,N_5864);
or U6946 (N_6946,N_5372,N_5473);
xor U6947 (N_6947,N_5155,N_5888);
nand U6948 (N_6948,N_5133,N_5602);
or U6949 (N_6949,N_5760,N_5248);
or U6950 (N_6950,N_5975,N_5406);
nand U6951 (N_6951,N_5377,N_5323);
and U6952 (N_6952,N_5582,N_5921);
xor U6953 (N_6953,N_5353,N_5205);
nand U6954 (N_6954,N_5532,N_5272);
and U6955 (N_6955,N_5862,N_5361);
xnor U6956 (N_6956,N_5410,N_5069);
and U6957 (N_6957,N_5750,N_5689);
or U6958 (N_6958,N_5326,N_5586);
or U6959 (N_6959,N_5898,N_5960);
nand U6960 (N_6960,N_5041,N_5978);
and U6961 (N_6961,N_5614,N_5779);
nand U6962 (N_6962,N_5124,N_5227);
nor U6963 (N_6963,N_5153,N_5248);
nor U6964 (N_6964,N_5834,N_5638);
xnor U6965 (N_6965,N_5061,N_5142);
and U6966 (N_6966,N_5402,N_5719);
and U6967 (N_6967,N_5084,N_5125);
or U6968 (N_6968,N_5384,N_5663);
xor U6969 (N_6969,N_5894,N_5559);
or U6970 (N_6970,N_5984,N_5478);
xor U6971 (N_6971,N_5922,N_5566);
or U6972 (N_6972,N_5526,N_5989);
or U6973 (N_6973,N_5732,N_5979);
and U6974 (N_6974,N_5278,N_5431);
nand U6975 (N_6975,N_5623,N_5820);
nor U6976 (N_6976,N_5546,N_5523);
nand U6977 (N_6977,N_5800,N_5117);
nor U6978 (N_6978,N_5524,N_5536);
nor U6979 (N_6979,N_5342,N_5072);
nor U6980 (N_6980,N_5204,N_5496);
nor U6981 (N_6981,N_5654,N_5928);
xor U6982 (N_6982,N_5487,N_5998);
nand U6983 (N_6983,N_5936,N_5583);
nor U6984 (N_6984,N_5246,N_5705);
or U6985 (N_6985,N_5026,N_5244);
nor U6986 (N_6986,N_5728,N_5839);
and U6987 (N_6987,N_5113,N_5825);
nand U6988 (N_6988,N_5172,N_5210);
nand U6989 (N_6989,N_5469,N_5140);
nand U6990 (N_6990,N_5019,N_5834);
nor U6991 (N_6991,N_5535,N_5580);
nor U6992 (N_6992,N_5309,N_5778);
or U6993 (N_6993,N_5930,N_5128);
nor U6994 (N_6994,N_5430,N_5784);
nor U6995 (N_6995,N_5224,N_5476);
nand U6996 (N_6996,N_5331,N_5831);
xnor U6997 (N_6997,N_5725,N_5879);
xor U6998 (N_6998,N_5385,N_5389);
and U6999 (N_6999,N_5872,N_5522);
nand U7000 (N_7000,N_6179,N_6505);
nor U7001 (N_7001,N_6522,N_6339);
and U7002 (N_7002,N_6013,N_6123);
and U7003 (N_7003,N_6661,N_6713);
xnor U7004 (N_7004,N_6251,N_6033);
xor U7005 (N_7005,N_6072,N_6605);
and U7006 (N_7006,N_6978,N_6308);
or U7007 (N_7007,N_6675,N_6940);
xor U7008 (N_7008,N_6706,N_6526);
or U7009 (N_7009,N_6521,N_6218);
xnor U7010 (N_7010,N_6088,N_6988);
nor U7011 (N_7011,N_6981,N_6135);
nand U7012 (N_7012,N_6823,N_6066);
or U7013 (N_7013,N_6780,N_6237);
nand U7014 (N_7014,N_6767,N_6461);
and U7015 (N_7015,N_6454,N_6480);
nor U7016 (N_7016,N_6821,N_6961);
nand U7017 (N_7017,N_6468,N_6854);
nor U7018 (N_7018,N_6220,N_6126);
nand U7019 (N_7019,N_6736,N_6843);
nand U7020 (N_7020,N_6330,N_6628);
nand U7021 (N_7021,N_6362,N_6720);
xnor U7022 (N_7022,N_6943,N_6465);
xnor U7023 (N_7023,N_6242,N_6015);
nor U7024 (N_7024,N_6653,N_6715);
xor U7025 (N_7025,N_6595,N_6097);
nor U7026 (N_7026,N_6450,N_6662);
nand U7027 (N_7027,N_6192,N_6846);
nand U7028 (N_7028,N_6495,N_6217);
xor U7029 (N_7029,N_6805,N_6773);
nor U7030 (N_7030,N_6031,N_6664);
xnor U7031 (N_7031,N_6162,N_6168);
or U7032 (N_7032,N_6674,N_6196);
nor U7033 (N_7033,N_6368,N_6555);
and U7034 (N_7034,N_6392,N_6474);
nand U7035 (N_7035,N_6875,N_6860);
nand U7036 (N_7036,N_6917,N_6876);
and U7037 (N_7037,N_6120,N_6371);
nor U7038 (N_7038,N_6083,N_6967);
or U7039 (N_7039,N_6409,N_6247);
nor U7040 (N_7040,N_6477,N_6898);
nand U7041 (N_7041,N_6905,N_6238);
and U7042 (N_7042,N_6446,N_6282);
nor U7043 (N_7043,N_6624,N_6222);
xor U7044 (N_7044,N_6858,N_6298);
or U7045 (N_7045,N_6908,N_6504);
or U7046 (N_7046,N_6143,N_6209);
nand U7047 (N_7047,N_6294,N_6401);
and U7048 (N_7048,N_6337,N_6829);
and U7049 (N_7049,N_6291,N_6267);
xnor U7050 (N_7050,N_6535,N_6991);
and U7051 (N_7051,N_6268,N_6863);
nand U7052 (N_7052,N_6701,N_6704);
nand U7053 (N_7053,N_6205,N_6751);
xor U7054 (N_7054,N_6197,N_6636);
xor U7055 (N_7055,N_6525,N_6946);
nand U7056 (N_7056,N_6417,N_6322);
nor U7057 (N_7057,N_6650,N_6885);
and U7058 (N_7058,N_6215,N_6941);
xor U7059 (N_7059,N_6746,N_6509);
xnor U7060 (N_7060,N_6319,N_6062);
and U7061 (N_7061,N_6486,N_6164);
nand U7062 (N_7062,N_6005,N_6629);
nor U7063 (N_7063,N_6129,N_6693);
xnor U7064 (N_7064,N_6317,N_6312);
or U7065 (N_7065,N_6663,N_6223);
xor U7066 (N_7066,N_6152,N_6467);
or U7067 (N_7067,N_6643,N_6797);
nor U7068 (N_7068,N_6093,N_6271);
and U7069 (N_7069,N_6012,N_6808);
or U7070 (N_7070,N_6657,N_6547);
and U7071 (N_7071,N_6916,N_6352);
and U7072 (N_7072,N_6149,N_6825);
nor U7073 (N_7073,N_6756,N_6104);
nand U7074 (N_7074,N_6793,N_6469);
nor U7075 (N_7075,N_6213,N_6175);
xor U7076 (N_7076,N_6951,N_6625);
or U7077 (N_7077,N_6040,N_6229);
and U7078 (N_7078,N_6029,N_6183);
and U7079 (N_7079,N_6707,N_6616);
nor U7080 (N_7080,N_6790,N_6838);
and U7081 (N_7081,N_6627,N_6889);
xor U7082 (N_7082,N_6512,N_6070);
nand U7083 (N_7083,N_6888,N_6831);
nor U7084 (N_7084,N_6906,N_6565);
xor U7085 (N_7085,N_6710,N_6970);
nand U7086 (N_7086,N_6911,N_6883);
nor U7087 (N_7087,N_6288,N_6189);
or U7088 (N_7088,N_6009,N_6749);
nand U7089 (N_7089,N_6199,N_6990);
or U7090 (N_7090,N_6195,N_6897);
xor U7091 (N_7091,N_6163,N_6191);
xor U7092 (N_7092,N_6491,N_6578);
nand U7093 (N_7093,N_6254,N_6110);
xnor U7094 (N_7094,N_6679,N_6383);
xor U7095 (N_7095,N_6021,N_6623);
nor U7096 (N_7096,N_6315,N_6000);
xnor U7097 (N_7097,N_6244,N_6051);
and U7098 (N_7098,N_6314,N_6779);
and U7099 (N_7099,N_6279,N_6249);
xnor U7100 (N_7100,N_6654,N_6646);
or U7101 (N_7101,N_6240,N_6777);
or U7102 (N_7102,N_6203,N_6476);
xnor U7103 (N_7103,N_6054,N_6923);
or U7104 (N_7104,N_6919,N_6552);
nor U7105 (N_7105,N_6792,N_6867);
or U7106 (N_7106,N_6166,N_6338);
or U7107 (N_7107,N_6640,N_6329);
or U7108 (N_7108,N_6904,N_6966);
and U7109 (N_7109,N_6484,N_6723);
and U7110 (N_7110,N_6599,N_6757);
or U7111 (N_7111,N_6499,N_6591);
xor U7112 (N_7112,N_6323,N_6676);
xnor U7113 (N_7113,N_6686,N_6007);
xor U7114 (N_7114,N_6171,N_6812);
or U7115 (N_7115,N_6327,N_6148);
nand U7116 (N_7116,N_6606,N_6376);
nand U7117 (N_7117,N_6065,N_6380);
nor U7118 (N_7118,N_6046,N_6553);
xnor U7119 (N_7119,N_6277,N_6245);
xor U7120 (N_7120,N_6730,N_6621);
nand U7121 (N_7121,N_6573,N_6581);
xor U7122 (N_7122,N_6566,N_6994);
or U7123 (N_7123,N_6395,N_6252);
or U7124 (N_7124,N_6313,N_6430);
or U7125 (N_7125,N_6370,N_6246);
nand U7126 (N_7126,N_6957,N_6109);
or U7127 (N_7127,N_6589,N_6464);
and U7128 (N_7128,N_6221,N_6765);
and U7129 (N_7129,N_6098,N_6369);
or U7130 (N_7130,N_6895,N_6788);
xnor U7131 (N_7131,N_6915,N_6677);
or U7132 (N_7132,N_6039,N_6969);
or U7133 (N_7133,N_6587,N_6343);
nand U7134 (N_7134,N_6443,N_6696);
and U7135 (N_7135,N_6037,N_6086);
xnor U7136 (N_7136,N_6320,N_6301);
nand U7137 (N_7137,N_6771,N_6048);
xnor U7138 (N_7138,N_6633,N_6520);
nor U7139 (N_7139,N_6125,N_6564);
and U7140 (N_7140,N_6456,N_6791);
nor U7141 (N_7141,N_6856,N_6794);
or U7142 (N_7142,N_6035,N_6059);
nand U7143 (N_7143,N_6708,N_6434);
xnor U7144 (N_7144,N_6665,N_6257);
nand U7145 (N_7145,N_6534,N_6324);
and U7146 (N_7146,N_6155,N_6726);
nor U7147 (N_7147,N_6878,N_6194);
xnor U7148 (N_7148,N_6731,N_6959);
and U7149 (N_7149,N_6333,N_6769);
or U7150 (N_7150,N_6427,N_6689);
nand U7151 (N_7151,N_6108,N_6714);
xor U7152 (N_7152,N_6334,N_6080);
nor U7153 (N_7153,N_6579,N_6722);
or U7154 (N_7154,N_6444,N_6106);
and U7155 (N_7155,N_6336,N_6099);
or U7156 (N_7156,N_6473,N_6851);
and U7157 (N_7157,N_6685,N_6810);
nand U7158 (N_7158,N_6735,N_6850);
or U7159 (N_7159,N_6198,N_6893);
nor U7160 (N_7160,N_6030,N_6502);
nor U7161 (N_7161,N_6006,N_6494);
and U7162 (N_7162,N_6741,N_6809);
xnor U7163 (N_7163,N_6248,N_6868);
nor U7164 (N_7164,N_6305,N_6140);
or U7165 (N_7165,N_6144,N_6702);
nor U7166 (N_7166,N_6847,N_6074);
nand U7167 (N_7167,N_6995,N_6820);
nand U7168 (N_7168,N_6881,N_6297);
or U7169 (N_7169,N_6842,N_6645);
xnor U7170 (N_7170,N_6986,N_6745);
nand U7171 (N_7171,N_6359,N_6023);
nand U7172 (N_7172,N_6281,N_6272);
nor U7173 (N_7173,N_6349,N_6394);
and U7174 (N_7174,N_6119,N_6105);
and U7175 (N_7175,N_6950,N_6382);
and U7176 (N_7176,N_6355,N_6864);
nor U7177 (N_7177,N_6052,N_6284);
nand U7178 (N_7178,N_6622,N_6413);
or U7179 (N_7179,N_6311,N_6452);
and U7180 (N_7180,N_6202,N_6415);
nand U7181 (N_7181,N_6920,N_6384);
and U7182 (N_7182,N_6912,N_6712);
xnor U7183 (N_7183,N_6445,N_6559);
or U7184 (N_7184,N_6471,N_6270);
and U7185 (N_7185,N_6658,N_6153);
nor U7186 (N_7186,N_6652,N_6803);
or U7187 (N_7187,N_6280,N_6239);
nor U7188 (N_7188,N_6835,N_6075);
or U7189 (N_7189,N_6848,N_6200);
or U7190 (N_7190,N_6416,N_6127);
and U7191 (N_7191,N_6342,N_6819);
nor U7192 (N_7192,N_6219,N_6607);
xor U7193 (N_7193,N_6344,N_6694);
nand U7194 (N_7194,N_6356,N_6768);
or U7195 (N_7195,N_6188,N_6892);
nand U7196 (N_7196,N_6930,N_6212);
xor U7197 (N_7197,N_6866,N_6763);
nor U7198 (N_7198,N_6309,N_6758);
nand U7199 (N_7199,N_6896,N_6531);
nor U7200 (N_7200,N_6551,N_6600);
nand U7201 (N_7201,N_6921,N_6659);
nor U7202 (N_7202,N_6177,N_6750);
nor U7203 (N_7203,N_6620,N_6304);
or U7204 (N_7204,N_6057,N_6615);
nand U7205 (N_7205,N_6441,N_6422);
or U7206 (N_7206,N_6691,N_6592);
nand U7207 (N_7207,N_6532,N_6403);
and U7208 (N_7208,N_6783,N_6700);
and U7209 (N_7209,N_6562,N_6576);
and U7210 (N_7210,N_6914,N_6488);
and U7211 (N_7211,N_6451,N_6873);
and U7212 (N_7212,N_6493,N_6373);
xnor U7213 (N_7213,N_6901,N_6572);
xor U7214 (N_7214,N_6487,N_6697);
xnor U7215 (N_7215,N_6554,N_6386);
or U7216 (N_7216,N_6610,N_6996);
nand U7217 (N_7217,N_6753,N_6455);
nand U7218 (N_7218,N_6258,N_6475);
and U7219 (N_7219,N_6001,N_6490);
nor U7220 (N_7220,N_6269,N_6236);
and U7221 (N_7221,N_6585,N_6972);
xnor U7222 (N_7222,N_6365,N_6945);
nor U7223 (N_7223,N_6782,N_6016);
or U7224 (N_7224,N_6293,N_6290);
or U7225 (N_7225,N_6283,N_6513);
or U7226 (N_7226,N_6241,N_6310);
or U7227 (N_7227,N_6909,N_6348);
nor U7228 (N_7228,N_6235,N_6784);
xor U7229 (N_7229,N_6299,N_6737);
or U7230 (N_7230,N_6557,N_6549);
or U7231 (N_7231,N_6594,N_6414);
or U7232 (N_7232,N_6569,N_6045);
nand U7233 (N_7233,N_6133,N_6038);
and U7234 (N_7234,N_6433,N_6385);
xnor U7235 (N_7235,N_6778,N_6147);
xor U7236 (N_7236,N_6924,N_6865);
nand U7237 (N_7237,N_6117,N_6956);
nor U7238 (N_7238,N_6346,N_6489);
nand U7239 (N_7239,N_6397,N_6316);
xor U7240 (N_7240,N_6067,N_6058);
and U7241 (N_7241,N_6377,N_6204);
or U7242 (N_7242,N_6260,N_6832);
xnor U7243 (N_7243,N_6890,N_6859);
or U7244 (N_7244,N_6262,N_6647);
and U7245 (N_7245,N_6887,N_6325);
xor U7246 (N_7246,N_6273,N_6849);
nor U7247 (N_7247,N_6224,N_6872);
nand U7248 (N_7248,N_6655,N_6903);
and U7249 (N_7249,N_6947,N_6225);
xor U7250 (N_7250,N_6457,N_6402);
nor U7251 (N_7251,N_6146,N_6632);
and U7252 (N_7252,N_6638,N_6011);
or U7253 (N_7253,N_6044,N_6335);
nand U7254 (N_7254,N_6598,N_6519);
nor U7255 (N_7255,N_6752,N_6186);
or U7256 (N_7256,N_6178,N_6295);
nand U7257 (N_7257,N_6609,N_6216);
and U7258 (N_7258,N_6560,N_6014);
or U7259 (N_7259,N_6453,N_6933);
or U7260 (N_7260,N_6910,N_6603);
nor U7261 (N_7261,N_6718,N_6458);
nor U7262 (N_7262,N_6176,N_6543);
and U7263 (N_7263,N_6228,N_6255);
and U7264 (N_7264,N_6800,N_6326);
and U7265 (N_7265,N_6078,N_6159);
or U7266 (N_7266,N_6150,N_6100);
xor U7267 (N_7267,N_6869,N_6024);
xor U7268 (N_7268,N_6507,N_6937);
and U7269 (N_7269,N_6743,N_6134);
nand U7270 (N_7270,N_6354,N_6678);
or U7271 (N_7271,N_6265,N_6321);
nand U7272 (N_7272,N_6094,N_6861);
nor U7273 (N_7273,N_6754,N_6425);
or U7274 (N_7274,N_6976,N_6460);
nand U7275 (N_7275,N_6503,N_6158);
xor U7276 (N_7276,N_6364,N_6174);
or U7277 (N_7277,N_6721,N_6410);
nand U7278 (N_7278,N_6498,N_6836);
nand U7279 (N_7279,N_6593,N_6300);
nand U7280 (N_7280,N_6463,N_6331);
xnor U7281 (N_7281,N_6739,N_6405);
nand U7282 (N_7282,N_6801,N_6366);
and U7283 (N_7283,N_6955,N_6799);
xor U7284 (N_7284,N_6227,N_6546);
nand U7285 (N_7285,N_6112,N_6411);
xor U7286 (N_7286,N_6630,N_6361);
or U7287 (N_7287,N_6396,N_6626);
and U7288 (N_7288,N_6785,N_6483);
and U7289 (N_7289,N_6608,N_6296);
nand U7290 (N_7290,N_6234,N_6518);
nand U7291 (N_7291,N_6979,N_6387);
and U7292 (N_7292,N_6567,N_6965);
and U7293 (N_7293,N_6447,N_6899);
nor U7294 (N_7294,N_6748,N_6528);
xnor U7295 (N_7295,N_6934,N_6759);
nor U7296 (N_7296,N_6285,N_6962);
nor U7297 (N_7297,N_6672,N_6478);
xor U7298 (N_7298,N_6656,N_6670);
nand U7299 (N_7299,N_6172,N_6649);
or U7300 (N_7300,N_6815,N_6727);
or U7301 (N_7301,N_6728,N_6182);
nor U7302 (N_7302,N_6137,N_6926);
nor U7303 (N_7303,N_6091,N_6840);
or U7304 (N_7304,N_6399,N_6442);
and U7305 (N_7305,N_6529,N_6264);
or U7306 (N_7306,N_6577,N_6938);
and U7307 (N_7307,N_6053,N_6210);
nand U7308 (N_7308,N_6724,N_6303);
xnor U7309 (N_7309,N_6187,N_6733);
nor U7310 (N_7310,N_6286,N_6485);
xnor U7311 (N_7311,N_6762,N_6406);
nor U7312 (N_7312,N_6027,N_6601);
nand U7313 (N_7313,N_6470,N_6772);
nand U7314 (N_7314,N_6918,N_6795);
xnor U7315 (N_7315,N_6827,N_6604);
and U7316 (N_7316,N_6041,N_6275);
nand U7317 (N_7317,N_6501,N_6660);
and U7318 (N_7318,N_6266,N_6524);
xor U7319 (N_7319,N_6536,N_6963);
nand U7320 (N_7320,N_6042,N_6548);
nor U7321 (N_7321,N_6612,N_6185);
nand U7322 (N_7322,N_6510,N_6673);
and U7323 (N_7323,N_6374,N_6684);
xor U7324 (N_7324,N_6449,N_6690);
xor U7325 (N_7325,N_6101,N_6230);
nand U7326 (N_7326,N_6989,N_6207);
xnor U7327 (N_7327,N_6145,N_6472);
nand U7328 (N_7328,N_6061,N_6424);
nor U7329 (N_7329,N_6390,N_6132);
nand U7330 (N_7330,N_6261,N_6975);
and U7331 (N_7331,N_6124,N_6913);
xor U7332 (N_7332,N_6538,N_6128);
nor U7333 (N_7333,N_6880,N_6419);
and U7334 (N_7334,N_6092,N_6738);
nand U7335 (N_7335,N_6987,N_6539);
or U7336 (N_7336,N_6992,N_6597);
and U7337 (N_7337,N_6681,N_6306);
and U7338 (N_7338,N_6250,N_6276);
nor U7339 (N_7339,N_6156,N_6618);
xnor U7340 (N_7340,N_6231,N_6043);
or U7341 (N_7341,N_6421,N_6429);
xnor U7342 (N_7342,N_6393,N_6774);
nand U7343 (N_7343,N_6818,N_6482);
nor U7344 (N_7344,N_6833,N_6165);
xnor U7345 (N_7345,N_6602,N_6004);
nor U7346 (N_7346,N_6882,N_6999);
or U7347 (N_7347,N_6292,N_6802);
nand U7348 (N_7348,N_6900,N_6206);
or U7349 (N_7349,N_6389,N_6492);
or U7350 (N_7350,N_6642,N_6523);
nand U7351 (N_7351,N_6611,N_6459);
nor U7352 (N_7352,N_6641,N_6617);
or U7353 (N_7353,N_6853,N_6407);
xnor U7354 (N_7354,N_6575,N_6563);
xnor U7355 (N_7355,N_6651,N_6826);
nor U7356 (N_7356,N_6755,N_6047);
nor U7357 (N_7357,N_6516,N_6614);
nand U7358 (N_7358,N_6026,N_6953);
and U7359 (N_7359,N_6340,N_6942);
or U7360 (N_7360,N_6077,N_6775);
nor U7361 (N_7361,N_6862,N_6180);
or U7362 (N_7362,N_6884,N_6232);
xor U7363 (N_7363,N_6351,N_6816);
nor U7364 (N_7364,N_6855,N_6839);
and U7365 (N_7365,N_6079,N_6050);
nor U7366 (N_7366,N_6069,N_6968);
xor U7367 (N_7367,N_6584,N_6997);
and U7368 (N_7368,N_6760,N_6017);
and U7369 (N_7369,N_6613,N_6060);
nor U7370 (N_7370,N_6687,N_6350);
or U7371 (N_7371,N_6139,N_6307);
or U7372 (N_7372,N_6466,N_6378);
nand U7373 (N_7373,N_6732,N_6318);
xnor U7374 (N_7374,N_6582,N_6122);
xor U7375 (N_7375,N_6977,N_6056);
nand U7376 (N_7376,N_6845,N_6003);
nand U7377 (N_7377,N_6208,N_6719);
and U7378 (N_7378,N_6438,N_6841);
nand U7379 (N_7379,N_6018,N_6734);
nand U7380 (N_7380,N_6857,N_6090);
xor U7381 (N_7381,N_6891,N_6391);
nor U7382 (N_7382,N_6766,N_6796);
or U7383 (N_7383,N_6436,N_6556);
and U7384 (N_7384,N_6644,N_6844);
and U7385 (N_7385,N_6824,N_6347);
or U7386 (N_7386,N_6682,N_6984);
nor U7387 (N_7387,N_6160,N_6786);
xor U7388 (N_7388,N_6637,N_6776);
xnor U7389 (N_7389,N_6983,N_6496);
and U7390 (N_7390,N_6639,N_6118);
or U7391 (N_7391,N_6302,N_6028);
xnor U7392 (N_7392,N_6063,N_6931);
nand U7393 (N_7393,N_6170,N_6558);
and U7394 (N_7394,N_6138,N_6729);
and U7395 (N_7395,N_6541,N_6328);
nor U7396 (N_7396,N_6811,N_6877);
nor U7397 (N_7397,N_6103,N_6341);
xor U7398 (N_7398,N_6064,N_6151);
nand U7399 (N_7399,N_6540,N_6571);
and U7400 (N_7400,N_6087,N_6437);
nor U7401 (N_7401,N_6462,N_6619);
nor U7402 (N_7402,N_6907,N_6952);
and U7403 (N_7403,N_6375,N_6142);
xor U7404 (N_7404,N_6974,N_6481);
nor U7405 (N_7405,N_6954,N_6113);
xor U7406 (N_7406,N_6927,N_6711);
xor U7407 (N_7407,N_6022,N_6211);
xnor U7408 (N_7408,N_6130,N_6002);
xor U7409 (N_7409,N_6932,N_6631);
xnor U7410 (N_7410,N_6894,N_6049);
nor U7411 (N_7411,N_6412,N_6479);
nand U7412 (N_7412,N_6680,N_6925);
and U7413 (N_7413,N_6367,N_6420);
xor U7414 (N_7414,N_6116,N_6744);
nor U7415 (N_7415,N_6717,N_6537);
and U7416 (N_7416,N_6993,N_6870);
nand U7417 (N_7417,N_6214,N_6161);
or U7418 (N_7418,N_6435,N_6233);
nand U7419 (N_7419,N_6527,N_6157);
and U7420 (N_7420,N_6596,N_6358);
nor U7421 (N_7421,N_6360,N_6440);
nand U7422 (N_7422,N_6287,N_6948);
nor U7423 (N_7423,N_6102,N_6431);
nand U7424 (N_7424,N_6274,N_6096);
xnor U7425 (N_7425,N_6226,N_6787);
xor U7426 (N_7426,N_6400,N_6964);
or U7427 (N_7427,N_6692,N_6770);
and U7428 (N_7428,N_6980,N_6439);
and U7429 (N_7429,N_6243,N_6852);
nand U7430 (N_7430,N_6111,N_6154);
and U7431 (N_7431,N_6036,N_6542);
xnor U7432 (N_7432,N_6879,N_6922);
xnor U7433 (N_7433,N_6278,N_6533);
and U7434 (N_7434,N_6259,N_6071);
or U7435 (N_7435,N_6971,N_6709);
nand U7436 (N_7436,N_6055,N_6789);
or U7437 (N_7437,N_6683,N_6034);
and U7438 (N_7438,N_6837,N_6363);
nand U7439 (N_7439,N_6583,N_6874);
or U7440 (N_7440,N_6173,N_6828);
nand U7441 (N_7441,N_6253,N_6570);
and U7442 (N_7442,N_6379,N_6184);
nor U7443 (N_7443,N_6671,N_6666);
and U7444 (N_7444,N_6497,N_6545);
nor U7445 (N_7445,N_6190,N_6114);
nor U7446 (N_7446,N_6372,N_6500);
nand U7447 (N_7447,N_6764,N_6949);
or U7448 (N_7448,N_6747,N_6982);
and U7449 (N_7449,N_6418,N_6648);
and U7450 (N_7450,N_6426,N_6668);
nor U7451 (N_7451,N_6740,N_6568);
nand U7452 (N_7452,N_6635,N_6806);
nand U7453 (N_7453,N_6669,N_6798);
and U7454 (N_7454,N_6193,N_6960);
and U7455 (N_7455,N_6761,N_6398);
xor U7456 (N_7456,N_6404,N_6506);
xnor U7457 (N_7457,N_6095,N_6936);
xnor U7458 (N_7458,N_6008,N_6357);
nand U7459 (N_7459,N_6725,N_6082);
and U7460 (N_7460,N_6167,N_6032);
nand U7461 (N_7461,N_6530,N_6985);
nor U7462 (N_7462,N_6073,N_6935);
xor U7463 (N_7463,N_6939,N_6634);
xor U7464 (N_7464,N_6508,N_6561);
and U7465 (N_7465,N_6263,N_6817);
xnor U7466 (N_7466,N_6814,N_6332);
nor U7467 (N_7467,N_6076,N_6871);
and U7468 (N_7468,N_6716,N_6010);
nand U7469 (N_7469,N_6448,N_6181);
xnor U7470 (N_7470,N_6998,N_6929);
or U7471 (N_7471,N_6742,N_6517);
nor U7472 (N_7472,N_6586,N_6201);
xnor U7473 (N_7473,N_6958,N_6699);
xor U7474 (N_7474,N_6511,N_6020);
or U7475 (N_7475,N_6514,N_6807);
nor U7476 (N_7476,N_6588,N_6973);
nor U7477 (N_7477,N_6136,N_6107);
nand U7478 (N_7478,N_6830,N_6580);
xnor U7479 (N_7479,N_6574,N_6822);
xor U7480 (N_7480,N_6085,N_6834);
and U7481 (N_7481,N_6813,N_6544);
nand U7482 (N_7482,N_6695,N_6025);
nor U7483 (N_7483,N_6169,N_6019);
and U7484 (N_7484,N_6408,N_6068);
or U7485 (N_7485,N_6289,N_6141);
or U7486 (N_7486,N_6084,N_6121);
xor U7487 (N_7487,N_6081,N_6423);
and U7488 (N_7488,N_6432,N_6590);
or U7489 (N_7489,N_6428,N_6928);
nor U7490 (N_7490,N_6353,N_6256);
nand U7491 (N_7491,N_6902,N_6089);
nand U7492 (N_7492,N_6703,N_6688);
xor U7493 (N_7493,N_6944,N_6698);
or U7494 (N_7494,N_6804,N_6388);
xnor U7495 (N_7495,N_6886,N_6705);
and U7496 (N_7496,N_6345,N_6550);
and U7497 (N_7497,N_6131,N_6381);
nand U7498 (N_7498,N_6115,N_6515);
nor U7499 (N_7499,N_6781,N_6667);
xor U7500 (N_7500,N_6645,N_6479);
and U7501 (N_7501,N_6905,N_6638);
or U7502 (N_7502,N_6782,N_6989);
and U7503 (N_7503,N_6841,N_6054);
xor U7504 (N_7504,N_6543,N_6325);
or U7505 (N_7505,N_6141,N_6976);
nor U7506 (N_7506,N_6064,N_6360);
and U7507 (N_7507,N_6380,N_6105);
and U7508 (N_7508,N_6584,N_6519);
and U7509 (N_7509,N_6033,N_6148);
xor U7510 (N_7510,N_6639,N_6007);
nand U7511 (N_7511,N_6548,N_6481);
nor U7512 (N_7512,N_6113,N_6651);
nand U7513 (N_7513,N_6996,N_6130);
xor U7514 (N_7514,N_6733,N_6399);
nor U7515 (N_7515,N_6517,N_6021);
nor U7516 (N_7516,N_6331,N_6156);
nor U7517 (N_7517,N_6350,N_6290);
nor U7518 (N_7518,N_6778,N_6131);
or U7519 (N_7519,N_6927,N_6769);
nor U7520 (N_7520,N_6234,N_6619);
nand U7521 (N_7521,N_6422,N_6384);
nor U7522 (N_7522,N_6999,N_6344);
nand U7523 (N_7523,N_6334,N_6803);
and U7524 (N_7524,N_6672,N_6165);
and U7525 (N_7525,N_6619,N_6709);
or U7526 (N_7526,N_6240,N_6500);
nand U7527 (N_7527,N_6436,N_6805);
and U7528 (N_7528,N_6514,N_6369);
xor U7529 (N_7529,N_6861,N_6479);
xnor U7530 (N_7530,N_6066,N_6134);
or U7531 (N_7531,N_6201,N_6512);
xnor U7532 (N_7532,N_6658,N_6293);
xnor U7533 (N_7533,N_6955,N_6782);
xor U7534 (N_7534,N_6486,N_6792);
nand U7535 (N_7535,N_6870,N_6723);
and U7536 (N_7536,N_6165,N_6658);
or U7537 (N_7537,N_6371,N_6106);
or U7538 (N_7538,N_6796,N_6027);
nor U7539 (N_7539,N_6696,N_6986);
and U7540 (N_7540,N_6263,N_6519);
or U7541 (N_7541,N_6164,N_6475);
nor U7542 (N_7542,N_6231,N_6298);
nor U7543 (N_7543,N_6156,N_6597);
or U7544 (N_7544,N_6649,N_6648);
xor U7545 (N_7545,N_6757,N_6346);
xor U7546 (N_7546,N_6506,N_6884);
or U7547 (N_7547,N_6896,N_6369);
nand U7548 (N_7548,N_6389,N_6225);
xor U7549 (N_7549,N_6322,N_6767);
nor U7550 (N_7550,N_6657,N_6412);
xnor U7551 (N_7551,N_6682,N_6195);
nor U7552 (N_7552,N_6303,N_6670);
nor U7553 (N_7553,N_6761,N_6212);
nor U7554 (N_7554,N_6769,N_6823);
or U7555 (N_7555,N_6423,N_6186);
or U7556 (N_7556,N_6622,N_6615);
xnor U7557 (N_7557,N_6399,N_6328);
nand U7558 (N_7558,N_6288,N_6163);
nor U7559 (N_7559,N_6850,N_6352);
nand U7560 (N_7560,N_6341,N_6426);
nand U7561 (N_7561,N_6193,N_6443);
xor U7562 (N_7562,N_6660,N_6730);
nand U7563 (N_7563,N_6887,N_6741);
or U7564 (N_7564,N_6393,N_6292);
nand U7565 (N_7565,N_6658,N_6750);
xor U7566 (N_7566,N_6095,N_6686);
nor U7567 (N_7567,N_6065,N_6095);
or U7568 (N_7568,N_6252,N_6264);
and U7569 (N_7569,N_6168,N_6631);
xnor U7570 (N_7570,N_6588,N_6281);
and U7571 (N_7571,N_6728,N_6266);
nand U7572 (N_7572,N_6193,N_6219);
nor U7573 (N_7573,N_6563,N_6766);
or U7574 (N_7574,N_6971,N_6026);
xor U7575 (N_7575,N_6175,N_6052);
xor U7576 (N_7576,N_6195,N_6935);
and U7577 (N_7577,N_6031,N_6248);
nor U7578 (N_7578,N_6259,N_6679);
or U7579 (N_7579,N_6393,N_6125);
nand U7580 (N_7580,N_6254,N_6361);
nand U7581 (N_7581,N_6445,N_6034);
and U7582 (N_7582,N_6890,N_6388);
xnor U7583 (N_7583,N_6534,N_6853);
xnor U7584 (N_7584,N_6785,N_6916);
and U7585 (N_7585,N_6055,N_6127);
or U7586 (N_7586,N_6595,N_6173);
and U7587 (N_7587,N_6773,N_6030);
and U7588 (N_7588,N_6088,N_6495);
and U7589 (N_7589,N_6794,N_6147);
or U7590 (N_7590,N_6097,N_6213);
nor U7591 (N_7591,N_6629,N_6579);
and U7592 (N_7592,N_6533,N_6843);
nor U7593 (N_7593,N_6104,N_6142);
nor U7594 (N_7594,N_6150,N_6408);
and U7595 (N_7595,N_6125,N_6124);
and U7596 (N_7596,N_6589,N_6873);
nand U7597 (N_7597,N_6149,N_6811);
or U7598 (N_7598,N_6017,N_6250);
or U7599 (N_7599,N_6838,N_6302);
or U7600 (N_7600,N_6133,N_6014);
and U7601 (N_7601,N_6455,N_6742);
and U7602 (N_7602,N_6053,N_6425);
or U7603 (N_7603,N_6216,N_6488);
or U7604 (N_7604,N_6870,N_6195);
and U7605 (N_7605,N_6809,N_6604);
xor U7606 (N_7606,N_6536,N_6556);
or U7607 (N_7607,N_6493,N_6782);
nand U7608 (N_7608,N_6751,N_6452);
nand U7609 (N_7609,N_6577,N_6987);
nand U7610 (N_7610,N_6619,N_6326);
and U7611 (N_7611,N_6273,N_6718);
xnor U7612 (N_7612,N_6137,N_6299);
xnor U7613 (N_7613,N_6198,N_6749);
nor U7614 (N_7614,N_6285,N_6721);
nor U7615 (N_7615,N_6466,N_6169);
xnor U7616 (N_7616,N_6576,N_6644);
or U7617 (N_7617,N_6231,N_6931);
nor U7618 (N_7618,N_6994,N_6469);
nor U7619 (N_7619,N_6558,N_6748);
or U7620 (N_7620,N_6008,N_6458);
nor U7621 (N_7621,N_6310,N_6921);
nand U7622 (N_7622,N_6991,N_6037);
nand U7623 (N_7623,N_6905,N_6533);
nor U7624 (N_7624,N_6840,N_6488);
xnor U7625 (N_7625,N_6212,N_6973);
and U7626 (N_7626,N_6594,N_6486);
and U7627 (N_7627,N_6336,N_6984);
nor U7628 (N_7628,N_6888,N_6893);
nand U7629 (N_7629,N_6041,N_6942);
nor U7630 (N_7630,N_6327,N_6492);
xnor U7631 (N_7631,N_6511,N_6840);
or U7632 (N_7632,N_6725,N_6222);
xnor U7633 (N_7633,N_6456,N_6342);
and U7634 (N_7634,N_6988,N_6506);
and U7635 (N_7635,N_6543,N_6034);
and U7636 (N_7636,N_6899,N_6914);
nor U7637 (N_7637,N_6022,N_6108);
xor U7638 (N_7638,N_6133,N_6522);
or U7639 (N_7639,N_6444,N_6756);
and U7640 (N_7640,N_6681,N_6013);
nor U7641 (N_7641,N_6348,N_6867);
nor U7642 (N_7642,N_6375,N_6416);
or U7643 (N_7643,N_6454,N_6271);
xor U7644 (N_7644,N_6325,N_6839);
xor U7645 (N_7645,N_6192,N_6483);
nand U7646 (N_7646,N_6208,N_6264);
and U7647 (N_7647,N_6167,N_6885);
nand U7648 (N_7648,N_6194,N_6808);
and U7649 (N_7649,N_6201,N_6898);
or U7650 (N_7650,N_6340,N_6174);
or U7651 (N_7651,N_6679,N_6730);
or U7652 (N_7652,N_6881,N_6322);
xor U7653 (N_7653,N_6917,N_6251);
xor U7654 (N_7654,N_6125,N_6835);
and U7655 (N_7655,N_6301,N_6089);
xnor U7656 (N_7656,N_6598,N_6368);
nor U7657 (N_7657,N_6134,N_6420);
nand U7658 (N_7658,N_6664,N_6137);
and U7659 (N_7659,N_6232,N_6105);
and U7660 (N_7660,N_6579,N_6841);
nor U7661 (N_7661,N_6631,N_6468);
nand U7662 (N_7662,N_6504,N_6427);
and U7663 (N_7663,N_6981,N_6390);
or U7664 (N_7664,N_6567,N_6829);
nand U7665 (N_7665,N_6116,N_6650);
xor U7666 (N_7666,N_6334,N_6002);
xor U7667 (N_7667,N_6997,N_6193);
or U7668 (N_7668,N_6602,N_6856);
nor U7669 (N_7669,N_6591,N_6076);
or U7670 (N_7670,N_6017,N_6477);
or U7671 (N_7671,N_6604,N_6243);
and U7672 (N_7672,N_6334,N_6113);
and U7673 (N_7673,N_6351,N_6121);
and U7674 (N_7674,N_6450,N_6729);
or U7675 (N_7675,N_6262,N_6069);
nor U7676 (N_7676,N_6704,N_6559);
nor U7677 (N_7677,N_6202,N_6393);
or U7678 (N_7678,N_6916,N_6590);
and U7679 (N_7679,N_6917,N_6487);
or U7680 (N_7680,N_6403,N_6392);
or U7681 (N_7681,N_6411,N_6740);
nor U7682 (N_7682,N_6317,N_6408);
xor U7683 (N_7683,N_6618,N_6382);
or U7684 (N_7684,N_6563,N_6348);
or U7685 (N_7685,N_6278,N_6849);
nand U7686 (N_7686,N_6173,N_6523);
nor U7687 (N_7687,N_6373,N_6914);
nor U7688 (N_7688,N_6652,N_6421);
or U7689 (N_7689,N_6033,N_6627);
nor U7690 (N_7690,N_6639,N_6665);
or U7691 (N_7691,N_6303,N_6283);
xnor U7692 (N_7692,N_6549,N_6435);
nand U7693 (N_7693,N_6190,N_6875);
or U7694 (N_7694,N_6598,N_6719);
and U7695 (N_7695,N_6568,N_6782);
or U7696 (N_7696,N_6219,N_6064);
nor U7697 (N_7697,N_6117,N_6055);
nand U7698 (N_7698,N_6943,N_6942);
nand U7699 (N_7699,N_6856,N_6307);
or U7700 (N_7700,N_6646,N_6479);
nand U7701 (N_7701,N_6968,N_6418);
nand U7702 (N_7702,N_6757,N_6746);
xnor U7703 (N_7703,N_6823,N_6993);
or U7704 (N_7704,N_6421,N_6570);
xnor U7705 (N_7705,N_6799,N_6722);
or U7706 (N_7706,N_6088,N_6193);
or U7707 (N_7707,N_6913,N_6191);
xnor U7708 (N_7708,N_6783,N_6438);
nor U7709 (N_7709,N_6726,N_6573);
and U7710 (N_7710,N_6024,N_6388);
xor U7711 (N_7711,N_6565,N_6061);
or U7712 (N_7712,N_6411,N_6177);
and U7713 (N_7713,N_6154,N_6858);
nor U7714 (N_7714,N_6330,N_6301);
or U7715 (N_7715,N_6630,N_6958);
xor U7716 (N_7716,N_6677,N_6923);
and U7717 (N_7717,N_6897,N_6355);
or U7718 (N_7718,N_6044,N_6446);
nor U7719 (N_7719,N_6141,N_6204);
and U7720 (N_7720,N_6727,N_6479);
xnor U7721 (N_7721,N_6492,N_6796);
nor U7722 (N_7722,N_6035,N_6600);
or U7723 (N_7723,N_6304,N_6795);
nor U7724 (N_7724,N_6982,N_6851);
or U7725 (N_7725,N_6137,N_6452);
or U7726 (N_7726,N_6354,N_6236);
xnor U7727 (N_7727,N_6352,N_6513);
xor U7728 (N_7728,N_6464,N_6501);
nor U7729 (N_7729,N_6936,N_6809);
nand U7730 (N_7730,N_6868,N_6975);
nand U7731 (N_7731,N_6554,N_6959);
nand U7732 (N_7732,N_6565,N_6183);
or U7733 (N_7733,N_6901,N_6090);
or U7734 (N_7734,N_6743,N_6157);
nand U7735 (N_7735,N_6008,N_6932);
xor U7736 (N_7736,N_6772,N_6106);
nor U7737 (N_7737,N_6123,N_6619);
xor U7738 (N_7738,N_6998,N_6593);
nor U7739 (N_7739,N_6878,N_6090);
and U7740 (N_7740,N_6485,N_6857);
nand U7741 (N_7741,N_6826,N_6231);
xnor U7742 (N_7742,N_6805,N_6958);
nor U7743 (N_7743,N_6075,N_6903);
or U7744 (N_7744,N_6724,N_6090);
and U7745 (N_7745,N_6902,N_6755);
nand U7746 (N_7746,N_6448,N_6439);
or U7747 (N_7747,N_6105,N_6887);
xnor U7748 (N_7748,N_6568,N_6741);
nor U7749 (N_7749,N_6023,N_6971);
nor U7750 (N_7750,N_6108,N_6777);
nand U7751 (N_7751,N_6253,N_6310);
xnor U7752 (N_7752,N_6393,N_6641);
and U7753 (N_7753,N_6999,N_6578);
and U7754 (N_7754,N_6535,N_6788);
nand U7755 (N_7755,N_6694,N_6167);
or U7756 (N_7756,N_6251,N_6029);
and U7757 (N_7757,N_6485,N_6575);
nor U7758 (N_7758,N_6656,N_6170);
and U7759 (N_7759,N_6292,N_6243);
nand U7760 (N_7760,N_6648,N_6703);
xor U7761 (N_7761,N_6946,N_6663);
nor U7762 (N_7762,N_6116,N_6270);
xor U7763 (N_7763,N_6585,N_6646);
xor U7764 (N_7764,N_6364,N_6847);
nand U7765 (N_7765,N_6263,N_6947);
nor U7766 (N_7766,N_6195,N_6448);
xnor U7767 (N_7767,N_6780,N_6627);
or U7768 (N_7768,N_6990,N_6073);
nand U7769 (N_7769,N_6151,N_6861);
xnor U7770 (N_7770,N_6317,N_6692);
or U7771 (N_7771,N_6334,N_6825);
and U7772 (N_7772,N_6588,N_6102);
and U7773 (N_7773,N_6017,N_6719);
and U7774 (N_7774,N_6679,N_6438);
xnor U7775 (N_7775,N_6756,N_6625);
and U7776 (N_7776,N_6784,N_6017);
xor U7777 (N_7777,N_6371,N_6961);
or U7778 (N_7778,N_6035,N_6296);
xnor U7779 (N_7779,N_6028,N_6927);
or U7780 (N_7780,N_6672,N_6034);
nor U7781 (N_7781,N_6213,N_6095);
or U7782 (N_7782,N_6482,N_6900);
or U7783 (N_7783,N_6455,N_6156);
and U7784 (N_7784,N_6409,N_6582);
nand U7785 (N_7785,N_6498,N_6445);
nor U7786 (N_7786,N_6314,N_6193);
nor U7787 (N_7787,N_6911,N_6762);
nor U7788 (N_7788,N_6735,N_6460);
and U7789 (N_7789,N_6944,N_6663);
xnor U7790 (N_7790,N_6442,N_6429);
and U7791 (N_7791,N_6973,N_6341);
or U7792 (N_7792,N_6204,N_6478);
nor U7793 (N_7793,N_6569,N_6458);
xnor U7794 (N_7794,N_6226,N_6170);
nor U7795 (N_7795,N_6770,N_6330);
nand U7796 (N_7796,N_6914,N_6401);
xnor U7797 (N_7797,N_6426,N_6995);
nand U7798 (N_7798,N_6615,N_6303);
or U7799 (N_7799,N_6780,N_6106);
nor U7800 (N_7800,N_6085,N_6622);
xor U7801 (N_7801,N_6027,N_6974);
nor U7802 (N_7802,N_6703,N_6789);
or U7803 (N_7803,N_6437,N_6105);
nand U7804 (N_7804,N_6427,N_6762);
nand U7805 (N_7805,N_6129,N_6511);
nor U7806 (N_7806,N_6468,N_6425);
xnor U7807 (N_7807,N_6410,N_6285);
nand U7808 (N_7808,N_6847,N_6033);
nor U7809 (N_7809,N_6910,N_6426);
nand U7810 (N_7810,N_6993,N_6603);
xnor U7811 (N_7811,N_6270,N_6510);
or U7812 (N_7812,N_6751,N_6841);
and U7813 (N_7813,N_6291,N_6429);
or U7814 (N_7814,N_6451,N_6164);
xnor U7815 (N_7815,N_6765,N_6525);
nand U7816 (N_7816,N_6889,N_6224);
nor U7817 (N_7817,N_6646,N_6212);
xnor U7818 (N_7818,N_6025,N_6133);
nor U7819 (N_7819,N_6907,N_6301);
xnor U7820 (N_7820,N_6630,N_6117);
xnor U7821 (N_7821,N_6601,N_6805);
xor U7822 (N_7822,N_6687,N_6050);
nand U7823 (N_7823,N_6541,N_6549);
nand U7824 (N_7824,N_6466,N_6240);
xnor U7825 (N_7825,N_6471,N_6904);
and U7826 (N_7826,N_6325,N_6642);
and U7827 (N_7827,N_6443,N_6083);
xnor U7828 (N_7828,N_6409,N_6771);
nand U7829 (N_7829,N_6152,N_6153);
nand U7830 (N_7830,N_6068,N_6083);
nand U7831 (N_7831,N_6524,N_6839);
xnor U7832 (N_7832,N_6118,N_6681);
xor U7833 (N_7833,N_6345,N_6284);
xor U7834 (N_7834,N_6968,N_6773);
and U7835 (N_7835,N_6898,N_6575);
or U7836 (N_7836,N_6436,N_6229);
or U7837 (N_7837,N_6454,N_6540);
xor U7838 (N_7838,N_6721,N_6320);
and U7839 (N_7839,N_6727,N_6077);
or U7840 (N_7840,N_6371,N_6364);
or U7841 (N_7841,N_6610,N_6211);
nor U7842 (N_7842,N_6595,N_6603);
nor U7843 (N_7843,N_6967,N_6228);
nor U7844 (N_7844,N_6347,N_6753);
nor U7845 (N_7845,N_6499,N_6059);
and U7846 (N_7846,N_6458,N_6352);
or U7847 (N_7847,N_6190,N_6957);
xor U7848 (N_7848,N_6868,N_6448);
and U7849 (N_7849,N_6135,N_6284);
nand U7850 (N_7850,N_6950,N_6175);
or U7851 (N_7851,N_6799,N_6331);
xnor U7852 (N_7852,N_6797,N_6732);
and U7853 (N_7853,N_6814,N_6992);
xor U7854 (N_7854,N_6368,N_6964);
nor U7855 (N_7855,N_6538,N_6651);
and U7856 (N_7856,N_6321,N_6713);
nor U7857 (N_7857,N_6914,N_6459);
xor U7858 (N_7858,N_6326,N_6820);
or U7859 (N_7859,N_6147,N_6653);
and U7860 (N_7860,N_6263,N_6772);
nand U7861 (N_7861,N_6048,N_6775);
and U7862 (N_7862,N_6780,N_6100);
nand U7863 (N_7863,N_6812,N_6169);
or U7864 (N_7864,N_6356,N_6912);
nor U7865 (N_7865,N_6236,N_6566);
nor U7866 (N_7866,N_6268,N_6046);
or U7867 (N_7867,N_6717,N_6650);
and U7868 (N_7868,N_6125,N_6396);
nand U7869 (N_7869,N_6401,N_6436);
nor U7870 (N_7870,N_6832,N_6793);
xnor U7871 (N_7871,N_6152,N_6936);
xor U7872 (N_7872,N_6520,N_6582);
or U7873 (N_7873,N_6608,N_6067);
xnor U7874 (N_7874,N_6255,N_6981);
or U7875 (N_7875,N_6078,N_6410);
nor U7876 (N_7876,N_6003,N_6998);
or U7877 (N_7877,N_6687,N_6890);
xnor U7878 (N_7878,N_6918,N_6282);
xor U7879 (N_7879,N_6543,N_6772);
xnor U7880 (N_7880,N_6281,N_6838);
xor U7881 (N_7881,N_6785,N_6170);
and U7882 (N_7882,N_6170,N_6478);
or U7883 (N_7883,N_6022,N_6041);
xor U7884 (N_7884,N_6904,N_6785);
or U7885 (N_7885,N_6598,N_6622);
and U7886 (N_7886,N_6378,N_6250);
and U7887 (N_7887,N_6156,N_6014);
nor U7888 (N_7888,N_6454,N_6984);
and U7889 (N_7889,N_6339,N_6203);
nand U7890 (N_7890,N_6930,N_6013);
xor U7891 (N_7891,N_6501,N_6809);
or U7892 (N_7892,N_6237,N_6485);
xnor U7893 (N_7893,N_6505,N_6922);
nor U7894 (N_7894,N_6909,N_6681);
or U7895 (N_7895,N_6877,N_6343);
or U7896 (N_7896,N_6617,N_6373);
nand U7897 (N_7897,N_6729,N_6371);
nand U7898 (N_7898,N_6746,N_6475);
nand U7899 (N_7899,N_6483,N_6660);
nand U7900 (N_7900,N_6135,N_6763);
and U7901 (N_7901,N_6187,N_6164);
or U7902 (N_7902,N_6093,N_6981);
xor U7903 (N_7903,N_6897,N_6495);
and U7904 (N_7904,N_6973,N_6015);
or U7905 (N_7905,N_6206,N_6581);
or U7906 (N_7906,N_6521,N_6328);
nor U7907 (N_7907,N_6004,N_6135);
nand U7908 (N_7908,N_6986,N_6748);
or U7909 (N_7909,N_6084,N_6203);
nor U7910 (N_7910,N_6254,N_6676);
xnor U7911 (N_7911,N_6917,N_6608);
or U7912 (N_7912,N_6720,N_6815);
nor U7913 (N_7913,N_6950,N_6822);
nor U7914 (N_7914,N_6713,N_6577);
and U7915 (N_7915,N_6870,N_6138);
or U7916 (N_7916,N_6272,N_6832);
nor U7917 (N_7917,N_6416,N_6849);
and U7918 (N_7918,N_6430,N_6966);
xnor U7919 (N_7919,N_6727,N_6766);
nand U7920 (N_7920,N_6246,N_6109);
nand U7921 (N_7921,N_6567,N_6352);
nand U7922 (N_7922,N_6654,N_6464);
or U7923 (N_7923,N_6202,N_6203);
xor U7924 (N_7924,N_6478,N_6301);
nand U7925 (N_7925,N_6919,N_6060);
xnor U7926 (N_7926,N_6620,N_6397);
xor U7927 (N_7927,N_6503,N_6685);
nand U7928 (N_7928,N_6603,N_6828);
nor U7929 (N_7929,N_6959,N_6856);
and U7930 (N_7930,N_6273,N_6711);
and U7931 (N_7931,N_6905,N_6883);
and U7932 (N_7932,N_6236,N_6014);
nand U7933 (N_7933,N_6483,N_6251);
nor U7934 (N_7934,N_6721,N_6751);
or U7935 (N_7935,N_6646,N_6567);
xor U7936 (N_7936,N_6077,N_6922);
nor U7937 (N_7937,N_6576,N_6131);
nand U7938 (N_7938,N_6579,N_6883);
nor U7939 (N_7939,N_6734,N_6616);
or U7940 (N_7940,N_6355,N_6279);
or U7941 (N_7941,N_6339,N_6652);
and U7942 (N_7942,N_6530,N_6302);
nor U7943 (N_7943,N_6113,N_6182);
or U7944 (N_7944,N_6974,N_6769);
and U7945 (N_7945,N_6215,N_6090);
nor U7946 (N_7946,N_6182,N_6502);
or U7947 (N_7947,N_6031,N_6220);
and U7948 (N_7948,N_6544,N_6268);
and U7949 (N_7949,N_6017,N_6179);
nor U7950 (N_7950,N_6982,N_6467);
and U7951 (N_7951,N_6948,N_6490);
and U7952 (N_7952,N_6165,N_6987);
and U7953 (N_7953,N_6761,N_6770);
and U7954 (N_7954,N_6239,N_6655);
nor U7955 (N_7955,N_6580,N_6930);
nand U7956 (N_7956,N_6125,N_6695);
nor U7957 (N_7957,N_6244,N_6377);
nand U7958 (N_7958,N_6526,N_6963);
xor U7959 (N_7959,N_6433,N_6337);
or U7960 (N_7960,N_6217,N_6261);
nand U7961 (N_7961,N_6475,N_6507);
nand U7962 (N_7962,N_6398,N_6770);
nand U7963 (N_7963,N_6227,N_6817);
xnor U7964 (N_7964,N_6990,N_6650);
xnor U7965 (N_7965,N_6846,N_6752);
nor U7966 (N_7966,N_6994,N_6128);
or U7967 (N_7967,N_6284,N_6786);
and U7968 (N_7968,N_6034,N_6313);
nor U7969 (N_7969,N_6783,N_6153);
or U7970 (N_7970,N_6472,N_6185);
xnor U7971 (N_7971,N_6186,N_6933);
and U7972 (N_7972,N_6165,N_6317);
or U7973 (N_7973,N_6039,N_6307);
nor U7974 (N_7974,N_6182,N_6123);
nand U7975 (N_7975,N_6491,N_6667);
xor U7976 (N_7976,N_6088,N_6989);
nand U7977 (N_7977,N_6861,N_6072);
nand U7978 (N_7978,N_6802,N_6064);
xnor U7979 (N_7979,N_6312,N_6338);
nor U7980 (N_7980,N_6531,N_6391);
nor U7981 (N_7981,N_6848,N_6796);
or U7982 (N_7982,N_6288,N_6204);
and U7983 (N_7983,N_6751,N_6657);
nor U7984 (N_7984,N_6947,N_6178);
and U7985 (N_7985,N_6547,N_6207);
nor U7986 (N_7986,N_6265,N_6454);
or U7987 (N_7987,N_6820,N_6900);
xor U7988 (N_7988,N_6590,N_6766);
or U7989 (N_7989,N_6720,N_6846);
or U7990 (N_7990,N_6357,N_6913);
and U7991 (N_7991,N_6224,N_6519);
nand U7992 (N_7992,N_6216,N_6152);
and U7993 (N_7993,N_6687,N_6783);
nand U7994 (N_7994,N_6074,N_6620);
and U7995 (N_7995,N_6486,N_6076);
nand U7996 (N_7996,N_6088,N_6408);
and U7997 (N_7997,N_6316,N_6925);
nand U7998 (N_7998,N_6064,N_6066);
nand U7999 (N_7999,N_6650,N_6150);
xnor U8000 (N_8000,N_7338,N_7337);
nand U8001 (N_8001,N_7404,N_7549);
xnor U8002 (N_8002,N_7039,N_7275);
nand U8003 (N_8003,N_7703,N_7194);
and U8004 (N_8004,N_7591,N_7653);
nand U8005 (N_8005,N_7684,N_7802);
nor U8006 (N_8006,N_7371,N_7765);
nand U8007 (N_8007,N_7285,N_7311);
or U8008 (N_8008,N_7236,N_7972);
xnor U8009 (N_8009,N_7139,N_7650);
and U8010 (N_8010,N_7135,N_7836);
nor U8011 (N_8011,N_7983,N_7682);
nand U8012 (N_8012,N_7152,N_7832);
and U8013 (N_8013,N_7671,N_7386);
nor U8014 (N_8014,N_7937,N_7730);
xor U8015 (N_8015,N_7146,N_7925);
nor U8016 (N_8016,N_7278,N_7843);
xor U8017 (N_8017,N_7379,N_7095);
and U8018 (N_8018,N_7279,N_7030);
nand U8019 (N_8019,N_7394,N_7190);
nor U8020 (N_8020,N_7222,N_7536);
and U8021 (N_8021,N_7686,N_7895);
or U8022 (N_8022,N_7851,N_7876);
nand U8023 (N_8023,N_7666,N_7077);
or U8024 (N_8024,N_7089,N_7216);
nor U8025 (N_8025,N_7313,N_7057);
xnor U8026 (N_8026,N_7729,N_7740);
nor U8027 (N_8027,N_7335,N_7233);
nor U8028 (N_8028,N_7797,N_7395);
nor U8029 (N_8029,N_7204,N_7389);
xor U8030 (N_8030,N_7980,N_7610);
or U8031 (N_8031,N_7559,N_7443);
or U8032 (N_8032,N_7970,N_7131);
xor U8033 (N_8033,N_7090,N_7072);
or U8034 (N_8034,N_7017,N_7618);
nand U8035 (N_8035,N_7526,N_7168);
xor U8036 (N_8036,N_7539,N_7396);
nand U8037 (N_8037,N_7174,N_7811);
nand U8038 (N_8038,N_7898,N_7791);
nor U8039 (N_8039,N_7491,N_7670);
nand U8040 (N_8040,N_7059,N_7008);
nand U8041 (N_8041,N_7128,N_7790);
nand U8042 (N_8042,N_7254,N_7614);
and U8043 (N_8043,N_7588,N_7122);
nand U8044 (N_8044,N_7622,N_7264);
or U8045 (N_8045,N_7325,N_7595);
xor U8046 (N_8046,N_7674,N_7697);
xor U8047 (N_8047,N_7213,N_7566);
nor U8048 (N_8048,N_7267,N_7497);
xor U8049 (N_8049,N_7268,N_7466);
xnor U8050 (N_8050,N_7628,N_7091);
or U8051 (N_8051,N_7367,N_7951);
nand U8052 (N_8052,N_7189,N_7726);
or U8053 (N_8053,N_7669,N_7166);
and U8054 (N_8054,N_7570,N_7855);
nor U8055 (N_8055,N_7508,N_7306);
and U8056 (N_8056,N_7144,N_7755);
nor U8057 (N_8057,N_7814,N_7783);
or U8058 (N_8058,N_7961,N_7002);
or U8059 (N_8059,N_7500,N_7935);
or U8060 (N_8060,N_7205,N_7431);
or U8061 (N_8061,N_7083,N_7971);
xnor U8062 (N_8062,N_7833,N_7110);
nand U8063 (N_8063,N_7635,N_7261);
nor U8064 (N_8064,N_7149,N_7303);
or U8065 (N_8065,N_7182,N_7237);
and U8066 (N_8066,N_7027,N_7123);
or U8067 (N_8067,N_7601,N_7247);
and U8068 (N_8068,N_7219,N_7307);
nand U8069 (N_8069,N_7619,N_7578);
nor U8070 (N_8070,N_7258,N_7116);
xor U8071 (N_8071,N_7270,N_7112);
or U8072 (N_8072,N_7555,N_7201);
nor U8073 (N_8073,N_7341,N_7630);
and U8074 (N_8074,N_7522,N_7217);
nand U8075 (N_8075,N_7659,N_7239);
or U8076 (N_8076,N_7881,N_7200);
xor U8077 (N_8077,N_7615,N_7286);
xnor U8078 (N_8078,N_7167,N_7999);
nor U8079 (N_8079,N_7828,N_7933);
nor U8080 (N_8080,N_7469,N_7043);
or U8081 (N_8081,N_7848,N_7481);
xor U8082 (N_8082,N_7033,N_7742);
nor U8083 (N_8083,N_7551,N_7314);
xor U8084 (N_8084,N_7556,N_7862);
nor U8085 (N_8085,N_7645,N_7774);
or U8086 (N_8086,N_7449,N_7022);
nor U8087 (N_8087,N_7102,N_7013);
xnor U8088 (N_8088,N_7098,N_7373);
and U8089 (N_8089,N_7963,N_7932);
and U8090 (N_8090,N_7798,N_7299);
and U8091 (N_8091,N_7710,N_7456);
and U8092 (N_8092,N_7639,N_7274);
nand U8093 (N_8093,N_7507,N_7447);
and U8094 (N_8094,N_7991,N_7725);
and U8095 (N_8095,N_7006,N_7973);
nand U8096 (N_8096,N_7067,N_7781);
and U8097 (N_8097,N_7667,N_7731);
xor U8098 (N_8098,N_7284,N_7520);
nor U8099 (N_8099,N_7966,N_7132);
and U8100 (N_8100,N_7967,N_7483);
xor U8101 (N_8101,N_7179,N_7606);
xnor U8102 (N_8102,N_7418,N_7020);
or U8103 (N_8103,N_7732,N_7575);
nand U8104 (N_8104,N_7332,N_7438);
nand U8105 (N_8105,N_7631,N_7356);
xor U8106 (N_8106,N_7221,N_7711);
nand U8107 (N_8107,N_7545,N_7119);
and U8108 (N_8108,N_7333,N_7212);
or U8109 (N_8109,N_7883,N_7871);
nand U8110 (N_8110,N_7459,N_7127);
nand U8111 (N_8111,N_7478,N_7530);
nand U8112 (N_8112,N_7885,N_7586);
xnor U8113 (N_8113,N_7572,N_7383);
xnor U8114 (N_8114,N_7207,N_7061);
nor U8115 (N_8115,N_7704,N_7318);
and U8116 (N_8116,N_7636,N_7272);
or U8117 (N_8117,N_7692,N_7965);
nand U8118 (N_8118,N_7251,N_7568);
or U8119 (N_8119,N_7501,N_7398);
xnor U8120 (N_8120,N_7060,N_7953);
and U8121 (N_8121,N_7440,N_7712);
or U8122 (N_8122,N_7365,N_7620);
nand U8123 (N_8123,N_7197,N_7256);
and U8124 (N_8124,N_7822,N_7206);
nand U8125 (N_8125,N_7596,N_7734);
nor U8126 (N_8126,N_7126,N_7849);
xor U8127 (N_8127,N_7745,N_7698);
xnor U8128 (N_8128,N_7915,N_7085);
nand U8129 (N_8129,N_7433,N_7467);
nor U8130 (N_8130,N_7019,N_7218);
nand U8131 (N_8131,N_7374,N_7576);
and U8132 (N_8132,N_7185,N_7052);
and U8133 (N_8133,N_7056,N_7942);
or U8134 (N_8134,N_7838,N_7042);
and U8135 (N_8135,N_7864,N_7954);
nor U8136 (N_8136,N_7529,N_7661);
and U8137 (N_8137,N_7416,N_7524);
nor U8138 (N_8138,N_7171,N_7273);
nand U8139 (N_8139,N_7762,N_7426);
nand U8140 (N_8140,N_7839,N_7489);
nand U8141 (N_8141,N_7191,N_7326);
and U8142 (N_8142,N_7600,N_7347);
or U8143 (N_8143,N_7423,N_7125);
and U8144 (N_8144,N_7114,N_7118);
nand U8145 (N_8145,N_7321,N_7805);
nor U8146 (N_8146,N_7892,N_7238);
nand U8147 (N_8147,N_7514,N_7796);
nand U8148 (N_8148,N_7888,N_7612);
and U8149 (N_8149,N_7176,N_7121);
nand U8150 (N_8150,N_7998,N_7437);
nand U8151 (N_8151,N_7384,N_7150);
nand U8152 (N_8152,N_7947,N_7164);
nand U8153 (N_8153,N_7241,N_7728);
or U8154 (N_8154,N_7457,N_7390);
or U8155 (N_8155,N_7768,N_7611);
nand U8156 (N_8156,N_7293,N_7535);
and U8157 (N_8157,N_7436,N_7608);
nor U8158 (N_8158,N_7700,N_7156);
or U8159 (N_8159,N_7751,N_7282);
or U8160 (N_8160,N_7941,N_7754);
or U8161 (N_8161,N_7801,N_7175);
xnor U8162 (N_8162,N_7415,N_7845);
nand U8163 (N_8163,N_7869,N_7603);
xnor U8164 (N_8164,N_7368,N_7914);
xor U8165 (N_8165,N_7472,N_7657);
and U8166 (N_8166,N_7081,N_7632);
or U8167 (N_8167,N_7353,N_7046);
or U8168 (N_8168,N_7070,N_7155);
xor U8169 (N_8169,N_7561,N_7547);
or U8170 (N_8170,N_7789,N_7548);
and U8171 (N_8171,N_7652,N_7761);
nor U8172 (N_8172,N_7880,N_7263);
nor U8173 (N_8173,N_7230,N_7111);
and U8174 (N_8174,N_7706,N_7370);
nand U8175 (N_8175,N_7658,N_7439);
nor U8176 (N_8176,N_7930,N_7253);
or U8177 (N_8177,N_7430,N_7360);
nor U8178 (N_8178,N_7224,N_7997);
or U8179 (N_8179,N_7492,N_7460);
or U8180 (N_8180,N_7872,N_7289);
or U8181 (N_8181,N_7688,N_7054);
nand U8182 (N_8182,N_7562,N_7651);
or U8183 (N_8183,N_7976,N_7104);
nand U8184 (N_8184,N_7494,N_7388);
nand U8185 (N_8185,N_7040,N_7151);
xor U8186 (N_8186,N_7598,N_7879);
and U8187 (N_8187,N_7908,N_7475);
or U8188 (N_8188,N_7000,N_7707);
or U8189 (N_8189,N_7228,N_7162);
or U8190 (N_8190,N_7778,N_7719);
or U8191 (N_8191,N_7032,N_7034);
nand U8192 (N_8192,N_7115,N_7567);
nor U8193 (N_8193,N_7560,N_7901);
or U8194 (N_8194,N_7451,N_7243);
nand U8195 (N_8195,N_7486,N_7249);
xnor U8196 (N_8196,N_7504,N_7777);
or U8197 (N_8197,N_7304,N_7994);
nor U8198 (N_8198,N_7375,N_7772);
and U8199 (N_8199,N_7775,N_7943);
nand U8200 (N_8200,N_7960,N_7737);
xnor U8201 (N_8201,N_7633,N_7904);
xor U8202 (N_8202,N_7830,N_7266);
xnor U8203 (N_8203,N_7533,N_7012);
nor U8204 (N_8204,N_7875,N_7782);
xor U8205 (N_8205,N_7184,N_7747);
nand U8206 (N_8206,N_7993,N_7767);
or U8207 (N_8207,N_7799,N_7294);
nor U8208 (N_8208,N_7290,N_7579);
and U8209 (N_8209,N_7495,N_7038);
and U8210 (N_8210,N_7288,N_7183);
nor U8211 (N_8211,N_7242,N_7084);
nor U8212 (N_8212,N_7844,N_7945);
xnor U8213 (N_8213,N_7235,N_7834);
and U8214 (N_8214,N_7865,N_7105);
nand U8215 (N_8215,N_7886,N_7434);
nor U8216 (N_8216,N_7982,N_7385);
nand U8217 (N_8217,N_7816,N_7257);
nand U8218 (N_8218,N_7410,N_7949);
nor U8219 (N_8219,N_7117,N_7137);
and U8220 (N_8220,N_7424,N_7563);
or U8221 (N_8221,N_7392,N_7784);
nand U8222 (N_8222,N_7071,N_7455);
nand U8223 (N_8223,N_7705,N_7690);
and U8224 (N_8224,N_7902,N_7234);
nor U8225 (N_8225,N_7157,N_7853);
and U8226 (N_8226,N_7382,N_7172);
nor U8227 (N_8227,N_7984,N_7452);
and U8228 (N_8228,N_7571,N_7014);
and U8229 (N_8229,N_7854,N_7764);
nor U8230 (N_8230,N_7316,N_7011);
or U8231 (N_8231,N_7987,N_7295);
xnor U8232 (N_8232,N_7401,N_7047);
nand U8233 (N_8233,N_7859,N_7330);
nand U8234 (N_8234,N_7557,N_7752);
and U8235 (N_8235,N_7897,N_7417);
and U8236 (N_8236,N_7153,N_7992);
and U8237 (N_8237,N_7372,N_7540);
nand U8238 (N_8238,N_7893,N_7795);
xor U8239 (N_8239,N_7887,N_7203);
nand U8240 (N_8240,N_7281,N_7169);
nand U8241 (N_8241,N_7969,N_7996);
nor U8242 (N_8242,N_7597,N_7470);
xor U8243 (N_8243,N_7718,N_7160);
nor U8244 (N_8244,N_7465,N_7148);
and U8245 (N_8245,N_7856,N_7036);
and U8246 (N_8246,N_7346,N_7884);
nand U8247 (N_8247,N_7924,N_7709);
or U8248 (N_8248,N_7532,N_7505);
nor U8249 (N_8249,N_7065,N_7894);
nor U8250 (N_8250,N_7178,N_7911);
nand U8251 (N_8251,N_7124,N_7988);
nand U8252 (N_8252,N_7340,N_7058);
nand U8253 (N_8253,N_7785,N_7106);
xnor U8254 (N_8254,N_7735,N_7513);
or U8255 (N_8255,N_7696,N_7616);
nand U8256 (N_8256,N_7521,N_7739);
nor U8257 (N_8257,N_7007,N_7021);
or U8258 (N_8258,N_7920,N_7818);
nand U8259 (N_8259,N_7344,N_7399);
and U8260 (N_8260,N_7581,N_7419);
and U8261 (N_8261,N_7005,N_7823);
nor U8262 (N_8262,N_7827,N_7644);
nand U8263 (N_8263,N_7870,N_7599);
xnor U8264 (N_8264,N_7051,N_7558);
or U8265 (N_8265,N_7621,N_7956);
nand U8266 (N_8266,N_7045,N_7035);
nor U8267 (N_8267,N_7411,N_7432);
nor U8268 (N_8268,N_7202,N_7946);
and U8269 (N_8269,N_7861,N_7262);
xnor U8270 (N_8270,N_7107,N_7917);
nor U8271 (N_8271,N_7287,N_7097);
or U8272 (N_8272,N_7354,N_7462);
and U8273 (N_8273,N_7769,N_7975);
nor U8274 (N_8274,N_7912,N_7758);
nand U8275 (N_8275,N_7076,N_7297);
xnor U8276 (N_8276,N_7713,N_7680);
nand U8277 (N_8277,N_7493,N_7477);
and U8278 (N_8278,N_7952,N_7271);
and U8279 (N_8279,N_7503,N_7627);
nor U8280 (N_8280,N_7406,N_7049);
or U8281 (N_8281,N_7453,N_7589);
and U8282 (N_8282,N_7582,N_7499);
nor U8283 (N_8283,N_7309,N_7677);
or U8284 (N_8284,N_7231,N_7868);
xnor U8285 (N_8285,N_7403,N_7334);
and U8286 (N_8286,N_7746,N_7794);
xor U8287 (N_8287,N_7319,N_7974);
or U8288 (N_8288,N_7420,N_7245);
nor U8289 (N_8289,N_7770,N_7177);
xor U8290 (N_8290,N_7874,N_7140);
nand U8291 (N_8291,N_7276,N_7594);
or U8292 (N_8292,N_7336,N_7929);
xnor U8293 (N_8293,N_7681,N_7847);
xnor U8294 (N_8294,N_7301,N_7479);
xor U8295 (N_8295,N_7683,N_7867);
and U8296 (N_8296,N_7348,N_7691);
xnor U8297 (N_8297,N_7638,N_7792);
and U8298 (N_8298,N_7074,N_7400);
nand U8299 (N_8299,N_7381,N_7302);
or U8300 (N_8300,N_7665,N_7041);
and U8301 (N_8301,N_7574,N_7078);
or U8302 (N_8302,N_7414,N_7749);
nor U8303 (N_8303,N_7429,N_7580);
and U8304 (N_8304,N_7850,N_7444);
and U8305 (N_8305,N_7656,N_7412);
nand U8306 (N_8306,N_7181,N_7938);
nand U8307 (N_8307,N_7248,N_7776);
or U8308 (N_8308,N_7722,N_7048);
or U8309 (N_8309,N_7685,N_7223);
and U8310 (N_8310,N_7468,N_7590);
nor U8311 (N_8311,N_7349,N_7625);
or U8312 (N_8312,N_7646,N_7094);
nand U8313 (N_8313,N_7748,N_7523);
nand U8314 (N_8314,N_7806,N_7023);
nand U8315 (N_8315,N_7981,N_7068);
nand U8316 (N_8316,N_7442,N_7130);
or U8317 (N_8317,N_7723,N_7721);
or U8318 (N_8318,N_7655,N_7905);
or U8319 (N_8319,N_7810,N_7339);
and U8320 (N_8320,N_7376,N_7458);
nor U8321 (N_8321,N_7446,N_7516);
xnor U8322 (N_8322,N_7787,N_7741);
and U8323 (N_8323,N_7528,N_7018);
nor U8324 (N_8324,N_7198,N_7583);
nor U8325 (N_8325,N_7957,N_7727);
xor U8326 (N_8326,N_7824,N_7990);
nand U8327 (N_8327,N_7485,N_7715);
xnor U8328 (N_8328,N_7858,N_7147);
nand U8329 (N_8329,N_7100,N_7793);
or U8330 (N_8330,N_7744,N_7195);
xnor U8331 (N_8331,N_7544,N_7968);
xnor U8332 (N_8332,N_7931,N_7812);
and U8333 (N_8333,N_7634,N_7369);
nor U8334 (N_8334,N_7129,N_7642);
xor U8335 (N_8335,N_7408,N_7617);
nand U8336 (N_8336,N_7866,N_7199);
xnor U8337 (N_8337,N_7808,N_7232);
and U8338 (N_8338,N_7250,N_7531);
nand U8339 (N_8339,N_7387,N_7154);
nand U8340 (N_8340,N_7565,N_7592);
nand U8341 (N_8341,N_7362,N_7327);
xnor U8342 (N_8342,N_7517,N_7577);
nor U8343 (N_8343,N_7675,N_7377);
xnor U8344 (N_8344,N_7649,N_7672);
xor U8345 (N_8345,N_7936,N_7890);
or U8346 (N_8346,N_7380,N_7629);
xnor U8347 (N_8347,N_7817,N_7978);
nor U8348 (N_8348,N_7800,N_7161);
nor U8349 (N_8349,N_7724,N_7063);
nor U8350 (N_8350,N_7743,N_7819);
nor U8351 (N_8351,N_7831,N_7480);
and U8352 (N_8352,N_7322,N_7214);
nand U8353 (N_8353,N_7538,N_7977);
or U8354 (N_8354,N_7320,N_7964);
nor U8355 (N_8355,N_7196,N_7702);
nor U8356 (N_8356,N_7210,N_7757);
nand U8357 (N_8357,N_7613,N_7720);
and U8358 (N_8358,N_7463,N_7676);
xor U8359 (N_8359,N_7053,N_7641);
nand U8360 (N_8360,N_7050,N_7317);
xor U8361 (N_8361,N_7693,N_7878);
or U8362 (N_8362,N_7552,N_7343);
or U8363 (N_8363,N_7986,N_7476);
xor U8364 (N_8364,N_7813,N_7873);
xor U8365 (N_8365,N_7413,N_7069);
xnor U8366 (N_8366,N_7010,N_7277);
nor U8367 (N_8367,N_7846,N_7393);
nand U8368 (N_8368,N_7525,N_7640);
and U8369 (N_8369,N_7510,N_7269);
or U8370 (N_8370,N_7860,N_7308);
nor U8371 (N_8371,N_7298,N_7515);
and U8372 (N_8372,N_7733,N_7989);
and U8373 (N_8373,N_7821,N_7291);
nor U8374 (N_8374,N_7995,N_7882);
nand U8375 (N_8375,N_7170,N_7009);
and U8376 (N_8376,N_7351,N_7402);
or U8377 (N_8377,N_7695,N_7918);
xor U8378 (N_8378,N_7427,N_7226);
or U8379 (N_8379,N_7923,N_7760);
and U8380 (N_8380,N_7328,N_7546);
xnor U8381 (N_8381,N_7029,N_7766);
nor U8382 (N_8382,N_7910,N_7073);
nor U8383 (N_8383,N_7461,N_7842);
nand U8384 (N_8384,N_7031,N_7227);
and U8385 (N_8385,N_7450,N_7209);
and U8386 (N_8386,N_7422,N_7738);
xnor U8387 (N_8387,N_7300,N_7584);
nor U8388 (N_8388,N_7096,N_7959);
nor U8389 (N_8389,N_7934,N_7877);
nor U8390 (N_8390,N_7717,N_7490);
and U8391 (N_8391,N_7134,N_7950);
and U8392 (N_8392,N_7701,N_7357);
and U8393 (N_8393,N_7143,N_7771);
nor U8394 (N_8394,N_7750,N_7948);
nor U8395 (N_8395,N_7407,N_7962);
or U8396 (N_8396,N_7891,N_7678);
nand U8397 (N_8397,N_7906,N_7165);
and U8398 (N_8398,N_7654,N_7927);
xnor U8399 (N_8399,N_7305,N_7448);
xnor U8400 (N_8400,N_7840,N_7225);
or U8401 (N_8401,N_7928,N_7315);
nor U8402 (N_8402,N_7679,N_7378);
xnor U8403 (N_8403,N_7240,N_7716);
nor U8404 (N_8404,N_7292,N_7896);
xor U8405 (N_8405,N_7044,N_7296);
xor U8406 (N_8406,N_7786,N_7807);
or U8407 (N_8407,N_7841,N_7086);
nor U8408 (N_8408,N_7331,N_7421);
xnor U8409 (N_8409,N_7425,N_7364);
xor U8410 (N_8410,N_7759,N_7173);
or U8411 (N_8411,N_7511,N_7926);
or U8412 (N_8412,N_7265,N_7913);
or U8413 (N_8413,N_7055,N_7820);
nor U8414 (N_8414,N_7604,N_7359);
nor U8415 (N_8415,N_7145,N_7099);
nand U8416 (N_8416,N_7863,N_7028);
and U8417 (N_8417,N_7687,N_7163);
or U8418 (N_8418,N_7773,N_7138);
and U8419 (N_8419,N_7133,N_7158);
xor U8420 (N_8420,N_7358,N_7916);
or U8421 (N_8421,N_7673,N_7648);
and U8422 (N_8422,N_7136,N_7985);
nor U8423 (N_8423,N_7829,N_7899);
nand U8424 (N_8424,N_7087,N_7889);
and U8425 (N_8425,N_7454,N_7944);
or U8426 (N_8426,N_7260,N_7668);
and U8427 (N_8427,N_7310,N_7405);
nor U8428 (N_8428,N_7736,N_7815);
and U8429 (N_8429,N_7512,N_7519);
nor U8430 (N_8430,N_7804,N_7474);
nor U8431 (N_8431,N_7763,N_7082);
or U8432 (N_8432,N_7391,N_7958);
xnor U8433 (N_8433,N_7255,N_7662);
or U8434 (N_8434,N_7498,N_7361);
nand U8435 (N_8435,N_7909,N_7602);
nor U8436 (N_8436,N_7192,N_7252);
and U8437 (N_8437,N_7626,N_7441);
and U8438 (N_8438,N_7496,N_7312);
or U8439 (N_8439,N_7837,N_7624);
or U8440 (N_8440,N_7229,N_7088);
or U8441 (N_8441,N_7428,N_7016);
nand U8442 (N_8442,N_7109,N_7756);
and U8443 (N_8443,N_7694,N_7825);
xnor U8444 (N_8444,N_7553,N_7593);
xor U8445 (N_8445,N_7664,N_7003);
nor U8446 (N_8446,N_7955,N_7780);
nor U8447 (N_8447,N_7092,N_7488);
nand U8448 (N_8448,N_7605,N_7001);
nand U8449 (N_8449,N_7788,N_7159);
xnor U8450 (N_8450,N_7919,N_7004);
and U8451 (N_8451,N_7506,N_7409);
nor U8452 (N_8452,N_7141,N_7075);
nor U8453 (N_8453,N_7120,N_7329);
nand U8454 (N_8454,N_7607,N_7093);
and U8455 (N_8455,N_7259,N_7643);
or U8456 (N_8456,N_7852,N_7623);
xor U8457 (N_8457,N_7907,N_7066);
and U8458 (N_8458,N_7903,N_7473);
and U8459 (N_8459,N_7324,N_7220);
and U8460 (N_8460,N_7509,N_7699);
xor U8461 (N_8461,N_7366,N_7283);
and U8462 (N_8462,N_7541,N_7355);
nor U8463 (N_8463,N_7024,N_7064);
and U8464 (N_8464,N_7564,N_7803);
and U8465 (N_8465,N_7482,N_7527);
xnor U8466 (N_8466,N_7835,N_7542);
nand U8467 (N_8467,N_7080,N_7663);
nor U8468 (N_8468,N_7714,N_7464);
nor U8469 (N_8469,N_7534,N_7826);
nand U8470 (N_8470,N_7689,N_7939);
or U8471 (N_8471,N_7979,N_7609);
nor U8472 (N_8472,N_7113,N_7637);
and U8473 (N_8473,N_7779,N_7108);
nand U8474 (N_8474,N_7350,N_7484);
or U8475 (N_8475,N_7026,N_7211);
or U8476 (N_8476,N_7940,N_7587);
nand U8477 (N_8477,N_7922,N_7537);
and U8478 (N_8478,N_7244,N_7037);
xnor U8479 (N_8479,N_7708,N_7208);
xnor U8480 (N_8480,N_7345,N_7015);
and U8481 (N_8481,N_7554,N_7397);
or U8482 (N_8482,N_7857,N_7550);
and U8483 (N_8483,N_7585,N_7363);
nor U8484 (N_8484,N_7573,N_7215);
nand U8485 (N_8485,N_7079,N_7180);
nor U8486 (N_8486,N_7569,N_7900);
nand U8487 (N_8487,N_7062,N_7647);
nand U8488 (N_8488,N_7188,N_7660);
xnor U8489 (N_8489,N_7025,N_7502);
nor U8490 (N_8490,N_7352,N_7543);
xor U8491 (N_8491,N_7487,N_7445);
or U8492 (N_8492,N_7342,N_7753);
nor U8493 (N_8493,N_7280,N_7921);
nor U8494 (N_8494,N_7323,N_7246);
nand U8495 (N_8495,N_7187,N_7193);
nor U8496 (N_8496,N_7471,N_7809);
or U8497 (N_8497,N_7186,N_7103);
xnor U8498 (N_8498,N_7101,N_7518);
and U8499 (N_8499,N_7435,N_7142);
nor U8500 (N_8500,N_7339,N_7920);
and U8501 (N_8501,N_7897,N_7477);
nand U8502 (N_8502,N_7927,N_7123);
or U8503 (N_8503,N_7120,N_7897);
or U8504 (N_8504,N_7492,N_7436);
nor U8505 (N_8505,N_7870,N_7347);
or U8506 (N_8506,N_7285,N_7313);
xor U8507 (N_8507,N_7504,N_7121);
and U8508 (N_8508,N_7863,N_7374);
xnor U8509 (N_8509,N_7619,N_7225);
or U8510 (N_8510,N_7769,N_7481);
nand U8511 (N_8511,N_7401,N_7109);
nor U8512 (N_8512,N_7163,N_7275);
nand U8513 (N_8513,N_7676,N_7772);
and U8514 (N_8514,N_7726,N_7103);
xor U8515 (N_8515,N_7747,N_7219);
and U8516 (N_8516,N_7632,N_7292);
xor U8517 (N_8517,N_7684,N_7996);
nor U8518 (N_8518,N_7279,N_7256);
nand U8519 (N_8519,N_7391,N_7695);
nand U8520 (N_8520,N_7153,N_7465);
nor U8521 (N_8521,N_7137,N_7251);
or U8522 (N_8522,N_7681,N_7839);
or U8523 (N_8523,N_7174,N_7920);
xnor U8524 (N_8524,N_7221,N_7222);
nand U8525 (N_8525,N_7682,N_7414);
and U8526 (N_8526,N_7125,N_7639);
or U8527 (N_8527,N_7503,N_7496);
nor U8528 (N_8528,N_7290,N_7765);
nor U8529 (N_8529,N_7992,N_7410);
nor U8530 (N_8530,N_7308,N_7244);
xor U8531 (N_8531,N_7252,N_7787);
or U8532 (N_8532,N_7260,N_7390);
and U8533 (N_8533,N_7628,N_7205);
nand U8534 (N_8534,N_7723,N_7948);
nand U8535 (N_8535,N_7664,N_7356);
nor U8536 (N_8536,N_7266,N_7369);
nor U8537 (N_8537,N_7598,N_7797);
and U8538 (N_8538,N_7164,N_7521);
nand U8539 (N_8539,N_7816,N_7247);
and U8540 (N_8540,N_7222,N_7447);
nand U8541 (N_8541,N_7532,N_7868);
xnor U8542 (N_8542,N_7181,N_7500);
nand U8543 (N_8543,N_7759,N_7842);
and U8544 (N_8544,N_7775,N_7054);
nor U8545 (N_8545,N_7692,N_7150);
and U8546 (N_8546,N_7263,N_7505);
and U8547 (N_8547,N_7287,N_7506);
nor U8548 (N_8548,N_7345,N_7802);
or U8549 (N_8549,N_7182,N_7492);
and U8550 (N_8550,N_7958,N_7198);
nor U8551 (N_8551,N_7615,N_7763);
xnor U8552 (N_8552,N_7169,N_7986);
nor U8553 (N_8553,N_7669,N_7990);
xnor U8554 (N_8554,N_7922,N_7110);
xnor U8555 (N_8555,N_7917,N_7675);
xor U8556 (N_8556,N_7772,N_7744);
nor U8557 (N_8557,N_7785,N_7729);
nand U8558 (N_8558,N_7818,N_7142);
nor U8559 (N_8559,N_7440,N_7635);
nor U8560 (N_8560,N_7262,N_7420);
or U8561 (N_8561,N_7125,N_7722);
xor U8562 (N_8562,N_7138,N_7700);
and U8563 (N_8563,N_7092,N_7198);
nand U8564 (N_8564,N_7406,N_7167);
nand U8565 (N_8565,N_7616,N_7598);
and U8566 (N_8566,N_7315,N_7055);
nor U8567 (N_8567,N_7730,N_7544);
or U8568 (N_8568,N_7315,N_7266);
and U8569 (N_8569,N_7055,N_7314);
and U8570 (N_8570,N_7065,N_7562);
and U8571 (N_8571,N_7703,N_7480);
nand U8572 (N_8572,N_7412,N_7052);
xnor U8573 (N_8573,N_7132,N_7103);
nand U8574 (N_8574,N_7147,N_7573);
xnor U8575 (N_8575,N_7958,N_7317);
xor U8576 (N_8576,N_7762,N_7169);
nand U8577 (N_8577,N_7689,N_7509);
nand U8578 (N_8578,N_7852,N_7594);
nor U8579 (N_8579,N_7764,N_7515);
or U8580 (N_8580,N_7029,N_7560);
xnor U8581 (N_8581,N_7539,N_7800);
nand U8582 (N_8582,N_7954,N_7497);
or U8583 (N_8583,N_7722,N_7160);
nor U8584 (N_8584,N_7616,N_7721);
nor U8585 (N_8585,N_7402,N_7867);
and U8586 (N_8586,N_7287,N_7525);
xnor U8587 (N_8587,N_7985,N_7578);
nor U8588 (N_8588,N_7844,N_7489);
xnor U8589 (N_8589,N_7148,N_7280);
xnor U8590 (N_8590,N_7266,N_7268);
or U8591 (N_8591,N_7723,N_7210);
or U8592 (N_8592,N_7953,N_7286);
or U8593 (N_8593,N_7885,N_7030);
or U8594 (N_8594,N_7634,N_7267);
nor U8595 (N_8595,N_7224,N_7598);
and U8596 (N_8596,N_7946,N_7966);
nand U8597 (N_8597,N_7545,N_7378);
nor U8598 (N_8598,N_7455,N_7266);
nand U8599 (N_8599,N_7802,N_7973);
and U8600 (N_8600,N_7057,N_7720);
or U8601 (N_8601,N_7511,N_7591);
and U8602 (N_8602,N_7165,N_7785);
xnor U8603 (N_8603,N_7838,N_7252);
or U8604 (N_8604,N_7612,N_7119);
xor U8605 (N_8605,N_7615,N_7738);
or U8606 (N_8606,N_7345,N_7798);
nand U8607 (N_8607,N_7857,N_7901);
nor U8608 (N_8608,N_7148,N_7799);
or U8609 (N_8609,N_7604,N_7650);
nor U8610 (N_8610,N_7762,N_7591);
nor U8611 (N_8611,N_7773,N_7666);
nand U8612 (N_8612,N_7185,N_7172);
xnor U8613 (N_8613,N_7195,N_7067);
nand U8614 (N_8614,N_7158,N_7390);
nor U8615 (N_8615,N_7937,N_7622);
nor U8616 (N_8616,N_7089,N_7347);
nor U8617 (N_8617,N_7768,N_7755);
xor U8618 (N_8618,N_7094,N_7551);
xor U8619 (N_8619,N_7892,N_7374);
or U8620 (N_8620,N_7122,N_7650);
or U8621 (N_8621,N_7327,N_7263);
and U8622 (N_8622,N_7645,N_7923);
xor U8623 (N_8623,N_7291,N_7399);
xnor U8624 (N_8624,N_7827,N_7417);
or U8625 (N_8625,N_7585,N_7775);
xnor U8626 (N_8626,N_7956,N_7346);
xor U8627 (N_8627,N_7777,N_7856);
nand U8628 (N_8628,N_7703,N_7464);
xnor U8629 (N_8629,N_7961,N_7484);
nor U8630 (N_8630,N_7234,N_7075);
nand U8631 (N_8631,N_7829,N_7617);
nor U8632 (N_8632,N_7662,N_7817);
nand U8633 (N_8633,N_7757,N_7947);
and U8634 (N_8634,N_7691,N_7408);
nand U8635 (N_8635,N_7601,N_7605);
or U8636 (N_8636,N_7334,N_7314);
nand U8637 (N_8637,N_7208,N_7612);
and U8638 (N_8638,N_7607,N_7155);
or U8639 (N_8639,N_7428,N_7632);
or U8640 (N_8640,N_7645,N_7734);
nor U8641 (N_8641,N_7794,N_7862);
nand U8642 (N_8642,N_7200,N_7512);
xnor U8643 (N_8643,N_7232,N_7024);
nand U8644 (N_8644,N_7450,N_7512);
nand U8645 (N_8645,N_7385,N_7853);
and U8646 (N_8646,N_7852,N_7134);
nand U8647 (N_8647,N_7369,N_7127);
nor U8648 (N_8648,N_7371,N_7845);
or U8649 (N_8649,N_7240,N_7809);
nand U8650 (N_8650,N_7725,N_7528);
or U8651 (N_8651,N_7572,N_7241);
and U8652 (N_8652,N_7017,N_7737);
nor U8653 (N_8653,N_7256,N_7523);
nand U8654 (N_8654,N_7917,N_7741);
nand U8655 (N_8655,N_7817,N_7571);
and U8656 (N_8656,N_7892,N_7009);
and U8657 (N_8657,N_7709,N_7784);
and U8658 (N_8658,N_7772,N_7356);
nor U8659 (N_8659,N_7148,N_7837);
and U8660 (N_8660,N_7990,N_7112);
and U8661 (N_8661,N_7215,N_7500);
nor U8662 (N_8662,N_7652,N_7567);
xnor U8663 (N_8663,N_7529,N_7134);
nand U8664 (N_8664,N_7706,N_7705);
xnor U8665 (N_8665,N_7448,N_7169);
xnor U8666 (N_8666,N_7115,N_7313);
nand U8667 (N_8667,N_7408,N_7308);
nor U8668 (N_8668,N_7501,N_7533);
nor U8669 (N_8669,N_7439,N_7563);
or U8670 (N_8670,N_7163,N_7156);
or U8671 (N_8671,N_7174,N_7205);
and U8672 (N_8672,N_7832,N_7403);
or U8673 (N_8673,N_7259,N_7258);
xnor U8674 (N_8674,N_7070,N_7311);
xnor U8675 (N_8675,N_7942,N_7051);
or U8676 (N_8676,N_7303,N_7773);
xor U8677 (N_8677,N_7870,N_7543);
and U8678 (N_8678,N_7944,N_7215);
nand U8679 (N_8679,N_7743,N_7439);
and U8680 (N_8680,N_7869,N_7025);
and U8681 (N_8681,N_7915,N_7937);
or U8682 (N_8682,N_7037,N_7939);
nand U8683 (N_8683,N_7395,N_7326);
or U8684 (N_8684,N_7130,N_7162);
or U8685 (N_8685,N_7307,N_7410);
nor U8686 (N_8686,N_7480,N_7660);
or U8687 (N_8687,N_7568,N_7076);
nor U8688 (N_8688,N_7689,N_7695);
nor U8689 (N_8689,N_7674,N_7787);
or U8690 (N_8690,N_7661,N_7109);
or U8691 (N_8691,N_7151,N_7414);
xor U8692 (N_8692,N_7390,N_7334);
nand U8693 (N_8693,N_7410,N_7215);
or U8694 (N_8694,N_7102,N_7977);
nand U8695 (N_8695,N_7642,N_7577);
nor U8696 (N_8696,N_7345,N_7661);
and U8697 (N_8697,N_7023,N_7060);
nand U8698 (N_8698,N_7613,N_7845);
xnor U8699 (N_8699,N_7245,N_7673);
nand U8700 (N_8700,N_7814,N_7989);
or U8701 (N_8701,N_7124,N_7047);
and U8702 (N_8702,N_7951,N_7702);
nand U8703 (N_8703,N_7226,N_7194);
nor U8704 (N_8704,N_7985,N_7609);
xnor U8705 (N_8705,N_7347,N_7578);
nand U8706 (N_8706,N_7723,N_7084);
nor U8707 (N_8707,N_7104,N_7200);
or U8708 (N_8708,N_7861,N_7055);
nor U8709 (N_8709,N_7099,N_7579);
or U8710 (N_8710,N_7757,N_7347);
and U8711 (N_8711,N_7828,N_7196);
and U8712 (N_8712,N_7108,N_7339);
nand U8713 (N_8713,N_7372,N_7480);
nand U8714 (N_8714,N_7517,N_7676);
nand U8715 (N_8715,N_7572,N_7678);
or U8716 (N_8716,N_7466,N_7967);
nor U8717 (N_8717,N_7148,N_7142);
nand U8718 (N_8718,N_7596,N_7455);
or U8719 (N_8719,N_7821,N_7493);
nand U8720 (N_8720,N_7590,N_7003);
or U8721 (N_8721,N_7246,N_7408);
and U8722 (N_8722,N_7780,N_7582);
xor U8723 (N_8723,N_7682,N_7779);
xnor U8724 (N_8724,N_7190,N_7705);
nand U8725 (N_8725,N_7638,N_7968);
or U8726 (N_8726,N_7217,N_7674);
nand U8727 (N_8727,N_7756,N_7916);
and U8728 (N_8728,N_7651,N_7216);
and U8729 (N_8729,N_7347,N_7996);
and U8730 (N_8730,N_7691,N_7870);
xnor U8731 (N_8731,N_7533,N_7885);
or U8732 (N_8732,N_7521,N_7264);
nor U8733 (N_8733,N_7336,N_7474);
nor U8734 (N_8734,N_7862,N_7978);
nand U8735 (N_8735,N_7868,N_7338);
xor U8736 (N_8736,N_7061,N_7224);
nand U8737 (N_8737,N_7311,N_7179);
and U8738 (N_8738,N_7269,N_7630);
xor U8739 (N_8739,N_7718,N_7244);
nor U8740 (N_8740,N_7071,N_7263);
and U8741 (N_8741,N_7249,N_7528);
and U8742 (N_8742,N_7119,N_7942);
and U8743 (N_8743,N_7850,N_7571);
nand U8744 (N_8744,N_7728,N_7710);
or U8745 (N_8745,N_7804,N_7857);
nor U8746 (N_8746,N_7811,N_7545);
nand U8747 (N_8747,N_7730,N_7326);
and U8748 (N_8748,N_7268,N_7844);
and U8749 (N_8749,N_7085,N_7595);
and U8750 (N_8750,N_7706,N_7890);
nand U8751 (N_8751,N_7089,N_7584);
or U8752 (N_8752,N_7186,N_7283);
xor U8753 (N_8753,N_7074,N_7069);
and U8754 (N_8754,N_7250,N_7619);
and U8755 (N_8755,N_7688,N_7342);
xor U8756 (N_8756,N_7102,N_7240);
or U8757 (N_8757,N_7770,N_7134);
xor U8758 (N_8758,N_7435,N_7233);
nor U8759 (N_8759,N_7692,N_7938);
or U8760 (N_8760,N_7451,N_7654);
or U8761 (N_8761,N_7590,N_7185);
and U8762 (N_8762,N_7245,N_7519);
and U8763 (N_8763,N_7638,N_7380);
xor U8764 (N_8764,N_7561,N_7891);
and U8765 (N_8765,N_7175,N_7971);
nand U8766 (N_8766,N_7525,N_7373);
or U8767 (N_8767,N_7355,N_7081);
nand U8768 (N_8768,N_7228,N_7115);
xor U8769 (N_8769,N_7113,N_7749);
nand U8770 (N_8770,N_7616,N_7144);
and U8771 (N_8771,N_7235,N_7054);
xnor U8772 (N_8772,N_7882,N_7375);
and U8773 (N_8773,N_7358,N_7373);
nor U8774 (N_8774,N_7477,N_7505);
and U8775 (N_8775,N_7993,N_7234);
or U8776 (N_8776,N_7337,N_7672);
xnor U8777 (N_8777,N_7611,N_7032);
nand U8778 (N_8778,N_7362,N_7245);
xnor U8779 (N_8779,N_7379,N_7796);
xor U8780 (N_8780,N_7385,N_7480);
or U8781 (N_8781,N_7075,N_7378);
or U8782 (N_8782,N_7758,N_7977);
and U8783 (N_8783,N_7597,N_7680);
nor U8784 (N_8784,N_7219,N_7354);
and U8785 (N_8785,N_7877,N_7792);
and U8786 (N_8786,N_7984,N_7332);
nand U8787 (N_8787,N_7053,N_7697);
or U8788 (N_8788,N_7569,N_7358);
nand U8789 (N_8789,N_7075,N_7920);
xnor U8790 (N_8790,N_7112,N_7625);
nand U8791 (N_8791,N_7747,N_7251);
and U8792 (N_8792,N_7201,N_7408);
and U8793 (N_8793,N_7944,N_7202);
xnor U8794 (N_8794,N_7836,N_7794);
nor U8795 (N_8795,N_7167,N_7091);
and U8796 (N_8796,N_7743,N_7356);
or U8797 (N_8797,N_7981,N_7913);
nand U8798 (N_8798,N_7537,N_7651);
nand U8799 (N_8799,N_7645,N_7714);
or U8800 (N_8800,N_7123,N_7351);
or U8801 (N_8801,N_7784,N_7583);
or U8802 (N_8802,N_7378,N_7163);
nand U8803 (N_8803,N_7571,N_7792);
or U8804 (N_8804,N_7143,N_7694);
nand U8805 (N_8805,N_7817,N_7417);
nand U8806 (N_8806,N_7882,N_7418);
or U8807 (N_8807,N_7315,N_7833);
nand U8808 (N_8808,N_7635,N_7632);
nor U8809 (N_8809,N_7381,N_7563);
nor U8810 (N_8810,N_7564,N_7387);
nand U8811 (N_8811,N_7889,N_7248);
or U8812 (N_8812,N_7051,N_7764);
and U8813 (N_8813,N_7266,N_7754);
xnor U8814 (N_8814,N_7523,N_7710);
xor U8815 (N_8815,N_7901,N_7347);
xnor U8816 (N_8816,N_7716,N_7973);
or U8817 (N_8817,N_7309,N_7993);
nor U8818 (N_8818,N_7077,N_7091);
or U8819 (N_8819,N_7459,N_7462);
nor U8820 (N_8820,N_7357,N_7984);
and U8821 (N_8821,N_7221,N_7208);
and U8822 (N_8822,N_7905,N_7604);
nand U8823 (N_8823,N_7124,N_7612);
and U8824 (N_8824,N_7961,N_7560);
xnor U8825 (N_8825,N_7702,N_7500);
or U8826 (N_8826,N_7832,N_7234);
or U8827 (N_8827,N_7436,N_7785);
or U8828 (N_8828,N_7008,N_7636);
xor U8829 (N_8829,N_7663,N_7079);
nand U8830 (N_8830,N_7040,N_7957);
or U8831 (N_8831,N_7034,N_7921);
nand U8832 (N_8832,N_7175,N_7428);
xnor U8833 (N_8833,N_7726,N_7127);
and U8834 (N_8834,N_7443,N_7609);
nand U8835 (N_8835,N_7082,N_7564);
nand U8836 (N_8836,N_7263,N_7144);
nand U8837 (N_8837,N_7238,N_7207);
nor U8838 (N_8838,N_7901,N_7819);
nor U8839 (N_8839,N_7913,N_7583);
xnor U8840 (N_8840,N_7961,N_7449);
nand U8841 (N_8841,N_7014,N_7655);
nor U8842 (N_8842,N_7693,N_7610);
and U8843 (N_8843,N_7503,N_7050);
nor U8844 (N_8844,N_7066,N_7966);
nand U8845 (N_8845,N_7894,N_7387);
or U8846 (N_8846,N_7692,N_7797);
xnor U8847 (N_8847,N_7166,N_7157);
or U8848 (N_8848,N_7238,N_7404);
and U8849 (N_8849,N_7214,N_7265);
nand U8850 (N_8850,N_7046,N_7406);
or U8851 (N_8851,N_7002,N_7061);
and U8852 (N_8852,N_7128,N_7955);
nor U8853 (N_8853,N_7945,N_7826);
nand U8854 (N_8854,N_7622,N_7932);
nand U8855 (N_8855,N_7180,N_7019);
nor U8856 (N_8856,N_7833,N_7113);
nor U8857 (N_8857,N_7905,N_7305);
nor U8858 (N_8858,N_7775,N_7445);
nor U8859 (N_8859,N_7988,N_7182);
and U8860 (N_8860,N_7716,N_7931);
xnor U8861 (N_8861,N_7581,N_7849);
xnor U8862 (N_8862,N_7881,N_7693);
nand U8863 (N_8863,N_7184,N_7426);
nor U8864 (N_8864,N_7659,N_7828);
or U8865 (N_8865,N_7745,N_7766);
nand U8866 (N_8866,N_7174,N_7719);
or U8867 (N_8867,N_7028,N_7055);
or U8868 (N_8868,N_7535,N_7688);
and U8869 (N_8869,N_7141,N_7177);
nor U8870 (N_8870,N_7425,N_7532);
xor U8871 (N_8871,N_7630,N_7223);
nand U8872 (N_8872,N_7375,N_7069);
nand U8873 (N_8873,N_7764,N_7740);
nand U8874 (N_8874,N_7360,N_7766);
nand U8875 (N_8875,N_7178,N_7298);
nor U8876 (N_8876,N_7691,N_7591);
nand U8877 (N_8877,N_7738,N_7156);
and U8878 (N_8878,N_7404,N_7333);
or U8879 (N_8879,N_7895,N_7243);
nand U8880 (N_8880,N_7626,N_7962);
nand U8881 (N_8881,N_7960,N_7430);
nand U8882 (N_8882,N_7679,N_7802);
and U8883 (N_8883,N_7295,N_7977);
nor U8884 (N_8884,N_7466,N_7103);
xnor U8885 (N_8885,N_7547,N_7584);
and U8886 (N_8886,N_7810,N_7950);
or U8887 (N_8887,N_7923,N_7121);
nand U8888 (N_8888,N_7954,N_7873);
nand U8889 (N_8889,N_7308,N_7176);
or U8890 (N_8890,N_7338,N_7679);
xor U8891 (N_8891,N_7274,N_7704);
or U8892 (N_8892,N_7933,N_7063);
or U8893 (N_8893,N_7713,N_7788);
and U8894 (N_8894,N_7403,N_7421);
and U8895 (N_8895,N_7085,N_7167);
and U8896 (N_8896,N_7241,N_7052);
or U8897 (N_8897,N_7255,N_7633);
nor U8898 (N_8898,N_7058,N_7958);
nand U8899 (N_8899,N_7913,N_7960);
and U8900 (N_8900,N_7508,N_7444);
and U8901 (N_8901,N_7851,N_7689);
nand U8902 (N_8902,N_7029,N_7743);
or U8903 (N_8903,N_7142,N_7673);
xnor U8904 (N_8904,N_7074,N_7383);
and U8905 (N_8905,N_7273,N_7168);
or U8906 (N_8906,N_7829,N_7447);
or U8907 (N_8907,N_7935,N_7075);
nor U8908 (N_8908,N_7423,N_7287);
xor U8909 (N_8909,N_7767,N_7650);
nand U8910 (N_8910,N_7256,N_7158);
xor U8911 (N_8911,N_7481,N_7107);
and U8912 (N_8912,N_7601,N_7694);
nand U8913 (N_8913,N_7093,N_7716);
nor U8914 (N_8914,N_7558,N_7602);
nand U8915 (N_8915,N_7020,N_7994);
nor U8916 (N_8916,N_7458,N_7745);
nor U8917 (N_8917,N_7254,N_7391);
and U8918 (N_8918,N_7904,N_7425);
or U8919 (N_8919,N_7860,N_7117);
nor U8920 (N_8920,N_7498,N_7325);
xnor U8921 (N_8921,N_7929,N_7927);
nor U8922 (N_8922,N_7690,N_7865);
or U8923 (N_8923,N_7157,N_7978);
or U8924 (N_8924,N_7008,N_7227);
and U8925 (N_8925,N_7978,N_7798);
or U8926 (N_8926,N_7378,N_7532);
nor U8927 (N_8927,N_7389,N_7134);
nor U8928 (N_8928,N_7956,N_7871);
nand U8929 (N_8929,N_7944,N_7329);
xnor U8930 (N_8930,N_7420,N_7810);
nor U8931 (N_8931,N_7065,N_7158);
xnor U8932 (N_8932,N_7147,N_7641);
nor U8933 (N_8933,N_7314,N_7412);
or U8934 (N_8934,N_7615,N_7558);
or U8935 (N_8935,N_7580,N_7629);
and U8936 (N_8936,N_7746,N_7369);
nor U8937 (N_8937,N_7216,N_7231);
xnor U8938 (N_8938,N_7595,N_7028);
or U8939 (N_8939,N_7786,N_7223);
nand U8940 (N_8940,N_7932,N_7525);
xnor U8941 (N_8941,N_7472,N_7782);
xnor U8942 (N_8942,N_7981,N_7674);
and U8943 (N_8943,N_7815,N_7483);
and U8944 (N_8944,N_7670,N_7847);
xor U8945 (N_8945,N_7969,N_7124);
and U8946 (N_8946,N_7668,N_7001);
and U8947 (N_8947,N_7792,N_7006);
xor U8948 (N_8948,N_7760,N_7269);
and U8949 (N_8949,N_7281,N_7422);
nand U8950 (N_8950,N_7835,N_7970);
nand U8951 (N_8951,N_7057,N_7620);
or U8952 (N_8952,N_7045,N_7916);
or U8953 (N_8953,N_7012,N_7586);
xor U8954 (N_8954,N_7900,N_7492);
nand U8955 (N_8955,N_7970,N_7572);
xor U8956 (N_8956,N_7862,N_7297);
and U8957 (N_8957,N_7239,N_7688);
and U8958 (N_8958,N_7240,N_7598);
xnor U8959 (N_8959,N_7459,N_7031);
nand U8960 (N_8960,N_7875,N_7236);
and U8961 (N_8961,N_7264,N_7563);
nor U8962 (N_8962,N_7462,N_7327);
and U8963 (N_8963,N_7387,N_7039);
nor U8964 (N_8964,N_7792,N_7323);
xnor U8965 (N_8965,N_7263,N_7899);
nand U8966 (N_8966,N_7886,N_7214);
nor U8967 (N_8967,N_7376,N_7294);
and U8968 (N_8968,N_7654,N_7377);
nor U8969 (N_8969,N_7711,N_7089);
nand U8970 (N_8970,N_7284,N_7434);
nor U8971 (N_8971,N_7069,N_7153);
or U8972 (N_8972,N_7955,N_7206);
and U8973 (N_8973,N_7011,N_7622);
nand U8974 (N_8974,N_7654,N_7976);
nor U8975 (N_8975,N_7299,N_7450);
xnor U8976 (N_8976,N_7369,N_7038);
xnor U8977 (N_8977,N_7118,N_7297);
nor U8978 (N_8978,N_7137,N_7510);
xor U8979 (N_8979,N_7501,N_7091);
or U8980 (N_8980,N_7396,N_7145);
nand U8981 (N_8981,N_7970,N_7244);
and U8982 (N_8982,N_7130,N_7550);
and U8983 (N_8983,N_7501,N_7074);
or U8984 (N_8984,N_7158,N_7699);
nand U8985 (N_8985,N_7183,N_7865);
nor U8986 (N_8986,N_7940,N_7210);
nor U8987 (N_8987,N_7159,N_7916);
nand U8988 (N_8988,N_7920,N_7227);
nor U8989 (N_8989,N_7419,N_7690);
xor U8990 (N_8990,N_7479,N_7657);
or U8991 (N_8991,N_7596,N_7442);
and U8992 (N_8992,N_7997,N_7198);
or U8993 (N_8993,N_7214,N_7173);
xnor U8994 (N_8994,N_7971,N_7673);
nor U8995 (N_8995,N_7252,N_7890);
or U8996 (N_8996,N_7947,N_7134);
and U8997 (N_8997,N_7747,N_7159);
nor U8998 (N_8998,N_7916,N_7820);
or U8999 (N_8999,N_7713,N_7609);
nand U9000 (N_9000,N_8455,N_8293);
nand U9001 (N_9001,N_8625,N_8702);
nand U9002 (N_9002,N_8492,N_8501);
xor U9003 (N_9003,N_8711,N_8729);
and U9004 (N_9004,N_8187,N_8669);
nor U9005 (N_9005,N_8125,N_8812);
and U9006 (N_9006,N_8986,N_8510);
xor U9007 (N_9007,N_8146,N_8860);
xor U9008 (N_9008,N_8328,N_8096);
and U9009 (N_9009,N_8880,N_8943);
nor U9010 (N_9010,N_8514,N_8129);
xor U9011 (N_9011,N_8322,N_8274);
nor U9012 (N_9012,N_8257,N_8407);
and U9013 (N_9013,N_8634,N_8984);
xnor U9014 (N_9014,N_8961,N_8798);
and U9015 (N_9015,N_8408,N_8589);
nor U9016 (N_9016,N_8268,N_8169);
xor U9017 (N_9017,N_8195,N_8043);
nor U9018 (N_9018,N_8562,N_8963);
xor U9019 (N_9019,N_8078,N_8520);
nor U9020 (N_9020,N_8672,N_8664);
nand U9021 (N_9021,N_8436,N_8130);
xor U9022 (N_9022,N_8049,N_8756);
nor U9023 (N_9023,N_8721,N_8347);
xor U9024 (N_9024,N_8720,N_8228);
and U9025 (N_9025,N_8114,N_8444);
nor U9026 (N_9026,N_8661,N_8369);
xnor U9027 (N_9027,N_8632,N_8240);
nand U9028 (N_9028,N_8512,N_8251);
nor U9029 (N_9029,N_8449,N_8784);
nor U9030 (N_9030,N_8184,N_8713);
xnor U9031 (N_9031,N_8331,N_8023);
nor U9032 (N_9032,N_8068,N_8121);
or U9033 (N_9033,N_8222,N_8133);
nand U9034 (N_9034,N_8806,N_8811);
nand U9035 (N_9035,N_8818,N_8925);
xnor U9036 (N_9036,N_8715,N_8662);
nor U9037 (N_9037,N_8103,N_8160);
nand U9038 (N_9038,N_8147,N_8016);
or U9039 (N_9039,N_8326,N_8092);
or U9040 (N_9040,N_8550,N_8522);
and U9041 (N_9041,N_8909,N_8760);
or U9042 (N_9042,N_8693,N_8728);
xnor U9043 (N_9043,N_8906,N_8137);
nand U9044 (N_9044,N_8248,N_8486);
nand U9045 (N_9045,N_8259,N_8588);
xor U9046 (N_9046,N_8979,N_8694);
xor U9047 (N_9047,N_8150,N_8519);
xnor U9048 (N_9048,N_8262,N_8992);
xor U9049 (N_9049,N_8610,N_8091);
nor U9050 (N_9050,N_8928,N_8143);
nand U9051 (N_9051,N_8463,N_8071);
nand U9052 (N_9052,N_8033,N_8960);
or U9053 (N_9053,N_8354,N_8592);
nor U9054 (N_9054,N_8215,N_8843);
or U9055 (N_9055,N_8095,N_8243);
nand U9056 (N_9056,N_8457,N_8573);
or U9057 (N_9057,N_8930,N_8586);
or U9058 (N_9058,N_8485,N_8738);
or U9059 (N_9059,N_8281,N_8036);
or U9060 (N_9060,N_8163,N_8288);
and U9061 (N_9061,N_8964,N_8168);
and U9062 (N_9062,N_8295,N_8052);
nand U9063 (N_9063,N_8236,N_8336);
or U9064 (N_9064,N_8265,N_8731);
xor U9065 (N_9065,N_8136,N_8997);
nand U9066 (N_9066,N_8681,N_8734);
nand U9067 (N_9067,N_8374,N_8406);
and U9068 (N_9068,N_8633,N_8099);
nand U9069 (N_9069,N_8749,N_8151);
xnor U9070 (N_9070,N_8403,N_8948);
and U9071 (N_9071,N_8161,N_8772);
xnor U9072 (N_9072,N_8080,N_8689);
or U9073 (N_9073,N_8093,N_8856);
and U9074 (N_9074,N_8500,N_8932);
xor U9075 (N_9075,N_8936,N_8207);
or U9076 (N_9076,N_8767,N_8356);
or U9077 (N_9077,N_8303,N_8175);
and U9078 (N_9078,N_8778,N_8552);
nand U9079 (N_9079,N_8167,N_8660);
or U9080 (N_9080,N_8947,N_8199);
xor U9081 (N_9081,N_8145,N_8282);
nor U9082 (N_9082,N_8088,N_8365);
xor U9083 (N_9083,N_8608,N_8206);
nand U9084 (N_9084,N_8885,N_8978);
xor U9085 (N_9085,N_8035,N_8927);
nor U9086 (N_9086,N_8431,N_8008);
nand U9087 (N_9087,N_8998,N_8312);
or U9088 (N_9088,N_8413,N_8679);
and U9089 (N_9089,N_8733,N_8718);
or U9090 (N_9090,N_8159,N_8613);
nand U9091 (N_9091,N_8626,N_8332);
xnor U9092 (N_9092,N_8044,N_8034);
xnor U9093 (N_9093,N_8793,N_8781);
nand U9094 (N_9094,N_8995,N_8646);
xor U9095 (N_9095,N_8657,N_8438);
nand U9096 (N_9096,N_8063,N_8824);
and U9097 (N_9097,N_8357,N_8323);
or U9098 (N_9098,N_8029,N_8275);
nand U9099 (N_9099,N_8764,N_8178);
nor U9100 (N_9100,N_8162,N_8518);
and U9101 (N_9101,N_8344,N_8920);
and U9102 (N_9102,N_8118,N_8046);
and U9103 (N_9103,N_8981,N_8405);
nor U9104 (N_9104,N_8391,N_8922);
and U9105 (N_9105,N_8081,N_8094);
or U9106 (N_9106,N_8242,N_8083);
nand U9107 (N_9107,N_8513,N_8667);
xnor U9108 (N_9108,N_8192,N_8075);
or U9109 (N_9109,N_8434,N_8830);
or U9110 (N_9110,N_8329,N_8845);
xor U9111 (N_9111,N_8805,N_8107);
xor U9112 (N_9112,N_8316,N_8591);
xor U9113 (N_9113,N_8226,N_8865);
nand U9114 (N_9114,N_8498,N_8571);
nor U9115 (N_9115,N_8676,N_8213);
nand U9116 (N_9116,N_8011,N_8367);
xor U9117 (N_9117,N_8604,N_8655);
nor U9118 (N_9118,N_8335,N_8266);
xnor U9119 (N_9119,N_8577,N_8284);
and U9120 (N_9120,N_8637,N_8358);
nand U9121 (N_9121,N_8801,N_8024);
nor U9122 (N_9122,N_8966,N_8901);
and U9123 (N_9123,N_8229,N_8690);
nand U9124 (N_9124,N_8197,N_8031);
nor U9125 (N_9125,N_8503,N_8467);
and U9126 (N_9126,N_8330,N_8461);
or U9127 (N_9127,N_8410,N_8051);
and U9128 (N_9128,N_8452,N_8460);
or U9129 (N_9129,N_8735,N_8343);
nand U9130 (N_9130,N_8447,N_8134);
or U9131 (N_9131,N_8258,N_8726);
xnor U9132 (N_9132,N_8196,N_8320);
nor U9133 (N_9133,N_8446,N_8070);
nand U9134 (N_9134,N_8556,N_8048);
xor U9135 (N_9135,N_8530,N_8314);
or U9136 (N_9136,N_8889,N_8013);
xor U9137 (N_9137,N_8509,N_8494);
nor U9138 (N_9138,N_8302,N_8837);
xor U9139 (N_9139,N_8705,N_8482);
nor U9140 (N_9140,N_8053,N_8983);
nand U9141 (N_9141,N_8506,N_8560);
and U9142 (N_9142,N_8601,N_8527);
nand U9143 (N_9143,N_8794,N_8808);
nor U9144 (N_9144,N_8952,N_8565);
and U9145 (N_9145,N_8618,N_8249);
and U9146 (N_9146,N_8290,N_8683);
nor U9147 (N_9147,N_8973,N_8116);
nor U9148 (N_9148,N_8531,N_8916);
nor U9149 (N_9149,N_8933,N_8473);
nand U9150 (N_9150,N_8766,N_8980);
or U9151 (N_9151,N_8027,N_8895);
xor U9152 (N_9152,N_8976,N_8832);
nor U9153 (N_9153,N_8021,N_8722);
nand U9154 (N_9154,N_8435,N_8006);
and U9155 (N_9155,N_8623,N_8292);
nand U9156 (N_9156,N_8624,N_8521);
xnor U9157 (N_9157,N_8792,N_8466);
nor U9158 (N_9158,N_8516,N_8703);
and U9159 (N_9159,N_8727,N_8084);
nand U9160 (N_9160,N_8595,N_8324);
nor U9161 (N_9161,N_8507,N_8777);
and U9162 (N_9162,N_8594,N_8924);
xor U9163 (N_9163,N_8174,N_8279);
xnor U9164 (N_9164,N_8969,N_8361);
and U9165 (N_9165,N_8650,N_8775);
or U9166 (N_9166,N_8014,N_8834);
nand U9167 (N_9167,N_8640,N_8779);
xnor U9168 (N_9168,N_8555,N_8350);
nand U9169 (N_9169,N_8119,N_8931);
nor U9170 (N_9170,N_8250,N_8934);
nor U9171 (N_9171,N_8086,N_8212);
nor U9172 (N_9172,N_8042,N_8656);
xor U9173 (N_9173,N_8993,N_8892);
nor U9174 (N_9174,N_8047,N_8607);
nor U9175 (N_9175,N_8180,N_8870);
xor U9176 (N_9176,N_8977,N_8581);
and U9177 (N_9177,N_8688,N_8788);
nand U9178 (N_9178,N_8989,N_8611);
nand U9179 (N_9179,N_8816,N_8959);
or U9180 (N_9180,N_8614,N_8897);
and U9181 (N_9181,N_8627,N_8907);
or U9182 (N_9182,N_8224,N_8419);
xor U9183 (N_9183,N_8123,N_8910);
nor U9184 (N_9184,N_8553,N_8575);
or U9185 (N_9185,N_8110,N_8642);
xnor U9186 (N_9186,N_8474,N_8493);
nand U9187 (N_9187,N_8797,N_8803);
and U9188 (N_9188,N_8183,N_8709);
and U9189 (N_9189,N_8790,N_8090);
and U9190 (N_9190,N_8317,N_8451);
nand U9191 (N_9191,N_8719,N_8082);
or U9192 (N_9192,N_8732,N_8990);
xor U9193 (N_9193,N_8040,N_8372);
nand U9194 (N_9194,N_8970,N_8489);
and U9195 (N_9195,N_8478,N_8508);
xnor U9196 (N_9196,N_8505,N_8165);
nor U9197 (N_9197,N_8415,N_8746);
nand U9198 (N_9198,N_8132,N_8201);
or U9199 (N_9199,N_8126,N_8872);
and U9200 (N_9200,N_8246,N_8205);
or U9201 (N_9201,N_8371,N_8422);
or U9202 (N_9202,N_8352,N_8386);
or U9203 (N_9203,N_8379,N_8346);
nor U9204 (N_9204,N_8437,N_8914);
and U9205 (N_9205,N_8341,N_8252);
or U9206 (N_9206,N_8349,N_8950);
and U9207 (N_9207,N_8537,N_8216);
nor U9208 (N_9208,N_8737,N_8138);
nor U9209 (N_9209,N_8334,N_8270);
nand U9210 (N_9210,N_8750,N_8076);
and U9211 (N_9211,N_8484,N_8769);
and U9212 (N_9212,N_8428,N_8390);
and U9213 (N_9213,N_8432,N_8267);
and U9214 (N_9214,N_8392,N_8987);
nor U9215 (N_9215,N_8840,N_8238);
nor U9216 (N_9216,N_8762,N_8652);
nor U9217 (N_9217,N_8533,N_8563);
nor U9218 (N_9218,N_8260,N_8574);
nor U9219 (N_9219,N_8389,N_8402);
xor U9220 (N_9220,N_8751,N_8115);
or U9221 (N_9221,N_8300,N_8225);
nor U9222 (N_9222,N_8409,N_8597);
nand U9223 (N_9223,N_8459,N_8450);
or U9224 (N_9224,N_8894,N_8230);
nand U9225 (N_9225,N_8638,N_8668);
xor U9226 (N_9226,N_8810,N_8758);
or U9227 (N_9227,N_8140,N_8898);
or U9228 (N_9228,N_8570,N_8915);
and U9229 (N_9229,N_8855,N_8218);
xnor U9230 (N_9230,N_8139,N_8665);
or U9231 (N_9231,N_8704,N_8158);
nand U9232 (N_9232,N_8965,N_8542);
nand U9233 (N_9233,N_8191,N_8888);
nand U9234 (N_9234,N_8237,N_8534);
nor U9235 (N_9235,N_8425,N_8429);
xnor U9236 (N_9236,N_8862,N_8340);
and U9237 (N_9237,N_8185,N_8838);
xnor U9238 (N_9238,N_8217,N_8972);
nand U9239 (N_9239,N_8325,N_8453);
nor U9240 (N_9240,N_8141,N_8214);
nand U9241 (N_9241,N_8182,N_8541);
and U9242 (N_9242,N_8710,N_8069);
nor U9243 (N_9243,N_8658,N_8113);
or U9244 (N_9244,N_8471,N_8800);
nand U9245 (N_9245,N_8748,N_8327);
nor U9246 (N_9246,N_8348,N_8686);
or U9247 (N_9247,N_8020,N_8698);
or U9248 (N_9248,N_8026,N_8653);
or U9249 (N_9249,N_8497,N_8120);
xor U9250 (N_9250,N_8062,N_8255);
xnor U9251 (N_9251,N_8397,N_8313);
xor U9252 (N_9252,N_8079,N_8787);
or U9253 (N_9253,N_8526,N_8421);
xnor U9254 (N_9254,N_8765,N_8401);
or U9255 (N_9255,N_8286,N_8414);
nor U9256 (N_9256,N_8942,N_8337);
xor U9257 (N_9257,N_8028,N_8476);
or U9258 (N_9258,N_8636,N_8622);
nand U9259 (N_9259,N_8572,N_8417);
and U9260 (N_9260,N_8100,N_8022);
xor U9261 (N_9261,N_8612,N_8564);
xnor U9262 (N_9262,N_8481,N_8770);
nand U9263 (N_9263,N_8321,N_8700);
xnor U9264 (N_9264,N_8420,N_8373);
nand U9265 (N_9265,N_8523,N_8831);
or U9266 (N_9266,N_8864,N_8842);
or U9267 (N_9267,N_8559,N_8905);
xnor U9268 (N_9268,N_8598,N_8863);
xnor U9269 (N_9269,N_8954,N_8558);
nor U9270 (N_9270,N_8566,N_8089);
and U9271 (N_9271,N_8495,N_8030);
nor U9272 (N_9272,N_8101,N_8861);
and U9273 (N_9273,N_8108,N_8768);
nand U9274 (N_9274,N_8621,N_8946);
or U9275 (N_9275,N_8227,N_8005);
nand U9276 (N_9276,N_8234,N_8850);
nor U9277 (N_9277,N_8283,N_8848);
and U9278 (N_9278,N_8730,N_8269);
nand U9279 (N_9279,N_8382,N_8561);
and U9280 (N_9280,N_8418,N_8362);
nand U9281 (N_9281,N_8487,N_8194);
and U9282 (N_9282,N_8189,N_8873);
xnor U9283 (N_9283,N_8469,N_8599);
and U9284 (N_9284,N_8568,N_8411);
xnor U9285 (N_9285,N_8551,N_8822);
xnor U9286 (N_9286,N_8456,N_8355);
nor U9287 (N_9287,N_8833,N_8651);
nand U9288 (N_9288,N_8783,N_8398);
nand U9289 (N_9289,N_8780,N_8529);
and U9290 (N_9290,N_8935,N_8917);
xnor U9291 (N_9291,N_8821,N_8789);
xnor U9292 (N_9292,N_8576,N_8839);
or U9293 (N_9293,N_8706,N_8799);
nor U9294 (N_9294,N_8585,N_8105);
xnor U9295 (N_9295,N_8368,N_8254);
xor U9296 (N_9296,N_8874,N_8241);
and U9297 (N_9297,N_8176,N_8817);
nand U9298 (N_9298,N_8433,N_8524);
or U9299 (N_9299,N_8996,N_8315);
or U9300 (N_9300,N_8659,N_8015);
nand U9301 (N_9301,N_8741,N_8219);
xnor U9302 (N_9302,N_8223,N_8142);
nand U9303 (N_9303,N_8815,N_8829);
and U9304 (N_9304,N_8232,N_8807);
or U9305 (N_9305,N_8605,N_8695);
and U9306 (N_9306,N_8804,N_8066);
xor U9307 (N_9307,N_8630,N_8654);
nand U9308 (N_9308,N_8745,N_8544);
or U9309 (N_9309,N_8464,N_8802);
nor U9310 (N_9310,N_8032,N_8380);
nand U9311 (N_9311,N_8525,N_8479);
and U9312 (N_9312,N_8554,N_8423);
or U9313 (N_9313,N_8543,N_8294);
xor U9314 (N_9314,N_8887,N_8763);
nor U9315 (N_9315,N_8825,N_8170);
xor U9316 (N_9316,N_8716,N_8913);
and U9317 (N_9317,N_8691,N_8809);
xor U9318 (N_9318,N_8603,N_8773);
nand U9319 (N_9319,N_8619,N_8424);
nand U9320 (N_9320,N_8221,N_8940);
or U9321 (N_9321,N_8871,N_8155);
nor U9322 (N_9322,N_8548,N_8412);
nor U9323 (N_9323,N_8853,N_8007);
or U9324 (N_9324,N_8173,N_8287);
nor U9325 (N_9325,N_8649,N_8579);
nand U9326 (N_9326,N_8009,N_8462);
xnor U9327 (N_9327,N_8220,N_8299);
nand U9328 (N_9328,N_8122,N_8955);
nand U9329 (N_9329,N_8128,N_8298);
xor U9330 (N_9330,N_8854,N_8231);
xnor U9331 (N_9331,N_8276,N_8515);
nand U9332 (N_9332,N_8465,N_8974);
nor U9333 (N_9333,N_8057,N_8306);
or U9334 (N_9334,N_8210,N_8430);
and U9335 (N_9335,N_8496,N_8426);
nand U9336 (N_9336,N_8442,N_8208);
nor U9337 (N_9337,N_8073,N_8580);
and U9338 (N_9338,N_8074,N_8304);
and U9339 (N_9339,N_8645,N_8037);
xnor U9340 (N_9340,N_8929,N_8439);
xor U9341 (N_9341,N_8038,N_8491);
xnor U9342 (N_9342,N_8823,N_8557);
nor U9343 (N_9343,N_8443,N_8743);
nor U9344 (N_9344,N_8814,N_8307);
or U9345 (N_9345,N_8752,N_8875);
and U9346 (N_9346,N_8985,N_8852);
xnor U9347 (N_9347,N_8866,N_8584);
xor U9348 (N_9348,N_8911,N_8319);
and U9349 (N_9349,N_8345,N_8578);
nand U9350 (N_9350,N_8893,N_8629);
and U9351 (N_9351,N_8360,N_8488);
nand U9352 (N_9352,N_8841,N_8097);
xnor U9353 (N_9353,N_8648,N_8697);
xor U9354 (N_9354,N_8958,N_8245);
nand U9355 (N_9355,N_8971,N_8416);
nor U9356 (N_9356,N_8725,N_8171);
xnor U9357 (N_9357,N_8918,N_8087);
xnor U9358 (N_9358,N_8593,N_8540);
or U9359 (N_9359,N_8851,N_8945);
nand U9360 (N_9360,N_8209,N_8342);
nor U9361 (N_9361,N_8261,N_8263);
and U9362 (N_9362,N_8050,N_8318);
xor U9363 (N_9363,N_8545,N_8253);
or U9364 (N_9364,N_8065,N_8826);
nand U9365 (N_9365,N_8297,N_8441);
nor U9366 (N_9366,N_8882,N_8363);
xnor U9367 (N_9367,N_8387,N_8127);
xor U9368 (N_9368,N_8289,N_8647);
or U9369 (N_9369,N_8061,N_8747);
nor U9370 (N_9370,N_8939,N_8724);
nand U9371 (N_9371,N_8333,N_8239);
or U9372 (N_9372,N_8117,N_8017);
and U9373 (N_9373,N_8754,N_8628);
xor U9374 (N_9374,N_8054,N_8394);
nand U9375 (N_9375,N_8277,N_8723);
or U9376 (N_9376,N_8502,N_8736);
xnor U9377 (N_9377,N_8609,N_8211);
nor U9378 (N_9378,N_8759,N_8285);
and U9379 (N_9379,N_8098,N_8708);
or U9380 (N_9380,N_8004,N_8532);
and U9381 (N_9381,N_8663,N_8152);
nand U9382 (N_9382,N_8166,N_8908);
and U9383 (N_9383,N_8511,N_8796);
nand U9384 (N_9384,N_8890,N_8353);
nand U9385 (N_9385,N_8366,N_8714);
nand U9386 (N_9386,N_8309,N_8280);
or U9387 (N_9387,N_8472,N_8926);
and U9388 (N_9388,N_8666,N_8968);
and U9389 (N_9389,N_8190,N_8549);
or U9390 (N_9390,N_8883,N_8962);
xor U9391 (N_9391,N_8153,N_8771);
or U9392 (N_9392,N_8002,N_8644);
xnor U9393 (N_9393,N_8782,N_8739);
nor U9394 (N_9394,N_8587,N_8235);
xnor U9395 (N_9395,N_8813,N_8154);
nand U9396 (N_9396,N_8202,N_8677);
nand U9397 (N_9397,N_8606,N_8836);
and U9398 (N_9398,N_8675,N_8085);
or U9399 (N_9399,N_8991,N_8041);
nor U9400 (N_9400,N_8753,N_8761);
xnor U9401 (N_9401,N_8396,N_8200);
nor U9402 (N_9402,N_8844,N_8000);
xnor U9403 (N_9403,N_8203,N_8381);
and U9404 (N_9404,N_8567,N_8018);
nor U9405 (N_9405,N_8899,N_8643);
or U9406 (N_9406,N_8827,N_8384);
nand U9407 (N_9407,N_8311,N_8602);
or U9408 (N_9408,N_8470,N_8858);
nor U9409 (N_9409,N_8359,N_8148);
and U9410 (N_9410,N_8308,N_8164);
nor U9411 (N_9411,N_8468,N_8059);
or U9412 (N_9412,N_8272,N_8448);
nor U9413 (N_9413,N_8835,N_8600);
xnor U9414 (N_9414,N_8849,N_8596);
nand U9415 (N_9415,N_8291,N_8937);
xnor U9416 (N_9416,N_8440,N_8135);
xor U9417 (N_9417,N_8956,N_8338);
or U9418 (N_9418,N_8064,N_8376);
nor U9419 (N_9419,N_8884,N_8699);
and U9420 (N_9420,N_8701,N_8301);
nor U9421 (N_9421,N_8941,N_8454);
nand U9422 (N_9422,N_8186,N_8427);
nor U9423 (N_9423,N_8635,N_8399);
nor U9424 (N_9424,N_8896,N_8535);
nand U9425 (N_9425,N_8538,N_8395);
and U9426 (N_9426,N_8177,N_8475);
or U9427 (N_9427,N_8999,N_8179);
xor U9428 (N_9428,N_8785,N_8483);
nor U9429 (N_9429,N_8383,N_8639);
xnor U9430 (N_9430,N_8003,N_8903);
or U9431 (N_9431,N_8058,N_8921);
and U9432 (N_9432,N_8204,N_8388);
xor U9433 (N_9433,N_8755,N_8846);
and U9434 (N_9434,N_8717,N_8687);
nor U9435 (N_9435,N_8919,N_8019);
xor U9436 (N_9436,N_8867,N_8377);
nand U9437 (N_9437,N_8902,N_8685);
and U9438 (N_9438,N_8504,N_8692);
nor U9439 (N_9439,N_8957,N_8539);
or U9440 (N_9440,N_8680,N_8536);
and U9441 (N_9441,N_8631,N_8517);
and U9442 (N_9442,N_8776,N_8445);
nor U9443 (N_9443,N_8857,N_8891);
nand U9444 (N_9444,N_8795,N_8616);
nor U9445 (N_9445,N_8944,N_8144);
and U9446 (N_9446,N_8244,N_8296);
xnor U9447 (N_9447,N_8982,N_8696);
nor U9448 (N_9448,N_8351,N_8271);
and U9449 (N_9449,N_8615,N_8673);
and U9450 (N_9450,N_8278,N_8923);
and U9451 (N_9451,N_8157,N_8247);
nor U9452 (N_9452,N_8879,N_8385);
or U9453 (N_9453,N_8378,N_8617);
or U9454 (N_9454,N_8975,N_8547);
xor U9455 (N_9455,N_8111,N_8106);
and U9456 (N_9456,N_8156,N_8869);
xnor U9457 (N_9457,N_8112,N_8364);
and U9458 (N_9458,N_8400,N_8757);
nand U9459 (N_9459,N_8868,N_8045);
nor U9460 (N_9460,N_8791,N_8499);
xnor U9461 (N_9461,N_8264,N_8273);
or U9462 (N_9462,N_8370,N_8994);
xor U9463 (N_9463,N_8786,N_8149);
and U9464 (N_9464,N_8740,N_8012);
nor U9465 (N_9465,N_8582,N_8109);
nor U9466 (N_9466,N_8967,N_8198);
nand U9467 (N_9467,N_8193,N_8181);
or U9468 (N_9468,N_8490,N_8819);
and U9469 (N_9469,N_8912,N_8712);
xor U9470 (N_9470,N_8641,N_8859);
nor U9471 (N_9471,N_8404,N_8876);
xor U9472 (N_9472,N_8707,N_8671);
xor U9473 (N_9473,N_8010,N_8077);
and U9474 (N_9474,N_8900,N_8393);
nor U9475 (N_9475,N_8678,N_8056);
nand U9476 (N_9476,N_8375,N_8477);
or U9477 (N_9477,N_8820,N_8886);
nor U9478 (N_9478,N_8256,N_8951);
nor U9479 (N_9479,N_8590,N_8774);
nand U9480 (N_9480,N_8124,N_8339);
and U9481 (N_9481,N_8172,N_8072);
nor U9482 (N_9482,N_8949,N_8480);
nor U9483 (N_9483,N_8233,N_8847);
xnor U9484 (N_9484,N_8001,N_8188);
nor U9485 (N_9485,N_8039,N_8938);
or U9486 (N_9486,N_8528,N_8674);
or U9487 (N_9487,N_8682,N_8988);
xor U9488 (N_9488,N_8878,N_8670);
or U9489 (N_9489,N_8828,N_8104);
nor U9490 (N_9490,N_8877,N_8742);
and U9491 (N_9491,N_8102,N_8744);
and U9492 (N_9492,N_8305,N_8569);
xor U9493 (N_9493,N_8131,N_8546);
xnor U9494 (N_9494,N_8025,N_8310);
and U9495 (N_9495,N_8583,N_8067);
xor U9496 (N_9496,N_8620,N_8684);
or U9497 (N_9497,N_8055,N_8953);
nand U9498 (N_9498,N_8881,N_8060);
nand U9499 (N_9499,N_8904,N_8458);
or U9500 (N_9500,N_8665,N_8449);
or U9501 (N_9501,N_8851,N_8342);
and U9502 (N_9502,N_8771,N_8295);
xor U9503 (N_9503,N_8636,N_8170);
xnor U9504 (N_9504,N_8042,N_8621);
or U9505 (N_9505,N_8506,N_8109);
xnor U9506 (N_9506,N_8463,N_8736);
or U9507 (N_9507,N_8394,N_8284);
or U9508 (N_9508,N_8252,N_8628);
nand U9509 (N_9509,N_8207,N_8574);
or U9510 (N_9510,N_8715,N_8951);
or U9511 (N_9511,N_8792,N_8033);
nand U9512 (N_9512,N_8646,N_8407);
xnor U9513 (N_9513,N_8117,N_8659);
nor U9514 (N_9514,N_8998,N_8559);
nor U9515 (N_9515,N_8387,N_8656);
or U9516 (N_9516,N_8973,N_8520);
nor U9517 (N_9517,N_8852,N_8429);
xor U9518 (N_9518,N_8996,N_8491);
xnor U9519 (N_9519,N_8823,N_8266);
nand U9520 (N_9520,N_8733,N_8806);
nor U9521 (N_9521,N_8505,N_8751);
xor U9522 (N_9522,N_8712,N_8228);
nand U9523 (N_9523,N_8573,N_8233);
xor U9524 (N_9524,N_8665,N_8841);
xnor U9525 (N_9525,N_8081,N_8767);
nor U9526 (N_9526,N_8789,N_8313);
or U9527 (N_9527,N_8878,N_8463);
xor U9528 (N_9528,N_8038,N_8904);
and U9529 (N_9529,N_8554,N_8716);
xor U9530 (N_9530,N_8505,N_8302);
nor U9531 (N_9531,N_8182,N_8721);
and U9532 (N_9532,N_8799,N_8701);
nand U9533 (N_9533,N_8713,N_8216);
nand U9534 (N_9534,N_8149,N_8672);
and U9535 (N_9535,N_8402,N_8919);
xor U9536 (N_9536,N_8870,N_8513);
xor U9537 (N_9537,N_8348,N_8127);
or U9538 (N_9538,N_8165,N_8871);
xor U9539 (N_9539,N_8741,N_8409);
nor U9540 (N_9540,N_8825,N_8600);
nand U9541 (N_9541,N_8527,N_8730);
nand U9542 (N_9542,N_8155,N_8277);
xnor U9543 (N_9543,N_8843,N_8999);
xnor U9544 (N_9544,N_8750,N_8855);
and U9545 (N_9545,N_8304,N_8779);
nand U9546 (N_9546,N_8085,N_8335);
and U9547 (N_9547,N_8698,N_8888);
xnor U9548 (N_9548,N_8045,N_8483);
nor U9549 (N_9549,N_8166,N_8273);
or U9550 (N_9550,N_8028,N_8186);
or U9551 (N_9551,N_8014,N_8449);
or U9552 (N_9552,N_8082,N_8507);
or U9553 (N_9553,N_8124,N_8971);
nand U9554 (N_9554,N_8863,N_8088);
or U9555 (N_9555,N_8802,N_8828);
nand U9556 (N_9556,N_8423,N_8533);
and U9557 (N_9557,N_8927,N_8928);
xor U9558 (N_9558,N_8058,N_8569);
xor U9559 (N_9559,N_8409,N_8187);
and U9560 (N_9560,N_8533,N_8431);
nand U9561 (N_9561,N_8382,N_8207);
nor U9562 (N_9562,N_8883,N_8879);
and U9563 (N_9563,N_8466,N_8631);
nand U9564 (N_9564,N_8809,N_8909);
or U9565 (N_9565,N_8533,N_8034);
nor U9566 (N_9566,N_8002,N_8843);
or U9567 (N_9567,N_8678,N_8523);
nor U9568 (N_9568,N_8652,N_8632);
and U9569 (N_9569,N_8177,N_8981);
nand U9570 (N_9570,N_8424,N_8036);
nor U9571 (N_9571,N_8650,N_8186);
nor U9572 (N_9572,N_8346,N_8689);
nand U9573 (N_9573,N_8188,N_8466);
xnor U9574 (N_9574,N_8135,N_8192);
nand U9575 (N_9575,N_8552,N_8690);
nor U9576 (N_9576,N_8371,N_8702);
xor U9577 (N_9577,N_8747,N_8927);
xor U9578 (N_9578,N_8109,N_8314);
nand U9579 (N_9579,N_8013,N_8234);
xor U9580 (N_9580,N_8204,N_8554);
nor U9581 (N_9581,N_8599,N_8687);
nor U9582 (N_9582,N_8515,N_8953);
nor U9583 (N_9583,N_8215,N_8580);
and U9584 (N_9584,N_8710,N_8070);
or U9585 (N_9585,N_8337,N_8556);
xor U9586 (N_9586,N_8748,N_8164);
xor U9587 (N_9587,N_8589,N_8650);
xnor U9588 (N_9588,N_8534,N_8881);
nand U9589 (N_9589,N_8433,N_8529);
and U9590 (N_9590,N_8121,N_8419);
nand U9591 (N_9591,N_8813,N_8832);
and U9592 (N_9592,N_8749,N_8252);
and U9593 (N_9593,N_8657,N_8529);
nor U9594 (N_9594,N_8471,N_8237);
and U9595 (N_9595,N_8483,N_8014);
xor U9596 (N_9596,N_8545,N_8143);
xnor U9597 (N_9597,N_8152,N_8531);
nand U9598 (N_9598,N_8497,N_8101);
nor U9599 (N_9599,N_8159,N_8296);
nand U9600 (N_9600,N_8851,N_8431);
xnor U9601 (N_9601,N_8221,N_8083);
and U9602 (N_9602,N_8300,N_8043);
nor U9603 (N_9603,N_8499,N_8842);
xnor U9604 (N_9604,N_8700,N_8188);
nand U9605 (N_9605,N_8811,N_8404);
nor U9606 (N_9606,N_8271,N_8605);
nand U9607 (N_9607,N_8756,N_8031);
or U9608 (N_9608,N_8860,N_8083);
nor U9609 (N_9609,N_8430,N_8328);
or U9610 (N_9610,N_8569,N_8846);
and U9611 (N_9611,N_8842,N_8717);
or U9612 (N_9612,N_8661,N_8278);
nand U9613 (N_9613,N_8738,N_8868);
xnor U9614 (N_9614,N_8878,N_8205);
nand U9615 (N_9615,N_8618,N_8736);
nand U9616 (N_9616,N_8166,N_8763);
and U9617 (N_9617,N_8445,N_8458);
nor U9618 (N_9618,N_8306,N_8908);
or U9619 (N_9619,N_8344,N_8046);
nand U9620 (N_9620,N_8756,N_8333);
or U9621 (N_9621,N_8902,N_8125);
and U9622 (N_9622,N_8006,N_8922);
and U9623 (N_9623,N_8687,N_8780);
and U9624 (N_9624,N_8154,N_8584);
or U9625 (N_9625,N_8600,N_8842);
nor U9626 (N_9626,N_8019,N_8416);
and U9627 (N_9627,N_8813,N_8448);
nand U9628 (N_9628,N_8258,N_8580);
nand U9629 (N_9629,N_8063,N_8564);
or U9630 (N_9630,N_8076,N_8276);
and U9631 (N_9631,N_8733,N_8675);
nand U9632 (N_9632,N_8075,N_8838);
xnor U9633 (N_9633,N_8119,N_8430);
nor U9634 (N_9634,N_8482,N_8623);
or U9635 (N_9635,N_8645,N_8188);
or U9636 (N_9636,N_8181,N_8689);
nand U9637 (N_9637,N_8087,N_8396);
xnor U9638 (N_9638,N_8009,N_8053);
nor U9639 (N_9639,N_8823,N_8902);
nor U9640 (N_9640,N_8150,N_8618);
nand U9641 (N_9641,N_8614,N_8770);
xor U9642 (N_9642,N_8791,N_8778);
xor U9643 (N_9643,N_8153,N_8468);
xnor U9644 (N_9644,N_8622,N_8089);
and U9645 (N_9645,N_8251,N_8104);
xor U9646 (N_9646,N_8459,N_8124);
or U9647 (N_9647,N_8033,N_8313);
xnor U9648 (N_9648,N_8781,N_8695);
xor U9649 (N_9649,N_8810,N_8075);
nand U9650 (N_9650,N_8972,N_8024);
xor U9651 (N_9651,N_8420,N_8064);
nand U9652 (N_9652,N_8946,N_8779);
nor U9653 (N_9653,N_8027,N_8335);
and U9654 (N_9654,N_8805,N_8286);
nor U9655 (N_9655,N_8354,N_8771);
xnor U9656 (N_9656,N_8212,N_8168);
nand U9657 (N_9657,N_8743,N_8147);
and U9658 (N_9658,N_8690,N_8344);
and U9659 (N_9659,N_8640,N_8480);
nand U9660 (N_9660,N_8503,N_8135);
or U9661 (N_9661,N_8138,N_8853);
and U9662 (N_9662,N_8534,N_8365);
and U9663 (N_9663,N_8691,N_8473);
or U9664 (N_9664,N_8862,N_8803);
and U9665 (N_9665,N_8162,N_8381);
or U9666 (N_9666,N_8099,N_8168);
nor U9667 (N_9667,N_8689,N_8205);
or U9668 (N_9668,N_8811,N_8371);
nor U9669 (N_9669,N_8723,N_8510);
and U9670 (N_9670,N_8260,N_8073);
and U9671 (N_9671,N_8675,N_8632);
nand U9672 (N_9672,N_8245,N_8091);
nand U9673 (N_9673,N_8396,N_8342);
nor U9674 (N_9674,N_8211,N_8392);
xor U9675 (N_9675,N_8765,N_8034);
or U9676 (N_9676,N_8152,N_8075);
xor U9677 (N_9677,N_8724,N_8793);
nand U9678 (N_9678,N_8275,N_8909);
and U9679 (N_9679,N_8977,N_8117);
nand U9680 (N_9680,N_8810,N_8046);
or U9681 (N_9681,N_8155,N_8355);
and U9682 (N_9682,N_8691,N_8853);
or U9683 (N_9683,N_8171,N_8447);
nor U9684 (N_9684,N_8917,N_8310);
or U9685 (N_9685,N_8036,N_8840);
xnor U9686 (N_9686,N_8774,N_8645);
or U9687 (N_9687,N_8342,N_8929);
or U9688 (N_9688,N_8057,N_8672);
or U9689 (N_9689,N_8488,N_8528);
xor U9690 (N_9690,N_8119,N_8681);
or U9691 (N_9691,N_8224,N_8312);
nor U9692 (N_9692,N_8920,N_8702);
and U9693 (N_9693,N_8650,N_8870);
nor U9694 (N_9694,N_8573,N_8711);
and U9695 (N_9695,N_8604,N_8707);
or U9696 (N_9696,N_8483,N_8901);
or U9697 (N_9697,N_8140,N_8114);
nand U9698 (N_9698,N_8240,N_8729);
or U9699 (N_9699,N_8355,N_8047);
nand U9700 (N_9700,N_8038,N_8982);
nor U9701 (N_9701,N_8279,N_8391);
xnor U9702 (N_9702,N_8514,N_8250);
or U9703 (N_9703,N_8376,N_8526);
or U9704 (N_9704,N_8854,N_8536);
or U9705 (N_9705,N_8505,N_8562);
and U9706 (N_9706,N_8084,N_8661);
and U9707 (N_9707,N_8991,N_8301);
nand U9708 (N_9708,N_8883,N_8453);
nor U9709 (N_9709,N_8734,N_8264);
nand U9710 (N_9710,N_8077,N_8382);
nand U9711 (N_9711,N_8905,N_8749);
nor U9712 (N_9712,N_8772,N_8988);
and U9713 (N_9713,N_8556,N_8615);
xor U9714 (N_9714,N_8869,N_8931);
nor U9715 (N_9715,N_8902,N_8494);
nor U9716 (N_9716,N_8367,N_8006);
xor U9717 (N_9717,N_8787,N_8985);
xor U9718 (N_9718,N_8614,N_8307);
or U9719 (N_9719,N_8574,N_8825);
and U9720 (N_9720,N_8159,N_8778);
nor U9721 (N_9721,N_8798,N_8029);
nand U9722 (N_9722,N_8757,N_8743);
nand U9723 (N_9723,N_8211,N_8482);
nor U9724 (N_9724,N_8627,N_8154);
xor U9725 (N_9725,N_8808,N_8844);
nor U9726 (N_9726,N_8989,N_8932);
nor U9727 (N_9727,N_8219,N_8959);
and U9728 (N_9728,N_8588,N_8832);
or U9729 (N_9729,N_8921,N_8480);
nand U9730 (N_9730,N_8894,N_8758);
nand U9731 (N_9731,N_8182,N_8426);
nand U9732 (N_9732,N_8695,N_8046);
or U9733 (N_9733,N_8679,N_8132);
or U9734 (N_9734,N_8490,N_8817);
nand U9735 (N_9735,N_8165,N_8584);
or U9736 (N_9736,N_8811,N_8331);
or U9737 (N_9737,N_8425,N_8126);
or U9738 (N_9738,N_8495,N_8652);
and U9739 (N_9739,N_8961,N_8323);
or U9740 (N_9740,N_8881,N_8940);
nor U9741 (N_9741,N_8016,N_8699);
nor U9742 (N_9742,N_8096,N_8484);
nand U9743 (N_9743,N_8127,N_8150);
nand U9744 (N_9744,N_8854,N_8671);
xor U9745 (N_9745,N_8356,N_8913);
xor U9746 (N_9746,N_8365,N_8716);
and U9747 (N_9747,N_8159,N_8548);
nor U9748 (N_9748,N_8607,N_8310);
or U9749 (N_9749,N_8717,N_8055);
and U9750 (N_9750,N_8674,N_8567);
nand U9751 (N_9751,N_8256,N_8313);
or U9752 (N_9752,N_8822,N_8220);
nor U9753 (N_9753,N_8864,N_8346);
or U9754 (N_9754,N_8453,N_8865);
and U9755 (N_9755,N_8044,N_8279);
nor U9756 (N_9756,N_8139,N_8303);
or U9757 (N_9757,N_8025,N_8689);
nor U9758 (N_9758,N_8875,N_8547);
nand U9759 (N_9759,N_8249,N_8814);
nand U9760 (N_9760,N_8099,N_8025);
nor U9761 (N_9761,N_8745,N_8608);
nor U9762 (N_9762,N_8976,N_8164);
or U9763 (N_9763,N_8514,N_8718);
xor U9764 (N_9764,N_8229,N_8030);
or U9765 (N_9765,N_8002,N_8557);
nor U9766 (N_9766,N_8309,N_8835);
xnor U9767 (N_9767,N_8088,N_8544);
and U9768 (N_9768,N_8852,N_8046);
xnor U9769 (N_9769,N_8622,N_8755);
nand U9770 (N_9770,N_8528,N_8994);
or U9771 (N_9771,N_8133,N_8892);
or U9772 (N_9772,N_8330,N_8234);
nand U9773 (N_9773,N_8750,N_8001);
or U9774 (N_9774,N_8349,N_8754);
nand U9775 (N_9775,N_8463,N_8107);
or U9776 (N_9776,N_8590,N_8159);
and U9777 (N_9777,N_8615,N_8142);
nand U9778 (N_9778,N_8380,N_8728);
xor U9779 (N_9779,N_8781,N_8848);
xor U9780 (N_9780,N_8992,N_8471);
nor U9781 (N_9781,N_8554,N_8603);
nand U9782 (N_9782,N_8575,N_8354);
nor U9783 (N_9783,N_8010,N_8562);
and U9784 (N_9784,N_8833,N_8581);
xnor U9785 (N_9785,N_8738,N_8754);
nor U9786 (N_9786,N_8437,N_8810);
nand U9787 (N_9787,N_8871,N_8472);
and U9788 (N_9788,N_8788,N_8714);
nand U9789 (N_9789,N_8792,N_8837);
and U9790 (N_9790,N_8287,N_8941);
xor U9791 (N_9791,N_8649,N_8791);
nand U9792 (N_9792,N_8383,N_8760);
xnor U9793 (N_9793,N_8573,N_8445);
nand U9794 (N_9794,N_8437,N_8766);
xnor U9795 (N_9795,N_8222,N_8527);
xnor U9796 (N_9796,N_8290,N_8963);
or U9797 (N_9797,N_8809,N_8075);
xor U9798 (N_9798,N_8236,N_8777);
nand U9799 (N_9799,N_8570,N_8386);
or U9800 (N_9800,N_8193,N_8200);
xor U9801 (N_9801,N_8250,N_8496);
xor U9802 (N_9802,N_8802,N_8628);
or U9803 (N_9803,N_8699,N_8633);
xor U9804 (N_9804,N_8618,N_8266);
nor U9805 (N_9805,N_8591,N_8455);
xor U9806 (N_9806,N_8647,N_8687);
nor U9807 (N_9807,N_8152,N_8529);
or U9808 (N_9808,N_8917,N_8182);
or U9809 (N_9809,N_8134,N_8286);
nor U9810 (N_9810,N_8973,N_8963);
and U9811 (N_9811,N_8246,N_8145);
or U9812 (N_9812,N_8026,N_8366);
nor U9813 (N_9813,N_8401,N_8743);
nand U9814 (N_9814,N_8987,N_8340);
and U9815 (N_9815,N_8080,N_8350);
xor U9816 (N_9816,N_8141,N_8102);
xor U9817 (N_9817,N_8610,N_8708);
xor U9818 (N_9818,N_8079,N_8184);
nand U9819 (N_9819,N_8863,N_8364);
xor U9820 (N_9820,N_8889,N_8632);
and U9821 (N_9821,N_8787,N_8939);
nor U9822 (N_9822,N_8481,N_8909);
and U9823 (N_9823,N_8236,N_8165);
or U9824 (N_9824,N_8024,N_8411);
nor U9825 (N_9825,N_8831,N_8453);
nand U9826 (N_9826,N_8064,N_8377);
nor U9827 (N_9827,N_8649,N_8822);
nand U9828 (N_9828,N_8782,N_8077);
and U9829 (N_9829,N_8609,N_8802);
and U9830 (N_9830,N_8314,N_8320);
and U9831 (N_9831,N_8447,N_8050);
xnor U9832 (N_9832,N_8314,N_8604);
nand U9833 (N_9833,N_8044,N_8136);
and U9834 (N_9834,N_8444,N_8277);
or U9835 (N_9835,N_8907,N_8333);
nand U9836 (N_9836,N_8989,N_8472);
and U9837 (N_9837,N_8846,N_8331);
and U9838 (N_9838,N_8743,N_8908);
nor U9839 (N_9839,N_8946,N_8935);
xor U9840 (N_9840,N_8740,N_8191);
xnor U9841 (N_9841,N_8674,N_8314);
xnor U9842 (N_9842,N_8131,N_8547);
xnor U9843 (N_9843,N_8220,N_8131);
nor U9844 (N_9844,N_8723,N_8633);
and U9845 (N_9845,N_8118,N_8742);
and U9846 (N_9846,N_8273,N_8506);
and U9847 (N_9847,N_8467,N_8061);
or U9848 (N_9848,N_8010,N_8026);
nor U9849 (N_9849,N_8203,N_8152);
nand U9850 (N_9850,N_8079,N_8472);
and U9851 (N_9851,N_8421,N_8247);
xnor U9852 (N_9852,N_8854,N_8142);
or U9853 (N_9853,N_8461,N_8223);
nor U9854 (N_9854,N_8655,N_8651);
nor U9855 (N_9855,N_8311,N_8390);
nor U9856 (N_9856,N_8694,N_8877);
nor U9857 (N_9857,N_8956,N_8900);
xnor U9858 (N_9858,N_8787,N_8916);
xnor U9859 (N_9859,N_8059,N_8499);
nor U9860 (N_9860,N_8872,N_8279);
nor U9861 (N_9861,N_8987,N_8196);
nand U9862 (N_9862,N_8024,N_8135);
xor U9863 (N_9863,N_8570,N_8872);
and U9864 (N_9864,N_8092,N_8403);
and U9865 (N_9865,N_8058,N_8004);
nor U9866 (N_9866,N_8643,N_8615);
and U9867 (N_9867,N_8530,N_8234);
or U9868 (N_9868,N_8458,N_8173);
xnor U9869 (N_9869,N_8841,N_8258);
and U9870 (N_9870,N_8565,N_8837);
nor U9871 (N_9871,N_8018,N_8308);
nor U9872 (N_9872,N_8623,N_8197);
nand U9873 (N_9873,N_8389,N_8104);
nand U9874 (N_9874,N_8826,N_8194);
or U9875 (N_9875,N_8575,N_8807);
or U9876 (N_9876,N_8073,N_8466);
or U9877 (N_9877,N_8360,N_8000);
nor U9878 (N_9878,N_8670,N_8658);
nand U9879 (N_9879,N_8038,N_8013);
or U9880 (N_9880,N_8794,N_8926);
nor U9881 (N_9881,N_8689,N_8939);
and U9882 (N_9882,N_8155,N_8951);
and U9883 (N_9883,N_8492,N_8405);
xnor U9884 (N_9884,N_8675,N_8299);
nand U9885 (N_9885,N_8089,N_8772);
nor U9886 (N_9886,N_8284,N_8246);
nand U9887 (N_9887,N_8306,N_8426);
nor U9888 (N_9888,N_8159,N_8410);
or U9889 (N_9889,N_8075,N_8335);
nand U9890 (N_9890,N_8811,N_8212);
xnor U9891 (N_9891,N_8195,N_8841);
nor U9892 (N_9892,N_8553,N_8289);
xnor U9893 (N_9893,N_8514,N_8698);
nor U9894 (N_9894,N_8194,N_8424);
nor U9895 (N_9895,N_8319,N_8765);
xnor U9896 (N_9896,N_8123,N_8296);
and U9897 (N_9897,N_8460,N_8081);
xnor U9898 (N_9898,N_8975,N_8132);
nor U9899 (N_9899,N_8189,N_8241);
xnor U9900 (N_9900,N_8850,N_8985);
nand U9901 (N_9901,N_8317,N_8777);
and U9902 (N_9902,N_8960,N_8615);
xnor U9903 (N_9903,N_8908,N_8619);
xor U9904 (N_9904,N_8624,N_8825);
or U9905 (N_9905,N_8325,N_8005);
or U9906 (N_9906,N_8035,N_8079);
and U9907 (N_9907,N_8736,N_8345);
xnor U9908 (N_9908,N_8569,N_8868);
nor U9909 (N_9909,N_8053,N_8288);
and U9910 (N_9910,N_8504,N_8284);
xnor U9911 (N_9911,N_8074,N_8916);
or U9912 (N_9912,N_8315,N_8138);
xnor U9913 (N_9913,N_8484,N_8853);
nor U9914 (N_9914,N_8864,N_8306);
or U9915 (N_9915,N_8157,N_8414);
nor U9916 (N_9916,N_8492,N_8789);
nand U9917 (N_9917,N_8469,N_8658);
and U9918 (N_9918,N_8914,N_8923);
and U9919 (N_9919,N_8269,N_8278);
and U9920 (N_9920,N_8813,N_8347);
xnor U9921 (N_9921,N_8048,N_8114);
nand U9922 (N_9922,N_8474,N_8381);
nand U9923 (N_9923,N_8474,N_8361);
or U9924 (N_9924,N_8327,N_8788);
nor U9925 (N_9925,N_8672,N_8323);
nand U9926 (N_9926,N_8072,N_8391);
nor U9927 (N_9927,N_8510,N_8631);
nand U9928 (N_9928,N_8083,N_8370);
and U9929 (N_9929,N_8463,N_8603);
nor U9930 (N_9930,N_8792,N_8530);
and U9931 (N_9931,N_8888,N_8996);
nand U9932 (N_9932,N_8626,N_8903);
nor U9933 (N_9933,N_8909,N_8013);
nor U9934 (N_9934,N_8906,N_8154);
xor U9935 (N_9935,N_8454,N_8425);
or U9936 (N_9936,N_8689,N_8621);
or U9937 (N_9937,N_8248,N_8073);
or U9938 (N_9938,N_8619,N_8131);
nand U9939 (N_9939,N_8545,N_8123);
and U9940 (N_9940,N_8937,N_8602);
xor U9941 (N_9941,N_8881,N_8929);
nand U9942 (N_9942,N_8020,N_8884);
nand U9943 (N_9943,N_8225,N_8093);
or U9944 (N_9944,N_8302,N_8311);
nand U9945 (N_9945,N_8383,N_8268);
and U9946 (N_9946,N_8608,N_8945);
nor U9947 (N_9947,N_8886,N_8748);
nand U9948 (N_9948,N_8393,N_8901);
nand U9949 (N_9949,N_8943,N_8327);
nand U9950 (N_9950,N_8679,N_8520);
xor U9951 (N_9951,N_8896,N_8206);
xnor U9952 (N_9952,N_8380,N_8354);
xnor U9953 (N_9953,N_8381,N_8690);
nor U9954 (N_9954,N_8161,N_8404);
nor U9955 (N_9955,N_8115,N_8763);
and U9956 (N_9956,N_8137,N_8405);
nand U9957 (N_9957,N_8643,N_8671);
xor U9958 (N_9958,N_8896,N_8080);
xnor U9959 (N_9959,N_8126,N_8348);
and U9960 (N_9960,N_8298,N_8408);
nand U9961 (N_9961,N_8327,N_8507);
and U9962 (N_9962,N_8187,N_8668);
and U9963 (N_9963,N_8778,N_8698);
nor U9964 (N_9964,N_8806,N_8787);
and U9965 (N_9965,N_8202,N_8999);
nand U9966 (N_9966,N_8535,N_8974);
nor U9967 (N_9967,N_8851,N_8693);
xor U9968 (N_9968,N_8655,N_8349);
nand U9969 (N_9969,N_8440,N_8504);
nand U9970 (N_9970,N_8364,N_8981);
nand U9971 (N_9971,N_8282,N_8976);
nand U9972 (N_9972,N_8784,N_8583);
nand U9973 (N_9973,N_8167,N_8138);
nor U9974 (N_9974,N_8707,N_8692);
xor U9975 (N_9975,N_8275,N_8884);
nor U9976 (N_9976,N_8665,N_8733);
xor U9977 (N_9977,N_8852,N_8367);
and U9978 (N_9978,N_8794,N_8976);
or U9979 (N_9979,N_8493,N_8991);
and U9980 (N_9980,N_8734,N_8496);
nand U9981 (N_9981,N_8884,N_8957);
and U9982 (N_9982,N_8611,N_8154);
and U9983 (N_9983,N_8819,N_8488);
nor U9984 (N_9984,N_8126,N_8198);
or U9985 (N_9985,N_8615,N_8565);
nor U9986 (N_9986,N_8189,N_8663);
nand U9987 (N_9987,N_8428,N_8985);
and U9988 (N_9988,N_8296,N_8116);
and U9989 (N_9989,N_8694,N_8078);
xnor U9990 (N_9990,N_8365,N_8005);
or U9991 (N_9991,N_8558,N_8038);
or U9992 (N_9992,N_8899,N_8005);
and U9993 (N_9993,N_8273,N_8641);
and U9994 (N_9994,N_8338,N_8441);
nand U9995 (N_9995,N_8980,N_8761);
and U9996 (N_9996,N_8343,N_8581);
xor U9997 (N_9997,N_8244,N_8599);
or U9998 (N_9998,N_8568,N_8189);
nand U9999 (N_9999,N_8167,N_8652);
nand U10000 (N_10000,N_9820,N_9937);
or U10001 (N_10001,N_9255,N_9051);
and U10002 (N_10002,N_9782,N_9398);
xor U10003 (N_10003,N_9703,N_9196);
nand U10004 (N_10004,N_9321,N_9179);
nand U10005 (N_10005,N_9263,N_9917);
or U10006 (N_10006,N_9974,N_9380);
or U10007 (N_10007,N_9879,N_9293);
and U10008 (N_10008,N_9150,N_9816);
nand U10009 (N_10009,N_9992,N_9824);
and U10010 (N_10010,N_9864,N_9546);
or U10011 (N_10011,N_9172,N_9658);
and U10012 (N_10012,N_9356,N_9166);
or U10013 (N_10013,N_9482,N_9827);
and U10014 (N_10014,N_9547,N_9696);
xor U10015 (N_10015,N_9279,N_9590);
or U10016 (N_10016,N_9564,N_9780);
nand U10017 (N_10017,N_9979,N_9897);
and U10018 (N_10018,N_9021,N_9553);
nand U10019 (N_10019,N_9659,N_9605);
or U10020 (N_10020,N_9272,N_9234);
nand U10021 (N_10021,N_9754,N_9834);
nand U10022 (N_10022,N_9884,N_9268);
xnor U10023 (N_10023,N_9448,N_9539);
xor U10024 (N_10024,N_9359,N_9372);
nand U10025 (N_10025,N_9521,N_9743);
nand U10026 (N_10026,N_9000,N_9475);
nor U10027 (N_10027,N_9235,N_9069);
nand U10028 (N_10028,N_9830,N_9241);
xor U10029 (N_10029,N_9560,N_9276);
or U10030 (N_10030,N_9669,N_9868);
xor U10031 (N_10031,N_9946,N_9443);
nor U10032 (N_10032,N_9706,N_9412);
or U10033 (N_10033,N_9516,N_9694);
or U10034 (N_10034,N_9245,N_9665);
and U10035 (N_10035,N_9154,N_9500);
or U10036 (N_10036,N_9143,N_9883);
nand U10037 (N_10037,N_9990,N_9677);
nand U10038 (N_10038,N_9987,N_9405);
nand U10039 (N_10039,N_9668,N_9673);
nand U10040 (N_10040,N_9977,N_9774);
or U10041 (N_10041,N_9488,N_9297);
nor U10042 (N_10042,N_9716,N_9116);
or U10043 (N_10043,N_9442,N_9700);
or U10044 (N_10044,N_9383,N_9175);
xnor U10045 (N_10045,N_9007,N_9544);
nand U10046 (N_10046,N_9271,N_9647);
nand U10047 (N_10047,N_9910,N_9818);
or U10048 (N_10048,N_9013,N_9455);
xor U10049 (N_10049,N_9115,N_9353);
xor U10050 (N_10050,N_9771,N_9996);
xnor U10051 (N_10051,N_9550,N_9760);
nand U10052 (N_10052,N_9980,N_9066);
or U10053 (N_10053,N_9316,N_9123);
or U10054 (N_10054,N_9233,N_9173);
nand U10055 (N_10055,N_9082,N_9178);
nor U10056 (N_10056,N_9765,N_9104);
or U10057 (N_10057,N_9653,N_9100);
xnor U10058 (N_10058,N_9549,N_9973);
and U10059 (N_10059,N_9872,N_9718);
and U10060 (N_10060,N_9918,N_9674);
nor U10061 (N_10061,N_9477,N_9167);
and U10062 (N_10062,N_9313,N_9367);
or U10063 (N_10063,N_9296,N_9587);
nand U10064 (N_10064,N_9707,N_9413);
or U10065 (N_10065,N_9147,N_9481);
nor U10066 (N_10066,N_9217,N_9062);
and U10067 (N_10067,N_9869,N_9772);
xnor U10068 (N_10068,N_9457,N_9230);
or U10069 (N_10069,N_9586,N_9859);
xnor U10070 (N_10070,N_9926,N_9400);
nor U10071 (N_10071,N_9833,N_9124);
nor U10072 (N_10072,N_9001,N_9844);
nand U10073 (N_10073,N_9324,N_9369);
nor U10074 (N_10074,N_9008,N_9803);
nand U10075 (N_10075,N_9155,N_9393);
nor U10076 (N_10076,N_9307,N_9038);
nand U10077 (N_10077,N_9458,N_9152);
nor U10078 (N_10078,N_9610,N_9159);
nand U10079 (N_10079,N_9030,N_9894);
xor U10080 (N_10080,N_9387,N_9170);
and U10081 (N_10081,N_9959,N_9683);
nand U10082 (N_10082,N_9936,N_9073);
xnor U10083 (N_10083,N_9893,N_9479);
nand U10084 (N_10084,N_9168,N_9319);
xor U10085 (N_10085,N_9414,N_9518);
nor U10086 (N_10086,N_9609,N_9841);
or U10087 (N_10087,N_9135,N_9314);
xor U10088 (N_10088,N_9212,N_9040);
xor U10089 (N_10089,N_9326,N_9078);
nor U10090 (N_10090,N_9111,N_9335);
nand U10091 (N_10091,N_9639,N_9410);
xor U10092 (N_10092,N_9077,N_9449);
xor U10093 (N_10093,N_9709,N_9507);
nor U10094 (N_10094,N_9595,N_9511);
and U10095 (N_10095,N_9289,N_9689);
and U10096 (N_10096,N_9381,N_9676);
and U10097 (N_10097,N_9645,N_9688);
or U10098 (N_10098,N_9982,N_9469);
xnor U10099 (N_10099,N_9731,N_9724);
or U10100 (N_10100,N_9885,N_9248);
or U10101 (N_10101,N_9403,N_9250);
nor U10102 (N_10102,N_9720,N_9513);
or U10103 (N_10103,N_9345,N_9064);
nor U10104 (N_10104,N_9127,N_9912);
and U10105 (N_10105,N_9985,N_9664);
xnor U10106 (N_10106,N_9984,N_9796);
and U10107 (N_10107,N_9598,N_9280);
or U10108 (N_10108,N_9141,N_9619);
and U10109 (N_10109,N_9913,N_9877);
xor U10110 (N_10110,N_9404,N_9563);
or U10111 (N_10111,N_9231,N_9121);
nand U10112 (N_10112,N_9532,N_9890);
nor U10113 (N_10113,N_9192,N_9228);
or U10114 (N_10114,N_9092,N_9510);
nor U10115 (N_10115,N_9744,N_9191);
nand U10116 (N_10116,N_9083,N_9714);
or U10117 (N_10117,N_9886,N_9266);
or U10118 (N_10118,N_9095,N_9540);
xor U10119 (N_10119,N_9294,N_9878);
nand U10120 (N_10120,N_9226,N_9079);
and U10121 (N_10121,N_9934,N_9764);
nand U10122 (N_10122,N_9584,N_9370);
nor U10123 (N_10123,N_9466,N_9363);
nand U10124 (N_10124,N_9227,N_9061);
and U10125 (N_10125,N_9811,N_9680);
nor U10126 (N_10126,N_9631,N_9867);
nand U10127 (N_10127,N_9474,N_9470);
or U10128 (N_10128,N_9330,N_9993);
nand U10129 (N_10129,N_9395,N_9144);
nor U10130 (N_10130,N_9295,N_9685);
and U10131 (N_10131,N_9735,N_9063);
xnor U10132 (N_10132,N_9920,N_9118);
nand U10133 (N_10133,N_9053,N_9134);
and U10134 (N_10134,N_9012,N_9922);
xor U10135 (N_10135,N_9569,N_9312);
or U10136 (N_10136,N_9298,N_9802);
and U10137 (N_10137,N_9804,N_9348);
nand U10138 (N_10138,N_9574,N_9267);
or U10139 (N_10139,N_9556,N_9328);
nor U10140 (N_10140,N_9637,N_9751);
or U10141 (N_10141,N_9286,N_9882);
nand U10142 (N_10142,N_9528,N_9336);
nor U10143 (N_10143,N_9965,N_9672);
and U10144 (N_10144,N_9374,N_9603);
or U10145 (N_10145,N_9219,N_9725);
and U10146 (N_10146,N_9512,N_9264);
xor U10147 (N_10147,N_9761,N_9309);
nor U10148 (N_10148,N_9997,N_9671);
xnor U10149 (N_10149,N_9087,N_9925);
nand U10150 (N_10150,N_9394,N_9342);
or U10151 (N_10151,N_9737,N_9025);
nand U10152 (N_10152,N_9060,N_9478);
nand U10153 (N_10153,N_9364,N_9107);
or U10154 (N_10154,N_9251,N_9853);
and U10155 (N_10155,N_9052,N_9006);
nand U10156 (N_10156,N_9432,N_9355);
nand U10157 (N_10157,N_9072,N_9242);
and U10158 (N_10158,N_9678,N_9325);
or U10159 (N_10159,N_9148,N_9520);
and U10160 (N_10160,N_9341,N_9583);
nand U10161 (N_10161,N_9682,N_9738);
xor U10162 (N_10162,N_9209,N_9205);
nand U10163 (N_10163,N_9055,N_9654);
and U10164 (N_10164,N_9514,N_9919);
xnor U10165 (N_10165,N_9005,N_9480);
xor U10166 (N_10166,N_9721,N_9182);
xnor U10167 (N_10167,N_9331,N_9870);
and U10168 (N_10168,N_9822,N_9852);
xor U10169 (N_10169,N_9746,N_9165);
xnor U10170 (N_10170,N_9787,N_9835);
nor U10171 (N_10171,N_9282,N_9401);
nor U10172 (N_10172,N_9952,N_9004);
and U10173 (N_10173,N_9770,N_9315);
or U10174 (N_10174,N_9068,N_9438);
nor U10175 (N_10175,N_9975,N_9281);
and U10176 (N_10176,N_9648,N_9211);
and U10177 (N_10177,N_9120,N_9184);
and U10178 (N_10178,N_9472,N_9164);
nor U10179 (N_10179,N_9875,N_9183);
and U10180 (N_10180,N_9909,N_9789);
or U10181 (N_10181,N_9577,N_9995);
xnor U10182 (N_10182,N_9200,N_9807);
nand U10183 (N_10183,N_9416,N_9881);
xor U10184 (N_10184,N_9146,N_9629);
nand U10185 (N_10185,N_9218,N_9453);
nor U10186 (N_10186,N_9785,N_9049);
nor U10187 (N_10187,N_9615,N_9594);
xor U10188 (N_10188,N_9138,N_9388);
nand U10189 (N_10189,N_9708,N_9578);
and U10190 (N_10190,N_9915,N_9174);
and U10191 (N_10191,N_9427,N_9950);
and U10192 (N_10192,N_9880,N_9652);
xnor U10193 (N_10193,N_9098,N_9794);
xnor U10194 (N_10194,N_9758,N_9541);
and U10195 (N_10195,N_9766,N_9411);
xnor U10196 (N_10196,N_9848,N_9932);
and U10197 (N_10197,N_9199,N_9283);
nand U10198 (N_10198,N_9260,N_9391);
xor U10199 (N_10199,N_9656,N_9810);
and U10200 (N_10200,N_9895,N_9084);
xnor U10201 (N_10201,N_9767,N_9221);
xor U10202 (N_10202,N_9128,N_9452);
and U10203 (N_10203,N_9132,N_9686);
xnor U10204 (N_10204,N_9499,N_9651);
and U10205 (N_10205,N_9091,N_9225);
xnor U10206 (N_10206,N_9429,N_9437);
or U10207 (N_10207,N_9028,N_9329);
nand U10208 (N_10208,N_9779,N_9642);
and U10209 (N_10209,N_9561,N_9426);
or U10210 (N_10210,N_9559,N_9597);
or U10211 (N_10211,N_9430,N_9311);
nor U10212 (N_10212,N_9037,N_9406);
and U10213 (N_10213,N_9889,N_9842);
nand U10214 (N_10214,N_9460,N_9243);
xnor U10215 (N_10215,N_9534,N_9846);
nand U10216 (N_10216,N_9015,N_9396);
and U10217 (N_10217,N_9828,N_9237);
or U10218 (N_10218,N_9142,N_9018);
nor U10219 (N_10219,N_9424,N_9206);
or U10220 (N_10220,N_9663,N_9467);
nand U10221 (N_10221,N_9357,N_9567);
or U10222 (N_10222,N_9445,N_9954);
and U10223 (N_10223,N_9566,N_9930);
or U10224 (N_10224,N_9014,N_9814);
and U10225 (N_10225,N_9726,N_9961);
or U10226 (N_10226,N_9836,N_9745);
or U10227 (N_10227,N_9131,N_9288);
nor U10228 (N_10228,N_9041,N_9047);
or U10229 (N_10229,N_9600,N_9957);
nor U10230 (N_10230,N_9854,N_9527);
or U10231 (N_10231,N_9058,N_9797);
and U10232 (N_10232,N_9627,N_9386);
nand U10233 (N_10233,N_9552,N_9284);
xnor U10234 (N_10234,N_9808,N_9964);
nand U10235 (N_10235,N_9033,N_9160);
or U10236 (N_10236,N_9011,N_9991);
nor U10237 (N_10237,N_9186,N_9622);
xor U10238 (N_10238,N_9130,N_9777);
or U10239 (N_10239,N_9291,N_9972);
xor U10240 (N_10240,N_9633,N_9273);
and U10241 (N_10241,N_9300,N_9695);
and U10242 (N_10242,N_9575,N_9752);
xor U10243 (N_10243,N_9749,N_9606);
nor U10244 (N_10244,N_9939,N_9464);
nand U10245 (N_10245,N_9838,N_9621);
nand U10246 (N_10246,N_9795,N_9801);
xnor U10247 (N_10247,N_9187,N_9046);
nor U10248 (N_10248,N_9888,N_9692);
or U10249 (N_10249,N_9819,N_9044);
or U10250 (N_10250,N_9378,N_9582);
and U10251 (N_10251,N_9215,N_9999);
nor U10252 (N_10252,N_9953,N_9277);
xor U10253 (N_10253,N_9149,N_9863);
or U10254 (N_10254,N_9866,N_9502);
or U10255 (N_10255,N_9258,N_9732);
or U10256 (N_10256,N_9232,N_9998);
nor U10257 (N_10257,N_9275,N_9246);
and U10258 (N_10258,N_9602,N_9496);
xor U10259 (N_10259,N_9632,N_9914);
nand U10260 (N_10260,N_9439,N_9831);
or U10261 (N_10261,N_9604,N_9776);
xnor U10262 (N_10262,N_9843,N_9809);
xor U10263 (N_10263,N_9176,N_9076);
or U10264 (N_10264,N_9322,N_9377);
xor U10265 (N_10265,N_9849,N_9945);
or U10266 (N_10266,N_9274,N_9417);
xor U10267 (N_10267,N_9431,N_9778);
nor U10268 (N_10268,N_9323,N_9265);
or U10269 (N_10269,N_9655,N_9628);
and U10270 (N_10270,N_9624,N_9533);
nor U10271 (N_10271,N_9887,N_9213);
nand U10272 (N_10272,N_9646,N_9487);
nor U10273 (N_10273,N_9662,N_9490);
xor U10274 (N_10274,N_9962,N_9379);
or U10275 (N_10275,N_9963,N_9723);
nor U10276 (N_10276,N_9856,N_9185);
nor U10277 (N_10277,N_9468,N_9224);
nor U10278 (N_10278,N_9074,N_9045);
and U10279 (N_10279,N_9090,N_9202);
or U10280 (N_10280,N_9681,N_9821);
and U10281 (N_10281,N_9420,N_9898);
nand U10282 (N_10282,N_9407,N_9489);
nand U10283 (N_10283,N_9684,N_9317);
and U10284 (N_10284,N_9944,N_9740);
or U10285 (N_10285,N_9085,N_9981);
xnor U10286 (N_10286,N_9545,N_9823);
xnor U10287 (N_10287,N_9641,N_9017);
nor U10288 (N_10288,N_9722,N_9382);
nor U10289 (N_10289,N_9059,N_9812);
and U10290 (N_10290,N_9554,N_9327);
xor U10291 (N_10291,N_9793,N_9376);
nor U10292 (N_10292,N_9599,N_9375);
or U10293 (N_10293,N_9781,N_9526);
nand U10294 (N_10294,N_9970,N_9441);
and U10295 (N_10295,N_9825,N_9911);
nand U10296 (N_10296,N_9171,N_9362);
or U10297 (N_10297,N_9713,N_9204);
and U10298 (N_10298,N_9110,N_9948);
xor U10299 (N_10299,N_9504,N_9903);
nor U10300 (N_10300,N_9601,N_9446);
xnor U10301 (N_10301,N_9422,N_9967);
or U10302 (N_10302,N_9784,N_9596);
or U10303 (N_10303,N_9103,N_9702);
nand U10304 (N_10304,N_9542,N_9197);
or U10305 (N_10305,N_9042,N_9303);
nor U10306 (N_10306,N_9334,N_9093);
nor U10307 (N_10307,N_9070,N_9137);
nor U10308 (N_10308,N_9613,N_9711);
nor U10309 (N_10309,N_9902,N_9865);
nor U10310 (N_10310,N_9239,N_9969);
xnor U10311 (N_10311,N_9366,N_9207);
nand U10312 (N_10312,N_9285,N_9717);
xor U10313 (N_10313,N_9792,N_9493);
xor U10314 (N_10314,N_9026,N_9290);
and U10315 (N_10315,N_9530,N_9238);
nor U10316 (N_10316,N_9687,N_9071);
nand U10317 (N_10317,N_9896,N_9436);
nor U10318 (N_10318,N_9690,N_9454);
nand U10319 (N_10319,N_9608,N_9741);
nor U10320 (N_10320,N_9180,N_9989);
nand U10321 (N_10321,N_9832,N_9057);
nand U10322 (N_10322,N_9096,N_9636);
or U10323 (N_10323,N_9065,N_9145);
xor U10324 (N_10324,N_9626,N_9177);
xnor U10325 (N_10325,N_9257,N_9506);
nor U10326 (N_10326,N_9693,N_9976);
nor U10327 (N_10327,N_9941,N_9113);
and U10328 (N_10328,N_9790,N_9572);
nand U10329 (N_10329,N_9840,N_9860);
xor U10330 (N_10330,N_9661,N_9960);
or U10331 (N_10331,N_9409,N_9891);
and U10332 (N_10332,N_9094,N_9733);
or U10333 (N_10333,N_9050,N_9508);
and U10334 (N_10334,N_9739,N_9390);
or U10335 (N_10335,N_9346,N_9032);
or U10336 (N_10336,N_9906,N_9108);
nand U10337 (N_10337,N_9947,N_9350);
nand U10338 (N_10338,N_9397,N_9483);
nand U10339 (N_10339,N_9201,N_9529);
nand U10340 (N_10340,N_9140,N_9451);
nand U10341 (N_10341,N_9270,N_9473);
and U10342 (N_10342,N_9054,N_9750);
nor U10343 (N_10343,N_9551,N_9861);
and U10344 (N_10344,N_9759,N_9340);
nand U10345 (N_10345,N_9592,N_9791);
xor U10346 (N_10346,N_9901,N_9900);
nor U10347 (N_10347,N_9162,N_9189);
nor U10348 (N_10348,N_9244,N_9612);
and U10349 (N_10349,N_9428,N_9119);
xnor U10350 (N_10350,N_9826,N_9299);
nand U10351 (N_10351,N_9009,N_9921);
nor U10352 (N_10352,N_9576,N_9773);
nor U10353 (N_10353,N_9614,N_9531);
xor U10354 (N_10354,N_9924,N_9099);
nand U10355 (N_10355,N_9871,N_9851);
and U10356 (N_10356,N_9434,N_9978);
or U10357 (N_10357,N_9968,N_9450);
and U10358 (N_10358,N_9568,N_9643);
and U10359 (N_10359,N_9798,N_9638);
nand U10360 (N_10360,N_9650,N_9847);
or U10361 (N_10361,N_9736,N_9813);
or U10362 (N_10362,N_9261,N_9193);
or U10363 (N_10363,N_9585,N_9928);
nand U10364 (N_10364,N_9892,N_9730);
nand U10365 (N_10365,N_9368,N_9617);
nor U10366 (N_10366,N_9611,N_9016);
nand U10367 (N_10367,N_9435,N_9169);
or U10368 (N_10368,N_9555,N_9710);
or U10369 (N_10369,N_9517,N_9343);
or U10370 (N_10370,N_9635,N_9701);
nand U10371 (N_10371,N_9019,N_9940);
nand U10372 (N_10372,N_9259,N_9775);
and U10373 (N_10373,N_9670,N_9347);
nand U10374 (N_10374,N_9523,N_9181);
nand U10375 (N_10375,N_9763,N_9579);
and U10376 (N_10376,N_9788,N_9558);
xor U10377 (N_10377,N_9462,N_9535);
xor U10378 (N_10378,N_9986,N_9679);
xnor U10379 (N_10379,N_9337,N_9106);
nand U10380 (N_10380,N_9931,N_9373);
nand U10381 (N_10381,N_9086,N_9850);
xnor U10382 (N_10382,N_9365,N_9262);
nor U10383 (N_10383,N_9188,N_9543);
xor U10384 (N_10384,N_9122,N_9565);
and U10385 (N_10385,N_9497,N_9158);
nand U10386 (N_10386,N_9208,N_9837);
nor U10387 (N_10387,N_9591,N_9461);
xnor U10388 (N_10388,N_9002,N_9151);
xor U10389 (N_10389,N_9229,N_9862);
nand U10390 (N_10390,N_9198,N_9515);
or U10391 (N_10391,N_9857,N_9415);
or U10392 (N_10392,N_9216,N_9908);
nand U10393 (N_10393,N_9024,N_9287);
nor U10394 (N_10394,N_9519,N_9756);
xnor U10395 (N_10395,N_9117,N_9942);
xnor U10396 (N_10396,N_9332,N_9027);
nor U10397 (N_10397,N_9114,N_9899);
nor U10398 (N_10398,N_9537,N_9503);
or U10399 (N_10399,N_9109,N_9361);
xor U10400 (N_10400,N_9035,N_9101);
and U10401 (N_10401,N_9573,N_9247);
nor U10402 (N_10402,N_9938,N_9222);
nand U10403 (N_10403,N_9753,N_9742);
and U10404 (N_10404,N_9492,N_9988);
or U10405 (N_10405,N_9634,N_9660);
xor U10406 (N_10406,N_9133,N_9728);
nor U10407 (N_10407,N_9252,N_9494);
xnor U10408 (N_10408,N_9081,N_9536);
and U10409 (N_10409,N_9194,N_9349);
xor U10410 (N_10410,N_9163,N_9214);
nor U10411 (N_10411,N_9943,N_9715);
nor U10412 (N_10412,N_9402,N_9010);
nor U10413 (N_10413,N_9338,N_9697);
nand U10414 (N_10414,N_9210,N_9333);
and U10415 (N_10415,N_9190,N_9022);
nand U10416 (N_10416,N_9593,N_9589);
or U10417 (N_10417,N_9029,N_9719);
nor U10418 (N_10418,N_9310,N_9048);
or U10419 (N_10419,N_9418,N_9799);
nand U10420 (N_10420,N_9949,N_9392);
nor U10421 (N_10421,N_9956,N_9983);
nor U10422 (N_10422,N_9419,N_9306);
or U10423 (N_10423,N_9916,N_9304);
xnor U10424 (N_10424,N_9845,N_9471);
nor U10425 (N_10425,N_9408,N_9548);
or U10426 (N_10426,N_9075,N_9620);
nor U10427 (N_10427,N_9240,N_9501);
nand U10428 (N_10428,N_9783,N_9236);
xor U10429 (N_10429,N_9389,N_9385);
nor U10430 (N_10430,N_9023,N_9089);
xnor U10431 (N_10431,N_9935,N_9675);
nor U10432 (N_10432,N_9195,N_9031);
xnor U10433 (N_10433,N_9136,N_9423);
nor U10434 (N_10434,N_9256,N_9640);
nand U10435 (N_10435,N_9344,N_9153);
or U10436 (N_10436,N_9768,N_9769);
nor U10437 (N_10437,N_9302,N_9657);
nor U10438 (N_10438,N_9581,N_9786);
or U10439 (N_10439,N_9360,N_9320);
and U10440 (N_10440,N_9484,N_9156);
nand U10441 (N_10441,N_9904,N_9649);
xor U10442 (N_10442,N_9126,N_9249);
or U10443 (N_10443,N_9139,N_9440);
xnor U10444 (N_10444,N_9056,N_9923);
xor U10445 (N_10445,N_9097,N_9459);
nor U10446 (N_10446,N_9399,N_9704);
and U10447 (N_10447,N_9444,N_9994);
nand U10448 (N_10448,N_9699,N_9278);
or U10449 (N_10449,N_9384,N_9088);
nor U10450 (N_10450,N_9485,N_9223);
nor U10451 (N_10451,N_9371,N_9644);
xnor U10452 (N_10452,N_9817,N_9958);
nand U10453 (N_10453,N_9666,N_9498);
xnor U10454 (N_10454,N_9829,N_9043);
nor U10455 (N_10455,N_9505,N_9800);
nor U10456 (N_10456,N_9815,N_9003);
nor U10457 (N_10457,N_9020,N_9757);
or U10458 (N_10458,N_9112,N_9433);
nand U10459 (N_10459,N_9705,N_9491);
nand U10460 (N_10460,N_9351,N_9301);
or U10461 (N_10461,N_9447,N_9855);
and U10462 (N_10462,N_9630,N_9269);
or U10463 (N_10463,N_9562,N_9618);
xor U10464 (N_10464,N_9524,N_9623);
nand U10465 (N_10465,N_9951,N_9352);
xor U10466 (N_10466,N_9067,N_9318);
nor U10467 (N_10467,N_9125,N_9425);
or U10468 (N_10468,N_9625,N_9580);
nand U10469 (N_10469,N_9305,N_9933);
nand U10470 (N_10470,N_9927,N_9698);
xnor U10471 (N_10471,N_9806,N_9308);
xor U10472 (N_10472,N_9161,N_9929);
nor U10473 (N_10473,N_9858,N_9762);
and U10474 (N_10474,N_9495,N_9557);
nor U10475 (N_10475,N_9876,N_9570);
xor U10476 (N_10476,N_9748,N_9955);
or U10477 (N_10477,N_9456,N_9421);
nand U10478 (N_10478,N_9966,N_9476);
or U10479 (N_10479,N_9691,N_9102);
or U10480 (N_10480,N_9253,N_9729);
or U10481 (N_10481,N_9727,N_9616);
xnor U10482 (N_10482,N_9873,N_9034);
or U10483 (N_10483,N_9712,N_9667);
nand U10484 (N_10484,N_9571,N_9220);
and U10485 (N_10485,N_9538,N_9805);
xor U10486 (N_10486,N_9465,N_9254);
and U10487 (N_10487,N_9522,N_9509);
and U10488 (N_10488,N_9354,N_9339);
or U10489 (N_10489,N_9129,N_9203);
or U10490 (N_10490,N_9080,N_9358);
nand U10491 (N_10491,N_9905,N_9525);
nand U10492 (N_10492,N_9907,N_9971);
and U10493 (N_10493,N_9747,N_9486);
or U10494 (N_10494,N_9039,N_9463);
nor U10495 (N_10495,N_9292,N_9588);
nor U10496 (N_10496,N_9607,N_9839);
nor U10497 (N_10497,N_9036,N_9755);
nand U10498 (N_10498,N_9105,N_9157);
xnor U10499 (N_10499,N_9734,N_9874);
xor U10500 (N_10500,N_9425,N_9953);
nand U10501 (N_10501,N_9514,N_9048);
nor U10502 (N_10502,N_9850,N_9782);
and U10503 (N_10503,N_9805,N_9822);
nand U10504 (N_10504,N_9781,N_9776);
nand U10505 (N_10505,N_9732,N_9255);
xor U10506 (N_10506,N_9169,N_9295);
xnor U10507 (N_10507,N_9387,N_9872);
and U10508 (N_10508,N_9445,N_9210);
nand U10509 (N_10509,N_9669,N_9780);
xnor U10510 (N_10510,N_9621,N_9366);
nor U10511 (N_10511,N_9127,N_9313);
or U10512 (N_10512,N_9152,N_9202);
nor U10513 (N_10513,N_9903,N_9121);
xnor U10514 (N_10514,N_9676,N_9876);
xor U10515 (N_10515,N_9628,N_9565);
nor U10516 (N_10516,N_9248,N_9235);
and U10517 (N_10517,N_9171,N_9126);
nand U10518 (N_10518,N_9646,N_9353);
or U10519 (N_10519,N_9591,N_9899);
and U10520 (N_10520,N_9389,N_9295);
or U10521 (N_10521,N_9765,N_9519);
or U10522 (N_10522,N_9885,N_9804);
xnor U10523 (N_10523,N_9336,N_9778);
nor U10524 (N_10524,N_9679,N_9901);
nand U10525 (N_10525,N_9460,N_9219);
and U10526 (N_10526,N_9785,N_9042);
xnor U10527 (N_10527,N_9738,N_9164);
xor U10528 (N_10528,N_9128,N_9378);
or U10529 (N_10529,N_9866,N_9686);
and U10530 (N_10530,N_9071,N_9001);
nor U10531 (N_10531,N_9691,N_9239);
nand U10532 (N_10532,N_9068,N_9923);
xnor U10533 (N_10533,N_9268,N_9052);
nand U10534 (N_10534,N_9165,N_9645);
and U10535 (N_10535,N_9362,N_9262);
xnor U10536 (N_10536,N_9366,N_9179);
nor U10537 (N_10537,N_9908,N_9992);
nand U10538 (N_10538,N_9634,N_9627);
nor U10539 (N_10539,N_9298,N_9541);
xnor U10540 (N_10540,N_9220,N_9048);
or U10541 (N_10541,N_9583,N_9729);
and U10542 (N_10542,N_9206,N_9150);
and U10543 (N_10543,N_9524,N_9658);
or U10544 (N_10544,N_9283,N_9961);
nand U10545 (N_10545,N_9759,N_9183);
xnor U10546 (N_10546,N_9677,N_9160);
nor U10547 (N_10547,N_9465,N_9982);
or U10548 (N_10548,N_9081,N_9874);
and U10549 (N_10549,N_9642,N_9931);
or U10550 (N_10550,N_9036,N_9581);
nor U10551 (N_10551,N_9222,N_9215);
xor U10552 (N_10552,N_9121,N_9908);
or U10553 (N_10553,N_9949,N_9325);
nand U10554 (N_10554,N_9019,N_9103);
nor U10555 (N_10555,N_9817,N_9637);
xor U10556 (N_10556,N_9304,N_9398);
nor U10557 (N_10557,N_9782,N_9647);
or U10558 (N_10558,N_9822,N_9093);
xor U10559 (N_10559,N_9556,N_9499);
or U10560 (N_10560,N_9778,N_9887);
and U10561 (N_10561,N_9508,N_9073);
or U10562 (N_10562,N_9583,N_9927);
nand U10563 (N_10563,N_9015,N_9432);
nor U10564 (N_10564,N_9577,N_9455);
xnor U10565 (N_10565,N_9249,N_9175);
and U10566 (N_10566,N_9187,N_9878);
nor U10567 (N_10567,N_9197,N_9108);
nor U10568 (N_10568,N_9361,N_9948);
xor U10569 (N_10569,N_9994,N_9610);
and U10570 (N_10570,N_9689,N_9929);
xor U10571 (N_10571,N_9734,N_9085);
or U10572 (N_10572,N_9067,N_9740);
nor U10573 (N_10573,N_9330,N_9910);
and U10574 (N_10574,N_9005,N_9002);
nand U10575 (N_10575,N_9547,N_9587);
xnor U10576 (N_10576,N_9346,N_9353);
xor U10577 (N_10577,N_9831,N_9023);
nor U10578 (N_10578,N_9955,N_9711);
nand U10579 (N_10579,N_9777,N_9425);
or U10580 (N_10580,N_9855,N_9337);
or U10581 (N_10581,N_9068,N_9805);
nor U10582 (N_10582,N_9098,N_9184);
nor U10583 (N_10583,N_9238,N_9398);
xor U10584 (N_10584,N_9953,N_9553);
nor U10585 (N_10585,N_9846,N_9575);
nor U10586 (N_10586,N_9868,N_9305);
and U10587 (N_10587,N_9932,N_9529);
or U10588 (N_10588,N_9864,N_9565);
nor U10589 (N_10589,N_9794,N_9448);
xnor U10590 (N_10590,N_9093,N_9389);
or U10591 (N_10591,N_9058,N_9326);
nand U10592 (N_10592,N_9357,N_9625);
nand U10593 (N_10593,N_9041,N_9722);
and U10594 (N_10594,N_9150,N_9507);
nor U10595 (N_10595,N_9313,N_9101);
and U10596 (N_10596,N_9601,N_9117);
and U10597 (N_10597,N_9880,N_9587);
and U10598 (N_10598,N_9694,N_9209);
xor U10599 (N_10599,N_9444,N_9579);
nand U10600 (N_10600,N_9388,N_9592);
nand U10601 (N_10601,N_9444,N_9424);
or U10602 (N_10602,N_9961,N_9618);
or U10603 (N_10603,N_9077,N_9297);
or U10604 (N_10604,N_9099,N_9168);
or U10605 (N_10605,N_9566,N_9151);
nor U10606 (N_10606,N_9496,N_9036);
nor U10607 (N_10607,N_9345,N_9288);
xnor U10608 (N_10608,N_9815,N_9098);
xnor U10609 (N_10609,N_9014,N_9504);
xnor U10610 (N_10610,N_9332,N_9299);
xor U10611 (N_10611,N_9940,N_9808);
xnor U10612 (N_10612,N_9994,N_9016);
nor U10613 (N_10613,N_9533,N_9573);
and U10614 (N_10614,N_9399,N_9881);
nand U10615 (N_10615,N_9295,N_9079);
and U10616 (N_10616,N_9777,N_9911);
nor U10617 (N_10617,N_9979,N_9047);
nor U10618 (N_10618,N_9673,N_9018);
nand U10619 (N_10619,N_9718,N_9320);
nor U10620 (N_10620,N_9643,N_9181);
nand U10621 (N_10621,N_9553,N_9118);
and U10622 (N_10622,N_9758,N_9261);
and U10623 (N_10623,N_9261,N_9851);
or U10624 (N_10624,N_9683,N_9378);
nand U10625 (N_10625,N_9553,N_9555);
or U10626 (N_10626,N_9232,N_9291);
and U10627 (N_10627,N_9178,N_9339);
or U10628 (N_10628,N_9172,N_9252);
xor U10629 (N_10629,N_9710,N_9463);
and U10630 (N_10630,N_9035,N_9733);
or U10631 (N_10631,N_9996,N_9641);
nand U10632 (N_10632,N_9304,N_9827);
xor U10633 (N_10633,N_9757,N_9904);
nor U10634 (N_10634,N_9171,N_9468);
nor U10635 (N_10635,N_9317,N_9864);
xnor U10636 (N_10636,N_9178,N_9789);
nor U10637 (N_10637,N_9613,N_9388);
xor U10638 (N_10638,N_9422,N_9968);
and U10639 (N_10639,N_9100,N_9922);
nand U10640 (N_10640,N_9282,N_9844);
or U10641 (N_10641,N_9413,N_9892);
nor U10642 (N_10642,N_9802,N_9437);
or U10643 (N_10643,N_9659,N_9789);
nor U10644 (N_10644,N_9666,N_9088);
xor U10645 (N_10645,N_9940,N_9467);
nor U10646 (N_10646,N_9723,N_9627);
xor U10647 (N_10647,N_9811,N_9031);
nand U10648 (N_10648,N_9322,N_9581);
nand U10649 (N_10649,N_9194,N_9816);
or U10650 (N_10650,N_9016,N_9949);
nand U10651 (N_10651,N_9630,N_9502);
nor U10652 (N_10652,N_9693,N_9689);
or U10653 (N_10653,N_9869,N_9022);
xnor U10654 (N_10654,N_9231,N_9624);
nor U10655 (N_10655,N_9558,N_9616);
and U10656 (N_10656,N_9072,N_9288);
nor U10657 (N_10657,N_9244,N_9700);
and U10658 (N_10658,N_9451,N_9684);
nor U10659 (N_10659,N_9841,N_9887);
or U10660 (N_10660,N_9021,N_9180);
and U10661 (N_10661,N_9637,N_9416);
or U10662 (N_10662,N_9427,N_9512);
or U10663 (N_10663,N_9918,N_9478);
nand U10664 (N_10664,N_9660,N_9197);
nand U10665 (N_10665,N_9828,N_9075);
nand U10666 (N_10666,N_9652,N_9008);
nor U10667 (N_10667,N_9706,N_9625);
nor U10668 (N_10668,N_9052,N_9735);
and U10669 (N_10669,N_9951,N_9367);
or U10670 (N_10670,N_9291,N_9367);
xnor U10671 (N_10671,N_9425,N_9906);
xnor U10672 (N_10672,N_9845,N_9272);
nand U10673 (N_10673,N_9855,N_9770);
or U10674 (N_10674,N_9452,N_9742);
or U10675 (N_10675,N_9049,N_9752);
and U10676 (N_10676,N_9048,N_9567);
nor U10677 (N_10677,N_9819,N_9327);
nand U10678 (N_10678,N_9037,N_9321);
and U10679 (N_10679,N_9030,N_9591);
and U10680 (N_10680,N_9027,N_9753);
xor U10681 (N_10681,N_9688,N_9562);
or U10682 (N_10682,N_9628,N_9076);
nor U10683 (N_10683,N_9275,N_9353);
or U10684 (N_10684,N_9315,N_9885);
nor U10685 (N_10685,N_9568,N_9761);
and U10686 (N_10686,N_9383,N_9768);
and U10687 (N_10687,N_9111,N_9101);
xor U10688 (N_10688,N_9409,N_9773);
and U10689 (N_10689,N_9692,N_9508);
or U10690 (N_10690,N_9123,N_9574);
nor U10691 (N_10691,N_9791,N_9829);
and U10692 (N_10692,N_9505,N_9430);
or U10693 (N_10693,N_9304,N_9585);
and U10694 (N_10694,N_9824,N_9040);
nor U10695 (N_10695,N_9085,N_9448);
nor U10696 (N_10696,N_9274,N_9954);
nand U10697 (N_10697,N_9220,N_9782);
nand U10698 (N_10698,N_9728,N_9843);
xor U10699 (N_10699,N_9186,N_9583);
xor U10700 (N_10700,N_9319,N_9927);
xnor U10701 (N_10701,N_9546,N_9062);
and U10702 (N_10702,N_9891,N_9920);
or U10703 (N_10703,N_9206,N_9136);
xnor U10704 (N_10704,N_9451,N_9676);
and U10705 (N_10705,N_9081,N_9884);
xnor U10706 (N_10706,N_9608,N_9086);
nor U10707 (N_10707,N_9064,N_9208);
xnor U10708 (N_10708,N_9461,N_9524);
nand U10709 (N_10709,N_9108,N_9589);
nor U10710 (N_10710,N_9663,N_9299);
nor U10711 (N_10711,N_9014,N_9930);
nand U10712 (N_10712,N_9975,N_9997);
xnor U10713 (N_10713,N_9368,N_9821);
nor U10714 (N_10714,N_9844,N_9112);
or U10715 (N_10715,N_9431,N_9181);
or U10716 (N_10716,N_9000,N_9969);
xor U10717 (N_10717,N_9726,N_9335);
nand U10718 (N_10718,N_9264,N_9226);
nor U10719 (N_10719,N_9797,N_9140);
nor U10720 (N_10720,N_9824,N_9501);
nor U10721 (N_10721,N_9207,N_9358);
xor U10722 (N_10722,N_9137,N_9383);
or U10723 (N_10723,N_9137,N_9318);
xor U10724 (N_10724,N_9242,N_9178);
xor U10725 (N_10725,N_9158,N_9260);
nand U10726 (N_10726,N_9370,N_9049);
nor U10727 (N_10727,N_9783,N_9591);
nor U10728 (N_10728,N_9292,N_9534);
nand U10729 (N_10729,N_9750,N_9083);
or U10730 (N_10730,N_9632,N_9547);
and U10731 (N_10731,N_9320,N_9404);
nor U10732 (N_10732,N_9205,N_9785);
or U10733 (N_10733,N_9254,N_9965);
nand U10734 (N_10734,N_9430,N_9557);
nand U10735 (N_10735,N_9066,N_9031);
or U10736 (N_10736,N_9268,N_9242);
and U10737 (N_10737,N_9360,N_9645);
xnor U10738 (N_10738,N_9525,N_9090);
or U10739 (N_10739,N_9496,N_9770);
nand U10740 (N_10740,N_9988,N_9810);
nor U10741 (N_10741,N_9829,N_9388);
or U10742 (N_10742,N_9972,N_9875);
or U10743 (N_10743,N_9835,N_9939);
xnor U10744 (N_10744,N_9257,N_9083);
or U10745 (N_10745,N_9428,N_9068);
nand U10746 (N_10746,N_9421,N_9744);
nor U10747 (N_10747,N_9276,N_9116);
nand U10748 (N_10748,N_9003,N_9207);
nor U10749 (N_10749,N_9197,N_9115);
nand U10750 (N_10750,N_9754,N_9008);
xnor U10751 (N_10751,N_9784,N_9722);
nor U10752 (N_10752,N_9115,N_9664);
and U10753 (N_10753,N_9290,N_9736);
and U10754 (N_10754,N_9619,N_9565);
nor U10755 (N_10755,N_9488,N_9755);
nor U10756 (N_10756,N_9208,N_9441);
and U10757 (N_10757,N_9412,N_9031);
and U10758 (N_10758,N_9086,N_9210);
nand U10759 (N_10759,N_9882,N_9113);
xor U10760 (N_10760,N_9754,N_9263);
or U10761 (N_10761,N_9982,N_9191);
nor U10762 (N_10762,N_9603,N_9574);
or U10763 (N_10763,N_9603,N_9062);
nand U10764 (N_10764,N_9154,N_9105);
nand U10765 (N_10765,N_9441,N_9981);
nor U10766 (N_10766,N_9242,N_9726);
nor U10767 (N_10767,N_9354,N_9536);
nand U10768 (N_10768,N_9574,N_9147);
nor U10769 (N_10769,N_9485,N_9518);
xnor U10770 (N_10770,N_9559,N_9408);
nand U10771 (N_10771,N_9685,N_9479);
nand U10772 (N_10772,N_9980,N_9018);
xor U10773 (N_10773,N_9442,N_9757);
or U10774 (N_10774,N_9186,N_9746);
and U10775 (N_10775,N_9708,N_9382);
or U10776 (N_10776,N_9954,N_9060);
xnor U10777 (N_10777,N_9738,N_9665);
or U10778 (N_10778,N_9230,N_9201);
or U10779 (N_10779,N_9083,N_9703);
nand U10780 (N_10780,N_9564,N_9967);
or U10781 (N_10781,N_9404,N_9811);
and U10782 (N_10782,N_9934,N_9216);
xor U10783 (N_10783,N_9239,N_9084);
or U10784 (N_10784,N_9424,N_9904);
xnor U10785 (N_10785,N_9738,N_9458);
nand U10786 (N_10786,N_9171,N_9331);
and U10787 (N_10787,N_9410,N_9171);
and U10788 (N_10788,N_9031,N_9688);
or U10789 (N_10789,N_9989,N_9939);
nor U10790 (N_10790,N_9336,N_9329);
and U10791 (N_10791,N_9443,N_9802);
nand U10792 (N_10792,N_9723,N_9739);
nand U10793 (N_10793,N_9200,N_9162);
nand U10794 (N_10794,N_9455,N_9161);
nand U10795 (N_10795,N_9692,N_9216);
xnor U10796 (N_10796,N_9463,N_9006);
xor U10797 (N_10797,N_9931,N_9724);
xor U10798 (N_10798,N_9399,N_9435);
and U10799 (N_10799,N_9511,N_9052);
xor U10800 (N_10800,N_9636,N_9498);
or U10801 (N_10801,N_9725,N_9808);
xnor U10802 (N_10802,N_9279,N_9034);
and U10803 (N_10803,N_9971,N_9191);
nand U10804 (N_10804,N_9308,N_9930);
xor U10805 (N_10805,N_9828,N_9248);
xor U10806 (N_10806,N_9005,N_9498);
and U10807 (N_10807,N_9290,N_9767);
nand U10808 (N_10808,N_9416,N_9009);
nand U10809 (N_10809,N_9531,N_9480);
xor U10810 (N_10810,N_9516,N_9491);
nand U10811 (N_10811,N_9376,N_9893);
nor U10812 (N_10812,N_9232,N_9710);
xnor U10813 (N_10813,N_9649,N_9842);
or U10814 (N_10814,N_9377,N_9616);
nand U10815 (N_10815,N_9933,N_9038);
xnor U10816 (N_10816,N_9055,N_9914);
nand U10817 (N_10817,N_9011,N_9054);
or U10818 (N_10818,N_9708,N_9997);
nor U10819 (N_10819,N_9245,N_9510);
nand U10820 (N_10820,N_9455,N_9802);
nor U10821 (N_10821,N_9789,N_9834);
nor U10822 (N_10822,N_9414,N_9433);
and U10823 (N_10823,N_9801,N_9225);
xor U10824 (N_10824,N_9115,N_9355);
and U10825 (N_10825,N_9970,N_9036);
or U10826 (N_10826,N_9799,N_9846);
nand U10827 (N_10827,N_9566,N_9526);
xor U10828 (N_10828,N_9644,N_9657);
xor U10829 (N_10829,N_9134,N_9592);
nand U10830 (N_10830,N_9252,N_9759);
nand U10831 (N_10831,N_9859,N_9007);
nor U10832 (N_10832,N_9804,N_9240);
nor U10833 (N_10833,N_9431,N_9849);
xnor U10834 (N_10834,N_9540,N_9791);
and U10835 (N_10835,N_9069,N_9961);
nor U10836 (N_10836,N_9941,N_9153);
and U10837 (N_10837,N_9171,N_9874);
xnor U10838 (N_10838,N_9209,N_9202);
or U10839 (N_10839,N_9665,N_9490);
and U10840 (N_10840,N_9717,N_9826);
and U10841 (N_10841,N_9419,N_9166);
xor U10842 (N_10842,N_9851,N_9835);
xnor U10843 (N_10843,N_9589,N_9156);
and U10844 (N_10844,N_9187,N_9103);
nor U10845 (N_10845,N_9296,N_9100);
xnor U10846 (N_10846,N_9999,N_9728);
and U10847 (N_10847,N_9219,N_9589);
nor U10848 (N_10848,N_9890,N_9410);
and U10849 (N_10849,N_9649,N_9626);
or U10850 (N_10850,N_9922,N_9236);
nand U10851 (N_10851,N_9681,N_9945);
nand U10852 (N_10852,N_9381,N_9440);
and U10853 (N_10853,N_9292,N_9638);
and U10854 (N_10854,N_9795,N_9960);
or U10855 (N_10855,N_9196,N_9920);
or U10856 (N_10856,N_9898,N_9312);
and U10857 (N_10857,N_9480,N_9290);
xor U10858 (N_10858,N_9769,N_9470);
or U10859 (N_10859,N_9834,N_9262);
nand U10860 (N_10860,N_9469,N_9076);
and U10861 (N_10861,N_9849,N_9125);
xor U10862 (N_10862,N_9956,N_9755);
xnor U10863 (N_10863,N_9496,N_9462);
xnor U10864 (N_10864,N_9450,N_9933);
nand U10865 (N_10865,N_9470,N_9735);
nand U10866 (N_10866,N_9911,N_9615);
xor U10867 (N_10867,N_9587,N_9119);
and U10868 (N_10868,N_9828,N_9092);
xor U10869 (N_10869,N_9507,N_9050);
nor U10870 (N_10870,N_9033,N_9811);
xnor U10871 (N_10871,N_9074,N_9125);
nand U10872 (N_10872,N_9265,N_9023);
xnor U10873 (N_10873,N_9902,N_9735);
and U10874 (N_10874,N_9238,N_9806);
xnor U10875 (N_10875,N_9807,N_9248);
or U10876 (N_10876,N_9710,N_9429);
or U10877 (N_10877,N_9517,N_9162);
xnor U10878 (N_10878,N_9007,N_9231);
and U10879 (N_10879,N_9090,N_9878);
and U10880 (N_10880,N_9267,N_9459);
nor U10881 (N_10881,N_9977,N_9810);
or U10882 (N_10882,N_9136,N_9104);
and U10883 (N_10883,N_9324,N_9400);
or U10884 (N_10884,N_9866,N_9338);
nand U10885 (N_10885,N_9545,N_9076);
and U10886 (N_10886,N_9844,N_9433);
nor U10887 (N_10887,N_9224,N_9559);
and U10888 (N_10888,N_9074,N_9779);
and U10889 (N_10889,N_9937,N_9248);
nand U10890 (N_10890,N_9225,N_9870);
or U10891 (N_10891,N_9021,N_9329);
nor U10892 (N_10892,N_9559,N_9843);
nor U10893 (N_10893,N_9511,N_9194);
and U10894 (N_10894,N_9258,N_9094);
nand U10895 (N_10895,N_9059,N_9410);
and U10896 (N_10896,N_9483,N_9261);
nor U10897 (N_10897,N_9264,N_9276);
or U10898 (N_10898,N_9613,N_9684);
or U10899 (N_10899,N_9267,N_9338);
nor U10900 (N_10900,N_9570,N_9055);
and U10901 (N_10901,N_9966,N_9364);
xor U10902 (N_10902,N_9724,N_9232);
and U10903 (N_10903,N_9100,N_9307);
and U10904 (N_10904,N_9833,N_9432);
or U10905 (N_10905,N_9188,N_9778);
nor U10906 (N_10906,N_9211,N_9275);
nand U10907 (N_10907,N_9284,N_9494);
nor U10908 (N_10908,N_9523,N_9017);
and U10909 (N_10909,N_9187,N_9058);
nor U10910 (N_10910,N_9497,N_9869);
or U10911 (N_10911,N_9296,N_9610);
nand U10912 (N_10912,N_9200,N_9622);
or U10913 (N_10913,N_9509,N_9793);
nand U10914 (N_10914,N_9986,N_9658);
or U10915 (N_10915,N_9900,N_9307);
nor U10916 (N_10916,N_9367,N_9855);
xnor U10917 (N_10917,N_9620,N_9793);
nand U10918 (N_10918,N_9264,N_9325);
nand U10919 (N_10919,N_9273,N_9815);
and U10920 (N_10920,N_9936,N_9074);
xor U10921 (N_10921,N_9168,N_9988);
or U10922 (N_10922,N_9779,N_9948);
nor U10923 (N_10923,N_9415,N_9955);
or U10924 (N_10924,N_9910,N_9695);
or U10925 (N_10925,N_9716,N_9921);
and U10926 (N_10926,N_9558,N_9549);
nor U10927 (N_10927,N_9300,N_9016);
and U10928 (N_10928,N_9601,N_9670);
or U10929 (N_10929,N_9651,N_9859);
and U10930 (N_10930,N_9206,N_9660);
nand U10931 (N_10931,N_9587,N_9136);
and U10932 (N_10932,N_9639,N_9620);
xor U10933 (N_10933,N_9404,N_9117);
or U10934 (N_10934,N_9537,N_9033);
xor U10935 (N_10935,N_9283,N_9474);
xor U10936 (N_10936,N_9879,N_9431);
or U10937 (N_10937,N_9298,N_9058);
nand U10938 (N_10938,N_9898,N_9335);
or U10939 (N_10939,N_9163,N_9735);
and U10940 (N_10940,N_9509,N_9045);
and U10941 (N_10941,N_9283,N_9761);
nand U10942 (N_10942,N_9947,N_9451);
nand U10943 (N_10943,N_9978,N_9329);
xor U10944 (N_10944,N_9518,N_9366);
nand U10945 (N_10945,N_9645,N_9484);
xor U10946 (N_10946,N_9872,N_9034);
or U10947 (N_10947,N_9462,N_9525);
xnor U10948 (N_10948,N_9931,N_9101);
or U10949 (N_10949,N_9820,N_9783);
or U10950 (N_10950,N_9708,N_9658);
xnor U10951 (N_10951,N_9597,N_9037);
nor U10952 (N_10952,N_9305,N_9928);
xnor U10953 (N_10953,N_9912,N_9294);
nor U10954 (N_10954,N_9715,N_9116);
and U10955 (N_10955,N_9726,N_9525);
xor U10956 (N_10956,N_9686,N_9701);
xnor U10957 (N_10957,N_9245,N_9025);
or U10958 (N_10958,N_9234,N_9746);
nand U10959 (N_10959,N_9061,N_9367);
and U10960 (N_10960,N_9748,N_9617);
nor U10961 (N_10961,N_9016,N_9376);
or U10962 (N_10962,N_9893,N_9702);
and U10963 (N_10963,N_9066,N_9367);
or U10964 (N_10964,N_9952,N_9440);
or U10965 (N_10965,N_9853,N_9013);
or U10966 (N_10966,N_9917,N_9154);
or U10967 (N_10967,N_9922,N_9194);
and U10968 (N_10968,N_9174,N_9252);
or U10969 (N_10969,N_9873,N_9570);
nor U10970 (N_10970,N_9011,N_9554);
and U10971 (N_10971,N_9103,N_9378);
nand U10972 (N_10972,N_9847,N_9797);
nand U10973 (N_10973,N_9289,N_9344);
or U10974 (N_10974,N_9408,N_9689);
nor U10975 (N_10975,N_9446,N_9740);
and U10976 (N_10976,N_9130,N_9525);
nand U10977 (N_10977,N_9312,N_9402);
nand U10978 (N_10978,N_9514,N_9462);
nor U10979 (N_10979,N_9009,N_9005);
nand U10980 (N_10980,N_9376,N_9588);
nand U10981 (N_10981,N_9200,N_9767);
or U10982 (N_10982,N_9043,N_9341);
nor U10983 (N_10983,N_9332,N_9156);
nor U10984 (N_10984,N_9398,N_9947);
xnor U10985 (N_10985,N_9507,N_9612);
and U10986 (N_10986,N_9367,N_9231);
and U10987 (N_10987,N_9645,N_9706);
nor U10988 (N_10988,N_9515,N_9865);
nor U10989 (N_10989,N_9925,N_9464);
nand U10990 (N_10990,N_9166,N_9486);
and U10991 (N_10991,N_9135,N_9040);
or U10992 (N_10992,N_9162,N_9550);
and U10993 (N_10993,N_9556,N_9651);
nor U10994 (N_10994,N_9840,N_9717);
and U10995 (N_10995,N_9537,N_9950);
and U10996 (N_10996,N_9928,N_9903);
xnor U10997 (N_10997,N_9659,N_9714);
xor U10998 (N_10998,N_9220,N_9381);
and U10999 (N_10999,N_9654,N_9491);
nand U11000 (N_11000,N_10943,N_10831);
or U11001 (N_11001,N_10161,N_10357);
and U11002 (N_11002,N_10698,N_10162);
nor U11003 (N_11003,N_10348,N_10886);
and U11004 (N_11004,N_10062,N_10879);
xor U11005 (N_11005,N_10141,N_10805);
xnor U11006 (N_11006,N_10350,N_10925);
nand U11007 (N_11007,N_10099,N_10036);
nand U11008 (N_11008,N_10351,N_10662);
or U11009 (N_11009,N_10987,N_10215);
nand U11010 (N_11010,N_10359,N_10221);
nand U11011 (N_11011,N_10848,N_10871);
xor U11012 (N_11012,N_10173,N_10420);
xor U11013 (N_11013,N_10236,N_10776);
xor U11014 (N_11014,N_10564,N_10815);
nor U11015 (N_11015,N_10619,N_10788);
or U11016 (N_11016,N_10074,N_10859);
nor U11017 (N_11017,N_10745,N_10755);
nor U11018 (N_11018,N_10884,N_10835);
nor U11019 (N_11019,N_10393,N_10344);
xnor U11020 (N_11020,N_10069,N_10136);
xor U11021 (N_11021,N_10550,N_10211);
nand U11022 (N_11022,N_10189,N_10433);
nand U11023 (N_11023,N_10511,N_10204);
and U11024 (N_11024,N_10363,N_10311);
or U11025 (N_11025,N_10981,N_10532);
nor U11026 (N_11026,N_10616,N_10440);
and U11027 (N_11027,N_10985,N_10458);
or U11028 (N_11028,N_10086,N_10728);
and U11029 (N_11029,N_10920,N_10515);
nor U11030 (N_11030,N_10414,N_10322);
and U11031 (N_11031,N_10463,N_10097);
and U11032 (N_11032,N_10064,N_10793);
or U11033 (N_11033,N_10775,N_10177);
xnor U11034 (N_11034,N_10536,N_10618);
and U11035 (N_11035,N_10449,N_10757);
or U11036 (N_11036,N_10356,N_10584);
or U11037 (N_11037,N_10464,N_10687);
nand U11038 (N_11038,N_10594,N_10644);
xor U11039 (N_11039,N_10545,N_10398);
nor U11040 (N_11040,N_10300,N_10767);
xor U11041 (N_11041,N_10736,N_10289);
nand U11042 (N_11042,N_10797,N_10499);
xor U11043 (N_11043,N_10885,N_10032);
nand U11044 (N_11044,N_10287,N_10002);
nand U11045 (N_11045,N_10600,N_10778);
nand U11046 (N_11046,N_10849,N_10853);
or U11047 (N_11047,N_10176,N_10780);
or U11048 (N_11048,N_10932,N_10593);
nor U11049 (N_11049,N_10281,N_10326);
xor U11050 (N_11050,N_10589,N_10347);
nor U11051 (N_11051,N_10954,N_10868);
or U11052 (N_11052,N_10073,N_10131);
xor U11053 (N_11053,N_10428,N_10994);
nand U11054 (N_11054,N_10270,N_10577);
nand U11055 (N_11055,N_10921,N_10934);
nor U11056 (N_11056,N_10025,N_10497);
nor U11057 (N_11057,N_10031,N_10956);
xnor U11058 (N_11058,N_10602,N_10517);
nand U11059 (N_11059,N_10383,N_10494);
nor U11060 (N_11060,N_10441,N_10333);
or U11061 (N_11061,N_10557,N_10199);
nor U11062 (N_11062,N_10685,N_10106);
and U11063 (N_11063,N_10486,N_10314);
nor U11064 (N_11064,N_10769,N_10731);
or U11065 (N_11065,N_10924,N_10462);
nor U11066 (N_11066,N_10178,N_10476);
nor U11067 (N_11067,N_10490,N_10659);
and U11068 (N_11068,N_10098,N_10562);
and U11069 (N_11069,N_10992,N_10008);
and U11070 (N_11070,N_10290,N_10092);
and U11071 (N_11071,N_10043,N_10958);
and U11072 (N_11072,N_10652,N_10792);
xor U11073 (N_11073,N_10371,N_10245);
xor U11074 (N_11074,N_10638,N_10259);
xnor U11075 (N_11075,N_10901,N_10139);
and U11076 (N_11076,N_10200,N_10624);
and U11077 (N_11077,N_10018,N_10291);
nor U11078 (N_11078,N_10172,N_10874);
nand U11079 (N_11079,N_10404,N_10096);
nor U11080 (N_11080,N_10896,N_10285);
xor U11081 (N_11081,N_10317,N_10844);
nor U11082 (N_11082,N_10058,N_10035);
or U11083 (N_11083,N_10389,N_10466);
xor U11084 (N_11084,N_10626,N_10621);
and U11085 (N_11085,N_10525,N_10524);
and U11086 (N_11086,N_10845,N_10278);
or U11087 (N_11087,N_10220,N_10916);
nand U11088 (N_11088,N_10045,N_10055);
xnor U11089 (N_11089,N_10372,N_10015);
and U11090 (N_11090,N_10858,N_10044);
nor U11091 (N_11091,N_10129,N_10457);
xor U11092 (N_11092,N_10774,N_10219);
xnor U11093 (N_11093,N_10202,N_10477);
nand U11094 (N_11094,N_10078,N_10487);
or U11095 (N_11095,N_10895,N_10764);
nand U11096 (N_11096,N_10455,N_10534);
and U11097 (N_11097,N_10654,N_10000);
or U11098 (N_11098,N_10700,N_10340);
nor U11099 (N_11099,N_10856,N_10324);
or U11100 (N_11100,N_10191,N_10334);
xnor U11101 (N_11101,N_10146,N_10240);
nand U11102 (N_11102,N_10005,N_10953);
xnor U11103 (N_11103,N_10242,N_10988);
nand U11104 (N_11104,N_10832,N_10979);
or U11105 (N_11105,N_10512,N_10699);
and U11106 (N_11106,N_10175,N_10996);
xor U11107 (N_11107,N_10902,N_10104);
xnor U11108 (N_11108,N_10418,N_10535);
and U11109 (N_11109,N_10928,N_10299);
nor U11110 (N_11110,N_10042,N_10459);
xnor U11111 (N_11111,N_10313,N_10120);
nor U11112 (N_11112,N_10822,N_10673);
nand U11113 (N_11113,N_10391,N_10234);
xnor U11114 (N_11114,N_10405,N_10377);
xnor U11115 (N_11115,N_10807,N_10452);
nor U11116 (N_11116,N_10142,N_10100);
and U11117 (N_11117,N_10130,N_10111);
and U11118 (N_11118,N_10740,N_10581);
nand U11119 (N_11119,N_10198,N_10152);
xor U11120 (N_11120,N_10663,N_10244);
xnor U11121 (N_11121,N_10110,N_10003);
and U11122 (N_11122,N_10810,N_10117);
nor U11123 (N_11123,N_10072,N_10272);
xor U11124 (N_11124,N_10900,N_10696);
nand U11125 (N_11125,N_10375,N_10158);
and U11126 (N_11126,N_10709,N_10399);
xor U11127 (N_11127,N_10516,N_10882);
or U11128 (N_11128,N_10783,N_10880);
or U11129 (N_11129,N_10303,N_10506);
and U11130 (N_11130,N_10020,N_10489);
xor U11131 (N_11131,N_10551,N_10495);
nand U11132 (N_11132,N_10688,N_10249);
and U11133 (N_11133,N_10226,N_10546);
nand U11134 (N_11134,N_10869,N_10770);
and U11135 (N_11135,N_10573,N_10331);
nand U11136 (N_11136,N_10316,N_10079);
xor U11137 (N_11137,N_10799,N_10505);
xor U11138 (N_11138,N_10364,N_10966);
nand U11139 (N_11139,N_10570,N_10125);
xor U11140 (N_11140,N_10867,N_10425);
xor U11141 (N_11141,N_10446,N_10250);
xor U11142 (N_11142,N_10268,N_10894);
xnor U11143 (N_11143,N_10530,N_10413);
nor U11144 (N_11144,N_10145,N_10187);
xor U11145 (N_11145,N_10637,N_10615);
nor U11146 (N_11146,N_10210,N_10075);
and U11147 (N_11147,N_10641,N_10430);
nor U11148 (N_11148,N_10473,N_10263);
nand U11149 (N_11149,N_10620,N_10697);
xnor U11150 (N_11150,N_10968,N_10837);
and U11151 (N_11151,N_10046,N_10862);
nand U11152 (N_11152,N_10491,N_10468);
and U11153 (N_11153,N_10059,N_10193);
nor U11154 (N_11154,N_10986,N_10328);
nor U11155 (N_11155,N_10784,N_10238);
nor U11156 (N_11156,N_10016,N_10857);
xnor U11157 (N_11157,N_10407,N_10197);
nor U11158 (N_11158,N_10386,N_10758);
or U11159 (N_11159,N_10355,N_10980);
and U11160 (N_11160,N_10049,N_10819);
xor U11161 (N_11161,N_10456,N_10684);
xnor U11162 (N_11162,N_10048,N_10261);
or U11163 (N_11163,N_10442,N_10646);
and U11164 (N_11164,N_10312,N_10601);
xnor U11165 (N_11165,N_10260,N_10686);
nor U11166 (N_11166,N_10645,N_10254);
and U11167 (N_11167,N_10415,N_10765);
nor U11168 (N_11168,N_10955,N_10742);
nand U11169 (N_11169,N_10960,N_10431);
nor U11170 (N_11170,N_10747,N_10575);
or U11171 (N_11171,N_10706,N_10115);
nor U11172 (N_11172,N_10450,N_10997);
nand U11173 (N_11173,N_10548,N_10520);
nor U11174 (N_11174,N_10631,N_10999);
or U11175 (N_11175,N_10174,N_10427);
or U11176 (N_11176,N_10338,N_10112);
nand U11177 (N_11177,N_10402,N_10453);
nand U11178 (N_11178,N_10563,N_10108);
xnor U11179 (N_11179,N_10066,N_10729);
and U11180 (N_11180,N_10056,N_10274);
xnor U11181 (N_11181,N_10649,N_10216);
nand U11182 (N_11182,N_10498,N_10039);
xor U11183 (N_11183,N_10022,N_10823);
nand U11184 (N_11184,N_10599,N_10743);
and U11185 (N_11185,N_10976,N_10623);
and U11186 (N_11186,N_10625,N_10277);
and U11187 (N_11187,N_10669,N_10258);
nand U11188 (N_11188,N_10472,N_10768);
and U11189 (N_11189,N_10243,N_10710);
and U11190 (N_11190,N_10713,N_10276);
nor U11191 (N_11191,N_10756,N_10082);
nor U11192 (N_11192,N_10318,N_10782);
and U11193 (N_11193,N_10689,N_10122);
nor U11194 (N_11194,N_10301,N_10021);
nand U11195 (N_11195,N_10384,N_10975);
and U11196 (N_11196,N_10423,N_10737);
nand U11197 (N_11197,N_10915,N_10722);
xor U11198 (N_11198,N_10116,N_10860);
nand U11199 (N_11199,N_10567,N_10478);
and U11200 (N_11200,N_10531,N_10762);
and U11201 (N_11201,N_10825,N_10692);
nand U11202 (N_11202,N_10041,N_10123);
xnor U11203 (N_11203,N_10292,N_10439);
xor U11204 (N_11204,N_10070,N_10801);
nand U11205 (N_11205,N_10503,N_10445);
nor U11206 (N_11206,N_10582,N_10339);
nor U11207 (N_11207,N_10488,N_10933);
or U11208 (N_11208,N_10962,N_10865);
nor U11209 (N_11209,N_10648,N_10561);
or U11210 (N_11210,N_10007,N_10169);
xor U11211 (N_11211,N_10566,N_10113);
or U11212 (N_11212,N_10940,N_10565);
nor U11213 (N_11213,N_10163,N_10772);
or U11214 (N_11214,N_10114,N_10872);
nor U11215 (N_11215,N_10461,N_10222);
or U11216 (N_11216,N_10948,N_10787);
and U11217 (N_11217,N_10381,N_10374);
nand U11218 (N_11218,N_10647,N_10961);
xnor U11219 (N_11219,N_10734,N_10887);
nor U11220 (N_11220,N_10542,N_10580);
nor U11221 (N_11221,N_10038,N_10057);
xor U11222 (N_11222,N_10855,N_10795);
and U11223 (N_11223,N_10027,N_10460);
and U11224 (N_11224,N_10556,N_10060);
nor U11225 (N_11225,N_10668,N_10089);
xor U11226 (N_11226,N_10369,N_10388);
xnor U11227 (N_11227,N_10540,N_10674);
and U11228 (N_11228,N_10320,N_10119);
and U11229 (N_11229,N_10101,N_10904);
and U11230 (N_11230,N_10410,N_10217);
or U11231 (N_11231,N_10998,N_10085);
and U11232 (N_11232,N_10063,N_10906);
and U11233 (N_11233,N_10727,N_10714);
and U11234 (N_11234,N_10135,N_10083);
and U11235 (N_11235,N_10401,N_10379);
and U11236 (N_11236,N_10675,N_10467);
nand U11237 (N_11237,N_10591,N_10306);
or U11238 (N_11238,N_10761,N_10804);
nand U11239 (N_11239,N_10352,N_10970);
xnor U11240 (N_11240,N_10485,N_10847);
or U11241 (N_11241,N_10409,N_10875);
nor U11242 (N_11242,N_10167,N_10617);
and U11243 (N_11243,N_10529,N_10429);
and U11244 (N_11244,N_10773,N_10387);
nor U11245 (N_11245,N_10814,N_10910);
and U11246 (N_11246,N_10877,N_10701);
nor U11247 (N_11247,N_10088,N_10206);
or U11248 (N_11248,N_10051,N_10752);
and U11249 (N_11249,N_10667,N_10500);
nand U11250 (N_11250,N_10155,N_10343);
nand U11251 (N_11251,N_10269,N_10241);
and U11252 (N_11252,N_10253,N_10733);
nor U11253 (N_11253,N_10481,N_10208);
nand U11254 (N_11254,N_10411,N_10978);
and U11255 (N_11255,N_10661,N_10597);
nor U11256 (N_11256,N_10385,N_10917);
and U11257 (N_11257,N_10811,N_10544);
xor U11258 (N_11258,N_10543,N_10518);
and U11259 (N_11259,N_10225,N_10212);
and U11260 (N_11260,N_10721,N_10907);
or U11261 (N_11261,N_10345,N_10337);
or U11262 (N_11262,N_10444,N_10033);
or U11263 (N_11263,N_10820,N_10930);
or U11264 (N_11264,N_10026,N_10507);
nand U11265 (N_11265,N_10090,N_10295);
nand U11266 (N_11266,N_10144,N_10315);
and U11267 (N_11267,N_10678,N_10977);
or U11268 (N_11268,N_10432,N_10680);
nor U11269 (N_11269,N_10982,N_10156);
nor U11270 (N_11270,N_10702,N_10818);
nor U11271 (N_11271,N_10660,N_10703);
nand U11272 (N_11272,N_10103,N_10942);
nor U11273 (N_11273,N_10179,N_10246);
and U11274 (N_11274,N_10671,N_10469);
and U11275 (N_11275,N_10346,N_10817);
and U11276 (N_11276,N_10170,N_10213);
or U11277 (N_11277,N_10124,N_10121);
xor U11278 (N_11278,N_10951,N_10666);
nor U11279 (N_11279,N_10627,N_10813);
or U11280 (N_11280,N_10188,N_10991);
nand U11281 (N_11281,N_10889,N_10195);
nor U11282 (N_11282,N_10012,N_10571);
nand U11283 (N_11283,N_10914,N_10358);
xnor U11284 (N_11284,N_10912,N_10255);
nor U11285 (N_11285,N_10830,N_10927);
nor U11286 (N_11286,N_10081,N_10382);
xnor U11287 (N_11287,N_10950,N_10808);
nor U11288 (N_11288,N_10650,N_10061);
or U11289 (N_11289,N_10585,N_10257);
nand U11290 (N_11290,N_10559,N_10077);
nor U11291 (N_11291,N_10102,N_10554);
and U11292 (N_11292,N_10911,N_10746);
nand U11293 (N_11293,N_10635,N_10194);
or U11294 (N_11294,N_10019,N_10093);
or U11295 (N_11295,N_10483,N_10523);
and U11296 (N_11296,N_10034,N_10040);
and U11297 (N_11297,N_10947,N_10403);
or U11298 (N_11298,N_10735,N_10368);
nor U11299 (N_11299,N_10555,N_10574);
nand U11300 (N_11300,N_10223,N_10612);
nor U11301 (N_11301,N_10154,N_10717);
or U11302 (N_11302,N_10267,N_10741);
and U11303 (N_11303,N_10610,N_10838);
xor U11304 (N_11304,N_10636,N_10604);
nor U11305 (N_11305,N_10839,N_10821);
xor U11306 (N_11306,N_10816,N_10944);
nand U11307 (N_11307,N_10547,N_10127);
xor U11308 (N_11308,N_10068,N_10993);
or U11309 (N_11309,N_10168,N_10959);
or U11310 (N_11310,N_10608,N_10852);
nand U11311 (N_11311,N_10651,N_10370);
nor U11312 (N_11312,N_10587,N_10024);
nand U11313 (N_11313,N_10185,N_10030);
xnor U11314 (N_11314,N_10286,N_10421);
and U11315 (N_11315,N_10094,N_10332);
nor U11316 (N_11316,N_10192,N_10938);
or U11317 (N_11317,N_10010,N_10247);
nor U11318 (N_11318,N_10630,N_10201);
and U11319 (N_11319,N_10378,N_10897);
and U11320 (N_11320,N_10160,N_10922);
xor U11321 (N_11321,N_10264,N_10873);
or U11322 (N_11322,N_10309,N_10723);
xor U11323 (N_11323,N_10796,N_10794);
xnor U11324 (N_11324,N_10308,N_10205);
nand U11325 (N_11325,N_10307,N_10798);
nor U11326 (N_11326,N_10899,N_10426);
or U11327 (N_11327,N_10186,N_10971);
and U11328 (N_11328,N_10084,N_10406);
xor U11329 (N_11329,N_10228,N_10539);
nand U11330 (N_11330,N_10480,N_10973);
nand U11331 (N_11331,N_10826,N_10560);
nor U11332 (N_11332,N_10329,N_10424);
or U11333 (N_11333,N_10779,N_10298);
and U11334 (N_11334,N_10164,N_10613);
and U11335 (N_11335,N_10157,N_10576);
nand U11336 (N_11336,N_10588,N_10964);
or U11337 (N_11337,N_10726,N_10622);
and U11338 (N_11338,N_10282,N_10229);
nor U11339 (N_11339,N_10454,N_10321);
and U11340 (N_11340,N_10800,N_10829);
or U11341 (N_11341,N_10840,N_10677);
xnor U11342 (N_11342,N_10294,N_10437);
or U11343 (N_11343,N_10558,N_10171);
nor U11344 (N_11344,N_10809,N_10676);
and U11345 (N_11345,N_10395,N_10908);
nor U11346 (N_11346,N_10080,N_10360);
nand U11347 (N_11347,N_10009,N_10732);
and U11348 (N_11348,N_10447,N_10209);
xnor U11349 (N_11349,N_10143,N_10004);
and U11350 (N_11350,N_10422,N_10715);
nand U11351 (N_11351,N_10704,N_10744);
and U11352 (N_11352,N_10288,N_10640);
nand U11353 (N_11353,N_10603,N_10750);
nor U11354 (N_11354,N_10541,N_10341);
nand U11355 (N_11355,N_10929,N_10695);
nand U11356 (N_11356,N_10140,N_10510);
xor U11357 (N_11357,N_10514,N_10790);
and U11358 (N_11358,N_10011,N_10974);
xor U11359 (N_11359,N_10777,N_10786);
xor U11360 (N_11360,N_10438,N_10076);
nand U11361 (N_11361,N_10293,N_10656);
xor U11362 (N_11362,N_10023,N_10946);
or U11363 (N_11363,N_10903,N_10936);
and U11364 (N_11364,N_10609,N_10785);
or U11365 (N_11365,N_10203,N_10578);
nand U11366 (N_11366,N_10711,N_10866);
or U11367 (N_11367,N_10720,N_10923);
and U11368 (N_11368,N_10716,N_10824);
or U11369 (N_11369,N_10147,N_10937);
or U11370 (N_11370,N_10682,N_10397);
nand U11371 (N_11371,N_10417,N_10771);
and U11372 (N_11372,N_10552,N_10931);
or U11373 (N_11373,N_10054,N_10605);
xor U11374 (N_11374,N_10569,N_10394);
nand U11375 (N_11375,N_10296,N_10501);
nand U11376 (N_11376,N_10607,N_10995);
nand U11377 (N_11377,N_10305,N_10724);
nor U11378 (N_11378,N_10248,N_10508);
and U11379 (N_11379,N_10606,N_10419);
nor U11380 (N_11380,N_10919,N_10284);
and U11381 (N_11381,N_10149,N_10166);
and U11382 (N_11382,N_10218,N_10583);
nand U11383 (N_11383,N_10017,N_10400);
nor U11384 (N_11384,N_10336,N_10470);
and U11385 (N_11385,N_10766,N_10071);
or U11386 (N_11386,N_10579,N_10367);
nand U11387 (N_11387,N_10230,N_10549);
and U11388 (N_11388,N_10319,N_10224);
nor U11389 (N_11389,N_10803,N_10707);
xnor U11390 (N_11390,N_10266,N_10361);
or U11391 (N_11391,N_10989,N_10893);
nand U11392 (N_11392,N_10841,N_10595);
and U11393 (N_11393,N_10196,N_10629);
xor U11394 (N_11394,N_10754,N_10392);
nor U11395 (N_11395,N_10091,N_10435);
nand U11396 (N_11396,N_10376,N_10888);
nor U11397 (N_11397,N_10683,N_10672);
nor U11398 (N_11398,N_10067,N_10492);
nor U11399 (N_11399,N_10693,N_10302);
nor U11400 (N_11400,N_10806,N_10504);
nand U11401 (N_11401,N_10365,N_10854);
and U11402 (N_11402,N_10759,N_10963);
nor U11403 (N_11403,N_10126,N_10969);
nor U11404 (N_11404,N_10132,N_10519);
and U11405 (N_11405,N_10232,N_10526);
and U11406 (N_11406,N_10107,N_10949);
nor U11407 (N_11407,N_10812,N_10926);
xor U11408 (N_11408,N_10527,N_10052);
nor U11409 (N_11409,N_10408,N_10941);
nand U11410 (N_11410,N_10753,N_10725);
nor U11411 (N_11411,N_10572,N_10751);
nor U11412 (N_11412,N_10628,N_10151);
nand U11413 (N_11413,N_10190,N_10691);
or U11414 (N_11414,N_10614,N_10690);
and U11415 (N_11415,N_10412,N_10029);
or U11416 (N_11416,N_10271,N_10967);
xnor U11417 (N_11417,N_10633,N_10180);
nor U11418 (N_11418,N_10863,N_10207);
nand U11419 (N_11419,N_10876,N_10836);
or U11420 (N_11420,N_10134,N_10730);
xor U11421 (N_11421,N_10353,N_10642);
or U11422 (N_11422,N_10065,N_10846);
nor U11423 (N_11423,N_10148,N_10050);
nor U11424 (N_11424,N_10279,N_10850);
nand U11425 (N_11425,N_10509,N_10482);
and U11426 (N_11426,N_10738,N_10828);
or U11427 (N_11427,N_10390,N_10237);
or U11428 (N_11428,N_10273,N_10833);
nand U11429 (N_11429,N_10013,N_10909);
and U11430 (N_11430,N_10434,N_10493);
or U11431 (N_11431,N_10006,N_10349);
or U11432 (N_11432,N_10883,N_10053);
xor U11433 (N_11433,N_10952,N_10513);
or U11434 (N_11434,N_10159,N_10611);
nor U11435 (N_11435,N_10150,N_10670);
or U11436 (N_11436,N_10598,N_10184);
nor U11437 (N_11437,N_10655,N_10990);
or U11438 (N_11438,N_10842,N_10262);
nor U11439 (N_11439,N_10323,N_10181);
or U11440 (N_11440,N_10763,N_10657);
nor U11441 (N_11441,N_10665,N_10479);
or U11442 (N_11442,N_10265,N_10905);
xor U11443 (N_11443,N_10643,N_10653);
nand U11444 (N_11444,N_10749,N_10105);
and U11445 (N_11445,N_10227,N_10984);
xor U11446 (N_11446,N_10165,N_10109);
and U11447 (N_11447,N_10128,N_10396);
or U11448 (N_11448,N_10416,N_10664);
xor U11449 (N_11449,N_10087,N_10708);
and U11450 (N_11450,N_10256,N_10335);
xnor U11451 (N_11451,N_10496,N_10471);
or U11452 (N_11452,N_10373,N_10451);
or U11453 (N_11453,N_10681,N_10153);
and U11454 (N_11454,N_10983,N_10330);
nand U11455 (N_11455,N_10632,N_10658);
or U11456 (N_11456,N_10639,N_10037);
nand U11457 (N_11457,N_10231,N_10537);
nand U11458 (N_11458,N_10138,N_10739);
and U11459 (N_11459,N_10843,N_10233);
nand U11460 (N_11460,N_10325,N_10133);
or U11461 (N_11461,N_10945,N_10235);
or U11462 (N_11462,N_10137,N_10528);
nand U11463 (N_11463,N_10448,N_10251);
nand U11464 (N_11464,N_10028,N_10436);
nand U11465 (N_11465,N_10297,N_10705);
xnor U11466 (N_11466,N_10719,N_10891);
and U11467 (N_11467,N_10957,N_10538);
and U11468 (N_11468,N_10590,N_10870);
or U11469 (N_11469,N_10342,N_10522);
and U11470 (N_11470,N_10864,N_10592);
nor U11471 (N_11471,N_10712,N_10118);
and U11472 (N_11472,N_10275,N_10327);
nor U11473 (N_11473,N_10748,N_10918);
nor U11474 (N_11474,N_10861,N_10475);
or U11475 (N_11475,N_10362,N_10802);
and U11476 (N_11476,N_10183,N_10310);
nor U11477 (N_11477,N_10878,N_10014);
and U11478 (N_11478,N_10047,N_10834);
xnor U11479 (N_11479,N_10596,N_10001);
and U11480 (N_11480,N_10304,N_10366);
or U11481 (N_11481,N_10252,N_10781);
nor U11482 (N_11482,N_10095,N_10972);
nand U11483 (N_11483,N_10892,N_10553);
nand U11484 (N_11484,N_10521,N_10214);
and U11485 (N_11485,N_10718,N_10791);
and U11486 (N_11486,N_10568,N_10851);
xor U11487 (N_11487,N_10484,N_10634);
nand U11488 (N_11488,N_10280,N_10881);
nand U11489 (N_11489,N_10465,N_10586);
xor U11490 (N_11490,N_10898,N_10502);
or U11491 (N_11491,N_10694,N_10965);
and U11492 (N_11492,N_10789,N_10533);
or U11493 (N_11493,N_10679,N_10283);
and U11494 (N_11494,N_10380,N_10354);
nand U11495 (N_11495,N_10239,N_10760);
and U11496 (N_11496,N_10182,N_10827);
nand U11497 (N_11497,N_10939,N_10935);
xor U11498 (N_11498,N_10913,N_10443);
and U11499 (N_11499,N_10474,N_10890);
or U11500 (N_11500,N_10471,N_10934);
nand U11501 (N_11501,N_10100,N_10697);
nor U11502 (N_11502,N_10131,N_10604);
nand U11503 (N_11503,N_10175,N_10567);
nand U11504 (N_11504,N_10225,N_10153);
xor U11505 (N_11505,N_10374,N_10835);
or U11506 (N_11506,N_10410,N_10758);
and U11507 (N_11507,N_10023,N_10625);
and U11508 (N_11508,N_10616,N_10056);
and U11509 (N_11509,N_10994,N_10797);
nor U11510 (N_11510,N_10828,N_10096);
and U11511 (N_11511,N_10464,N_10400);
and U11512 (N_11512,N_10558,N_10741);
nand U11513 (N_11513,N_10266,N_10348);
nand U11514 (N_11514,N_10427,N_10659);
and U11515 (N_11515,N_10891,N_10734);
xnor U11516 (N_11516,N_10973,N_10145);
xor U11517 (N_11517,N_10677,N_10890);
nor U11518 (N_11518,N_10295,N_10602);
or U11519 (N_11519,N_10442,N_10929);
nand U11520 (N_11520,N_10591,N_10492);
xor U11521 (N_11521,N_10001,N_10724);
and U11522 (N_11522,N_10001,N_10676);
nand U11523 (N_11523,N_10399,N_10044);
or U11524 (N_11524,N_10002,N_10847);
nand U11525 (N_11525,N_10256,N_10943);
xnor U11526 (N_11526,N_10814,N_10534);
or U11527 (N_11527,N_10340,N_10132);
nor U11528 (N_11528,N_10193,N_10125);
or U11529 (N_11529,N_10395,N_10525);
nand U11530 (N_11530,N_10687,N_10851);
nor U11531 (N_11531,N_10962,N_10202);
xor U11532 (N_11532,N_10891,N_10804);
xnor U11533 (N_11533,N_10001,N_10848);
and U11534 (N_11534,N_10247,N_10668);
or U11535 (N_11535,N_10688,N_10421);
nand U11536 (N_11536,N_10218,N_10403);
xor U11537 (N_11537,N_10843,N_10781);
and U11538 (N_11538,N_10723,N_10854);
and U11539 (N_11539,N_10057,N_10559);
nand U11540 (N_11540,N_10761,N_10368);
xnor U11541 (N_11541,N_10085,N_10076);
and U11542 (N_11542,N_10333,N_10019);
xnor U11543 (N_11543,N_10707,N_10664);
nand U11544 (N_11544,N_10714,N_10823);
xnor U11545 (N_11545,N_10383,N_10279);
or U11546 (N_11546,N_10501,N_10740);
nand U11547 (N_11547,N_10450,N_10806);
xnor U11548 (N_11548,N_10625,N_10804);
or U11549 (N_11549,N_10007,N_10732);
xnor U11550 (N_11550,N_10571,N_10727);
nor U11551 (N_11551,N_10395,N_10954);
nor U11552 (N_11552,N_10124,N_10838);
or U11553 (N_11553,N_10025,N_10874);
and U11554 (N_11554,N_10908,N_10149);
nor U11555 (N_11555,N_10009,N_10149);
nand U11556 (N_11556,N_10805,N_10201);
xor U11557 (N_11557,N_10058,N_10887);
nor U11558 (N_11558,N_10367,N_10192);
nor U11559 (N_11559,N_10248,N_10592);
xor U11560 (N_11560,N_10616,N_10165);
xnor U11561 (N_11561,N_10800,N_10356);
nor U11562 (N_11562,N_10601,N_10429);
nand U11563 (N_11563,N_10873,N_10860);
nand U11564 (N_11564,N_10402,N_10141);
xor U11565 (N_11565,N_10652,N_10599);
xnor U11566 (N_11566,N_10744,N_10313);
and U11567 (N_11567,N_10105,N_10666);
nor U11568 (N_11568,N_10849,N_10896);
xor U11569 (N_11569,N_10768,N_10531);
or U11570 (N_11570,N_10062,N_10725);
and U11571 (N_11571,N_10777,N_10118);
xor U11572 (N_11572,N_10932,N_10998);
nand U11573 (N_11573,N_10849,N_10674);
and U11574 (N_11574,N_10158,N_10153);
nor U11575 (N_11575,N_10594,N_10755);
or U11576 (N_11576,N_10336,N_10176);
or U11577 (N_11577,N_10075,N_10775);
or U11578 (N_11578,N_10200,N_10768);
nand U11579 (N_11579,N_10943,N_10761);
or U11580 (N_11580,N_10513,N_10445);
and U11581 (N_11581,N_10430,N_10406);
nand U11582 (N_11582,N_10459,N_10311);
or U11583 (N_11583,N_10348,N_10050);
xnor U11584 (N_11584,N_10142,N_10295);
or U11585 (N_11585,N_10513,N_10005);
nand U11586 (N_11586,N_10020,N_10233);
xnor U11587 (N_11587,N_10964,N_10353);
nand U11588 (N_11588,N_10350,N_10280);
xnor U11589 (N_11589,N_10110,N_10717);
or U11590 (N_11590,N_10826,N_10724);
nor U11591 (N_11591,N_10140,N_10465);
nor U11592 (N_11592,N_10255,N_10823);
nor U11593 (N_11593,N_10767,N_10105);
nand U11594 (N_11594,N_10344,N_10164);
or U11595 (N_11595,N_10155,N_10101);
nor U11596 (N_11596,N_10217,N_10382);
nor U11597 (N_11597,N_10961,N_10871);
and U11598 (N_11598,N_10523,N_10953);
or U11599 (N_11599,N_10330,N_10213);
xor U11600 (N_11600,N_10223,N_10454);
nand U11601 (N_11601,N_10620,N_10197);
xor U11602 (N_11602,N_10891,N_10042);
or U11603 (N_11603,N_10498,N_10066);
xor U11604 (N_11604,N_10666,N_10228);
nor U11605 (N_11605,N_10991,N_10587);
or U11606 (N_11606,N_10365,N_10174);
nand U11607 (N_11607,N_10760,N_10217);
nor U11608 (N_11608,N_10691,N_10708);
and U11609 (N_11609,N_10694,N_10671);
nor U11610 (N_11610,N_10814,N_10571);
or U11611 (N_11611,N_10843,N_10423);
nor U11612 (N_11612,N_10401,N_10510);
xor U11613 (N_11613,N_10739,N_10905);
and U11614 (N_11614,N_10865,N_10239);
and U11615 (N_11615,N_10007,N_10392);
and U11616 (N_11616,N_10326,N_10386);
nand U11617 (N_11617,N_10992,N_10436);
nand U11618 (N_11618,N_10386,N_10278);
or U11619 (N_11619,N_10568,N_10219);
xnor U11620 (N_11620,N_10116,N_10601);
and U11621 (N_11621,N_10557,N_10510);
xor U11622 (N_11622,N_10951,N_10081);
and U11623 (N_11623,N_10863,N_10267);
xor U11624 (N_11624,N_10968,N_10396);
xor U11625 (N_11625,N_10339,N_10770);
nor U11626 (N_11626,N_10462,N_10121);
and U11627 (N_11627,N_10399,N_10131);
or U11628 (N_11628,N_10695,N_10020);
or U11629 (N_11629,N_10575,N_10948);
nor U11630 (N_11630,N_10571,N_10802);
xor U11631 (N_11631,N_10564,N_10972);
and U11632 (N_11632,N_10157,N_10938);
nand U11633 (N_11633,N_10430,N_10193);
nor U11634 (N_11634,N_10139,N_10919);
and U11635 (N_11635,N_10563,N_10506);
nor U11636 (N_11636,N_10785,N_10593);
xnor U11637 (N_11637,N_10636,N_10243);
and U11638 (N_11638,N_10806,N_10068);
nor U11639 (N_11639,N_10056,N_10136);
nor U11640 (N_11640,N_10442,N_10922);
xor U11641 (N_11641,N_10308,N_10248);
and U11642 (N_11642,N_10621,N_10293);
xnor U11643 (N_11643,N_10778,N_10129);
xor U11644 (N_11644,N_10446,N_10732);
xnor U11645 (N_11645,N_10828,N_10636);
and U11646 (N_11646,N_10136,N_10327);
nand U11647 (N_11647,N_10240,N_10522);
xnor U11648 (N_11648,N_10268,N_10907);
and U11649 (N_11649,N_10198,N_10957);
and U11650 (N_11650,N_10019,N_10257);
xnor U11651 (N_11651,N_10364,N_10248);
and U11652 (N_11652,N_10384,N_10162);
nor U11653 (N_11653,N_10184,N_10900);
nor U11654 (N_11654,N_10444,N_10708);
or U11655 (N_11655,N_10507,N_10193);
nand U11656 (N_11656,N_10550,N_10036);
or U11657 (N_11657,N_10977,N_10857);
or U11658 (N_11658,N_10316,N_10602);
nor U11659 (N_11659,N_10775,N_10407);
or U11660 (N_11660,N_10963,N_10882);
and U11661 (N_11661,N_10440,N_10990);
and U11662 (N_11662,N_10722,N_10161);
or U11663 (N_11663,N_10440,N_10655);
and U11664 (N_11664,N_10530,N_10183);
nor U11665 (N_11665,N_10915,N_10694);
xor U11666 (N_11666,N_10246,N_10144);
or U11667 (N_11667,N_10830,N_10355);
or U11668 (N_11668,N_10583,N_10084);
nor U11669 (N_11669,N_10949,N_10289);
and U11670 (N_11670,N_10987,N_10334);
nor U11671 (N_11671,N_10399,N_10693);
or U11672 (N_11672,N_10365,N_10605);
nand U11673 (N_11673,N_10674,N_10054);
and U11674 (N_11674,N_10445,N_10825);
xor U11675 (N_11675,N_10620,N_10895);
nor U11676 (N_11676,N_10378,N_10801);
nor U11677 (N_11677,N_10002,N_10361);
xor U11678 (N_11678,N_10100,N_10438);
nand U11679 (N_11679,N_10294,N_10226);
nor U11680 (N_11680,N_10686,N_10024);
nand U11681 (N_11681,N_10407,N_10368);
xor U11682 (N_11682,N_10567,N_10785);
nor U11683 (N_11683,N_10452,N_10086);
nor U11684 (N_11684,N_10075,N_10474);
xor U11685 (N_11685,N_10452,N_10982);
xnor U11686 (N_11686,N_10735,N_10849);
or U11687 (N_11687,N_10544,N_10678);
or U11688 (N_11688,N_10009,N_10779);
or U11689 (N_11689,N_10314,N_10565);
nor U11690 (N_11690,N_10329,N_10981);
or U11691 (N_11691,N_10109,N_10481);
nand U11692 (N_11692,N_10578,N_10439);
and U11693 (N_11693,N_10593,N_10270);
or U11694 (N_11694,N_10160,N_10254);
xnor U11695 (N_11695,N_10388,N_10339);
and U11696 (N_11696,N_10245,N_10091);
nand U11697 (N_11697,N_10010,N_10492);
xor U11698 (N_11698,N_10049,N_10880);
nor U11699 (N_11699,N_10926,N_10426);
and U11700 (N_11700,N_10133,N_10022);
or U11701 (N_11701,N_10458,N_10652);
or U11702 (N_11702,N_10146,N_10139);
and U11703 (N_11703,N_10149,N_10763);
or U11704 (N_11704,N_10108,N_10348);
nand U11705 (N_11705,N_10420,N_10287);
or U11706 (N_11706,N_10528,N_10123);
nor U11707 (N_11707,N_10831,N_10676);
and U11708 (N_11708,N_10795,N_10033);
nand U11709 (N_11709,N_10804,N_10861);
nor U11710 (N_11710,N_10587,N_10307);
nor U11711 (N_11711,N_10951,N_10501);
nor U11712 (N_11712,N_10533,N_10785);
nor U11713 (N_11713,N_10637,N_10569);
nor U11714 (N_11714,N_10740,N_10777);
and U11715 (N_11715,N_10877,N_10489);
xor U11716 (N_11716,N_10522,N_10826);
nand U11717 (N_11717,N_10739,N_10780);
or U11718 (N_11718,N_10062,N_10264);
or U11719 (N_11719,N_10810,N_10326);
and U11720 (N_11720,N_10129,N_10565);
xnor U11721 (N_11721,N_10229,N_10303);
and U11722 (N_11722,N_10189,N_10833);
xor U11723 (N_11723,N_10034,N_10290);
nor U11724 (N_11724,N_10933,N_10071);
and U11725 (N_11725,N_10587,N_10224);
and U11726 (N_11726,N_10031,N_10689);
nor U11727 (N_11727,N_10431,N_10551);
or U11728 (N_11728,N_10989,N_10947);
nor U11729 (N_11729,N_10223,N_10996);
nor U11730 (N_11730,N_10374,N_10025);
or U11731 (N_11731,N_10404,N_10525);
nand U11732 (N_11732,N_10676,N_10079);
xor U11733 (N_11733,N_10284,N_10876);
or U11734 (N_11734,N_10051,N_10337);
and U11735 (N_11735,N_10867,N_10180);
nor U11736 (N_11736,N_10813,N_10279);
or U11737 (N_11737,N_10777,N_10628);
nand U11738 (N_11738,N_10665,N_10624);
or U11739 (N_11739,N_10343,N_10030);
nand U11740 (N_11740,N_10459,N_10392);
nand U11741 (N_11741,N_10171,N_10019);
or U11742 (N_11742,N_10443,N_10049);
nand U11743 (N_11743,N_10938,N_10849);
or U11744 (N_11744,N_10008,N_10370);
or U11745 (N_11745,N_10573,N_10749);
xnor U11746 (N_11746,N_10295,N_10403);
or U11747 (N_11747,N_10314,N_10962);
and U11748 (N_11748,N_10986,N_10477);
xnor U11749 (N_11749,N_10007,N_10695);
nor U11750 (N_11750,N_10594,N_10226);
nor U11751 (N_11751,N_10291,N_10651);
nand U11752 (N_11752,N_10138,N_10025);
or U11753 (N_11753,N_10891,N_10715);
nand U11754 (N_11754,N_10995,N_10065);
xnor U11755 (N_11755,N_10297,N_10129);
nor U11756 (N_11756,N_10716,N_10806);
and U11757 (N_11757,N_10500,N_10101);
xor U11758 (N_11758,N_10455,N_10791);
and U11759 (N_11759,N_10931,N_10934);
nand U11760 (N_11760,N_10995,N_10507);
xnor U11761 (N_11761,N_10206,N_10553);
nand U11762 (N_11762,N_10107,N_10724);
or U11763 (N_11763,N_10591,N_10392);
nand U11764 (N_11764,N_10042,N_10225);
nand U11765 (N_11765,N_10725,N_10902);
or U11766 (N_11766,N_10955,N_10731);
xor U11767 (N_11767,N_10429,N_10908);
xor U11768 (N_11768,N_10970,N_10319);
xor U11769 (N_11769,N_10032,N_10051);
and U11770 (N_11770,N_10065,N_10315);
nor U11771 (N_11771,N_10810,N_10197);
nand U11772 (N_11772,N_10635,N_10012);
nor U11773 (N_11773,N_10054,N_10236);
nand U11774 (N_11774,N_10850,N_10511);
xnor U11775 (N_11775,N_10724,N_10337);
or U11776 (N_11776,N_10181,N_10454);
and U11777 (N_11777,N_10557,N_10705);
nand U11778 (N_11778,N_10734,N_10391);
and U11779 (N_11779,N_10274,N_10060);
and U11780 (N_11780,N_10823,N_10758);
nand U11781 (N_11781,N_10681,N_10849);
or U11782 (N_11782,N_10503,N_10074);
and U11783 (N_11783,N_10048,N_10614);
or U11784 (N_11784,N_10780,N_10605);
nand U11785 (N_11785,N_10823,N_10225);
nor U11786 (N_11786,N_10903,N_10459);
and U11787 (N_11787,N_10759,N_10531);
xor U11788 (N_11788,N_10701,N_10367);
xnor U11789 (N_11789,N_10027,N_10898);
or U11790 (N_11790,N_10454,N_10241);
and U11791 (N_11791,N_10892,N_10785);
nand U11792 (N_11792,N_10753,N_10551);
nand U11793 (N_11793,N_10899,N_10449);
or U11794 (N_11794,N_10673,N_10126);
nand U11795 (N_11795,N_10761,N_10082);
or U11796 (N_11796,N_10206,N_10017);
nor U11797 (N_11797,N_10979,N_10060);
and U11798 (N_11798,N_10649,N_10302);
and U11799 (N_11799,N_10772,N_10979);
xor U11800 (N_11800,N_10883,N_10911);
xor U11801 (N_11801,N_10104,N_10918);
xnor U11802 (N_11802,N_10507,N_10151);
xnor U11803 (N_11803,N_10138,N_10987);
nor U11804 (N_11804,N_10337,N_10108);
xnor U11805 (N_11805,N_10611,N_10161);
or U11806 (N_11806,N_10708,N_10818);
or U11807 (N_11807,N_10863,N_10747);
nand U11808 (N_11808,N_10304,N_10830);
xnor U11809 (N_11809,N_10627,N_10341);
and U11810 (N_11810,N_10969,N_10456);
or U11811 (N_11811,N_10067,N_10555);
or U11812 (N_11812,N_10716,N_10197);
nand U11813 (N_11813,N_10065,N_10904);
nand U11814 (N_11814,N_10042,N_10169);
or U11815 (N_11815,N_10590,N_10610);
xnor U11816 (N_11816,N_10150,N_10324);
or U11817 (N_11817,N_10249,N_10580);
nor U11818 (N_11818,N_10373,N_10855);
nor U11819 (N_11819,N_10585,N_10668);
or U11820 (N_11820,N_10078,N_10759);
xnor U11821 (N_11821,N_10384,N_10761);
nor U11822 (N_11822,N_10182,N_10778);
nor U11823 (N_11823,N_10380,N_10897);
nand U11824 (N_11824,N_10783,N_10919);
and U11825 (N_11825,N_10324,N_10358);
nand U11826 (N_11826,N_10376,N_10203);
nor U11827 (N_11827,N_10164,N_10072);
and U11828 (N_11828,N_10134,N_10139);
and U11829 (N_11829,N_10681,N_10310);
nor U11830 (N_11830,N_10610,N_10531);
nor U11831 (N_11831,N_10515,N_10468);
xnor U11832 (N_11832,N_10457,N_10144);
and U11833 (N_11833,N_10678,N_10748);
nand U11834 (N_11834,N_10171,N_10239);
xor U11835 (N_11835,N_10534,N_10845);
and U11836 (N_11836,N_10078,N_10409);
nand U11837 (N_11837,N_10112,N_10612);
nor U11838 (N_11838,N_10658,N_10791);
nor U11839 (N_11839,N_10350,N_10950);
nand U11840 (N_11840,N_10151,N_10269);
and U11841 (N_11841,N_10907,N_10010);
nand U11842 (N_11842,N_10853,N_10181);
nand U11843 (N_11843,N_10998,N_10999);
nand U11844 (N_11844,N_10866,N_10869);
or U11845 (N_11845,N_10805,N_10812);
or U11846 (N_11846,N_10344,N_10118);
nor U11847 (N_11847,N_10271,N_10531);
or U11848 (N_11848,N_10244,N_10547);
and U11849 (N_11849,N_10636,N_10940);
xnor U11850 (N_11850,N_10410,N_10549);
or U11851 (N_11851,N_10330,N_10730);
xnor U11852 (N_11852,N_10255,N_10017);
nand U11853 (N_11853,N_10850,N_10193);
or U11854 (N_11854,N_10053,N_10477);
nor U11855 (N_11855,N_10676,N_10455);
xnor U11856 (N_11856,N_10603,N_10412);
and U11857 (N_11857,N_10026,N_10695);
nor U11858 (N_11858,N_10650,N_10032);
nor U11859 (N_11859,N_10139,N_10137);
nor U11860 (N_11860,N_10004,N_10989);
nand U11861 (N_11861,N_10612,N_10403);
nor U11862 (N_11862,N_10678,N_10448);
nor U11863 (N_11863,N_10365,N_10841);
and U11864 (N_11864,N_10457,N_10861);
nand U11865 (N_11865,N_10446,N_10731);
and U11866 (N_11866,N_10532,N_10217);
nor U11867 (N_11867,N_10402,N_10473);
or U11868 (N_11868,N_10453,N_10021);
nor U11869 (N_11869,N_10827,N_10768);
nand U11870 (N_11870,N_10689,N_10824);
or U11871 (N_11871,N_10686,N_10477);
nand U11872 (N_11872,N_10234,N_10572);
nor U11873 (N_11873,N_10777,N_10211);
nand U11874 (N_11874,N_10568,N_10459);
nand U11875 (N_11875,N_10771,N_10894);
nand U11876 (N_11876,N_10530,N_10490);
nor U11877 (N_11877,N_10622,N_10463);
and U11878 (N_11878,N_10032,N_10835);
or U11879 (N_11879,N_10916,N_10997);
or U11880 (N_11880,N_10903,N_10715);
xor U11881 (N_11881,N_10431,N_10029);
xor U11882 (N_11882,N_10679,N_10144);
xnor U11883 (N_11883,N_10963,N_10210);
xor U11884 (N_11884,N_10693,N_10592);
xnor U11885 (N_11885,N_10495,N_10614);
or U11886 (N_11886,N_10115,N_10412);
or U11887 (N_11887,N_10166,N_10845);
and U11888 (N_11888,N_10684,N_10418);
nor U11889 (N_11889,N_10041,N_10085);
xnor U11890 (N_11890,N_10719,N_10790);
nor U11891 (N_11891,N_10876,N_10902);
or U11892 (N_11892,N_10560,N_10090);
xor U11893 (N_11893,N_10306,N_10330);
and U11894 (N_11894,N_10394,N_10438);
nor U11895 (N_11895,N_10195,N_10936);
and U11896 (N_11896,N_10365,N_10303);
nor U11897 (N_11897,N_10598,N_10257);
nor U11898 (N_11898,N_10331,N_10897);
xor U11899 (N_11899,N_10292,N_10464);
xor U11900 (N_11900,N_10584,N_10177);
nand U11901 (N_11901,N_10250,N_10040);
or U11902 (N_11902,N_10055,N_10866);
nor U11903 (N_11903,N_10113,N_10017);
nor U11904 (N_11904,N_10761,N_10772);
nor U11905 (N_11905,N_10625,N_10121);
nand U11906 (N_11906,N_10917,N_10715);
and U11907 (N_11907,N_10292,N_10645);
or U11908 (N_11908,N_10627,N_10498);
xnor U11909 (N_11909,N_10093,N_10836);
or U11910 (N_11910,N_10852,N_10583);
and U11911 (N_11911,N_10016,N_10050);
nor U11912 (N_11912,N_10266,N_10029);
xnor U11913 (N_11913,N_10886,N_10512);
or U11914 (N_11914,N_10246,N_10941);
or U11915 (N_11915,N_10594,N_10308);
and U11916 (N_11916,N_10892,N_10706);
nor U11917 (N_11917,N_10805,N_10106);
xor U11918 (N_11918,N_10082,N_10655);
or U11919 (N_11919,N_10011,N_10411);
and U11920 (N_11920,N_10646,N_10522);
xor U11921 (N_11921,N_10765,N_10207);
nand U11922 (N_11922,N_10754,N_10946);
or U11923 (N_11923,N_10176,N_10753);
xnor U11924 (N_11924,N_10765,N_10656);
and U11925 (N_11925,N_10722,N_10901);
nand U11926 (N_11926,N_10559,N_10802);
and U11927 (N_11927,N_10019,N_10206);
xor U11928 (N_11928,N_10818,N_10568);
nand U11929 (N_11929,N_10892,N_10671);
xnor U11930 (N_11930,N_10257,N_10811);
and U11931 (N_11931,N_10172,N_10134);
xor U11932 (N_11932,N_10457,N_10524);
or U11933 (N_11933,N_10646,N_10592);
or U11934 (N_11934,N_10992,N_10408);
xnor U11935 (N_11935,N_10437,N_10122);
or U11936 (N_11936,N_10060,N_10653);
nor U11937 (N_11937,N_10140,N_10215);
nor U11938 (N_11938,N_10580,N_10377);
and U11939 (N_11939,N_10217,N_10718);
nand U11940 (N_11940,N_10988,N_10584);
nand U11941 (N_11941,N_10409,N_10259);
nor U11942 (N_11942,N_10456,N_10343);
or U11943 (N_11943,N_10149,N_10370);
nand U11944 (N_11944,N_10359,N_10443);
nand U11945 (N_11945,N_10159,N_10796);
nand U11946 (N_11946,N_10375,N_10775);
xor U11947 (N_11947,N_10914,N_10748);
nor U11948 (N_11948,N_10023,N_10816);
xnor U11949 (N_11949,N_10775,N_10122);
and U11950 (N_11950,N_10847,N_10742);
and U11951 (N_11951,N_10342,N_10040);
or U11952 (N_11952,N_10194,N_10715);
nor U11953 (N_11953,N_10808,N_10057);
nand U11954 (N_11954,N_10237,N_10501);
nand U11955 (N_11955,N_10617,N_10220);
nand U11956 (N_11956,N_10409,N_10188);
and U11957 (N_11957,N_10643,N_10770);
xor U11958 (N_11958,N_10114,N_10342);
xor U11959 (N_11959,N_10354,N_10920);
nand U11960 (N_11960,N_10885,N_10902);
or U11961 (N_11961,N_10370,N_10885);
nor U11962 (N_11962,N_10506,N_10178);
xnor U11963 (N_11963,N_10655,N_10827);
and U11964 (N_11964,N_10097,N_10435);
xor U11965 (N_11965,N_10624,N_10130);
and U11966 (N_11966,N_10284,N_10340);
nor U11967 (N_11967,N_10066,N_10994);
or U11968 (N_11968,N_10590,N_10810);
and U11969 (N_11969,N_10512,N_10755);
xnor U11970 (N_11970,N_10741,N_10972);
xnor U11971 (N_11971,N_10079,N_10490);
nor U11972 (N_11972,N_10489,N_10324);
nor U11973 (N_11973,N_10521,N_10145);
and U11974 (N_11974,N_10917,N_10598);
nor U11975 (N_11975,N_10123,N_10605);
nor U11976 (N_11976,N_10076,N_10500);
nor U11977 (N_11977,N_10719,N_10020);
or U11978 (N_11978,N_10514,N_10359);
and U11979 (N_11979,N_10592,N_10093);
or U11980 (N_11980,N_10630,N_10055);
xor U11981 (N_11981,N_10624,N_10753);
and U11982 (N_11982,N_10970,N_10020);
nor U11983 (N_11983,N_10153,N_10976);
nand U11984 (N_11984,N_10121,N_10764);
xnor U11985 (N_11985,N_10448,N_10077);
and U11986 (N_11986,N_10742,N_10669);
and U11987 (N_11987,N_10096,N_10347);
and U11988 (N_11988,N_10489,N_10323);
xnor U11989 (N_11989,N_10319,N_10375);
xnor U11990 (N_11990,N_10825,N_10644);
xor U11991 (N_11991,N_10849,N_10605);
and U11992 (N_11992,N_10242,N_10883);
xor U11993 (N_11993,N_10038,N_10487);
and U11994 (N_11994,N_10894,N_10316);
nand U11995 (N_11995,N_10557,N_10091);
and U11996 (N_11996,N_10184,N_10141);
nor U11997 (N_11997,N_10304,N_10696);
or U11998 (N_11998,N_10881,N_10686);
nand U11999 (N_11999,N_10362,N_10381);
nor U12000 (N_12000,N_11031,N_11956);
xnor U12001 (N_12001,N_11378,N_11477);
xnor U12002 (N_12002,N_11740,N_11311);
xnor U12003 (N_12003,N_11738,N_11763);
or U12004 (N_12004,N_11504,N_11985);
or U12005 (N_12005,N_11360,N_11458);
nand U12006 (N_12006,N_11082,N_11330);
nand U12007 (N_12007,N_11780,N_11196);
nand U12008 (N_12008,N_11578,N_11306);
or U12009 (N_12009,N_11284,N_11423);
nand U12010 (N_12010,N_11735,N_11960);
nor U12011 (N_12011,N_11747,N_11524);
nor U12012 (N_12012,N_11730,N_11705);
nand U12013 (N_12013,N_11745,N_11255);
nor U12014 (N_12014,N_11115,N_11681);
xnor U12015 (N_12015,N_11077,N_11123);
nand U12016 (N_12016,N_11021,N_11023);
xnor U12017 (N_12017,N_11512,N_11973);
nor U12018 (N_12018,N_11538,N_11979);
nor U12019 (N_12019,N_11888,N_11913);
nor U12020 (N_12020,N_11319,N_11907);
and U12021 (N_12021,N_11584,N_11204);
or U12022 (N_12022,N_11310,N_11739);
or U12023 (N_12023,N_11700,N_11778);
or U12024 (N_12024,N_11962,N_11889);
xnor U12025 (N_12025,N_11006,N_11808);
or U12026 (N_12026,N_11500,N_11384);
or U12027 (N_12027,N_11851,N_11085);
nand U12028 (N_12028,N_11975,N_11124);
xnor U12029 (N_12029,N_11569,N_11086);
or U12030 (N_12030,N_11722,N_11886);
nand U12031 (N_12031,N_11874,N_11797);
or U12032 (N_12032,N_11998,N_11663);
nor U12033 (N_12033,N_11025,N_11243);
and U12034 (N_12034,N_11020,N_11698);
or U12035 (N_12035,N_11048,N_11910);
and U12036 (N_12036,N_11993,N_11265);
or U12037 (N_12037,N_11782,N_11826);
and U12038 (N_12038,N_11142,N_11665);
xor U12039 (N_12039,N_11566,N_11228);
and U12040 (N_12040,N_11746,N_11001);
nor U12041 (N_12041,N_11338,N_11097);
nand U12042 (N_12042,N_11644,N_11661);
nor U12043 (N_12043,N_11550,N_11211);
nand U12044 (N_12044,N_11534,N_11028);
nand U12045 (N_12045,N_11220,N_11218);
or U12046 (N_12046,N_11003,N_11453);
nand U12047 (N_12047,N_11468,N_11564);
nand U12048 (N_12048,N_11685,N_11260);
or U12049 (N_12049,N_11729,N_11995);
nor U12050 (N_12050,N_11125,N_11779);
nor U12051 (N_12051,N_11672,N_11891);
xnor U12052 (N_12052,N_11965,N_11688);
xor U12053 (N_12053,N_11827,N_11883);
or U12054 (N_12054,N_11143,N_11164);
and U12055 (N_12055,N_11075,N_11475);
or U12056 (N_12056,N_11622,N_11425);
nand U12057 (N_12057,N_11497,N_11377);
xnor U12058 (N_12058,N_11406,N_11270);
or U12059 (N_12059,N_11596,N_11288);
and U12060 (N_12060,N_11600,N_11420);
or U12061 (N_12061,N_11172,N_11620);
nand U12062 (N_12062,N_11022,N_11556);
xnor U12063 (N_12063,N_11083,N_11103);
and U12064 (N_12064,N_11060,N_11868);
xnor U12065 (N_12065,N_11855,N_11011);
nor U12066 (N_12066,N_11929,N_11442);
and U12067 (N_12067,N_11231,N_11343);
nand U12068 (N_12068,N_11232,N_11182);
xor U12069 (N_12069,N_11947,N_11293);
nor U12070 (N_12070,N_11754,N_11119);
xnor U12071 (N_12071,N_11731,N_11503);
nand U12072 (N_12072,N_11071,N_11176);
nand U12073 (N_12073,N_11836,N_11224);
nand U12074 (N_12074,N_11638,N_11005);
nor U12075 (N_12075,N_11169,N_11852);
xnor U12076 (N_12076,N_11771,N_11667);
nand U12077 (N_12077,N_11752,N_11461);
nor U12078 (N_12078,N_11187,N_11253);
xnor U12079 (N_12079,N_11056,N_11290);
and U12080 (N_12080,N_11530,N_11004);
nor U12081 (N_12081,N_11646,N_11273);
xnor U12082 (N_12082,N_11967,N_11794);
nor U12083 (N_12083,N_11767,N_11699);
xor U12084 (N_12084,N_11470,N_11058);
xor U12085 (N_12085,N_11183,N_11893);
nor U12086 (N_12086,N_11203,N_11146);
nand U12087 (N_12087,N_11510,N_11828);
xor U12088 (N_12088,N_11340,N_11178);
xnor U12089 (N_12089,N_11509,N_11536);
xnor U12090 (N_12090,N_11271,N_11400);
xnor U12091 (N_12091,N_11895,N_11350);
or U12092 (N_12092,N_11236,N_11331);
and U12093 (N_12093,N_11549,N_11925);
or U12094 (N_12094,N_11456,N_11894);
nor U12095 (N_12095,N_11132,N_11519);
nor U12096 (N_12096,N_11944,N_11079);
or U12097 (N_12097,N_11065,N_11820);
xnor U12098 (N_12098,N_11171,N_11399);
or U12099 (N_12099,N_11501,N_11155);
nor U12100 (N_12100,N_11434,N_11626);
xor U12101 (N_12101,N_11026,N_11133);
or U12102 (N_12102,N_11084,N_11815);
or U12103 (N_12103,N_11440,N_11842);
or U12104 (N_12104,N_11508,N_11354);
or U12105 (N_12105,N_11368,N_11007);
and U12106 (N_12106,N_11990,N_11315);
nand U12107 (N_12107,N_11351,N_11678);
xor U12108 (N_12108,N_11958,N_11099);
xor U12109 (N_12109,N_11034,N_11230);
and U12110 (N_12110,N_11019,N_11559);
or U12111 (N_12111,N_11674,N_11721);
nor U12112 (N_12112,N_11609,N_11843);
nor U12113 (N_12113,N_11135,N_11636);
xor U12114 (N_12114,N_11690,N_11267);
nor U12115 (N_12115,N_11447,N_11599);
xnor U12116 (N_12116,N_11612,N_11551);
xor U12117 (N_12117,N_11094,N_11717);
xor U12118 (N_12118,N_11691,N_11353);
or U12119 (N_12119,N_11937,N_11884);
xor U12120 (N_12120,N_11489,N_11844);
and U12121 (N_12121,N_11777,N_11408);
nor U12122 (N_12122,N_11972,N_11585);
nand U12123 (N_12123,N_11106,N_11159);
nor U12124 (N_12124,N_11128,N_11571);
or U12125 (N_12125,N_11055,N_11981);
and U12126 (N_12126,N_11484,N_11292);
xor U12127 (N_12127,N_11824,N_11069);
xor U12128 (N_12128,N_11464,N_11113);
or U12129 (N_12129,N_11445,N_11249);
nand U12130 (N_12130,N_11539,N_11526);
nor U12131 (N_12131,N_11673,N_11364);
and U12132 (N_12132,N_11162,N_11093);
nor U12133 (N_12133,N_11064,N_11225);
and U12134 (N_12134,N_11810,N_11396);
nor U12135 (N_12135,N_11591,N_11219);
and U12136 (N_12136,N_11733,N_11529);
xnor U12137 (N_12137,N_11819,N_11194);
and U12138 (N_12138,N_11753,N_11185);
nand U12139 (N_12139,N_11649,N_11713);
nand U12140 (N_12140,N_11511,N_11344);
xor U12141 (N_12141,N_11057,N_11522);
or U12142 (N_12142,N_11502,N_11439);
or U12143 (N_12143,N_11710,N_11269);
or U12144 (N_12144,N_11562,N_11383);
or U12145 (N_12145,N_11275,N_11983);
nand U12146 (N_12146,N_11321,N_11516);
xnor U12147 (N_12147,N_11297,N_11567);
xnor U12148 (N_12148,N_11853,N_11602);
and U12149 (N_12149,N_11210,N_11948);
and U12150 (N_12150,N_11848,N_11553);
nand U12151 (N_12151,N_11773,N_11333);
xnor U12152 (N_12152,N_11216,N_11309);
nand U12153 (N_12153,N_11117,N_11481);
nor U12154 (N_12154,N_11168,N_11296);
and U12155 (N_12155,N_11866,N_11165);
nand U12156 (N_12156,N_11490,N_11643);
or U12157 (N_12157,N_11433,N_11581);
or U12158 (N_12158,N_11882,N_11601);
and U12159 (N_12159,N_11463,N_11558);
or U12160 (N_12160,N_11573,N_11801);
or U12161 (N_12161,N_11281,N_11443);
nor U12162 (N_12162,N_11769,N_11109);
and U12163 (N_12163,N_11614,N_11095);
nand U12164 (N_12164,N_11968,N_11587);
nor U12165 (N_12165,N_11438,N_11316);
nor U12166 (N_12166,N_11802,N_11561);
and U12167 (N_12167,N_11467,N_11372);
or U12168 (N_12168,N_11978,N_11719);
nand U12169 (N_12169,N_11630,N_11786);
and U12170 (N_12170,N_11419,N_11637);
nor U12171 (N_12171,N_11362,N_11394);
nor U12172 (N_12172,N_11525,N_11544);
xnor U12173 (N_12173,N_11042,N_11588);
xor U12174 (N_12174,N_11335,N_11098);
nand U12175 (N_12175,N_11254,N_11590);
nor U12176 (N_12176,N_11061,N_11865);
and U12177 (N_12177,N_11989,N_11954);
and U12178 (N_12178,N_11625,N_11088);
nand U12179 (N_12179,N_11762,N_11613);
and U12180 (N_12180,N_11302,N_11137);
or U12181 (N_12181,N_11352,N_11565);
or U12182 (N_12182,N_11469,N_11078);
and U12183 (N_12183,N_11361,N_11715);
nor U12184 (N_12184,N_11336,N_11633);
nand U12185 (N_12185,N_11862,N_11671);
xor U12186 (N_12186,N_11935,N_11675);
nor U12187 (N_12187,N_11970,N_11543);
nor U12188 (N_12188,N_11493,N_11939);
xor U12189 (N_12189,N_11422,N_11984);
or U12190 (N_12190,N_11341,N_11540);
nor U12191 (N_12191,N_11669,N_11631);
and U12192 (N_12192,N_11732,N_11592);
nand U12193 (N_12193,N_11473,N_11560);
and U12194 (N_12194,N_11045,N_11193);
nor U12195 (N_12195,N_11043,N_11010);
and U12196 (N_12196,N_11314,N_11287);
or U12197 (N_12197,N_11918,N_11190);
xor U12198 (N_12198,N_11724,N_11547);
xor U12199 (N_12199,N_11689,N_11009);
nand U12200 (N_12200,N_11148,N_11217);
and U12201 (N_12201,N_11506,N_11157);
nand U12202 (N_12202,N_11834,N_11505);
or U12203 (N_12203,N_11282,N_11881);
nand U12204 (N_12204,N_11312,N_11385);
or U12205 (N_12205,N_11476,N_11652);
nor U12206 (N_12206,N_11908,N_11520);
nor U12207 (N_12207,N_11024,N_11161);
nand U12208 (N_12208,N_11850,N_11904);
or U12209 (N_12209,N_11897,N_11900);
or U12210 (N_12210,N_11285,N_11527);
nand U12211 (N_12211,N_11393,N_11847);
or U12212 (N_12212,N_11240,N_11403);
nand U12213 (N_12213,N_11381,N_11821);
nand U12214 (N_12214,N_11427,N_11572);
and U12215 (N_12215,N_11101,N_11370);
or U12216 (N_12216,N_11658,N_11655);
nand U12217 (N_12217,N_11140,N_11577);
or U12218 (N_12218,N_11632,N_11846);
nand U12219 (N_12219,N_11479,N_11666);
nand U12220 (N_12220,N_11931,N_11814);
and U12221 (N_12221,N_11062,N_11971);
and U12222 (N_12222,N_11709,N_11790);
or U12223 (N_12223,N_11987,N_11038);
xor U12224 (N_12224,N_11415,N_11213);
nand U12225 (N_12225,N_11407,N_11090);
or U12226 (N_12226,N_11059,N_11728);
nor U12227 (N_12227,N_11914,N_11879);
nand U12228 (N_12228,N_11387,N_11076);
xnor U12229 (N_12229,N_11934,N_11483);
xnor U12230 (N_12230,N_11327,N_11205);
xor U12231 (N_12231,N_11430,N_11300);
nand U12232 (N_12232,N_11180,N_11744);
nand U12233 (N_12233,N_11037,N_11706);
and U12234 (N_12234,N_11320,N_11092);
nand U12235 (N_12235,N_11455,N_11405);
nand U12236 (N_12236,N_11039,N_11154);
nand U12237 (N_12237,N_11365,N_11857);
or U12238 (N_12238,N_11545,N_11864);
nand U12239 (N_12239,N_11197,N_11743);
or U12240 (N_12240,N_11212,N_11390);
or U12241 (N_12241,N_11936,N_11029);
nor U12242 (N_12242,N_11807,N_11460);
nor U12243 (N_12243,N_11261,N_11653);
and U12244 (N_12244,N_11849,N_11208);
or U12245 (N_12245,N_11869,N_11334);
or U12246 (N_12246,N_11299,N_11959);
nor U12247 (N_12247,N_11391,N_11957);
or U12248 (N_12248,N_11694,N_11478);
xnor U12249 (N_12249,N_11923,N_11920);
xnor U12250 (N_12250,N_11662,N_11980);
nor U12251 (N_12251,N_11604,N_11809);
xnor U12252 (N_12252,N_11933,N_11811);
and U12253 (N_12253,N_11768,N_11494);
nand U12254 (N_12254,N_11416,N_11648);
nor U12255 (N_12255,N_11756,N_11992);
and U12256 (N_12256,N_11452,N_11668);
xnor U12257 (N_12257,N_11829,N_11774);
or U12258 (N_12258,N_11791,N_11051);
xor U12259 (N_12259,N_11521,N_11757);
and U12260 (N_12260,N_11872,N_11887);
or U12261 (N_12261,N_11835,N_11186);
and U12262 (N_12262,N_11635,N_11242);
xnor U12263 (N_12263,N_11431,N_11091);
and U12264 (N_12264,N_11696,N_11451);
nand U12265 (N_12265,N_11389,N_11053);
xnor U12266 (N_12266,N_11823,N_11147);
and U12267 (N_12267,N_11418,N_11191);
nand U12268 (N_12268,N_11603,N_11693);
and U12269 (N_12269,N_11486,N_11676);
or U12270 (N_12270,N_11170,N_11942);
and U12271 (N_12271,N_11775,N_11533);
and U12272 (N_12272,N_11660,N_11474);
nor U12273 (N_12273,N_11301,N_11324);
xnor U12274 (N_12274,N_11426,N_11153);
nor U12275 (N_12275,N_11495,N_11656);
nand U12276 (N_12276,N_11692,N_11044);
nand U12277 (N_12277,N_11030,N_11040);
nand U12278 (N_12278,N_11174,N_11804);
xor U12279 (N_12279,N_11226,N_11749);
nand U12280 (N_12280,N_11244,N_11683);
xnor U12281 (N_12281,N_11491,N_11582);
and U12282 (N_12282,N_11748,N_11594);
nand U12283 (N_12283,N_11272,N_11304);
or U12284 (N_12284,N_11742,N_11050);
nor U12285 (N_12285,N_11152,N_11195);
xor U12286 (N_12286,N_11465,N_11912);
and U12287 (N_12287,N_11818,N_11949);
nor U12288 (N_12288,N_11803,N_11876);
xor U12289 (N_12289,N_11200,N_11008);
and U12290 (N_12290,N_11120,N_11554);
and U12291 (N_12291,N_11812,N_11969);
or U12292 (N_12292,N_11513,N_11018);
xnor U12293 (N_12293,N_11395,N_11121);
or U12294 (N_12294,N_11623,N_11974);
xnor U12295 (N_12295,N_11404,N_11515);
nor U12296 (N_12296,N_11682,N_11122);
and U12297 (N_12297,N_11448,N_11861);
and U12298 (N_12298,N_11898,N_11016);
xor U12299 (N_12299,N_11239,N_11496);
and U12300 (N_12300,N_11664,N_11369);
or U12301 (N_12301,N_11347,N_11758);
nor U12302 (N_12302,N_11449,N_11118);
nor U12303 (N_12303,N_11063,N_11928);
xor U12304 (N_12304,N_11245,N_11707);
nand U12305 (N_12305,N_11107,N_11997);
nand U12306 (N_12306,N_11878,N_11645);
and U12307 (N_12307,N_11392,N_11313);
nor U12308 (N_12308,N_11988,N_11607);
xor U12309 (N_12309,N_11875,N_11175);
and U12310 (N_12310,N_11295,N_11902);
nor U12311 (N_12311,N_11617,N_11563);
nand U12312 (N_12312,N_11574,N_11346);
or U12313 (N_12313,N_11687,N_11555);
or U12314 (N_12314,N_11570,N_11237);
or U12315 (N_12315,N_11289,N_11579);
nand U12316 (N_12316,N_11332,N_11776);
or U12317 (N_12317,N_11677,N_11339);
xnor U12318 (N_12318,N_11318,N_11257);
and U12319 (N_12319,N_11785,N_11799);
nand U12320 (N_12320,N_11518,N_11150);
nor U12321 (N_12321,N_11279,N_11052);
xor U12322 (N_12322,N_11201,N_11532);
nand U12323 (N_12323,N_11256,N_11736);
xor U12324 (N_12324,N_11627,N_11624);
xor U12325 (N_12325,N_11945,N_11414);
xnor U12326 (N_12326,N_11189,N_11386);
xor U12327 (N_12327,N_11568,N_11615);
or U12328 (N_12328,N_11890,N_11375);
nor U12329 (N_12329,N_11013,N_11116);
or U12330 (N_12330,N_11618,N_11999);
xnor U12331 (N_12331,N_11033,N_11839);
and U12332 (N_12332,N_11789,N_11922);
nand U12333 (N_12333,N_11342,N_11184);
nor U12334 (N_12334,N_11382,N_11946);
or U12335 (N_12335,N_11374,N_11634);
and U12336 (N_12336,N_11488,N_11940);
and U12337 (N_12337,N_11163,N_11723);
or U12338 (N_12338,N_11130,N_11134);
nor U12339 (N_12339,N_11877,N_11996);
nand U12340 (N_12340,N_11517,N_11358);
or U12341 (N_12341,N_11840,N_11457);
or U12342 (N_12342,N_11616,N_11411);
nor U12343 (N_12343,N_11294,N_11198);
and U12344 (N_12344,N_11552,N_11428);
or U12345 (N_12345,N_11982,N_11199);
nand U12346 (N_12346,N_11366,N_11348);
and U12347 (N_12347,N_11054,N_11081);
xnor U12348 (N_12348,N_11177,N_11074);
or U12349 (N_12349,N_11277,N_11961);
or U12350 (N_12350,N_11325,N_11017);
nor U12351 (N_12351,N_11480,N_11298);
or U12352 (N_12352,N_11867,N_11950);
nor U12353 (N_12353,N_11535,N_11067);
xor U12354 (N_12354,N_11697,N_11783);
xor U12355 (N_12355,N_11233,N_11087);
or U12356 (N_12356,N_11498,N_11266);
and U12357 (N_12357,N_11472,N_11714);
nand U12358 (N_12358,N_11932,N_11976);
nor U12359 (N_12359,N_11138,N_11830);
xor U12360 (N_12360,N_11576,N_11305);
or U12361 (N_12361,N_11307,N_11379);
nor U12362 (N_12362,N_11605,N_11167);
nor U12363 (N_12363,N_11432,N_11557);
or U12364 (N_12364,N_11126,N_11859);
or U12365 (N_12365,N_11583,N_11703);
and U12366 (N_12366,N_11214,N_11854);
and U12367 (N_12367,N_11450,N_11207);
nand U12368 (N_12368,N_11800,N_11640);
and U12369 (N_12369,N_11308,N_11899);
nand U12370 (N_12370,N_11924,N_11816);
or U12371 (N_12371,N_11755,N_11611);
xor U12372 (N_12372,N_11892,N_11049);
nand U12373 (N_12373,N_11328,N_11838);
nand U12374 (N_12374,N_11421,N_11337);
nand U12375 (N_12375,N_11072,N_11047);
and U12376 (N_12376,N_11514,N_11188);
or U12377 (N_12377,N_11291,N_11485);
xor U12378 (N_12378,N_11014,N_11542);
nor U12379 (N_12379,N_11329,N_11817);
and U12380 (N_12380,N_11227,N_11371);
nor U12381 (N_12381,N_11238,N_11955);
nand U12382 (N_12382,N_11909,N_11482);
nor U12383 (N_12383,N_11994,N_11258);
or U12384 (N_12384,N_11750,N_11679);
or U12385 (N_12385,N_11725,N_11398);
and U12386 (N_12386,N_11259,N_11454);
nand U12387 (N_12387,N_11856,N_11487);
or U12388 (N_12388,N_11492,N_11252);
and U12389 (N_12389,N_11606,N_11248);
or U12390 (N_12390,N_11102,N_11651);
nand U12391 (N_12391,N_11073,N_11435);
nand U12392 (N_12392,N_11951,N_11160);
and U12393 (N_12393,N_11066,N_11792);
or U12394 (N_12394,N_11129,N_11278);
and U12395 (N_12395,N_11206,N_11772);
or U12396 (N_12396,N_11359,N_11127);
and U12397 (N_12397,N_11111,N_11659);
nor U12398 (N_12398,N_11112,N_11356);
and U12399 (N_12399,N_11684,N_11952);
or U12400 (N_12400,N_11917,N_11471);
xnor U12401 (N_12401,N_11642,N_11446);
and U12402 (N_12402,N_11250,N_11926);
nor U12403 (N_12403,N_11149,N_11032);
or U12404 (N_12404,N_11537,N_11268);
and U12405 (N_12405,N_11144,N_11795);
nor U12406 (N_12406,N_11586,N_11264);
nand U12407 (N_12407,N_11376,N_11100);
nand U12408 (N_12408,N_11873,N_11041);
nor U12409 (N_12409,N_11104,N_11179);
and U12410 (N_12410,N_11303,N_11858);
and U12411 (N_12411,N_11765,N_11734);
xor U12412 (N_12412,N_11680,N_11380);
xor U12413 (N_12413,N_11905,N_11546);
nor U12414 (N_12414,N_11650,N_11880);
xnor U12415 (N_12415,N_11412,N_11720);
and U12416 (N_12416,N_11927,N_11708);
nor U12417 (N_12417,N_11263,N_11388);
xor U12418 (N_12418,N_11209,N_11367);
nand U12419 (N_12419,N_11871,N_11145);
nor U12420 (N_12420,N_11915,N_11941);
and U12421 (N_12421,N_11241,N_11760);
nor U12422 (N_12422,N_11963,N_11202);
or U12423 (N_12423,N_11046,N_11089);
nand U12424 (N_12424,N_11991,N_11695);
or U12425 (N_12425,N_11441,N_11276);
xnor U12426 (N_12426,N_11741,N_11896);
nand U12427 (N_12427,N_11528,N_11373);
and U12428 (N_12428,N_11788,N_11608);
xnor U12429 (N_12429,N_11286,N_11466);
or U12430 (N_12430,N_11110,N_11507);
nand U12431 (N_12431,N_11322,N_11413);
and U12432 (N_12432,N_11357,N_11628);
nor U12433 (N_12433,N_11531,N_11262);
nand U12434 (N_12434,N_11911,N_11841);
and U12435 (N_12435,N_11787,N_11580);
or U12436 (N_12436,N_11349,N_11424);
nand U12437 (N_12437,N_11247,N_11919);
or U12438 (N_12438,N_11712,N_11727);
nand U12439 (N_12439,N_11444,N_11657);
or U12440 (N_12440,N_11136,N_11686);
or U12441 (N_12441,N_11108,N_11813);
and U12442 (N_12442,N_11761,N_11610);
nor U12443 (N_12443,N_11766,N_11986);
nor U12444 (N_12444,N_11166,N_11639);
xnor U12445 (N_12445,N_11015,N_11012);
nor U12446 (N_12446,N_11977,N_11141);
nor U12447 (N_12447,N_11223,N_11921);
and U12448 (N_12448,N_11966,N_11598);
or U12449 (N_12449,N_11726,N_11139);
xnor U12450 (N_12450,N_11901,N_11173);
and U12451 (N_12451,N_11323,N_11181);
nand U12452 (N_12452,N_11784,N_11436);
xnor U12453 (N_12453,N_11845,N_11462);
nand U12454 (N_12454,N_11930,N_11870);
nor U12455 (N_12455,N_11621,N_11832);
nor U12456 (N_12456,N_11903,N_11629);
xnor U12457 (N_12457,N_11229,N_11080);
or U12458 (N_12458,N_11409,N_11770);
nor U12459 (N_12459,N_11096,N_11363);
nand U12460 (N_12460,N_11906,N_11718);
xnor U12461 (N_12461,N_11222,N_11670);
nand U12462 (N_12462,N_11943,N_11831);
xnor U12463 (N_12463,N_11796,N_11781);
and U12464 (N_12464,N_11751,N_11711);
nand U12465 (N_12465,N_11002,N_11158);
or U12466 (N_12466,N_11068,N_11251);
nor U12467 (N_12467,N_11597,N_11595);
xor U12468 (N_12468,N_11541,N_11716);
nand U12469 (N_12469,N_11548,N_11860);
nand U12470 (N_12470,N_11793,N_11402);
or U12471 (N_12471,N_11589,N_11317);
xnor U12472 (N_12472,N_11523,N_11221);
nor U12473 (N_12473,N_11035,N_11964);
and U12474 (N_12474,N_11953,N_11885);
nand U12475 (N_12475,N_11070,N_11759);
nand U12476 (N_12476,N_11283,N_11105);
or U12477 (N_12477,N_11417,N_11437);
nand U12478 (N_12478,N_11764,N_11355);
nor U12479 (N_12479,N_11215,N_11156);
and U12480 (N_12480,N_11837,N_11701);
xor U12481 (N_12481,N_11274,N_11641);
and U12482 (N_12482,N_11036,N_11151);
nor U12483 (N_12483,N_11410,N_11863);
or U12484 (N_12484,N_11619,N_11575);
or U12485 (N_12485,N_11825,N_11401);
and U12486 (N_12486,N_11345,N_11192);
xor U12487 (N_12487,N_11131,N_11805);
nor U12488 (N_12488,N_11654,N_11822);
nand U12489 (N_12489,N_11798,N_11647);
nor U12490 (N_12490,N_11000,N_11397);
nor U12491 (N_12491,N_11806,N_11916);
and U12492 (N_12492,N_11234,N_11235);
nor U12493 (N_12493,N_11429,N_11702);
nand U12494 (N_12494,N_11326,N_11246);
nand U12495 (N_12495,N_11280,N_11499);
nor U12496 (N_12496,N_11833,N_11027);
or U12497 (N_12497,N_11593,N_11737);
xnor U12498 (N_12498,N_11114,N_11459);
xnor U12499 (N_12499,N_11938,N_11704);
and U12500 (N_12500,N_11412,N_11047);
xor U12501 (N_12501,N_11459,N_11678);
xnor U12502 (N_12502,N_11237,N_11587);
and U12503 (N_12503,N_11646,N_11111);
nor U12504 (N_12504,N_11513,N_11439);
or U12505 (N_12505,N_11379,N_11724);
xnor U12506 (N_12506,N_11998,N_11973);
xnor U12507 (N_12507,N_11674,N_11856);
or U12508 (N_12508,N_11428,N_11403);
nor U12509 (N_12509,N_11730,N_11525);
or U12510 (N_12510,N_11969,N_11355);
nor U12511 (N_12511,N_11395,N_11993);
nand U12512 (N_12512,N_11260,N_11777);
and U12513 (N_12513,N_11430,N_11751);
nor U12514 (N_12514,N_11773,N_11116);
or U12515 (N_12515,N_11786,N_11468);
or U12516 (N_12516,N_11447,N_11717);
nand U12517 (N_12517,N_11026,N_11825);
or U12518 (N_12518,N_11582,N_11226);
and U12519 (N_12519,N_11306,N_11326);
or U12520 (N_12520,N_11185,N_11924);
nand U12521 (N_12521,N_11756,N_11249);
and U12522 (N_12522,N_11452,N_11450);
nor U12523 (N_12523,N_11089,N_11042);
xor U12524 (N_12524,N_11280,N_11760);
and U12525 (N_12525,N_11697,N_11836);
and U12526 (N_12526,N_11455,N_11038);
nand U12527 (N_12527,N_11256,N_11635);
nor U12528 (N_12528,N_11845,N_11530);
nand U12529 (N_12529,N_11974,N_11033);
xnor U12530 (N_12530,N_11317,N_11249);
xor U12531 (N_12531,N_11888,N_11739);
and U12532 (N_12532,N_11957,N_11669);
or U12533 (N_12533,N_11088,N_11402);
or U12534 (N_12534,N_11771,N_11747);
or U12535 (N_12535,N_11141,N_11593);
nand U12536 (N_12536,N_11973,N_11434);
nor U12537 (N_12537,N_11847,N_11000);
xnor U12538 (N_12538,N_11700,N_11839);
and U12539 (N_12539,N_11940,N_11906);
xor U12540 (N_12540,N_11304,N_11867);
nand U12541 (N_12541,N_11448,N_11839);
or U12542 (N_12542,N_11180,N_11201);
nor U12543 (N_12543,N_11517,N_11880);
and U12544 (N_12544,N_11714,N_11626);
or U12545 (N_12545,N_11805,N_11808);
nand U12546 (N_12546,N_11062,N_11673);
xor U12547 (N_12547,N_11953,N_11321);
or U12548 (N_12548,N_11993,N_11215);
nand U12549 (N_12549,N_11878,N_11850);
nand U12550 (N_12550,N_11934,N_11996);
nor U12551 (N_12551,N_11976,N_11606);
nand U12552 (N_12552,N_11642,N_11270);
xnor U12553 (N_12553,N_11267,N_11742);
xnor U12554 (N_12554,N_11935,N_11742);
xor U12555 (N_12555,N_11872,N_11754);
xor U12556 (N_12556,N_11812,N_11335);
or U12557 (N_12557,N_11300,N_11900);
nor U12558 (N_12558,N_11301,N_11921);
nand U12559 (N_12559,N_11970,N_11801);
nor U12560 (N_12560,N_11625,N_11143);
and U12561 (N_12561,N_11859,N_11489);
or U12562 (N_12562,N_11540,N_11321);
xnor U12563 (N_12563,N_11722,N_11893);
and U12564 (N_12564,N_11415,N_11744);
and U12565 (N_12565,N_11390,N_11451);
nor U12566 (N_12566,N_11632,N_11952);
or U12567 (N_12567,N_11871,N_11751);
xor U12568 (N_12568,N_11650,N_11072);
nor U12569 (N_12569,N_11753,N_11166);
or U12570 (N_12570,N_11080,N_11133);
nor U12571 (N_12571,N_11595,N_11550);
and U12572 (N_12572,N_11652,N_11641);
nand U12573 (N_12573,N_11842,N_11928);
or U12574 (N_12574,N_11127,N_11837);
nor U12575 (N_12575,N_11731,N_11838);
or U12576 (N_12576,N_11855,N_11802);
or U12577 (N_12577,N_11680,N_11758);
nor U12578 (N_12578,N_11842,N_11156);
nand U12579 (N_12579,N_11362,N_11194);
xor U12580 (N_12580,N_11487,N_11323);
nor U12581 (N_12581,N_11341,N_11372);
nand U12582 (N_12582,N_11874,N_11954);
xnor U12583 (N_12583,N_11801,N_11737);
nand U12584 (N_12584,N_11812,N_11532);
or U12585 (N_12585,N_11561,N_11843);
and U12586 (N_12586,N_11133,N_11296);
and U12587 (N_12587,N_11473,N_11357);
or U12588 (N_12588,N_11910,N_11033);
nor U12589 (N_12589,N_11552,N_11112);
xor U12590 (N_12590,N_11936,N_11538);
xor U12591 (N_12591,N_11396,N_11267);
or U12592 (N_12592,N_11094,N_11750);
or U12593 (N_12593,N_11942,N_11492);
nor U12594 (N_12594,N_11999,N_11007);
nor U12595 (N_12595,N_11635,N_11605);
nand U12596 (N_12596,N_11862,N_11570);
xor U12597 (N_12597,N_11938,N_11709);
or U12598 (N_12598,N_11611,N_11661);
nor U12599 (N_12599,N_11678,N_11730);
and U12600 (N_12600,N_11290,N_11787);
and U12601 (N_12601,N_11096,N_11097);
and U12602 (N_12602,N_11247,N_11619);
nand U12603 (N_12603,N_11619,N_11698);
and U12604 (N_12604,N_11195,N_11184);
or U12605 (N_12605,N_11109,N_11392);
nor U12606 (N_12606,N_11363,N_11291);
xnor U12607 (N_12607,N_11542,N_11060);
xor U12608 (N_12608,N_11582,N_11039);
nor U12609 (N_12609,N_11634,N_11160);
and U12610 (N_12610,N_11149,N_11219);
xor U12611 (N_12611,N_11749,N_11969);
xor U12612 (N_12612,N_11758,N_11941);
and U12613 (N_12613,N_11405,N_11350);
nand U12614 (N_12614,N_11841,N_11642);
and U12615 (N_12615,N_11775,N_11732);
nor U12616 (N_12616,N_11790,N_11685);
and U12617 (N_12617,N_11627,N_11310);
and U12618 (N_12618,N_11130,N_11100);
and U12619 (N_12619,N_11316,N_11965);
or U12620 (N_12620,N_11353,N_11562);
nand U12621 (N_12621,N_11362,N_11337);
nand U12622 (N_12622,N_11581,N_11015);
nor U12623 (N_12623,N_11852,N_11611);
nor U12624 (N_12624,N_11884,N_11792);
nor U12625 (N_12625,N_11085,N_11264);
nor U12626 (N_12626,N_11692,N_11053);
nand U12627 (N_12627,N_11193,N_11507);
xnor U12628 (N_12628,N_11552,N_11085);
and U12629 (N_12629,N_11777,N_11470);
nor U12630 (N_12630,N_11047,N_11769);
xor U12631 (N_12631,N_11403,N_11784);
xnor U12632 (N_12632,N_11457,N_11068);
or U12633 (N_12633,N_11012,N_11709);
nor U12634 (N_12634,N_11985,N_11512);
xnor U12635 (N_12635,N_11187,N_11622);
xor U12636 (N_12636,N_11098,N_11533);
nor U12637 (N_12637,N_11526,N_11840);
nand U12638 (N_12638,N_11994,N_11365);
nor U12639 (N_12639,N_11539,N_11883);
or U12640 (N_12640,N_11409,N_11852);
xnor U12641 (N_12641,N_11375,N_11424);
or U12642 (N_12642,N_11030,N_11763);
nand U12643 (N_12643,N_11676,N_11100);
xnor U12644 (N_12644,N_11595,N_11647);
xor U12645 (N_12645,N_11417,N_11883);
xnor U12646 (N_12646,N_11000,N_11759);
or U12647 (N_12647,N_11115,N_11919);
xnor U12648 (N_12648,N_11109,N_11250);
and U12649 (N_12649,N_11667,N_11568);
or U12650 (N_12650,N_11127,N_11449);
or U12651 (N_12651,N_11315,N_11072);
and U12652 (N_12652,N_11842,N_11862);
or U12653 (N_12653,N_11954,N_11234);
or U12654 (N_12654,N_11217,N_11594);
nand U12655 (N_12655,N_11604,N_11312);
or U12656 (N_12656,N_11608,N_11064);
nor U12657 (N_12657,N_11274,N_11911);
or U12658 (N_12658,N_11336,N_11341);
and U12659 (N_12659,N_11852,N_11112);
xnor U12660 (N_12660,N_11772,N_11006);
nor U12661 (N_12661,N_11623,N_11968);
xnor U12662 (N_12662,N_11218,N_11872);
xor U12663 (N_12663,N_11772,N_11278);
xor U12664 (N_12664,N_11185,N_11331);
and U12665 (N_12665,N_11180,N_11227);
nor U12666 (N_12666,N_11340,N_11028);
nor U12667 (N_12667,N_11867,N_11619);
nor U12668 (N_12668,N_11171,N_11937);
or U12669 (N_12669,N_11091,N_11846);
or U12670 (N_12670,N_11821,N_11831);
nor U12671 (N_12671,N_11751,N_11336);
or U12672 (N_12672,N_11056,N_11383);
nor U12673 (N_12673,N_11326,N_11462);
or U12674 (N_12674,N_11594,N_11612);
nand U12675 (N_12675,N_11308,N_11495);
nand U12676 (N_12676,N_11798,N_11878);
and U12677 (N_12677,N_11809,N_11573);
or U12678 (N_12678,N_11407,N_11432);
or U12679 (N_12679,N_11442,N_11214);
xnor U12680 (N_12680,N_11522,N_11126);
nand U12681 (N_12681,N_11910,N_11271);
xnor U12682 (N_12682,N_11726,N_11663);
nand U12683 (N_12683,N_11186,N_11455);
nand U12684 (N_12684,N_11681,N_11665);
xor U12685 (N_12685,N_11062,N_11951);
and U12686 (N_12686,N_11160,N_11633);
nand U12687 (N_12687,N_11248,N_11802);
and U12688 (N_12688,N_11488,N_11212);
nand U12689 (N_12689,N_11050,N_11292);
and U12690 (N_12690,N_11200,N_11436);
xnor U12691 (N_12691,N_11864,N_11602);
and U12692 (N_12692,N_11168,N_11098);
or U12693 (N_12693,N_11705,N_11200);
and U12694 (N_12694,N_11595,N_11646);
and U12695 (N_12695,N_11041,N_11322);
nand U12696 (N_12696,N_11216,N_11278);
or U12697 (N_12697,N_11055,N_11576);
nor U12698 (N_12698,N_11281,N_11192);
nor U12699 (N_12699,N_11072,N_11298);
nand U12700 (N_12700,N_11402,N_11274);
xor U12701 (N_12701,N_11970,N_11696);
nand U12702 (N_12702,N_11794,N_11278);
nor U12703 (N_12703,N_11300,N_11663);
xnor U12704 (N_12704,N_11903,N_11031);
nand U12705 (N_12705,N_11727,N_11177);
and U12706 (N_12706,N_11948,N_11792);
xor U12707 (N_12707,N_11513,N_11456);
nand U12708 (N_12708,N_11140,N_11478);
or U12709 (N_12709,N_11797,N_11141);
xnor U12710 (N_12710,N_11330,N_11005);
or U12711 (N_12711,N_11150,N_11774);
nand U12712 (N_12712,N_11133,N_11271);
or U12713 (N_12713,N_11753,N_11580);
and U12714 (N_12714,N_11030,N_11503);
nor U12715 (N_12715,N_11889,N_11225);
nand U12716 (N_12716,N_11965,N_11045);
or U12717 (N_12717,N_11936,N_11898);
nand U12718 (N_12718,N_11668,N_11601);
nor U12719 (N_12719,N_11125,N_11536);
nor U12720 (N_12720,N_11619,N_11535);
or U12721 (N_12721,N_11732,N_11298);
and U12722 (N_12722,N_11223,N_11362);
and U12723 (N_12723,N_11315,N_11407);
or U12724 (N_12724,N_11636,N_11884);
or U12725 (N_12725,N_11366,N_11403);
nor U12726 (N_12726,N_11140,N_11755);
or U12727 (N_12727,N_11798,N_11891);
xnor U12728 (N_12728,N_11011,N_11573);
and U12729 (N_12729,N_11144,N_11078);
nor U12730 (N_12730,N_11606,N_11423);
nor U12731 (N_12731,N_11169,N_11736);
nor U12732 (N_12732,N_11504,N_11881);
and U12733 (N_12733,N_11402,N_11019);
xnor U12734 (N_12734,N_11120,N_11114);
nand U12735 (N_12735,N_11494,N_11928);
nand U12736 (N_12736,N_11482,N_11457);
xnor U12737 (N_12737,N_11469,N_11742);
nand U12738 (N_12738,N_11495,N_11192);
nor U12739 (N_12739,N_11535,N_11122);
xor U12740 (N_12740,N_11367,N_11675);
nand U12741 (N_12741,N_11673,N_11183);
nor U12742 (N_12742,N_11978,N_11154);
nor U12743 (N_12743,N_11293,N_11331);
and U12744 (N_12744,N_11391,N_11958);
nand U12745 (N_12745,N_11174,N_11047);
xnor U12746 (N_12746,N_11781,N_11365);
nor U12747 (N_12747,N_11625,N_11877);
and U12748 (N_12748,N_11601,N_11590);
or U12749 (N_12749,N_11730,N_11807);
xnor U12750 (N_12750,N_11928,N_11189);
xor U12751 (N_12751,N_11219,N_11403);
or U12752 (N_12752,N_11694,N_11487);
xnor U12753 (N_12753,N_11460,N_11483);
nand U12754 (N_12754,N_11874,N_11220);
and U12755 (N_12755,N_11305,N_11034);
and U12756 (N_12756,N_11633,N_11393);
and U12757 (N_12757,N_11071,N_11213);
nor U12758 (N_12758,N_11164,N_11527);
xor U12759 (N_12759,N_11232,N_11344);
nor U12760 (N_12760,N_11452,N_11980);
nor U12761 (N_12761,N_11654,N_11811);
nand U12762 (N_12762,N_11946,N_11230);
or U12763 (N_12763,N_11863,N_11287);
or U12764 (N_12764,N_11107,N_11664);
and U12765 (N_12765,N_11911,N_11951);
and U12766 (N_12766,N_11607,N_11173);
and U12767 (N_12767,N_11575,N_11933);
or U12768 (N_12768,N_11239,N_11351);
nand U12769 (N_12769,N_11839,N_11727);
nor U12770 (N_12770,N_11356,N_11681);
or U12771 (N_12771,N_11915,N_11317);
xor U12772 (N_12772,N_11174,N_11562);
and U12773 (N_12773,N_11023,N_11321);
xnor U12774 (N_12774,N_11518,N_11195);
xor U12775 (N_12775,N_11450,N_11730);
or U12776 (N_12776,N_11820,N_11610);
nor U12777 (N_12777,N_11583,N_11835);
nand U12778 (N_12778,N_11046,N_11364);
and U12779 (N_12779,N_11010,N_11964);
or U12780 (N_12780,N_11853,N_11793);
xor U12781 (N_12781,N_11539,N_11605);
or U12782 (N_12782,N_11175,N_11798);
and U12783 (N_12783,N_11725,N_11280);
xnor U12784 (N_12784,N_11296,N_11419);
nand U12785 (N_12785,N_11386,N_11652);
nor U12786 (N_12786,N_11606,N_11719);
xor U12787 (N_12787,N_11882,N_11618);
or U12788 (N_12788,N_11645,N_11580);
or U12789 (N_12789,N_11811,N_11307);
nand U12790 (N_12790,N_11643,N_11936);
and U12791 (N_12791,N_11845,N_11933);
xor U12792 (N_12792,N_11804,N_11705);
nor U12793 (N_12793,N_11477,N_11606);
and U12794 (N_12794,N_11184,N_11672);
and U12795 (N_12795,N_11482,N_11037);
and U12796 (N_12796,N_11582,N_11253);
and U12797 (N_12797,N_11263,N_11331);
xnor U12798 (N_12798,N_11260,N_11948);
nor U12799 (N_12799,N_11944,N_11707);
xnor U12800 (N_12800,N_11405,N_11048);
nor U12801 (N_12801,N_11975,N_11052);
nand U12802 (N_12802,N_11852,N_11760);
nor U12803 (N_12803,N_11924,N_11762);
nor U12804 (N_12804,N_11824,N_11107);
xor U12805 (N_12805,N_11069,N_11365);
nor U12806 (N_12806,N_11217,N_11037);
nand U12807 (N_12807,N_11109,N_11974);
nand U12808 (N_12808,N_11925,N_11713);
and U12809 (N_12809,N_11363,N_11815);
nand U12810 (N_12810,N_11624,N_11185);
and U12811 (N_12811,N_11760,N_11679);
or U12812 (N_12812,N_11181,N_11523);
or U12813 (N_12813,N_11852,N_11324);
xnor U12814 (N_12814,N_11441,N_11285);
and U12815 (N_12815,N_11099,N_11289);
xor U12816 (N_12816,N_11119,N_11761);
and U12817 (N_12817,N_11283,N_11243);
nor U12818 (N_12818,N_11367,N_11866);
and U12819 (N_12819,N_11551,N_11166);
nand U12820 (N_12820,N_11009,N_11948);
nand U12821 (N_12821,N_11074,N_11969);
xor U12822 (N_12822,N_11140,N_11767);
nand U12823 (N_12823,N_11018,N_11686);
nor U12824 (N_12824,N_11088,N_11311);
and U12825 (N_12825,N_11393,N_11299);
nor U12826 (N_12826,N_11180,N_11033);
xnor U12827 (N_12827,N_11447,N_11304);
xnor U12828 (N_12828,N_11039,N_11295);
xor U12829 (N_12829,N_11774,N_11480);
nand U12830 (N_12830,N_11436,N_11162);
xor U12831 (N_12831,N_11093,N_11720);
or U12832 (N_12832,N_11591,N_11012);
nand U12833 (N_12833,N_11515,N_11541);
nor U12834 (N_12834,N_11463,N_11618);
nand U12835 (N_12835,N_11125,N_11118);
or U12836 (N_12836,N_11294,N_11330);
xnor U12837 (N_12837,N_11386,N_11684);
nand U12838 (N_12838,N_11817,N_11565);
xor U12839 (N_12839,N_11012,N_11866);
and U12840 (N_12840,N_11874,N_11811);
and U12841 (N_12841,N_11011,N_11218);
or U12842 (N_12842,N_11495,N_11693);
nand U12843 (N_12843,N_11782,N_11911);
xnor U12844 (N_12844,N_11550,N_11639);
nor U12845 (N_12845,N_11223,N_11682);
or U12846 (N_12846,N_11558,N_11562);
nand U12847 (N_12847,N_11570,N_11985);
or U12848 (N_12848,N_11211,N_11791);
xnor U12849 (N_12849,N_11523,N_11022);
and U12850 (N_12850,N_11856,N_11476);
nand U12851 (N_12851,N_11205,N_11262);
nor U12852 (N_12852,N_11358,N_11450);
or U12853 (N_12853,N_11819,N_11273);
nand U12854 (N_12854,N_11082,N_11834);
xor U12855 (N_12855,N_11006,N_11230);
or U12856 (N_12856,N_11677,N_11501);
or U12857 (N_12857,N_11113,N_11188);
and U12858 (N_12858,N_11019,N_11894);
xnor U12859 (N_12859,N_11480,N_11127);
nor U12860 (N_12860,N_11635,N_11803);
and U12861 (N_12861,N_11894,N_11403);
and U12862 (N_12862,N_11995,N_11403);
nor U12863 (N_12863,N_11561,N_11519);
nor U12864 (N_12864,N_11209,N_11564);
nor U12865 (N_12865,N_11705,N_11445);
and U12866 (N_12866,N_11715,N_11638);
xor U12867 (N_12867,N_11743,N_11049);
nand U12868 (N_12868,N_11329,N_11608);
nand U12869 (N_12869,N_11922,N_11614);
nor U12870 (N_12870,N_11227,N_11555);
and U12871 (N_12871,N_11697,N_11960);
and U12872 (N_12872,N_11458,N_11324);
and U12873 (N_12873,N_11533,N_11226);
or U12874 (N_12874,N_11671,N_11591);
nor U12875 (N_12875,N_11429,N_11742);
nand U12876 (N_12876,N_11415,N_11430);
nand U12877 (N_12877,N_11941,N_11740);
nor U12878 (N_12878,N_11680,N_11677);
and U12879 (N_12879,N_11478,N_11983);
nor U12880 (N_12880,N_11994,N_11694);
or U12881 (N_12881,N_11043,N_11743);
xnor U12882 (N_12882,N_11830,N_11951);
nor U12883 (N_12883,N_11189,N_11088);
or U12884 (N_12884,N_11135,N_11950);
nand U12885 (N_12885,N_11370,N_11455);
xnor U12886 (N_12886,N_11993,N_11485);
nand U12887 (N_12887,N_11597,N_11387);
nor U12888 (N_12888,N_11279,N_11672);
and U12889 (N_12889,N_11016,N_11726);
or U12890 (N_12890,N_11468,N_11993);
xor U12891 (N_12891,N_11230,N_11197);
and U12892 (N_12892,N_11537,N_11094);
xnor U12893 (N_12893,N_11890,N_11464);
xnor U12894 (N_12894,N_11892,N_11844);
nor U12895 (N_12895,N_11737,N_11290);
and U12896 (N_12896,N_11899,N_11802);
nor U12897 (N_12897,N_11799,N_11082);
and U12898 (N_12898,N_11917,N_11291);
nand U12899 (N_12899,N_11353,N_11663);
nor U12900 (N_12900,N_11412,N_11804);
nor U12901 (N_12901,N_11995,N_11419);
and U12902 (N_12902,N_11531,N_11442);
nand U12903 (N_12903,N_11757,N_11606);
nor U12904 (N_12904,N_11003,N_11314);
nor U12905 (N_12905,N_11537,N_11788);
nor U12906 (N_12906,N_11415,N_11482);
nor U12907 (N_12907,N_11341,N_11822);
nor U12908 (N_12908,N_11062,N_11818);
nor U12909 (N_12909,N_11001,N_11111);
or U12910 (N_12910,N_11446,N_11038);
xor U12911 (N_12911,N_11885,N_11760);
and U12912 (N_12912,N_11577,N_11642);
xor U12913 (N_12913,N_11719,N_11694);
or U12914 (N_12914,N_11433,N_11586);
nand U12915 (N_12915,N_11530,N_11431);
or U12916 (N_12916,N_11928,N_11445);
nor U12917 (N_12917,N_11727,N_11342);
nor U12918 (N_12918,N_11080,N_11142);
or U12919 (N_12919,N_11523,N_11922);
nand U12920 (N_12920,N_11685,N_11346);
and U12921 (N_12921,N_11094,N_11295);
nand U12922 (N_12922,N_11776,N_11853);
nand U12923 (N_12923,N_11374,N_11919);
nor U12924 (N_12924,N_11295,N_11416);
or U12925 (N_12925,N_11362,N_11612);
and U12926 (N_12926,N_11801,N_11694);
nand U12927 (N_12927,N_11908,N_11527);
and U12928 (N_12928,N_11634,N_11051);
nand U12929 (N_12929,N_11243,N_11429);
nand U12930 (N_12930,N_11810,N_11984);
xor U12931 (N_12931,N_11404,N_11697);
xnor U12932 (N_12932,N_11530,N_11410);
nor U12933 (N_12933,N_11229,N_11557);
nand U12934 (N_12934,N_11292,N_11815);
xor U12935 (N_12935,N_11222,N_11838);
nand U12936 (N_12936,N_11599,N_11865);
nand U12937 (N_12937,N_11267,N_11926);
nor U12938 (N_12938,N_11711,N_11335);
xor U12939 (N_12939,N_11690,N_11076);
nand U12940 (N_12940,N_11712,N_11974);
xor U12941 (N_12941,N_11285,N_11962);
and U12942 (N_12942,N_11285,N_11996);
and U12943 (N_12943,N_11081,N_11204);
xor U12944 (N_12944,N_11561,N_11971);
or U12945 (N_12945,N_11629,N_11432);
xor U12946 (N_12946,N_11311,N_11572);
and U12947 (N_12947,N_11869,N_11621);
nand U12948 (N_12948,N_11587,N_11129);
xnor U12949 (N_12949,N_11062,N_11726);
nor U12950 (N_12950,N_11221,N_11395);
xnor U12951 (N_12951,N_11832,N_11374);
xnor U12952 (N_12952,N_11877,N_11647);
and U12953 (N_12953,N_11350,N_11854);
and U12954 (N_12954,N_11872,N_11612);
xnor U12955 (N_12955,N_11132,N_11390);
nor U12956 (N_12956,N_11294,N_11425);
and U12957 (N_12957,N_11158,N_11426);
or U12958 (N_12958,N_11244,N_11055);
or U12959 (N_12959,N_11262,N_11364);
and U12960 (N_12960,N_11868,N_11462);
xnor U12961 (N_12961,N_11056,N_11030);
xor U12962 (N_12962,N_11063,N_11673);
xor U12963 (N_12963,N_11259,N_11145);
and U12964 (N_12964,N_11970,N_11306);
or U12965 (N_12965,N_11706,N_11297);
and U12966 (N_12966,N_11805,N_11220);
nand U12967 (N_12967,N_11376,N_11372);
and U12968 (N_12968,N_11285,N_11444);
or U12969 (N_12969,N_11431,N_11820);
nor U12970 (N_12970,N_11744,N_11998);
or U12971 (N_12971,N_11863,N_11513);
and U12972 (N_12972,N_11734,N_11236);
and U12973 (N_12973,N_11392,N_11270);
nand U12974 (N_12974,N_11137,N_11824);
and U12975 (N_12975,N_11374,N_11623);
nand U12976 (N_12976,N_11724,N_11864);
nand U12977 (N_12977,N_11529,N_11973);
or U12978 (N_12978,N_11002,N_11286);
and U12979 (N_12979,N_11531,N_11413);
and U12980 (N_12980,N_11922,N_11602);
and U12981 (N_12981,N_11903,N_11009);
and U12982 (N_12982,N_11646,N_11158);
xor U12983 (N_12983,N_11867,N_11236);
nand U12984 (N_12984,N_11010,N_11327);
nand U12985 (N_12985,N_11513,N_11406);
xnor U12986 (N_12986,N_11840,N_11242);
or U12987 (N_12987,N_11633,N_11978);
xnor U12988 (N_12988,N_11386,N_11614);
and U12989 (N_12989,N_11502,N_11196);
xor U12990 (N_12990,N_11095,N_11677);
xor U12991 (N_12991,N_11547,N_11387);
nor U12992 (N_12992,N_11843,N_11029);
or U12993 (N_12993,N_11468,N_11601);
or U12994 (N_12994,N_11309,N_11245);
nor U12995 (N_12995,N_11875,N_11652);
nor U12996 (N_12996,N_11039,N_11647);
and U12997 (N_12997,N_11708,N_11652);
nor U12998 (N_12998,N_11627,N_11612);
nor U12999 (N_12999,N_11488,N_11425);
or U13000 (N_13000,N_12625,N_12772);
or U13001 (N_13001,N_12368,N_12822);
nand U13002 (N_13002,N_12582,N_12282);
xor U13003 (N_13003,N_12130,N_12457);
and U13004 (N_13004,N_12838,N_12225);
and U13005 (N_13005,N_12219,N_12409);
xnor U13006 (N_13006,N_12761,N_12996);
nand U13007 (N_13007,N_12333,N_12026);
nor U13008 (N_13008,N_12759,N_12231);
nand U13009 (N_13009,N_12245,N_12849);
or U13010 (N_13010,N_12117,N_12399);
xor U13011 (N_13011,N_12114,N_12186);
or U13012 (N_13012,N_12581,N_12795);
or U13013 (N_13013,N_12813,N_12145);
nand U13014 (N_13014,N_12535,N_12745);
nand U13015 (N_13015,N_12052,N_12785);
xnor U13016 (N_13016,N_12687,N_12251);
xnor U13017 (N_13017,N_12847,N_12275);
nand U13018 (N_13018,N_12736,N_12043);
nor U13019 (N_13019,N_12608,N_12104);
nor U13020 (N_13020,N_12442,N_12132);
xor U13021 (N_13021,N_12390,N_12141);
or U13022 (N_13022,N_12283,N_12890);
nand U13023 (N_13023,N_12916,N_12893);
nand U13024 (N_13024,N_12209,N_12600);
or U13025 (N_13025,N_12048,N_12447);
and U13026 (N_13026,N_12035,N_12841);
xnor U13027 (N_13027,N_12748,N_12196);
nor U13028 (N_13028,N_12153,N_12458);
or U13029 (N_13029,N_12329,N_12110);
and U13030 (N_13030,N_12467,N_12797);
and U13031 (N_13031,N_12870,N_12798);
nor U13032 (N_13032,N_12638,N_12911);
xor U13033 (N_13033,N_12900,N_12183);
xor U13034 (N_13034,N_12489,N_12370);
nor U13035 (N_13035,N_12299,N_12803);
nor U13036 (N_13036,N_12904,N_12669);
xnor U13037 (N_13037,N_12987,N_12311);
nor U13038 (N_13038,N_12357,N_12871);
or U13039 (N_13039,N_12363,N_12902);
xnor U13040 (N_13040,N_12895,N_12391);
or U13041 (N_13041,N_12405,N_12671);
xor U13042 (N_13042,N_12242,N_12906);
and U13043 (N_13043,N_12273,N_12212);
or U13044 (N_13044,N_12081,N_12989);
or U13045 (N_13045,N_12665,N_12596);
nand U13046 (N_13046,N_12852,N_12019);
nand U13047 (N_13047,N_12905,N_12091);
and U13048 (N_13048,N_12738,N_12339);
and U13049 (N_13049,N_12940,N_12147);
nand U13050 (N_13050,N_12783,N_12878);
and U13051 (N_13051,N_12599,N_12611);
and U13052 (N_13052,N_12025,N_12042);
nor U13053 (N_13053,N_12965,N_12078);
xnor U13054 (N_13054,N_12359,N_12695);
xor U13055 (N_13055,N_12994,N_12888);
xor U13056 (N_13056,N_12478,N_12526);
or U13057 (N_13057,N_12630,N_12731);
nor U13058 (N_13058,N_12481,N_12606);
and U13059 (N_13059,N_12627,N_12848);
nor U13060 (N_13060,N_12885,N_12438);
and U13061 (N_13061,N_12869,N_12144);
nand U13062 (N_13062,N_12677,N_12154);
xnor U13063 (N_13063,N_12933,N_12971);
and U13064 (N_13064,N_12187,N_12594);
nand U13065 (N_13065,N_12127,N_12663);
or U13066 (N_13066,N_12693,N_12790);
nand U13067 (N_13067,N_12022,N_12376);
nand U13068 (N_13068,N_12810,N_12898);
nand U13069 (N_13069,N_12604,N_12876);
nor U13070 (N_13070,N_12754,N_12716);
nor U13071 (N_13071,N_12650,N_12845);
or U13072 (N_13072,N_12168,N_12455);
nor U13073 (N_13073,N_12942,N_12562);
and U13074 (N_13074,N_12515,N_12367);
nor U13075 (N_13075,N_12372,N_12805);
xnor U13076 (N_13076,N_12784,N_12986);
nand U13077 (N_13077,N_12249,N_12020);
and U13078 (N_13078,N_12944,N_12527);
nor U13079 (N_13079,N_12158,N_12935);
xnor U13080 (N_13080,N_12381,N_12646);
nand U13081 (N_13081,N_12583,N_12016);
xnor U13082 (N_13082,N_12003,N_12598);
xnor U13083 (N_13083,N_12278,N_12434);
or U13084 (N_13084,N_12142,N_12241);
and U13085 (N_13085,N_12758,N_12248);
or U13086 (N_13086,N_12193,N_12921);
nor U13087 (N_13087,N_12685,N_12364);
nand U13088 (N_13088,N_12176,N_12571);
nand U13089 (N_13089,N_12725,N_12943);
xor U13090 (N_13090,N_12733,N_12766);
nand U13091 (N_13091,N_12877,N_12688);
and U13092 (N_13092,N_12773,N_12129);
xnor U13093 (N_13093,N_12471,N_12559);
nor U13094 (N_13094,N_12444,N_12675);
and U13095 (N_13095,N_12879,N_12403);
nand U13096 (N_13096,N_12382,N_12206);
xor U13097 (N_13097,N_12366,N_12844);
or U13098 (N_13098,N_12238,N_12338);
nor U13099 (N_13099,N_12528,N_12284);
nand U13100 (N_13100,N_12757,N_12433);
nor U13101 (N_13101,N_12556,N_12605);
and U13102 (N_13102,N_12224,N_12373);
nand U13103 (N_13103,N_12085,N_12239);
and U13104 (N_13104,N_12446,N_12120);
nand U13105 (N_13105,N_12937,N_12723);
xnor U13106 (N_13106,N_12941,N_12769);
and U13107 (N_13107,N_12440,N_12652);
xnor U13108 (N_13108,N_12839,N_12896);
xor U13109 (N_13109,N_12930,N_12667);
xnor U13110 (N_13110,N_12353,N_12384);
nand U13111 (N_13111,N_12522,N_12518);
or U13112 (N_13112,N_12086,N_12701);
xor U13113 (N_13113,N_12636,N_12756);
and U13114 (N_13114,N_12782,N_12710);
nand U13115 (N_13115,N_12083,N_12791);
nor U13116 (N_13116,N_12073,N_12912);
and U13117 (N_13117,N_12228,N_12326);
nor U13118 (N_13118,N_12149,N_12683);
nor U13119 (N_13119,N_12220,N_12770);
nor U13120 (N_13120,N_12165,N_12549);
or U13121 (N_13121,N_12775,N_12272);
nand U13122 (N_13122,N_12613,N_12512);
and U13123 (N_13123,N_12684,N_12058);
or U13124 (N_13124,N_12680,N_12076);
or U13125 (N_13125,N_12614,N_12946);
nand U13126 (N_13126,N_12097,N_12497);
or U13127 (N_13127,N_12018,N_12059);
xor U13128 (N_13128,N_12387,N_12846);
xor U13129 (N_13129,N_12253,N_12629);
and U13130 (N_13130,N_12448,N_12369);
and U13131 (N_13131,N_12265,N_12974);
and U13132 (N_13132,N_12516,N_12169);
nand U13133 (N_13133,N_12074,N_12578);
nor U13134 (N_13134,N_12166,N_12577);
or U13135 (N_13135,N_12771,N_12015);
xnor U13136 (N_13136,N_12707,N_12880);
nor U13137 (N_13137,N_12654,N_12028);
or U13138 (N_13138,N_12816,N_12826);
nand U13139 (N_13139,N_12011,N_12696);
xor U13140 (N_13140,N_12294,N_12925);
nor U13141 (N_13141,N_12576,N_12626);
and U13142 (N_13142,N_12909,N_12881);
nor U13143 (N_13143,N_12715,N_12044);
xor U13144 (N_13144,N_12427,N_12737);
nand U13145 (N_13145,N_12714,N_12198);
xor U13146 (N_13146,N_12408,N_12860);
nor U13147 (N_13147,N_12386,N_12708);
and U13148 (N_13148,N_12213,N_12050);
xnor U13149 (N_13149,N_12831,N_12226);
nand U13150 (N_13150,N_12595,N_12936);
nor U13151 (N_13151,N_12465,N_12252);
xor U13152 (N_13152,N_12395,N_12227);
nand U13153 (N_13153,N_12874,N_12155);
and U13154 (N_13154,N_12079,N_12645);
nor U13155 (N_13155,N_12919,N_12205);
nor U13156 (N_13156,N_12317,N_12109);
and U13157 (N_13157,N_12229,N_12620);
and U13158 (N_13158,N_12362,N_12678);
and U13159 (N_13159,N_12108,N_12005);
nor U13160 (N_13160,N_12195,N_12873);
nor U13161 (N_13161,N_12393,N_12235);
and U13162 (N_13162,N_12069,N_12118);
and U13163 (N_13163,N_12825,N_12705);
or U13164 (N_13164,N_12853,N_12146);
nor U13165 (N_13165,N_12740,N_12607);
nand U13166 (N_13166,N_12800,N_12344);
nor U13167 (N_13167,N_12815,N_12063);
xnor U13168 (N_13168,N_12419,N_12123);
nand U13169 (N_13169,N_12126,N_12060);
nor U13170 (N_13170,N_12938,N_12106);
or U13171 (N_13171,N_12428,N_12172);
nand U13172 (N_13172,N_12140,N_12612);
xnor U13173 (N_13173,N_12601,N_12309);
and U13174 (N_13174,N_12466,N_12922);
and U13175 (N_13175,N_12832,N_12891);
xnor U13176 (N_13176,N_12477,N_12643);
and U13177 (N_13177,N_12222,N_12441);
xor U13178 (N_13178,N_12482,N_12009);
and U13179 (N_13179,N_12570,N_12762);
nor U13180 (N_13180,N_12546,N_12411);
nor U13181 (N_13181,N_12306,N_12305);
or U13182 (N_13182,N_12013,N_12637);
nand U13183 (N_13183,N_12981,N_12519);
and U13184 (N_13184,N_12875,N_12973);
or U13185 (N_13185,N_12978,N_12959);
and U13186 (N_13186,N_12463,N_12640);
nand U13187 (N_13187,N_12732,N_12237);
and U13188 (N_13188,N_12819,N_12289);
and U13189 (N_13189,N_12586,N_12647);
or U13190 (N_13190,N_12713,N_12365);
or U13191 (N_13191,N_12950,N_12014);
nor U13192 (N_13192,N_12415,N_12077);
xor U13193 (N_13193,N_12297,N_12180);
xnor U13194 (N_13194,N_12926,N_12915);
nor U13195 (N_13195,N_12483,N_12164);
nor U13196 (N_13196,N_12036,N_12812);
nand U13197 (N_13197,N_12223,N_12356);
and U13198 (N_13198,N_12982,N_12719);
or U13199 (N_13199,N_12301,N_12274);
or U13200 (N_13200,N_12194,N_12547);
or U13201 (N_13201,N_12181,N_12006);
xnor U13202 (N_13202,N_12510,N_12349);
or U13203 (N_13203,N_12388,N_12383);
or U13204 (N_13204,N_12722,N_12045);
xnor U13205 (N_13205,N_12616,N_12966);
or U13206 (N_13206,N_12103,N_12037);
nand U13207 (N_13207,N_12892,N_12068);
and U13208 (N_13208,N_12240,N_12778);
nand U13209 (N_13209,N_12210,N_12975);
nand U13210 (N_13210,N_12823,N_12287);
nor U13211 (N_13211,N_12254,N_12484);
and U13212 (N_13212,N_12479,N_12644);
and U13213 (N_13213,N_12692,N_12413);
or U13214 (N_13214,N_12184,N_12953);
xnor U13215 (N_13215,N_12247,N_12332);
and U13216 (N_13216,N_12967,N_12883);
and U13217 (N_13217,N_12843,N_12163);
nand U13218 (N_13218,N_12351,N_12323);
nor U13219 (N_13219,N_12592,N_12550);
or U13220 (N_13220,N_12749,N_12295);
or U13221 (N_13221,N_12956,N_12285);
nor U13222 (N_13222,N_12500,N_12691);
nand U13223 (N_13223,N_12504,N_12334);
xor U13224 (N_13224,N_12742,N_12065);
nand U13225 (N_13225,N_12866,N_12779);
xnor U13226 (N_13226,N_12730,N_12894);
xor U13227 (N_13227,N_12589,N_12536);
nor U13228 (N_13228,N_12410,N_12088);
nor U13229 (N_13229,N_12098,N_12752);
or U13230 (N_13230,N_12591,N_12682);
xor U13231 (N_13231,N_12539,N_12100);
nor U13232 (N_13232,N_12859,N_12506);
and U13233 (N_13233,N_12218,N_12668);
and U13234 (N_13234,N_12173,N_12379);
nor U13235 (N_13235,N_12192,N_12143);
xor U13236 (N_13236,N_12089,N_12914);
and U13237 (N_13237,N_12579,N_12360);
nand U13238 (N_13238,N_12821,N_12835);
nand U13239 (N_13239,N_12121,N_12699);
and U13240 (N_13240,N_12452,N_12190);
nand U13241 (N_13241,N_12266,N_12062);
nor U13242 (N_13242,N_12331,N_12315);
xnor U13243 (N_13243,N_12070,N_12468);
xnor U13244 (N_13244,N_12469,N_12177);
or U13245 (N_13245,N_12789,N_12928);
nor U13246 (N_13246,N_12107,N_12000);
xnor U13247 (N_13247,N_12017,N_12407);
nor U13248 (N_13248,N_12765,N_12361);
and U13249 (N_13249,N_12216,N_12348);
or U13250 (N_13250,N_12138,N_12156);
xnor U13251 (N_13251,N_12801,N_12174);
and U13252 (N_13252,N_12179,N_12416);
or U13253 (N_13253,N_12533,N_12189);
and U13254 (N_13254,N_12969,N_12777);
or U13255 (N_13255,N_12985,N_12087);
xnor U13256 (N_13256,N_12486,N_12342);
nand U13257 (N_13257,N_12603,N_12041);
nor U13258 (N_13258,N_12991,N_12199);
and U13259 (N_13259,N_12431,N_12633);
xor U13260 (N_13260,N_12712,N_12917);
nor U13261 (N_13261,N_12865,N_12498);
nor U13262 (N_13262,N_12857,N_12054);
nand U13263 (N_13263,N_12350,N_12378);
or U13264 (N_13264,N_12717,N_12207);
or U13265 (N_13265,N_12259,N_12246);
xor U13266 (N_13266,N_12686,N_12105);
nand U13267 (N_13267,N_12521,N_12552);
nand U13268 (N_13268,N_12659,N_12221);
nor U13269 (N_13269,N_12868,N_12032);
nor U13270 (N_13270,N_12728,N_12056);
xor U13271 (N_13271,N_12122,N_12711);
or U13272 (N_13272,N_12963,N_12945);
xnor U13273 (N_13273,N_12739,N_12182);
nor U13274 (N_13274,N_12072,N_12341);
xor U13275 (N_13275,N_12744,N_12281);
and U13276 (N_13276,N_12188,N_12008);
nand U13277 (N_13277,N_12160,N_12939);
xor U13278 (N_13278,N_12672,N_12340);
and U13279 (N_13279,N_12622,N_12624);
nor U13280 (N_13280,N_12631,N_12664);
nor U13281 (N_13281,N_12330,N_12377);
or U13282 (N_13282,N_12234,N_12354);
nand U13283 (N_13283,N_12760,N_12907);
and U13284 (N_13284,N_12319,N_12543);
nand U13285 (N_13285,N_12995,N_12850);
nor U13286 (N_13286,N_12566,N_12093);
and U13287 (N_13287,N_12047,N_12394);
xor U13288 (N_13288,N_12300,N_12304);
nor U13289 (N_13289,N_12538,N_12726);
xnor U13290 (N_13290,N_12027,N_12551);
or U13291 (N_13291,N_12298,N_12437);
xor U13292 (N_13292,N_12290,N_12530);
nor U13293 (N_13293,N_12806,N_12660);
xnor U13294 (N_13294,N_12727,N_12488);
xnor U13295 (N_13295,N_12337,N_12288);
xnor U13296 (N_13296,N_12430,N_12662);
nor U13297 (N_13297,N_12700,N_12886);
nand U13298 (N_13298,N_12802,N_12268);
and U13299 (N_13299,N_12615,N_12374);
xor U13300 (N_13300,N_12057,N_12657);
and U13301 (N_13301,N_12542,N_12096);
nor U13302 (N_13302,N_12743,N_12574);
or U13303 (N_13303,N_12824,N_12414);
nor U13304 (N_13304,N_12460,N_12970);
xor U13305 (N_13305,N_12398,N_12040);
nor U13306 (N_13306,N_12634,N_12236);
nor U13307 (N_13307,N_12116,N_12913);
or U13308 (N_13308,N_12794,N_12617);
nor U13309 (N_13309,N_12112,N_12046);
xor U13310 (N_13310,N_12406,N_12150);
and U13311 (N_13311,N_12724,N_12055);
and U13312 (N_13312,N_12352,N_12523);
nor U13313 (N_13313,N_12670,N_12541);
nor U13314 (N_13314,N_12320,N_12421);
nor U13315 (N_13315,N_12520,N_12264);
and U13316 (N_13316,N_12658,N_12402);
nor U13317 (N_13317,N_12211,N_12961);
nand U13318 (N_13318,N_12704,N_12830);
xor U13319 (N_13319,N_12066,N_12954);
nor U13320 (N_13320,N_12292,N_12464);
xnor U13321 (N_13321,N_12828,N_12609);
or U13322 (N_13322,N_12260,N_12661);
nor U13323 (N_13323,N_12404,N_12327);
and U13324 (N_13324,N_12854,N_12651);
nand U13325 (N_13325,N_12799,N_12811);
or U13326 (N_13326,N_12544,N_12313);
and U13327 (N_13327,N_12261,N_12053);
or U13328 (N_13328,N_12918,N_12010);
and U13329 (N_13329,N_12979,N_12064);
or U13330 (N_13330,N_12532,N_12593);
xor U13331 (N_13331,N_12157,N_12030);
xnor U13332 (N_13332,N_12271,N_12729);
nand U13333 (N_13333,N_12610,N_12628);
xor U13334 (N_13334,N_12563,N_12308);
and U13335 (N_13335,N_12417,N_12972);
nor U13336 (N_13336,N_12316,N_12021);
or U13337 (N_13337,N_12555,N_12508);
or U13338 (N_13338,N_12741,N_12310);
and U13339 (N_13339,N_12621,N_12099);
and U13340 (N_13340,N_12690,N_12851);
and U13341 (N_13341,N_12012,N_12929);
nor U13342 (N_13342,N_12947,N_12572);
xor U13343 (N_13343,N_12286,N_12540);
nand U13344 (N_13344,N_12561,N_12033);
nand U13345 (N_13345,N_12133,N_12152);
nand U13346 (N_13346,N_12703,N_12951);
nand U13347 (N_13347,N_12128,N_12554);
xnor U13348 (N_13348,N_12007,N_12768);
or U13349 (N_13349,N_12920,N_12780);
xnor U13350 (N_13350,N_12461,N_12649);
nand U13351 (N_13351,N_12597,N_12474);
xor U13352 (N_13352,N_12346,N_12666);
and U13353 (N_13353,N_12380,N_12502);
nor U13354 (N_13354,N_12899,N_12517);
and U13355 (N_13355,N_12202,N_12618);
or U13356 (N_13356,N_12347,N_12204);
nor U13357 (N_13357,N_12302,N_12197);
or U13358 (N_13358,N_12889,N_12923);
xnor U13359 (N_13359,N_12641,N_12175);
or U13360 (N_13360,N_12071,N_12746);
nor U13361 (N_13361,N_12702,N_12296);
nand U13362 (N_13362,N_12964,N_12855);
xnor U13363 (N_13363,N_12734,N_12709);
nor U13364 (N_13364,N_12080,N_12924);
nand U13365 (N_13365,N_12276,N_12511);
xor U13366 (N_13366,N_12485,N_12375);
or U13367 (N_13367,N_12639,N_12655);
or U13368 (N_13368,N_12400,N_12793);
nor U13369 (N_13369,N_12401,N_12092);
nand U13370 (N_13370,N_12113,N_12840);
nor U13371 (N_13371,N_12753,N_12927);
and U13372 (N_13372,N_12827,N_12689);
and U13373 (N_13373,N_12952,N_12392);
and U13374 (N_13374,N_12997,N_12834);
and U13375 (N_13375,N_12135,N_12884);
or U13376 (N_13376,N_12720,N_12931);
nor U13377 (N_13377,N_12755,N_12396);
nand U13378 (N_13378,N_12514,N_12990);
nor U13379 (N_13379,N_12524,N_12257);
xor U13380 (N_13380,N_12312,N_12861);
nor U13381 (N_13381,N_12882,N_12587);
and U13382 (N_13382,N_12124,N_12082);
or U13383 (N_13383,N_12580,N_12420);
nand U13384 (N_13384,N_12335,N_12679);
or U13385 (N_13385,N_12034,N_12001);
nand U13386 (N_13386,N_12809,N_12178);
nand U13387 (N_13387,N_12503,N_12602);
xor U13388 (N_13388,N_12293,N_12075);
nor U13389 (N_13389,N_12837,N_12314);
nand U13390 (N_13390,N_12718,N_12004);
xor U13391 (N_13391,N_12462,N_12998);
nand U13392 (N_13392,N_12322,N_12255);
nand U13393 (N_13393,N_12324,N_12422);
nand U13394 (N_13394,N_12932,N_12233);
nor U13395 (N_13395,N_12094,N_12694);
nor U13396 (N_13396,N_12872,N_12786);
nor U13397 (N_13397,N_12119,N_12796);
nor U13398 (N_13398,N_12307,N_12575);
xor U13399 (N_13399,N_12787,N_12358);
nand U13400 (N_13400,N_12808,N_12449);
nand U13401 (N_13401,N_12499,N_12792);
or U13402 (N_13402,N_12553,N_12897);
nand U13403 (N_13403,N_12167,N_12788);
and U13404 (N_13404,N_12336,N_12325);
xor U13405 (N_13405,N_12564,N_12051);
nor U13406 (N_13406,N_12653,N_12429);
xor U13407 (N_13407,N_12476,N_12084);
or U13408 (N_13408,N_12318,N_12049);
nor U13409 (N_13409,N_12545,N_12244);
nor U13410 (N_13410,N_12493,N_12529);
or U13411 (N_13411,N_12858,N_12161);
or U13412 (N_13412,N_12781,N_12136);
and U13413 (N_13413,N_12303,N_12454);
and U13414 (N_13414,N_12389,N_12584);
nor U13415 (N_13415,N_12491,N_12472);
xor U13416 (N_13416,N_12151,N_12492);
nand U13417 (N_13417,N_12090,N_12115);
xnor U13418 (N_13418,N_12676,N_12901);
or U13419 (N_13419,N_12480,N_12818);
xor U13420 (N_13420,N_12201,N_12002);
or U13421 (N_13421,N_12548,N_12993);
nor U13422 (N_13422,N_12807,N_12345);
or U13423 (N_13423,N_12038,N_12908);
xor U13424 (N_13424,N_12134,N_12321);
xnor U13425 (N_13425,N_12988,N_12567);
and U13426 (N_13426,N_12568,N_12513);
or U13427 (N_13427,N_12698,N_12980);
or U13428 (N_13428,N_12148,N_12820);
nand U13429 (N_13429,N_12557,N_12162);
nand U13430 (N_13430,N_12425,N_12208);
nand U13431 (N_13431,N_12473,N_12565);
xnor U13432 (N_13432,N_12948,N_12185);
or U13433 (N_13433,N_12450,N_12426);
nand U13434 (N_13434,N_12588,N_12200);
nor U13435 (N_13435,N_12962,N_12501);
nand U13436 (N_13436,N_12735,N_12230);
nand U13437 (N_13437,N_12217,N_12635);
and U13438 (N_13438,N_12355,N_12804);
nor U13439 (N_13439,N_12418,N_12423);
nand U13440 (N_13440,N_12291,N_12864);
or U13441 (N_13441,N_12102,N_12910);
or U13442 (N_13442,N_12537,N_12459);
xor U13443 (N_13443,N_12280,N_12023);
nand U13444 (N_13444,N_12619,N_12039);
xnor U13445 (N_13445,N_12256,N_12842);
nand U13446 (N_13446,N_12496,N_12270);
nand U13447 (N_13447,N_12955,N_12642);
and U13448 (N_13448,N_12095,N_12934);
or U13449 (N_13449,N_12475,N_12867);
nor U13450 (N_13450,N_12125,N_12451);
nor U13451 (N_13451,N_12470,N_12992);
xnor U13452 (N_13452,N_12191,N_12887);
xor U13453 (N_13453,N_12585,N_12432);
xor U13454 (N_13454,N_12328,N_12397);
nor U13455 (N_13455,N_12697,N_12763);
nand U13456 (N_13456,N_12067,N_12774);
nand U13457 (N_13457,N_12814,N_12531);
xor U13458 (N_13458,N_12817,N_12984);
nand U13459 (N_13459,N_12024,N_12385);
and U13460 (N_13460,N_12590,N_12767);
nor U13461 (N_13461,N_12750,N_12436);
or U13462 (N_13462,N_12439,N_12829);
or U13463 (N_13463,N_12279,N_12856);
nor U13464 (N_13464,N_12560,N_12957);
or U13465 (N_13465,N_12495,N_12776);
nand U13466 (N_13466,N_12031,N_12487);
nand U13467 (N_13467,N_12999,N_12747);
or U13468 (N_13468,N_12833,N_12214);
nand U13469 (N_13469,N_12456,N_12269);
nand U13470 (N_13470,N_12203,N_12490);
nor U13471 (N_13471,N_12509,N_12764);
or U13472 (N_13472,N_12243,N_12507);
and U13473 (N_13473,N_12958,N_12632);
or U13474 (N_13474,N_12412,N_12648);
nor U13475 (N_13475,N_12534,N_12262);
and U13476 (N_13476,N_12836,N_12977);
nand U13477 (N_13477,N_12371,N_12721);
or U13478 (N_13478,N_12558,N_12960);
or U13479 (N_13479,N_12424,N_12258);
nand U13480 (N_13480,N_12139,N_12061);
xnor U13481 (N_13481,N_12171,N_12569);
or U13482 (N_13482,N_12983,N_12505);
nand U13483 (N_13483,N_12976,N_12137);
xnor U13484 (N_13484,N_12525,N_12751);
nand U13485 (N_13485,N_12111,N_12131);
nor U13486 (N_13486,N_12232,N_12343);
nand U13487 (N_13487,N_12903,N_12863);
nand U13488 (N_13488,N_12159,N_12681);
nor U13489 (N_13489,N_12623,N_12101);
xnor U13490 (N_13490,N_12573,N_12263);
and U13491 (N_13491,N_12673,N_12706);
or U13492 (N_13492,N_12949,N_12277);
nand U13493 (N_13493,N_12170,N_12250);
nor U13494 (N_13494,N_12267,N_12968);
nor U13495 (N_13495,N_12453,N_12674);
nor U13496 (N_13496,N_12029,N_12445);
nand U13497 (N_13497,N_12656,N_12862);
or U13498 (N_13498,N_12215,N_12443);
nand U13499 (N_13499,N_12494,N_12435);
nor U13500 (N_13500,N_12957,N_12837);
xor U13501 (N_13501,N_12139,N_12680);
xnor U13502 (N_13502,N_12620,N_12648);
nor U13503 (N_13503,N_12050,N_12700);
or U13504 (N_13504,N_12361,N_12676);
xnor U13505 (N_13505,N_12860,N_12050);
nor U13506 (N_13506,N_12630,N_12101);
xor U13507 (N_13507,N_12783,N_12333);
and U13508 (N_13508,N_12878,N_12599);
nand U13509 (N_13509,N_12153,N_12716);
nand U13510 (N_13510,N_12669,N_12363);
xor U13511 (N_13511,N_12067,N_12491);
or U13512 (N_13512,N_12734,N_12143);
or U13513 (N_13513,N_12314,N_12291);
and U13514 (N_13514,N_12162,N_12499);
nor U13515 (N_13515,N_12379,N_12513);
or U13516 (N_13516,N_12985,N_12305);
and U13517 (N_13517,N_12215,N_12816);
xor U13518 (N_13518,N_12015,N_12131);
nand U13519 (N_13519,N_12468,N_12093);
nand U13520 (N_13520,N_12284,N_12841);
nand U13521 (N_13521,N_12036,N_12198);
or U13522 (N_13522,N_12492,N_12941);
or U13523 (N_13523,N_12049,N_12545);
or U13524 (N_13524,N_12418,N_12449);
and U13525 (N_13525,N_12134,N_12910);
nor U13526 (N_13526,N_12713,N_12879);
nand U13527 (N_13527,N_12266,N_12759);
xor U13528 (N_13528,N_12416,N_12704);
or U13529 (N_13529,N_12255,N_12958);
xnor U13530 (N_13530,N_12858,N_12801);
xnor U13531 (N_13531,N_12812,N_12174);
or U13532 (N_13532,N_12045,N_12572);
xnor U13533 (N_13533,N_12975,N_12301);
or U13534 (N_13534,N_12275,N_12973);
or U13535 (N_13535,N_12458,N_12420);
nor U13536 (N_13536,N_12211,N_12826);
or U13537 (N_13537,N_12320,N_12462);
and U13538 (N_13538,N_12763,N_12742);
xnor U13539 (N_13539,N_12220,N_12350);
xor U13540 (N_13540,N_12594,N_12613);
nand U13541 (N_13541,N_12165,N_12151);
nor U13542 (N_13542,N_12048,N_12153);
nor U13543 (N_13543,N_12936,N_12120);
nor U13544 (N_13544,N_12956,N_12842);
and U13545 (N_13545,N_12360,N_12066);
or U13546 (N_13546,N_12423,N_12491);
and U13547 (N_13547,N_12431,N_12580);
and U13548 (N_13548,N_12885,N_12290);
xnor U13549 (N_13549,N_12438,N_12384);
or U13550 (N_13550,N_12089,N_12909);
nand U13551 (N_13551,N_12213,N_12165);
or U13552 (N_13552,N_12874,N_12354);
xnor U13553 (N_13553,N_12150,N_12635);
xnor U13554 (N_13554,N_12994,N_12455);
nand U13555 (N_13555,N_12000,N_12384);
or U13556 (N_13556,N_12289,N_12221);
and U13557 (N_13557,N_12535,N_12396);
nand U13558 (N_13558,N_12575,N_12506);
and U13559 (N_13559,N_12720,N_12618);
xnor U13560 (N_13560,N_12558,N_12455);
nand U13561 (N_13561,N_12610,N_12684);
nand U13562 (N_13562,N_12528,N_12135);
and U13563 (N_13563,N_12009,N_12557);
xor U13564 (N_13564,N_12306,N_12745);
xor U13565 (N_13565,N_12455,N_12344);
xnor U13566 (N_13566,N_12656,N_12689);
xor U13567 (N_13567,N_12219,N_12778);
or U13568 (N_13568,N_12005,N_12069);
xor U13569 (N_13569,N_12790,N_12614);
and U13570 (N_13570,N_12321,N_12136);
xnor U13571 (N_13571,N_12359,N_12235);
nand U13572 (N_13572,N_12564,N_12174);
nor U13573 (N_13573,N_12177,N_12590);
or U13574 (N_13574,N_12919,N_12716);
and U13575 (N_13575,N_12968,N_12942);
and U13576 (N_13576,N_12331,N_12239);
or U13577 (N_13577,N_12471,N_12270);
nor U13578 (N_13578,N_12048,N_12058);
nor U13579 (N_13579,N_12078,N_12394);
and U13580 (N_13580,N_12857,N_12320);
nand U13581 (N_13581,N_12797,N_12550);
nor U13582 (N_13582,N_12761,N_12431);
and U13583 (N_13583,N_12563,N_12813);
nor U13584 (N_13584,N_12978,N_12068);
xnor U13585 (N_13585,N_12730,N_12695);
nand U13586 (N_13586,N_12739,N_12469);
and U13587 (N_13587,N_12510,N_12830);
nor U13588 (N_13588,N_12699,N_12791);
nor U13589 (N_13589,N_12476,N_12538);
or U13590 (N_13590,N_12923,N_12792);
nand U13591 (N_13591,N_12601,N_12044);
or U13592 (N_13592,N_12752,N_12877);
xor U13593 (N_13593,N_12481,N_12583);
or U13594 (N_13594,N_12538,N_12306);
and U13595 (N_13595,N_12735,N_12109);
and U13596 (N_13596,N_12695,N_12134);
nand U13597 (N_13597,N_12409,N_12286);
and U13598 (N_13598,N_12977,N_12795);
and U13599 (N_13599,N_12739,N_12780);
or U13600 (N_13600,N_12546,N_12953);
nor U13601 (N_13601,N_12365,N_12368);
nand U13602 (N_13602,N_12572,N_12384);
xnor U13603 (N_13603,N_12773,N_12153);
xnor U13604 (N_13604,N_12549,N_12910);
nand U13605 (N_13605,N_12356,N_12750);
nand U13606 (N_13606,N_12904,N_12778);
or U13607 (N_13607,N_12889,N_12457);
xor U13608 (N_13608,N_12006,N_12590);
or U13609 (N_13609,N_12946,N_12828);
nand U13610 (N_13610,N_12164,N_12504);
nand U13611 (N_13611,N_12480,N_12248);
or U13612 (N_13612,N_12469,N_12374);
nor U13613 (N_13613,N_12508,N_12031);
nor U13614 (N_13614,N_12392,N_12692);
nand U13615 (N_13615,N_12929,N_12740);
xnor U13616 (N_13616,N_12281,N_12236);
nor U13617 (N_13617,N_12198,N_12831);
nor U13618 (N_13618,N_12995,N_12413);
xnor U13619 (N_13619,N_12282,N_12313);
and U13620 (N_13620,N_12526,N_12525);
xor U13621 (N_13621,N_12239,N_12120);
or U13622 (N_13622,N_12763,N_12906);
or U13623 (N_13623,N_12600,N_12696);
xnor U13624 (N_13624,N_12625,N_12063);
xor U13625 (N_13625,N_12927,N_12559);
and U13626 (N_13626,N_12783,N_12938);
or U13627 (N_13627,N_12926,N_12301);
and U13628 (N_13628,N_12332,N_12106);
xnor U13629 (N_13629,N_12440,N_12276);
and U13630 (N_13630,N_12122,N_12652);
nor U13631 (N_13631,N_12825,N_12775);
xor U13632 (N_13632,N_12494,N_12324);
or U13633 (N_13633,N_12937,N_12705);
xor U13634 (N_13634,N_12958,N_12097);
xor U13635 (N_13635,N_12108,N_12821);
or U13636 (N_13636,N_12635,N_12373);
nor U13637 (N_13637,N_12452,N_12343);
and U13638 (N_13638,N_12914,N_12365);
nand U13639 (N_13639,N_12910,N_12019);
nor U13640 (N_13640,N_12981,N_12916);
or U13641 (N_13641,N_12702,N_12225);
nor U13642 (N_13642,N_12429,N_12976);
nor U13643 (N_13643,N_12688,N_12754);
xor U13644 (N_13644,N_12016,N_12396);
xnor U13645 (N_13645,N_12470,N_12214);
nor U13646 (N_13646,N_12328,N_12520);
or U13647 (N_13647,N_12071,N_12853);
nor U13648 (N_13648,N_12845,N_12713);
or U13649 (N_13649,N_12283,N_12734);
or U13650 (N_13650,N_12463,N_12973);
xnor U13651 (N_13651,N_12300,N_12575);
and U13652 (N_13652,N_12424,N_12363);
nand U13653 (N_13653,N_12299,N_12337);
xnor U13654 (N_13654,N_12090,N_12048);
and U13655 (N_13655,N_12565,N_12846);
and U13656 (N_13656,N_12354,N_12400);
or U13657 (N_13657,N_12474,N_12233);
and U13658 (N_13658,N_12293,N_12510);
nand U13659 (N_13659,N_12808,N_12342);
nand U13660 (N_13660,N_12409,N_12332);
or U13661 (N_13661,N_12647,N_12099);
xor U13662 (N_13662,N_12942,N_12615);
nand U13663 (N_13663,N_12461,N_12381);
nor U13664 (N_13664,N_12224,N_12190);
nand U13665 (N_13665,N_12134,N_12804);
and U13666 (N_13666,N_12047,N_12722);
nor U13667 (N_13667,N_12667,N_12170);
and U13668 (N_13668,N_12112,N_12667);
and U13669 (N_13669,N_12182,N_12189);
xor U13670 (N_13670,N_12797,N_12004);
nand U13671 (N_13671,N_12254,N_12344);
xnor U13672 (N_13672,N_12309,N_12823);
nand U13673 (N_13673,N_12162,N_12935);
and U13674 (N_13674,N_12899,N_12829);
or U13675 (N_13675,N_12043,N_12012);
or U13676 (N_13676,N_12213,N_12793);
nand U13677 (N_13677,N_12923,N_12613);
or U13678 (N_13678,N_12061,N_12275);
nor U13679 (N_13679,N_12839,N_12060);
xnor U13680 (N_13680,N_12326,N_12515);
nor U13681 (N_13681,N_12179,N_12195);
nand U13682 (N_13682,N_12358,N_12029);
nor U13683 (N_13683,N_12959,N_12932);
nand U13684 (N_13684,N_12828,N_12139);
xor U13685 (N_13685,N_12142,N_12757);
or U13686 (N_13686,N_12280,N_12050);
xor U13687 (N_13687,N_12481,N_12504);
xor U13688 (N_13688,N_12736,N_12780);
nor U13689 (N_13689,N_12418,N_12733);
xor U13690 (N_13690,N_12571,N_12974);
xor U13691 (N_13691,N_12959,N_12893);
and U13692 (N_13692,N_12522,N_12941);
nor U13693 (N_13693,N_12792,N_12726);
and U13694 (N_13694,N_12722,N_12455);
nor U13695 (N_13695,N_12817,N_12254);
xnor U13696 (N_13696,N_12148,N_12131);
nor U13697 (N_13697,N_12884,N_12968);
nand U13698 (N_13698,N_12525,N_12036);
nor U13699 (N_13699,N_12844,N_12697);
xnor U13700 (N_13700,N_12052,N_12960);
or U13701 (N_13701,N_12813,N_12722);
xnor U13702 (N_13702,N_12962,N_12664);
nor U13703 (N_13703,N_12606,N_12754);
or U13704 (N_13704,N_12870,N_12406);
nand U13705 (N_13705,N_12422,N_12546);
nor U13706 (N_13706,N_12258,N_12720);
xnor U13707 (N_13707,N_12354,N_12986);
xnor U13708 (N_13708,N_12376,N_12470);
xnor U13709 (N_13709,N_12708,N_12338);
or U13710 (N_13710,N_12249,N_12475);
nor U13711 (N_13711,N_12359,N_12834);
or U13712 (N_13712,N_12213,N_12327);
nor U13713 (N_13713,N_12228,N_12556);
xor U13714 (N_13714,N_12296,N_12286);
and U13715 (N_13715,N_12735,N_12051);
or U13716 (N_13716,N_12933,N_12917);
or U13717 (N_13717,N_12374,N_12946);
nand U13718 (N_13718,N_12252,N_12498);
and U13719 (N_13719,N_12027,N_12447);
xor U13720 (N_13720,N_12257,N_12683);
xnor U13721 (N_13721,N_12244,N_12732);
nand U13722 (N_13722,N_12698,N_12266);
xnor U13723 (N_13723,N_12286,N_12900);
or U13724 (N_13724,N_12115,N_12409);
or U13725 (N_13725,N_12837,N_12506);
nor U13726 (N_13726,N_12018,N_12779);
or U13727 (N_13727,N_12256,N_12679);
nor U13728 (N_13728,N_12295,N_12188);
and U13729 (N_13729,N_12399,N_12485);
xnor U13730 (N_13730,N_12626,N_12846);
nand U13731 (N_13731,N_12502,N_12538);
and U13732 (N_13732,N_12448,N_12254);
nand U13733 (N_13733,N_12755,N_12536);
and U13734 (N_13734,N_12217,N_12991);
nor U13735 (N_13735,N_12048,N_12284);
nand U13736 (N_13736,N_12019,N_12009);
and U13737 (N_13737,N_12230,N_12348);
or U13738 (N_13738,N_12781,N_12525);
nor U13739 (N_13739,N_12066,N_12570);
nand U13740 (N_13740,N_12723,N_12384);
nor U13741 (N_13741,N_12598,N_12481);
xnor U13742 (N_13742,N_12472,N_12717);
nand U13743 (N_13743,N_12864,N_12234);
and U13744 (N_13744,N_12561,N_12337);
or U13745 (N_13745,N_12475,N_12760);
nand U13746 (N_13746,N_12770,N_12015);
and U13747 (N_13747,N_12618,N_12387);
nor U13748 (N_13748,N_12375,N_12040);
xor U13749 (N_13749,N_12765,N_12440);
or U13750 (N_13750,N_12971,N_12925);
or U13751 (N_13751,N_12831,N_12482);
xor U13752 (N_13752,N_12632,N_12560);
nor U13753 (N_13753,N_12726,N_12148);
xnor U13754 (N_13754,N_12103,N_12555);
nand U13755 (N_13755,N_12302,N_12464);
nor U13756 (N_13756,N_12383,N_12438);
xor U13757 (N_13757,N_12244,N_12423);
and U13758 (N_13758,N_12510,N_12268);
nor U13759 (N_13759,N_12305,N_12668);
and U13760 (N_13760,N_12159,N_12138);
nand U13761 (N_13761,N_12918,N_12502);
or U13762 (N_13762,N_12911,N_12836);
xnor U13763 (N_13763,N_12480,N_12395);
xnor U13764 (N_13764,N_12362,N_12097);
nor U13765 (N_13765,N_12278,N_12411);
nor U13766 (N_13766,N_12991,N_12791);
nand U13767 (N_13767,N_12901,N_12007);
xor U13768 (N_13768,N_12827,N_12726);
and U13769 (N_13769,N_12076,N_12313);
xnor U13770 (N_13770,N_12798,N_12467);
xor U13771 (N_13771,N_12512,N_12539);
xor U13772 (N_13772,N_12567,N_12195);
nor U13773 (N_13773,N_12772,N_12163);
xor U13774 (N_13774,N_12723,N_12831);
xnor U13775 (N_13775,N_12173,N_12028);
nand U13776 (N_13776,N_12489,N_12518);
xnor U13777 (N_13777,N_12866,N_12347);
and U13778 (N_13778,N_12924,N_12138);
or U13779 (N_13779,N_12135,N_12554);
nor U13780 (N_13780,N_12268,N_12758);
nand U13781 (N_13781,N_12677,N_12602);
and U13782 (N_13782,N_12053,N_12038);
nor U13783 (N_13783,N_12356,N_12875);
nor U13784 (N_13784,N_12334,N_12213);
nor U13785 (N_13785,N_12388,N_12378);
nand U13786 (N_13786,N_12747,N_12239);
nand U13787 (N_13787,N_12094,N_12299);
nand U13788 (N_13788,N_12464,N_12901);
or U13789 (N_13789,N_12066,N_12277);
and U13790 (N_13790,N_12021,N_12698);
nor U13791 (N_13791,N_12821,N_12161);
and U13792 (N_13792,N_12362,N_12831);
or U13793 (N_13793,N_12346,N_12840);
and U13794 (N_13794,N_12820,N_12452);
and U13795 (N_13795,N_12069,N_12555);
nor U13796 (N_13796,N_12326,N_12110);
and U13797 (N_13797,N_12433,N_12443);
or U13798 (N_13798,N_12031,N_12488);
or U13799 (N_13799,N_12971,N_12363);
or U13800 (N_13800,N_12200,N_12289);
nor U13801 (N_13801,N_12800,N_12549);
xor U13802 (N_13802,N_12133,N_12014);
nor U13803 (N_13803,N_12560,N_12784);
nor U13804 (N_13804,N_12390,N_12760);
nor U13805 (N_13805,N_12567,N_12268);
xor U13806 (N_13806,N_12262,N_12501);
nor U13807 (N_13807,N_12934,N_12716);
nand U13808 (N_13808,N_12320,N_12163);
or U13809 (N_13809,N_12252,N_12239);
xor U13810 (N_13810,N_12901,N_12490);
or U13811 (N_13811,N_12457,N_12445);
nand U13812 (N_13812,N_12156,N_12883);
or U13813 (N_13813,N_12181,N_12354);
nor U13814 (N_13814,N_12845,N_12102);
or U13815 (N_13815,N_12352,N_12690);
xnor U13816 (N_13816,N_12772,N_12881);
and U13817 (N_13817,N_12841,N_12781);
or U13818 (N_13818,N_12678,N_12960);
nand U13819 (N_13819,N_12400,N_12648);
and U13820 (N_13820,N_12548,N_12752);
nand U13821 (N_13821,N_12768,N_12659);
and U13822 (N_13822,N_12324,N_12461);
nand U13823 (N_13823,N_12845,N_12198);
nand U13824 (N_13824,N_12958,N_12573);
nand U13825 (N_13825,N_12709,N_12325);
nor U13826 (N_13826,N_12539,N_12091);
and U13827 (N_13827,N_12235,N_12445);
nor U13828 (N_13828,N_12885,N_12287);
and U13829 (N_13829,N_12521,N_12510);
or U13830 (N_13830,N_12211,N_12478);
xor U13831 (N_13831,N_12773,N_12250);
or U13832 (N_13832,N_12271,N_12383);
and U13833 (N_13833,N_12449,N_12922);
and U13834 (N_13834,N_12636,N_12110);
nand U13835 (N_13835,N_12787,N_12650);
nor U13836 (N_13836,N_12798,N_12464);
nor U13837 (N_13837,N_12659,N_12616);
xor U13838 (N_13838,N_12269,N_12032);
xor U13839 (N_13839,N_12835,N_12246);
or U13840 (N_13840,N_12377,N_12418);
nor U13841 (N_13841,N_12127,N_12209);
and U13842 (N_13842,N_12284,N_12320);
nor U13843 (N_13843,N_12352,N_12060);
nor U13844 (N_13844,N_12114,N_12803);
xnor U13845 (N_13845,N_12512,N_12514);
and U13846 (N_13846,N_12227,N_12467);
or U13847 (N_13847,N_12378,N_12428);
or U13848 (N_13848,N_12697,N_12987);
and U13849 (N_13849,N_12372,N_12498);
and U13850 (N_13850,N_12639,N_12921);
xor U13851 (N_13851,N_12022,N_12400);
nor U13852 (N_13852,N_12836,N_12468);
nor U13853 (N_13853,N_12022,N_12943);
and U13854 (N_13854,N_12889,N_12202);
nor U13855 (N_13855,N_12222,N_12480);
nand U13856 (N_13856,N_12721,N_12043);
and U13857 (N_13857,N_12363,N_12941);
nand U13858 (N_13858,N_12562,N_12624);
nand U13859 (N_13859,N_12043,N_12541);
and U13860 (N_13860,N_12542,N_12221);
or U13861 (N_13861,N_12589,N_12510);
or U13862 (N_13862,N_12897,N_12352);
nor U13863 (N_13863,N_12305,N_12842);
nor U13864 (N_13864,N_12985,N_12481);
xor U13865 (N_13865,N_12277,N_12417);
or U13866 (N_13866,N_12479,N_12757);
or U13867 (N_13867,N_12017,N_12351);
and U13868 (N_13868,N_12253,N_12252);
and U13869 (N_13869,N_12990,N_12295);
and U13870 (N_13870,N_12025,N_12743);
xor U13871 (N_13871,N_12564,N_12258);
xnor U13872 (N_13872,N_12040,N_12640);
or U13873 (N_13873,N_12070,N_12974);
or U13874 (N_13874,N_12653,N_12350);
or U13875 (N_13875,N_12880,N_12212);
nor U13876 (N_13876,N_12015,N_12161);
and U13877 (N_13877,N_12248,N_12915);
xnor U13878 (N_13878,N_12681,N_12796);
nand U13879 (N_13879,N_12792,N_12752);
nor U13880 (N_13880,N_12746,N_12172);
xnor U13881 (N_13881,N_12931,N_12722);
nor U13882 (N_13882,N_12341,N_12491);
nor U13883 (N_13883,N_12753,N_12208);
and U13884 (N_13884,N_12435,N_12146);
and U13885 (N_13885,N_12714,N_12109);
and U13886 (N_13886,N_12005,N_12756);
xor U13887 (N_13887,N_12654,N_12053);
or U13888 (N_13888,N_12539,N_12863);
or U13889 (N_13889,N_12740,N_12475);
nor U13890 (N_13890,N_12616,N_12308);
nor U13891 (N_13891,N_12047,N_12172);
nand U13892 (N_13892,N_12719,N_12579);
or U13893 (N_13893,N_12604,N_12196);
nand U13894 (N_13894,N_12272,N_12163);
nor U13895 (N_13895,N_12332,N_12972);
xor U13896 (N_13896,N_12385,N_12511);
and U13897 (N_13897,N_12395,N_12925);
xor U13898 (N_13898,N_12552,N_12786);
nor U13899 (N_13899,N_12490,N_12454);
and U13900 (N_13900,N_12192,N_12442);
nand U13901 (N_13901,N_12398,N_12695);
or U13902 (N_13902,N_12069,N_12007);
xor U13903 (N_13903,N_12528,N_12378);
nand U13904 (N_13904,N_12086,N_12361);
nor U13905 (N_13905,N_12610,N_12928);
and U13906 (N_13906,N_12633,N_12510);
nor U13907 (N_13907,N_12039,N_12987);
and U13908 (N_13908,N_12743,N_12584);
or U13909 (N_13909,N_12644,N_12365);
and U13910 (N_13910,N_12058,N_12755);
or U13911 (N_13911,N_12947,N_12185);
nand U13912 (N_13912,N_12935,N_12813);
and U13913 (N_13913,N_12668,N_12487);
nor U13914 (N_13914,N_12315,N_12023);
or U13915 (N_13915,N_12814,N_12521);
and U13916 (N_13916,N_12656,N_12848);
nand U13917 (N_13917,N_12858,N_12787);
nand U13918 (N_13918,N_12977,N_12357);
and U13919 (N_13919,N_12978,N_12469);
nand U13920 (N_13920,N_12051,N_12755);
nor U13921 (N_13921,N_12787,N_12490);
or U13922 (N_13922,N_12249,N_12741);
and U13923 (N_13923,N_12437,N_12970);
nor U13924 (N_13924,N_12156,N_12500);
nand U13925 (N_13925,N_12369,N_12624);
nor U13926 (N_13926,N_12051,N_12315);
and U13927 (N_13927,N_12472,N_12569);
and U13928 (N_13928,N_12724,N_12132);
nand U13929 (N_13929,N_12696,N_12527);
or U13930 (N_13930,N_12155,N_12808);
nand U13931 (N_13931,N_12083,N_12166);
xnor U13932 (N_13932,N_12616,N_12513);
nand U13933 (N_13933,N_12195,N_12845);
nor U13934 (N_13934,N_12178,N_12879);
xor U13935 (N_13935,N_12797,N_12460);
or U13936 (N_13936,N_12827,N_12991);
or U13937 (N_13937,N_12846,N_12533);
or U13938 (N_13938,N_12965,N_12311);
and U13939 (N_13939,N_12576,N_12341);
and U13940 (N_13940,N_12934,N_12540);
nand U13941 (N_13941,N_12798,N_12764);
xnor U13942 (N_13942,N_12626,N_12754);
and U13943 (N_13943,N_12439,N_12256);
nand U13944 (N_13944,N_12744,N_12737);
nor U13945 (N_13945,N_12481,N_12696);
nand U13946 (N_13946,N_12447,N_12431);
xnor U13947 (N_13947,N_12675,N_12640);
and U13948 (N_13948,N_12791,N_12684);
nor U13949 (N_13949,N_12412,N_12842);
nand U13950 (N_13950,N_12183,N_12742);
or U13951 (N_13951,N_12296,N_12728);
or U13952 (N_13952,N_12727,N_12898);
and U13953 (N_13953,N_12488,N_12426);
and U13954 (N_13954,N_12399,N_12634);
or U13955 (N_13955,N_12739,N_12249);
and U13956 (N_13956,N_12002,N_12012);
nand U13957 (N_13957,N_12376,N_12027);
nand U13958 (N_13958,N_12648,N_12538);
or U13959 (N_13959,N_12770,N_12834);
xor U13960 (N_13960,N_12879,N_12756);
nand U13961 (N_13961,N_12493,N_12896);
xor U13962 (N_13962,N_12835,N_12273);
nor U13963 (N_13963,N_12407,N_12076);
xor U13964 (N_13964,N_12593,N_12878);
xor U13965 (N_13965,N_12558,N_12397);
and U13966 (N_13966,N_12457,N_12779);
or U13967 (N_13967,N_12390,N_12991);
nand U13968 (N_13968,N_12569,N_12546);
nor U13969 (N_13969,N_12897,N_12769);
nand U13970 (N_13970,N_12470,N_12761);
nand U13971 (N_13971,N_12389,N_12632);
or U13972 (N_13972,N_12939,N_12479);
and U13973 (N_13973,N_12542,N_12795);
and U13974 (N_13974,N_12320,N_12456);
xnor U13975 (N_13975,N_12103,N_12216);
nor U13976 (N_13976,N_12969,N_12842);
nor U13977 (N_13977,N_12141,N_12257);
xor U13978 (N_13978,N_12926,N_12536);
xnor U13979 (N_13979,N_12624,N_12311);
and U13980 (N_13980,N_12549,N_12473);
or U13981 (N_13981,N_12358,N_12604);
or U13982 (N_13982,N_12060,N_12616);
or U13983 (N_13983,N_12060,N_12045);
nand U13984 (N_13984,N_12227,N_12842);
and U13985 (N_13985,N_12863,N_12993);
or U13986 (N_13986,N_12941,N_12434);
or U13987 (N_13987,N_12215,N_12515);
nand U13988 (N_13988,N_12231,N_12111);
and U13989 (N_13989,N_12584,N_12026);
xor U13990 (N_13990,N_12852,N_12108);
and U13991 (N_13991,N_12452,N_12904);
or U13992 (N_13992,N_12215,N_12701);
nor U13993 (N_13993,N_12310,N_12822);
nand U13994 (N_13994,N_12943,N_12009);
nor U13995 (N_13995,N_12158,N_12777);
and U13996 (N_13996,N_12491,N_12820);
nand U13997 (N_13997,N_12650,N_12640);
xor U13998 (N_13998,N_12822,N_12600);
or U13999 (N_13999,N_12772,N_12263);
xor U14000 (N_14000,N_13190,N_13113);
nor U14001 (N_14001,N_13672,N_13577);
nor U14002 (N_14002,N_13624,N_13952);
xor U14003 (N_14003,N_13681,N_13739);
nand U14004 (N_14004,N_13000,N_13518);
xnor U14005 (N_14005,N_13875,N_13640);
nor U14006 (N_14006,N_13993,N_13852);
and U14007 (N_14007,N_13399,N_13830);
and U14008 (N_14008,N_13569,N_13509);
nand U14009 (N_14009,N_13460,N_13213);
and U14010 (N_14010,N_13598,N_13345);
xor U14011 (N_14011,N_13006,N_13408);
or U14012 (N_14012,N_13118,N_13825);
nand U14013 (N_14013,N_13948,N_13103);
and U14014 (N_14014,N_13706,N_13058);
nand U14015 (N_14015,N_13230,N_13140);
nand U14016 (N_14016,N_13304,N_13588);
and U14017 (N_14017,N_13652,N_13034);
nand U14018 (N_14018,N_13774,N_13650);
nand U14019 (N_14019,N_13777,N_13620);
xnor U14020 (N_14020,N_13032,N_13425);
xnor U14021 (N_14021,N_13307,N_13347);
or U14022 (N_14022,N_13222,N_13963);
nand U14023 (N_14023,N_13236,N_13584);
and U14024 (N_14024,N_13075,N_13506);
xnor U14025 (N_14025,N_13623,N_13242);
and U14026 (N_14026,N_13269,N_13836);
xnor U14027 (N_14027,N_13607,N_13265);
xnor U14028 (N_14028,N_13651,N_13784);
or U14029 (N_14029,N_13478,N_13004);
xor U14030 (N_14030,N_13386,N_13497);
and U14031 (N_14031,N_13746,N_13821);
nand U14032 (N_14032,N_13332,N_13532);
nor U14033 (N_14033,N_13363,N_13889);
nor U14034 (N_14034,N_13750,N_13763);
xor U14035 (N_14035,N_13978,N_13248);
nand U14036 (N_14036,N_13559,N_13091);
nor U14037 (N_14037,N_13234,N_13790);
xnor U14038 (N_14038,N_13418,N_13301);
nor U14039 (N_14039,N_13964,N_13522);
nand U14040 (N_14040,N_13106,N_13197);
or U14041 (N_14041,N_13144,N_13052);
and U14042 (N_14042,N_13011,N_13877);
xor U14043 (N_14043,N_13828,N_13949);
or U14044 (N_14044,N_13547,N_13918);
or U14045 (N_14045,N_13759,N_13531);
nand U14046 (N_14046,N_13002,N_13170);
xor U14047 (N_14047,N_13558,N_13528);
nor U14048 (N_14048,N_13553,N_13226);
or U14049 (N_14049,N_13663,N_13811);
xnor U14050 (N_14050,N_13153,N_13896);
and U14051 (N_14051,N_13074,N_13675);
xnor U14052 (N_14052,N_13917,N_13289);
or U14053 (N_14053,N_13986,N_13618);
xor U14054 (N_14054,N_13054,N_13717);
xnor U14055 (N_14055,N_13406,N_13127);
nor U14056 (N_14056,N_13692,N_13676);
nand U14057 (N_14057,N_13606,N_13600);
nand U14058 (N_14058,N_13229,N_13449);
nand U14059 (N_14059,N_13057,N_13589);
xor U14060 (N_14060,N_13070,N_13177);
or U14061 (N_14061,N_13669,N_13521);
and U14062 (N_14062,N_13326,N_13429);
nand U14063 (N_14063,N_13239,N_13255);
xnor U14064 (N_14064,N_13491,N_13945);
xnor U14065 (N_14065,N_13366,N_13719);
nand U14066 (N_14066,N_13446,N_13130);
nor U14067 (N_14067,N_13101,N_13319);
and U14068 (N_14068,N_13609,N_13415);
and U14069 (N_14069,N_13880,N_13299);
and U14070 (N_14070,N_13235,N_13227);
nor U14071 (N_14071,N_13359,N_13554);
nor U14072 (N_14072,N_13555,N_13857);
and U14073 (N_14073,N_13966,N_13556);
xnor U14074 (N_14074,N_13303,N_13733);
or U14075 (N_14075,N_13368,N_13817);
or U14076 (N_14076,N_13925,N_13349);
nand U14077 (N_14077,N_13404,N_13832);
and U14078 (N_14078,N_13803,N_13295);
xnor U14079 (N_14079,N_13934,N_13040);
and U14080 (N_14080,N_13346,N_13022);
or U14081 (N_14081,N_13268,N_13357);
nand U14082 (N_14082,N_13284,N_13954);
and U14083 (N_14083,N_13796,N_13597);
nand U14084 (N_14084,N_13145,N_13036);
and U14085 (N_14085,N_13988,N_13968);
nand U14086 (N_14086,N_13693,N_13016);
and U14087 (N_14087,N_13341,N_13695);
or U14088 (N_14088,N_13690,N_13160);
or U14089 (N_14089,N_13174,N_13715);
nand U14090 (N_14090,N_13855,N_13178);
nor U14091 (N_14091,N_13822,N_13231);
nand U14092 (N_14092,N_13493,N_13383);
and U14093 (N_14093,N_13646,N_13061);
or U14094 (N_14094,N_13604,N_13742);
nand U14095 (N_14095,N_13537,N_13807);
xor U14096 (N_14096,N_13550,N_13453);
nor U14097 (N_14097,N_13534,N_13691);
nor U14098 (N_14098,N_13973,N_13310);
nand U14099 (N_14099,N_13309,N_13541);
nand U14100 (N_14100,N_13328,N_13315);
and U14101 (N_14101,N_13564,N_13495);
or U14102 (N_14102,N_13258,N_13276);
nor U14103 (N_14103,N_13581,N_13906);
and U14104 (N_14104,N_13439,N_13867);
nor U14105 (N_14105,N_13560,N_13254);
and U14106 (N_14106,N_13616,N_13320);
nand U14107 (N_14107,N_13898,N_13352);
or U14108 (N_14108,N_13731,N_13043);
nor U14109 (N_14109,N_13189,N_13996);
and U14110 (N_14110,N_13335,N_13205);
nand U14111 (N_14111,N_13382,N_13947);
nor U14112 (N_14112,N_13270,N_13612);
nand U14113 (N_14113,N_13162,N_13393);
xnor U14114 (N_14114,N_13500,N_13049);
nor U14115 (N_14115,N_13987,N_13394);
xor U14116 (N_14116,N_13789,N_13240);
nand U14117 (N_14117,N_13501,N_13012);
xor U14118 (N_14118,N_13378,N_13751);
nor U14119 (N_14119,N_13067,N_13102);
and U14120 (N_14120,N_13452,N_13907);
or U14121 (N_14121,N_13208,N_13869);
and U14122 (N_14122,N_13180,N_13353);
nand U14123 (N_14123,N_13264,N_13519);
xor U14124 (N_14124,N_13440,N_13462);
or U14125 (N_14125,N_13782,N_13024);
or U14126 (N_14126,N_13355,N_13908);
or U14127 (N_14127,N_13225,N_13956);
and U14128 (N_14128,N_13527,N_13922);
xnor U14129 (N_14129,N_13095,N_13021);
and U14130 (N_14130,N_13743,N_13929);
nand U14131 (N_14131,N_13193,N_13961);
xor U14132 (N_14132,N_13568,N_13364);
nand U14133 (N_14133,N_13882,N_13188);
nand U14134 (N_14134,N_13017,N_13904);
and U14135 (N_14135,N_13970,N_13591);
nand U14136 (N_14136,N_13163,N_13712);
xnor U14137 (N_14137,N_13697,N_13463);
and U14138 (N_14138,N_13228,N_13068);
and U14139 (N_14139,N_13080,N_13562);
xor U14140 (N_14140,N_13432,N_13812);
and U14141 (N_14141,N_13336,N_13979);
xnor U14142 (N_14142,N_13123,N_13707);
nand U14143 (N_14143,N_13985,N_13090);
xnor U14144 (N_14144,N_13826,N_13769);
nor U14145 (N_14145,N_13206,N_13277);
and U14146 (N_14146,N_13147,N_13930);
xnor U14147 (N_14147,N_13157,N_13635);
nand U14148 (N_14148,N_13139,N_13696);
xor U14149 (N_14149,N_13909,N_13078);
nand U14150 (N_14150,N_13905,N_13659);
xor U14151 (N_14151,N_13250,N_13232);
and U14152 (N_14152,N_13121,N_13056);
nor U14153 (N_14153,N_13370,N_13658);
nor U14154 (N_14154,N_13813,N_13686);
or U14155 (N_14155,N_13483,N_13152);
and U14156 (N_14156,N_13146,N_13486);
and U14157 (N_14157,N_13776,N_13698);
nand U14158 (N_14158,N_13998,N_13736);
xor U14159 (N_14159,N_13324,N_13728);
xnor U14160 (N_14160,N_13735,N_13990);
nand U14161 (N_14161,N_13350,N_13786);
or U14162 (N_14162,N_13194,N_13586);
nand U14163 (N_14163,N_13876,N_13410);
nor U14164 (N_14164,N_13437,N_13809);
nand U14165 (N_14165,N_13246,N_13535);
nor U14166 (N_14166,N_13561,N_13983);
nor U14167 (N_14167,N_13414,N_13861);
nor U14168 (N_14168,N_13662,N_13096);
or U14169 (N_14169,N_13244,N_13883);
and U14170 (N_14170,N_13247,N_13260);
or U14171 (N_14171,N_13885,N_13371);
xor U14172 (N_14172,N_13647,N_13316);
nand U14173 (N_14173,N_13020,N_13816);
or U14174 (N_14174,N_13259,N_13575);
xnor U14175 (N_14175,N_13085,N_13331);
xor U14176 (N_14176,N_13843,N_13594);
xnor U14177 (N_14177,N_13902,N_13063);
nand U14178 (N_14178,N_13721,N_13942);
xor U14179 (N_14179,N_13262,N_13007);
xnor U14180 (N_14180,N_13872,N_13860);
nor U14181 (N_14181,N_13281,N_13788);
nor U14182 (N_14182,N_13940,N_13279);
or U14183 (N_14183,N_13187,N_13451);
and U14184 (N_14184,N_13175,N_13421);
nand U14185 (N_14185,N_13957,N_13156);
and U14186 (N_14186,N_13967,N_13685);
or U14187 (N_14187,N_13120,N_13724);
xor U14188 (N_14188,N_13155,N_13076);
and U14189 (N_14189,N_13916,N_13142);
nand U14190 (N_14190,N_13039,N_13614);
and U14191 (N_14191,N_13955,N_13610);
nor U14192 (N_14192,N_13204,N_13426);
nand U14193 (N_14193,N_13543,N_13413);
and U14194 (N_14194,N_13720,N_13975);
or U14195 (N_14195,N_13464,N_13098);
xnor U14196 (N_14196,N_13536,N_13253);
xnor U14197 (N_14197,N_13504,N_13533);
xnor U14198 (N_14198,N_13482,N_13116);
nand U14199 (N_14199,N_13741,N_13673);
or U14200 (N_14200,N_13141,N_13680);
nor U14201 (N_14201,N_13725,N_13411);
nor U14202 (N_14202,N_13395,N_13823);
and U14203 (N_14203,N_13848,N_13333);
or U14204 (N_14204,N_13548,N_13218);
nor U14205 (N_14205,N_13283,N_13932);
or U14206 (N_14206,N_13664,N_13377);
or U14207 (N_14207,N_13780,N_13005);
and U14208 (N_14208,N_13291,N_13864);
nand U14209 (N_14209,N_13570,N_13312);
xor U14210 (N_14210,N_13571,N_13029);
nor U14211 (N_14211,N_13919,N_13081);
or U14212 (N_14212,N_13512,N_13599);
and U14213 (N_14213,N_13787,N_13565);
xnor U14214 (N_14214,N_13196,N_13065);
or U14215 (N_14215,N_13069,N_13845);
xor U14216 (N_14216,N_13734,N_13847);
nor U14217 (N_14217,N_13164,N_13376);
or U14218 (N_14218,N_13455,N_13465);
or U14219 (N_14219,N_13801,N_13911);
nand U14220 (N_14220,N_13709,N_13980);
nand U14221 (N_14221,N_13540,N_13526);
or U14222 (N_14222,N_13573,N_13633);
or U14223 (N_14223,N_13999,N_13358);
nor U14224 (N_14224,N_13766,N_13820);
nand U14225 (N_14225,N_13682,N_13271);
nor U14226 (N_14226,N_13708,N_13631);
nor U14227 (N_14227,N_13417,N_13913);
or U14228 (N_14228,N_13977,N_13110);
or U14229 (N_14229,N_13765,N_13965);
nand U14230 (N_14230,N_13938,N_13479);
xnor U14231 (N_14231,N_13396,N_13549);
nor U14232 (N_14232,N_13398,N_13064);
and U14233 (N_14233,N_13468,N_13859);
and U14234 (N_14234,N_13539,N_13764);
nor U14235 (N_14235,N_13023,N_13994);
nand U14236 (N_14236,N_13829,N_13133);
nor U14237 (N_14237,N_13516,N_13771);
xor U14238 (N_14238,N_13819,N_13237);
xnor U14239 (N_14239,N_13292,N_13037);
xor U14240 (N_14240,N_13470,N_13329);
and U14241 (N_14241,N_13031,N_13617);
or U14242 (N_14242,N_13995,N_13566);
and U14243 (N_14243,N_13492,N_13935);
nor U14244 (N_14244,N_13420,N_13792);
nand U14245 (N_14245,N_13360,N_13959);
nand U14246 (N_14246,N_13732,N_13317);
or U14247 (N_14247,N_13436,N_13891);
xor U14248 (N_14248,N_13740,N_13808);
xnor U14249 (N_14249,N_13428,N_13125);
xor U14250 (N_14250,N_13062,N_13373);
or U14251 (N_14251,N_13634,N_13579);
nand U14252 (N_14252,N_13901,N_13109);
and U14253 (N_14253,N_13627,N_13387);
xor U14254 (N_14254,N_13487,N_13356);
xnor U14255 (N_14255,N_13888,N_13221);
nand U14256 (N_14256,N_13195,N_13783);
nand U14257 (N_14257,N_13611,N_13033);
nand U14258 (N_14258,N_13161,N_13545);
xnor U14259 (N_14259,N_13214,N_13870);
and U14260 (N_14260,N_13171,N_13198);
or U14261 (N_14261,N_13969,N_13167);
nand U14262 (N_14262,N_13173,N_13334);
or U14263 (N_14263,N_13791,N_13321);
or U14264 (N_14264,N_13001,N_13592);
nand U14265 (N_14265,N_13050,N_13055);
xnor U14266 (N_14266,N_13895,N_13722);
nand U14267 (N_14267,N_13752,N_13835);
nor U14268 (N_14268,N_13687,N_13924);
nor U14269 (N_14269,N_13014,N_13060);
or U14270 (N_14270,N_13636,N_13168);
xnor U14271 (N_14271,N_13149,N_13827);
and U14272 (N_14272,N_13991,N_13768);
or U14273 (N_14273,N_13758,N_13119);
and U14274 (N_14274,N_13878,N_13107);
xor U14275 (N_14275,N_13511,N_13525);
and U14276 (N_14276,N_13210,N_13914);
or U14277 (N_14277,N_13059,N_13422);
or U14278 (N_14278,N_13677,N_13494);
and U14279 (N_14279,N_13475,N_13223);
nor U14280 (N_14280,N_13181,N_13311);
nor U14281 (N_14281,N_13596,N_13441);
nand U14282 (N_14282,N_13053,N_13100);
nor U14283 (N_14283,N_13344,N_13389);
or U14284 (N_14284,N_13434,N_13183);
xnor U14285 (N_14285,N_13297,N_13866);
nor U14286 (N_14286,N_13762,N_13089);
and U14287 (N_14287,N_13245,N_13490);
nand U14288 (N_14288,N_13684,N_13288);
or U14289 (N_14289,N_13143,N_13151);
or U14290 (N_14290,N_13045,N_13314);
xor U14291 (N_14291,N_13132,N_13282);
nand U14292 (N_14292,N_13115,N_13520);
or U14293 (N_14293,N_13122,N_13354);
nor U14294 (N_14294,N_13481,N_13302);
nor U14295 (N_14295,N_13503,N_13154);
nor U14296 (N_14296,N_13351,N_13412);
or U14297 (N_14297,N_13392,N_13854);
nor U14298 (N_14298,N_13038,N_13688);
nor U14299 (N_14299,N_13800,N_13461);
or U14300 (N_14300,N_13894,N_13900);
and U14301 (N_14301,N_13703,N_13756);
nor U14302 (N_14302,N_13042,N_13233);
or U14303 (N_14303,N_13480,N_13445);
xor U14304 (N_14304,N_13749,N_13694);
nor U14305 (N_14305,N_13273,N_13515);
and U14306 (N_14306,N_13833,N_13200);
nor U14307 (N_14307,N_13099,N_13252);
and U14308 (N_14308,N_13844,N_13590);
or U14309 (N_14309,N_13323,N_13019);
and U14310 (N_14310,N_13711,N_13873);
nand U14311 (N_14311,N_13622,N_13216);
nand U14312 (N_14312,N_13632,N_13915);
or U14313 (N_14313,N_13931,N_13340);
xnor U14314 (N_14314,N_13958,N_13362);
nor U14315 (N_14315,N_13815,N_13191);
and U14316 (N_14316,N_13397,N_13111);
xor U14317 (N_14317,N_13524,N_13179);
nand U14318 (N_14318,N_13427,N_13760);
or U14319 (N_14319,N_13793,N_13256);
and U14320 (N_14320,N_13542,N_13087);
or U14321 (N_14321,N_13086,N_13619);
nand U14322 (N_14322,N_13484,N_13071);
or U14323 (N_14323,N_13795,N_13984);
or U14324 (N_14324,N_13073,N_13308);
and U14325 (N_14325,N_13215,N_13159);
or U14326 (N_14326,N_13642,N_13249);
and U14327 (N_14327,N_13653,N_13313);
and U14328 (N_14328,N_13003,N_13390);
or U14329 (N_14329,N_13846,N_13300);
xor U14330 (N_14330,N_13294,N_13567);
nor U14331 (N_14331,N_13266,N_13613);
nor U14332 (N_14332,N_13498,N_13135);
or U14333 (N_14333,N_13286,N_13804);
or U14334 (N_14334,N_13699,N_13375);
xnor U14335 (N_14335,N_13903,N_13407);
nor U14336 (N_14336,N_13009,N_13856);
nand U14337 (N_14337,N_13778,N_13476);
nand U14338 (N_14338,N_13972,N_13775);
and U14339 (N_14339,N_13148,N_13327);
and U14340 (N_14340,N_13257,N_13028);
and U14341 (N_14341,N_13946,N_13094);
nand U14342 (N_14342,N_13941,N_13459);
and U14343 (N_14343,N_13423,N_13131);
or U14344 (N_14344,N_13637,N_13048);
nor U14345 (N_14345,N_13450,N_13272);
nand U14346 (N_14346,N_13517,N_13010);
or U14347 (N_14347,N_13380,N_13219);
nand U14348 (N_14348,N_13084,N_13409);
nand U14349 (N_14349,N_13890,N_13608);
nor U14350 (N_14350,N_13137,N_13220);
xor U14351 (N_14351,N_13665,N_13278);
xor U14352 (N_14352,N_13670,N_13656);
and U14353 (N_14353,N_13603,N_13723);
nor U14354 (N_14354,N_13097,N_13251);
or U14355 (N_14355,N_13667,N_13374);
xnor U14356 (N_14356,N_13176,N_13051);
xnor U14357 (N_14357,N_13472,N_13887);
nor U14358 (N_14358,N_13834,N_13473);
and U14359 (N_14359,N_13514,N_13367);
nand U14360 (N_14360,N_13971,N_13079);
or U14361 (N_14361,N_13884,N_13595);
and U14362 (N_14362,N_13150,N_13530);
xnor U14363 (N_14363,N_13339,N_13761);
nor U14364 (N_14364,N_13391,N_13689);
or U14365 (N_14365,N_13726,N_13438);
nor U14366 (N_14366,N_13402,N_13874);
or U14367 (N_14367,N_13082,N_13285);
xor U14368 (N_14368,N_13296,N_13660);
and U14369 (N_14369,N_13136,N_13138);
nor U14370 (N_14370,N_13641,N_13199);
or U14371 (N_14371,N_13405,N_13092);
xor U14372 (N_14372,N_13342,N_13126);
xnor U14373 (N_14373,N_13865,N_13505);
nor U14374 (N_14374,N_13112,N_13802);
nand U14375 (N_14375,N_13114,N_13117);
nor U14376 (N_14376,N_13644,N_13893);
nand U14377 (N_14377,N_13657,N_13325);
nand U14378 (N_14378,N_13551,N_13818);
xnor U14379 (N_14379,N_13605,N_13025);
nor U14380 (N_14380,N_13951,N_13066);
xnor U14381 (N_14381,N_13943,N_13625);
and U14382 (N_14382,N_13628,N_13241);
or U14383 (N_14383,N_13753,N_13431);
xor U14384 (N_14384,N_13185,N_13529);
xor U14385 (N_14385,N_13757,N_13477);
xor U14386 (N_14386,N_13654,N_13920);
and U14387 (N_14387,N_13008,N_13496);
or U14388 (N_14388,N_13474,N_13928);
nand U14389 (N_14389,N_13824,N_13361);
nand U14390 (N_14390,N_13997,N_13794);
nand U14391 (N_14391,N_13679,N_13343);
nor U14392 (N_14392,N_13671,N_13655);
or U14393 (N_14393,N_13379,N_13621);
nand U14394 (N_14394,N_13458,N_13912);
xnor U14395 (N_14395,N_13744,N_13466);
nand U14396 (N_14396,N_13950,N_13737);
nand U14397 (N_14397,N_13580,N_13730);
nor U14398 (N_14398,N_13702,N_13444);
nand U14399 (N_14399,N_13601,N_13372);
and U14400 (N_14400,N_13837,N_13202);
nand U14401 (N_14401,N_13849,N_13810);
xnor U14402 (N_14402,N_13108,N_13018);
nand U14403 (N_14403,N_13544,N_13892);
xor U14404 (N_14404,N_13926,N_13937);
nor U14405 (N_14405,N_13330,N_13727);
or U14406 (N_14406,N_13471,N_13212);
or U14407 (N_14407,N_13443,N_13585);
nor U14408 (N_14408,N_13469,N_13899);
nor U14409 (N_14409,N_13209,N_13203);
or U14410 (N_14410,N_13638,N_13661);
xnor U14411 (N_14411,N_13124,N_13798);
xor U14412 (N_14412,N_13169,N_13044);
nand U14413 (N_14413,N_13083,N_13416);
and U14414 (N_14414,N_13649,N_13243);
or U14415 (N_14415,N_13933,N_13862);
nor U14416 (N_14416,N_13369,N_13805);
nand U14417 (N_14417,N_13104,N_13668);
xor U14418 (N_14418,N_13629,N_13026);
nand U14419 (N_14419,N_13072,N_13338);
nand U14420 (N_14420,N_13563,N_13700);
and U14421 (N_14421,N_13552,N_13489);
nand U14422 (N_14422,N_13293,N_13921);
xor U14423 (N_14423,N_13639,N_13306);
and U14424 (N_14424,N_13593,N_13401);
and U14425 (N_14425,N_13842,N_13546);
or U14426 (N_14426,N_13318,N_13701);
and U14427 (N_14427,N_13863,N_13615);
nor U14428 (N_14428,N_13337,N_13508);
and U14429 (N_14429,N_13838,N_13280);
or U14430 (N_14430,N_13851,N_13274);
or U14431 (N_14431,N_13814,N_13871);
or U14432 (N_14432,N_13348,N_13944);
nor U14433 (N_14433,N_13738,N_13513);
xor U14434 (N_14434,N_13645,N_13523);
xor U14435 (N_14435,N_13981,N_13172);
or U14436 (N_14436,N_13910,N_13046);
and U14437 (N_14437,N_13041,N_13578);
xnor U14438 (N_14438,N_13704,N_13030);
nor U14439 (N_14439,N_13035,N_13841);
and U14440 (N_14440,N_13158,N_13705);
and U14441 (N_14441,N_13365,N_13485);
and U14442 (N_14442,N_13201,N_13976);
nor U14443 (N_14443,N_13879,N_13457);
or U14444 (N_14444,N_13134,N_13587);
xor U14445 (N_14445,N_13224,N_13077);
nor U14446 (N_14446,N_13027,N_13992);
nor U14447 (N_14447,N_13982,N_13454);
nor U14448 (N_14448,N_13047,N_13488);
xnor U14449 (N_14449,N_13186,N_13275);
xnor U14450 (N_14450,N_13710,N_13433);
xor U14451 (N_14451,N_13419,N_13088);
and U14452 (N_14452,N_13674,N_13298);
xor U14453 (N_14453,N_13868,N_13806);
nand U14454 (N_14454,N_13583,N_13381);
nand U14455 (N_14455,N_13729,N_13238);
xor U14456 (N_14456,N_13850,N_13630);
nand U14457 (N_14457,N_13538,N_13602);
xor U14458 (N_14458,N_13683,N_13557);
and U14459 (N_14459,N_13960,N_13714);
nand U14460 (N_14460,N_13974,N_13166);
and U14461 (N_14461,N_13442,N_13384);
nand U14462 (N_14462,N_13853,N_13456);
nor U14463 (N_14463,N_13385,N_13927);
and U14464 (N_14464,N_13207,N_13448);
nor U14465 (N_14465,N_13267,N_13713);
or U14466 (N_14466,N_13263,N_13388);
and U14467 (N_14467,N_13962,N_13499);
and U14468 (N_14468,N_13858,N_13797);
xor U14469 (N_14469,N_13447,N_13953);
nand U14470 (N_14470,N_13840,N_13290);
nor U14471 (N_14471,N_13897,N_13424);
and U14472 (N_14472,N_13322,N_13093);
or U14473 (N_14473,N_13767,N_13748);
and U14474 (N_14474,N_13881,N_13400);
nor U14475 (N_14475,N_13502,N_13770);
xor U14476 (N_14476,N_13105,N_13666);
or U14477 (N_14477,N_13772,N_13716);
nor U14478 (N_14478,N_13182,N_13643);
nor U14479 (N_14479,N_13936,N_13403);
xor U14480 (N_14480,N_13015,N_13165);
nor U14481 (N_14481,N_13192,N_13754);
xnor U14482 (N_14482,N_13129,N_13755);
xnor U14483 (N_14483,N_13572,N_13507);
or U14484 (N_14484,N_13781,N_13217);
xnor U14485 (N_14485,N_13747,N_13430);
xnor U14486 (N_14486,N_13574,N_13510);
nor U14487 (N_14487,N_13773,N_13261);
xor U14488 (N_14488,N_13211,N_13626);
xnor U14489 (N_14489,N_13745,N_13305);
nor U14490 (N_14490,N_13886,N_13839);
or U14491 (N_14491,N_13989,N_13184);
nand U14492 (N_14492,N_13923,N_13582);
or U14493 (N_14493,N_13648,N_13779);
and U14494 (N_14494,N_13287,N_13435);
and U14495 (N_14495,N_13939,N_13831);
nor U14496 (N_14496,N_13799,N_13013);
nand U14497 (N_14497,N_13128,N_13467);
nand U14498 (N_14498,N_13576,N_13678);
nand U14499 (N_14499,N_13785,N_13718);
or U14500 (N_14500,N_13862,N_13516);
or U14501 (N_14501,N_13687,N_13987);
and U14502 (N_14502,N_13163,N_13107);
nand U14503 (N_14503,N_13662,N_13482);
nor U14504 (N_14504,N_13535,N_13711);
and U14505 (N_14505,N_13736,N_13234);
and U14506 (N_14506,N_13901,N_13344);
nor U14507 (N_14507,N_13547,N_13688);
xor U14508 (N_14508,N_13715,N_13711);
xnor U14509 (N_14509,N_13780,N_13711);
nor U14510 (N_14510,N_13966,N_13786);
and U14511 (N_14511,N_13464,N_13591);
or U14512 (N_14512,N_13268,N_13330);
nor U14513 (N_14513,N_13472,N_13627);
nor U14514 (N_14514,N_13113,N_13971);
nand U14515 (N_14515,N_13639,N_13608);
xor U14516 (N_14516,N_13347,N_13676);
xor U14517 (N_14517,N_13686,N_13843);
or U14518 (N_14518,N_13696,N_13834);
or U14519 (N_14519,N_13520,N_13522);
and U14520 (N_14520,N_13552,N_13099);
nand U14521 (N_14521,N_13584,N_13063);
xor U14522 (N_14522,N_13514,N_13328);
nand U14523 (N_14523,N_13400,N_13529);
or U14524 (N_14524,N_13329,N_13709);
xnor U14525 (N_14525,N_13929,N_13554);
xor U14526 (N_14526,N_13617,N_13226);
nand U14527 (N_14527,N_13325,N_13233);
xor U14528 (N_14528,N_13375,N_13407);
or U14529 (N_14529,N_13668,N_13328);
xnor U14530 (N_14530,N_13056,N_13597);
nand U14531 (N_14531,N_13930,N_13451);
and U14532 (N_14532,N_13757,N_13720);
and U14533 (N_14533,N_13229,N_13218);
or U14534 (N_14534,N_13472,N_13393);
and U14535 (N_14535,N_13870,N_13566);
nor U14536 (N_14536,N_13275,N_13988);
and U14537 (N_14537,N_13782,N_13701);
xnor U14538 (N_14538,N_13023,N_13880);
nand U14539 (N_14539,N_13717,N_13895);
nand U14540 (N_14540,N_13050,N_13127);
xnor U14541 (N_14541,N_13969,N_13503);
xnor U14542 (N_14542,N_13659,N_13980);
xnor U14543 (N_14543,N_13035,N_13847);
nor U14544 (N_14544,N_13599,N_13552);
nand U14545 (N_14545,N_13687,N_13598);
xor U14546 (N_14546,N_13013,N_13951);
xnor U14547 (N_14547,N_13966,N_13171);
or U14548 (N_14548,N_13570,N_13229);
or U14549 (N_14549,N_13925,N_13557);
and U14550 (N_14550,N_13128,N_13556);
xnor U14551 (N_14551,N_13362,N_13306);
nor U14552 (N_14552,N_13445,N_13502);
nor U14553 (N_14553,N_13888,N_13255);
nor U14554 (N_14554,N_13645,N_13570);
nor U14555 (N_14555,N_13984,N_13898);
or U14556 (N_14556,N_13229,N_13935);
or U14557 (N_14557,N_13411,N_13655);
and U14558 (N_14558,N_13659,N_13700);
nor U14559 (N_14559,N_13694,N_13456);
and U14560 (N_14560,N_13618,N_13364);
nand U14561 (N_14561,N_13790,N_13566);
nand U14562 (N_14562,N_13434,N_13229);
or U14563 (N_14563,N_13975,N_13404);
or U14564 (N_14564,N_13923,N_13000);
nand U14565 (N_14565,N_13783,N_13922);
nor U14566 (N_14566,N_13372,N_13414);
and U14567 (N_14567,N_13968,N_13805);
nand U14568 (N_14568,N_13889,N_13296);
and U14569 (N_14569,N_13890,N_13636);
xnor U14570 (N_14570,N_13421,N_13000);
nor U14571 (N_14571,N_13553,N_13722);
xor U14572 (N_14572,N_13675,N_13676);
or U14573 (N_14573,N_13968,N_13906);
nand U14574 (N_14574,N_13195,N_13211);
or U14575 (N_14575,N_13858,N_13216);
or U14576 (N_14576,N_13085,N_13409);
nand U14577 (N_14577,N_13537,N_13026);
nand U14578 (N_14578,N_13613,N_13467);
or U14579 (N_14579,N_13541,N_13189);
and U14580 (N_14580,N_13328,N_13701);
xnor U14581 (N_14581,N_13631,N_13220);
and U14582 (N_14582,N_13734,N_13567);
nand U14583 (N_14583,N_13875,N_13099);
or U14584 (N_14584,N_13830,N_13417);
or U14585 (N_14585,N_13433,N_13978);
or U14586 (N_14586,N_13015,N_13447);
and U14587 (N_14587,N_13544,N_13198);
nand U14588 (N_14588,N_13852,N_13211);
and U14589 (N_14589,N_13000,N_13753);
and U14590 (N_14590,N_13994,N_13368);
nor U14591 (N_14591,N_13904,N_13808);
or U14592 (N_14592,N_13559,N_13686);
xnor U14593 (N_14593,N_13883,N_13498);
nor U14594 (N_14594,N_13251,N_13297);
nand U14595 (N_14595,N_13009,N_13473);
xnor U14596 (N_14596,N_13145,N_13222);
and U14597 (N_14597,N_13115,N_13601);
nor U14598 (N_14598,N_13701,N_13432);
xnor U14599 (N_14599,N_13650,N_13864);
nor U14600 (N_14600,N_13888,N_13671);
xnor U14601 (N_14601,N_13938,N_13634);
nor U14602 (N_14602,N_13591,N_13290);
or U14603 (N_14603,N_13964,N_13588);
and U14604 (N_14604,N_13890,N_13353);
and U14605 (N_14605,N_13006,N_13382);
xor U14606 (N_14606,N_13711,N_13549);
nor U14607 (N_14607,N_13714,N_13116);
or U14608 (N_14608,N_13901,N_13208);
or U14609 (N_14609,N_13393,N_13831);
nor U14610 (N_14610,N_13626,N_13280);
nand U14611 (N_14611,N_13464,N_13070);
nor U14612 (N_14612,N_13221,N_13163);
or U14613 (N_14613,N_13707,N_13722);
xnor U14614 (N_14614,N_13979,N_13736);
nand U14615 (N_14615,N_13473,N_13780);
xor U14616 (N_14616,N_13644,N_13863);
xor U14617 (N_14617,N_13058,N_13636);
xnor U14618 (N_14618,N_13808,N_13507);
and U14619 (N_14619,N_13883,N_13001);
or U14620 (N_14620,N_13601,N_13008);
xnor U14621 (N_14621,N_13168,N_13639);
xor U14622 (N_14622,N_13592,N_13832);
nand U14623 (N_14623,N_13230,N_13663);
nand U14624 (N_14624,N_13440,N_13898);
xnor U14625 (N_14625,N_13449,N_13138);
xnor U14626 (N_14626,N_13209,N_13796);
or U14627 (N_14627,N_13482,N_13065);
and U14628 (N_14628,N_13599,N_13158);
and U14629 (N_14629,N_13737,N_13768);
xor U14630 (N_14630,N_13412,N_13662);
nand U14631 (N_14631,N_13059,N_13471);
nand U14632 (N_14632,N_13686,N_13215);
xnor U14633 (N_14633,N_13824,N_13171);
or U14634 (N_14634,N_13802,N_13261);
xor U14635 (N_14635,N_13871,N_13418);
or U14636 (N_14636,N_13473,N_13921);
xor U14637 (N_14637,N_13201,N_13623);
nor U14638 (N_14638,N_13691,N_13268);
xnor U14639 (N_14639,N_13276,N_13189);
and U14640 (N_14640,N_13265,N_13023);
xnor U14641 (N_14641,N_13164,N_13765);
nor U14642 (N_14642,N_13324,N_13261);
nand U14643 (N_14643,N_13085,N_13857);
or U14644 (N_14644,N_13192,N_13577);
or U14645 (N_14645,N_13708,N_13393);
nor U14646 (N_14646,N_13820,N_13242);
nand U14647 (N_14647,N_13610,N_13276);
and U14648 (N_14648,N_13962,N_13833);
or U14649 (N_14649,N_13094,N_13175);
nor U14650 (N_14650,N_13292,N_13644);
and U14651 (N_14651,N_13072,N_13269);
nor U14652 (N_14652,N_13029,N_13475);
xnor U14653 (N_14653,N_13926,N_13337);
nor U14654 (N_14654,N_13772,N_13944);
and U14655 (N_14655,N_13388,N_13805);
or U14656 (N_14656,N_13413,N_13130);
and U14657 (N_14657,N_13731,N_13615);
or U14658 (N_14658,N_13924,N_13447);
xnor U14659 (N_14659,N_13424,N_13733);
nand U14660 (N_14660,N_13757,N_13891);
nor U14661 (N_14661,N_13195,N_13753);
and U14662 (N_14662,N_13796,N_13120);
nor U14663 (N_14663,N_13846,N_13236);
nor U14664 (N_14664,N_13375,N_13400);
nor U14665 (N_14665,N_13113,N_13640);
or U14666 (N_14666,N_13937,N_13975);
xor U14667 (N_14667,N_13911,N_13661);
nor U14668 (N_14668,N_13069,N_13591);
nor U14669 (N_14669,N_13727,N_13139);
xnor U14670 (N_14670,N_13515,N_13424);
and U14671 (N_14671,N_13869,N_13028);
or U14672 (N_14672,N_13640,N_13955);
xor U14673 (N_14673,N_13149,N_13905);
xor U14674 (N_14674,N_13978,N_13243);
xor U14675 (N_14675,N_13525,N_13518);
nor U14676 (N_14676,N_13917,N_13830);
nand U14677 (N_14677,N_13604,N_13403);
or U14678 (N_14678,N_13824,N_13509);
xnor U14679 (N_14679,N_13081,N_13452);
nor U14680 (N_14680,N_13565,N_13824);
xnor U14681 (N_14681,N_13570,N_13592);
nand U14682 (N_14682,N_13714,N_13393);
xnor U14683 (N_14683,N_13353,N_13136);
and U14684 (N_14684,N_13795,N_13161);
xor U14685 (N_14685,N_13697,N_13518);
or U14686 (N_14686,N_13361,N_13771);
or U14687 (N_14687,N_13385,N_13834);
xor U14688 (N_14688,N_13009,N_13569);
nor U14689 (N_14689,N_13287,N_13068);
and U14690 (N_14690,N_13713,N_13287);
xor U14691 (N_14691,N_13491,N_13595);
or U14692 (N_14692,N_13645,N_13364);
or U14693 (N_14693,N_13056,N_13304);
and U14694 (N_14694,N_13003,N_13601);
and U14695 (N_14695,N_13781,N_13664);
nand U14696 (N_14696,N_13295,N_13421);
xnor U14697 (N_14697,N_13662,N_13880);
nand U14698 (N_14698,N_13664,N_13366);
or U14699 (N_14699,N_13952,N_13693);
or U14700 (N_14700,N_13814,N_13791);
and U14701 (N_14701,N_13294,N_13461);
and U14702 (N_14702,N_13841,N_13695);
and U14703 (N_14703,N_13529,N_13726);
and U14704 (N_14704,N_13327,N_13718);
xor U14705 (N_14705,N_13100,N_13223);
nand U14706 (N_14706,N_13414,N_13032);
xnor U14707 (N_14707,N_13737,N_13498);
nand U14708 (N_14708,N_13101,N_13805);
nor U14709 (N_14709,N_13646,N_13712);
xnor U14710 (N_14710,N_13713,N_13528);
nor U14711 (N_14711,N_13710,N_13521);
nand U14712 (N_14712,N_13991,N_13470);
or U14713 (N_14713,N_13416,N_13313);
nand U14714 (N_14714,N_13387,N_13895);
or U14715 (N_14715,N_13545,N_13132);
and U14716 (N_14716,N_13306,N_13399);
xor U14717 (N_14717,N_13189,N_13847);
nand U14718 (N_14718,N_13513,N_13015);
xor U14719 (N_14719,N_13606,N_13052);
or U14720 (N_14720,N_13101,N_13738);
nor U14721 (N_14721,N_13463,N_13760);
xnor U14722 (N_14722,N_13335,N_13820);
nand U14723 (N_14723,N_13248,N_13460);
nand U14724 (N_14724,N_13897,N_13958);
and U14725 (N_14725,N_13780,N_13422);
and U14726 (N_14726,N_13945,N_13199);
nand U14727 (N_14727,N_13779,N_13301);
and U14728 (N_14728,N_13824,N_13906);
xnor U14729 (N_14729,N_13868,N_13652);
and U14730 (N_14730,N_13460,N_13276);
xnor U14731 (N_14731,N_13830,N_13664);
nor U14732 (N_14732,N_13844,N_13936);
xor U14733 (N_14733,N_13066,N_13801);
or U14734 (N_14734,N_13016,N_13040);
nor U14735 (N_14735,N_13755,N_13122);
and U14736 (N_14736,N_13967,N_13189);
or U14737 (N_14737,N_13931,N_13345);
and U14738 (N_14738,N_13884,N_13526);
nor U14739 (N_14739,N_13754,N_13677);
nand U14740 (N_14740,N_13554,N_13857);
nor U14741 (N_14741,N_13968,N_13117);
nand U14742 (N_14742,N_13076,N_13941);
nor U14743 (N_14743,N_13779,N_13323);
or U14744 (N_14744,N_13737,N_13605);
nor U14745 (N_14745,N_13189,N_13198);
xnor U14746 (N_14746,N_13379,N_13993);
or U14747 (N_14747,N_13816,N_13149);
nand U14748 (N_14748,N_13226,N_13947);
nand U14749 (N_14749,N_13084,N_13880);
xor U14750 (N_14750,N_13985,N_13822);
or U14751 (N_14751,N_13474,N_13231);
or U14752 (N_14752,N_13632,N_13354);
or U14753 (N_14753,N_13486,N_13326);
nand U14754 (N_14754,N_13480,N_13774);
and U14755 (N_14755,N_13870,N_13415);
nand U14756 (N_14756,N_13306,N_13118);
nor U14757 (N_14757,N_13002,N_13924);
or U14758 (N_14758,N_13583,N_13406);
or U14759 (N_14759,N_13208,N_13771);
nor U14760 (N_14760,N_13646,N_13287);
and U14761 (N_14761,N_13057,N_13966);
xor U14762 (N_14762,N_13603,N_13995);
nand U14763 (N_14763,N_13433,N_13923);
nor U14764 (N_14764,N_13201,N_13212);
nor U14765 (N_14765,N_13078,N_13239);
nand U14766 (N_14766,N_13679,N_13673);
nand U14767 (N_14767,N_13364,N_13373);
nand U14768 (N_14768,N_13146,N_13713);
and U14769 (N_14769,N_13386,N_13519);
xor U14770 (N_14770,N_13875,N_13832);
nor U14771 (N_14771,N_13761,N_13193);
xnor U14772 (N_14772,N_13969,N_13055);
nor U14773 (N_14773,N_13238,N_13561);
nor U14774 (N_14774,N_13529,N_13431);
and U14775 (N_14775,N_13302,N_13142);
xor U14776 (N_14776,N_13119,N_13848);
nor U14777 (N_14777,N_13923,N_13244);
or U14778 (N_14778,N_13422,N_13875);
xor U14779 (N_14779,N_13131,N_13114);
xnor U14780 (N_14780,N_13228,N_13794);
or U14781 (N_14781,N_13182,N_13611);
or U14782 (N_14782,N_13652,N_13221);
or U14783 (N_14783,N_13668,N_13640);
nand U14784 (N_14784,N_13469,N_13381);
or U14785 (N_14785,N_13643,N_13401);
nand U14786 (N_14786,N_13433,N_13319);
nand U14787 (N_14787,N_13593,N_13915);
nand U14788 (N_14788,N_13927,N_13265);
or U14789 (N_14789,N_13066,N_13275);
or U14790 (N_14790,N_13293,N_13044);
or U14791 (N_14791,N_13745,N_13242);
or U14792 (N_14792,N_13759,N_13866);
nor U14793 (N_14793,N_13556,N_13969);
or U14794 (N_14794,N_13428,N_13599);
or U14795 (N_14795,N_13406,N_13399);
or U14796 (N_14796,N_13885,N_13121);
xnor U14797 (N_14797,N_13318,N_13434);
nor U14798 (N_14798,N_13286,N_13215);
and U14799 (N_14799,N_13745,N_13985);
xor U14800 (N_14800,N_13285,N_13234);
nand U14801 (N_14801,N_13139,N_13562);
nor U14802 (N_14802,N_13433,N_13911);
nand U14803 (N_14803,N_13698,N_13228);
xor U14804 (N_14804,N_13505,N_13939);
nor U14805 (N_14805,N_13232,N_13028);
nor U14806 (N_14806,N_13641,N_13351);
xnor U14807 (N_14807,N_13130,N_13369);
xnor U14808 (N_14808,N_13995,N_13845);
nor U14809 (N_14809,N_13447,N_13468);
nand U14810 (N_14810,N_13709,N_13185);
or U14811 (N_14811,N_13298,N_13642);
nand U14812 (N_14812,N_13076,N_13433);
nand U14813 (N_14813,N_13948,N_13427);
or U14814 (N_14814,N_13717,N_13787);
and U14815 (N_14815,N_13234,N_13777);
xor U14816 (N_14816,N_13235,N_13336);
xnor U14817 (N_14817,N_13447,N_13421);
xnor U14818 (N_14818,N_13600,N_13040);
nor U14819 (N_14819,N_13083,N_13691);
nor U14820 (N_14820,N_13024,N_13658);
and U14821 (N_14821,N_13059,N_13208);
xnor U14822 (N_14822,N_13312,N_13455);
nand U14823 (N_14823,N_13949,N_13181);
xor U14824 (N_14824,N_13698,N_13063);
xor U14825 (N_14825,N_13520,N_13538);
nor U14826 (N_14826,N_13266,N_13338);
and U14827 (N_14827,N_13100,N_13421);
nand U14828 (N_14828,N_13067,N_13969);
or U14829 (N_14829,N_13255,N_13868);
or U14830 (N_14830,N_13010,N_13736);
nor U14831 (N_14831,N_13245,N_13069);
and U14832 (N_14832,N_13151,N_13565);
and U14833 (N_14833,N_13072,N_13775);
and U14834 (N_14834,N_13854,N_13547);
xor U14835 (N_14835,N_13524,N_13956);
xor U14836 (N_14836,N_13389,N_13219);
nand U14837 (N_14837,N_13938,N_13675);
nor U14838 (N_14838,N_13321,N_13398);
or U14839 (N_14839,N_13083,N_13758);
nor U14840 (N_14840,N_13773,N_13502);
nand U14841 (N_14841,N_13296,N_13781);
xor U14842 (N_14842,N_13472,N_13710);
nor U14843 (N_14843,N_13527,N_13214);
xor U14844 (N_14844,N_13308,N_13568);
xnor U14845 (N_14845,N_13229,N_13781);
and U14846 (N_14846,N_13805,N_13957);
or U14847 (N_14847,N_13238,N_13405);
or U14848 (N_14848,N_13076,N_13915);
xor U14849 (N_14849,N_13444,N_13097);
or U14850 (N_14850,N_13729,N_13049);
nand U14851 (N_14851,N_13976,N_13874);
and U14852 (N_14852,N_13447,N_13920);
or U14853 (N_14853,N_13031,N_13538);
or U14854 (N_14854,N_13701,N_13989);
nor U14855 (N_14855,N_13705,N_13323);
xnor U14856 (N_14856,N_13224,N_13155);
nand U14857 (N_14857,N_13032,N_13949);
nor U14858 (N_14858,N_13353,N_13748);
nor U14859 (N_14859,N_13247,N_13370);
nor U14860 (N_14860,N_13243,N_13407);
nand U14861 (N_14861,N_13844,N_13791);
or U14862 (N_14862,N_13387,N_13868);
nor U14863 (N_14863,N_13111,N_13811);
xor U14864 (N_14864,N_13164,N_13797);
xor U14865 (N_14865,N_13846,N_13200);
nand U14866 (N_14866,N_13949,N_13438);
and U14867 (N_14867,N_13077,N_13113);
or U14868 (N_14868,N_13956,N_13970);
xor U14869 (N_14869,N_13159,N_13110);
nor U14870 (N_14870,N_13318,N_13114);
or U14871 (N_14871,N_13056,N_13175);
nand U14872 (N_14872,N_13546,N_13320);
xnor U14873 (N_14873,N_13094,N_13654);
and U14874 (N_14874,N_13404,N_13387);
and U14875 (N_14875,N_13461,N_13791);
nand U14876 (N_14876,N_13266,N_13412);
and U14877 (N_14877,N_13280,N_13353);
and U14878 (N_14878,N_13754,N_13770);
xor U14879 (N_14879,N_13811,N_13268);
or U14880 (N_14880,N_13336,N_13973);
xnor U14881 (N_14881,N_13088,N_13322);
nand U14882 (N_14882,N_13222,N_13446);
nand U14883 (N_14883,N_13479,N_13166);
or U14884 (N_14884,N_13906,N_13372);
nand U14885 (N_14885,N_13997,N_13669);
and U14886 (N_14886,N_13006,N_13466);
and U14887 (N_14887,N_13866,N_13320);
xnor U14888 (N_14888,N_13337,N_13921);
xnor U14889 (N_14889,N_13804,N_13809);
and U14890 (N_14890,N_13874,N_13531);
xor U14891 (N_14891,N_13277,N_13270);
or U14892 (N_14892,N_13332,N_13140);
and U14893 (N_14893,N_13938,N_13955);
xnor U14894 (N_14894,N_13701,N_13735);
nor U14895 (N_14895,N_13095,N_13854);
and U14896 (N_14896,N_13035,N_13029);
xor U14897 (N_14897,N_13966,N_13169);
and U14898 (N_14898,N_13483,N_13039);
and U14899 (N_14899,N_13468,N_13491);
xnor U14900 (N_14900,N_13866,N_13098);
xor U14901 (N_14901,N_13313,N_13097);
nand U14902 (N_14902,N_13928,N_13884);
and U14903 (N_14903,N_13219,N_13246);
nor U14904 (N_14904,N_13107,N_13858);
or U14905 (N_14905,N_13608,N_13580);
or U14906 (N_14906,N_13999,N_13095);
or U14907 (N_14907,N_13929,N_13366);
or U14908 (N_14908,N_13914,N_13998);
and U14909 (N_14909,N_13540,N_13476);
nor U14910 (N_14910,N_13015,N_13449);
xor U14911 (N_14911,N_13556,N_13588);
nor U14912 (N_14912,N_13163,N_13296);
nand U14913 (N_14913,N_13697,N_13390);
xor U14914 (N_14914,N_13184,N_13626);
nand U14915 (N_14915,N_13414,N_13075);
and U14916 (N_14916,N_13006,N_13528);
nand U14917 (N_14917,N_13792,N_13465);
and U14918 (N_14918,N_13713,N_13117);
or U14919 (N_14919,N_13428,N_13116);
or U14920 (N_14920,N_13340,N_13091);
nor U14921 (N_14921,N_13010,N_13215);
or U14922 (N_14922,N_13182,N_13544);
or U14923 (N_14923,N_13091,N_13353);
nand U14924 (N_14924,N_13677,N_13827);
nand U14925 (N_14925,N_13436,N_13614);
nand U14926 (N_14926,N_13487,N_13963);
or U14927 (N_14927,N_13573,N_13346);
nand U14928 (N_14928,N_13790,N_13230);
or U14929 (N_14929,N_13908,N_13668);
and U14930 (N_14930,N_13709,N_13841);
nand U14931 (N_14931,N_13830,N_13180);
nand U14932 (N_14932,N_13739,N_13797);
nand U14933 (N_14933,N_13045,N_13034);
nor U14934 (N_14934,N_13344,N_13494);
xor U14935 (N_14935,N_13006,N_13928);
nand U14936 (N_14936,N_13137,N_13375);
xor U14937 (N_14937,N_13832,N_13302);
nor U14938 (N_14938,N_13928,N_13778);
or U14939 (N_14939,N_13864,N_13951);
nand U14940 (N_14940,N_13446,N_13657);
nor U14941 (N_14941,N_13942,N_13981);
and U14942 (N_14942,N_13870,N_13890);
or U14943 (N_14943,N_13463,N_13185);
and U14944 (N_14944,N_13942,N_13402);
nand U14945 (N_14945,N_13162,N_13262);
nor U14946 (N_14946,N_13146,N_13720);
nor U14947 (N_14947,N_13124,N_13814);
nand U14948 (N_14948,N_13089,N_13204);
nor U14949 (N_14949,N_13249,N_13021);
nand U14950 (N_14950,N_13218,N_13957);
nor U14951 (N_14951,N_13268,N_13113);
nand U14952 (N_14952,N_13389,N_13590);
nor U14953 (N_14953,N_13171,N_13139);
or U14954 (N_14954,N_13606,N_13602);
and U14955 (N_14955,N_13764,N_13104);
and U14956 (N_14956,N_13812,N_13808);
xnor U14957 (N_14957,N_13628,N_13091);
nand U14958 (N_14958,N_13025,N_13313);
or U14959 (N_14959,N_13549,N_13980);
xor U14960 (N_14960,N_13854,N_13387);
nor U14961 (N_14961,N_13024,N_13244);
nand U14962 (N_14962,N_13584,N_13031);
nand U14963 (N_14963,N_13965,N_13096);
and U14964 (N_14964,N_13508,N_13465);
nor U14965 (N_14965,N_13953,N_13270);
nand U14966 (N_14966,N_13658,N_13423);
nand U14967 (N_14967,N_13741,N_13327);
nand U14968 (N_14968,N_13795,N_13688);
nor U14969 (N_14969,N_13709,N_13109);
xnor U14970 (N_14970,N_13440,N_13745);
and U14971 (N_14971,N_13368,N_13276);
nor U14972 (N_14972,N_13237,N_13401);
nand U14973 (N_14973,N_13132,N_13239);
and U14974 (N_14974,N_13231,N_13391);
xor U14975 (N_14975,N_13891,N_13819);
xor U14976 (N_14976,N_13779,N_13900);
or U14977 (N_14977,N_13893,N_13734);
nor U14978 (N_14978,N_13604,N_13234);
xor U14979 (N_14979,N_13318,N_13969);
nor U14980 (N_14980,N_13255,N_13477);
or U14981 (N_14981,N_13055,N_13407);
or U14982 (N_14982,N_13357,N_13061);
nor U14983 (N_14983,N_13298,N_13100);
nand U14984 (N_14984,N_13292,N_13512);
and U14985 (N_14985,N_13581,N_13469);
nor U14986 (N_14986,N_13923,N_13838);
nor U14987 (N_14987,N_13028,N_13551);
and U14988 (N_14988,N_13730,N_13870);
nor U14989 (N_14989,N_13296,N_13585);
xnor U14990 (N_14990,N_13828,N_13205);
nor U14991 (N_14991,N_13706,N_13120);
or U14992 (N_14992,N_13846,N_13258);
or U14993 (N_14993,N_13744,N_13452);
nand U14994 (N_14994,N_13017,N_13928);
nand U14995 (N_14995,N_13170,N_13096);
nor U14996 (N_14996,N_13893,N_13326);
or U14997 (N_14997,N_13523,N_13952);
nor U14998 (N_14998,N_13988,N_13739);
or U14999 (N_14999,N_13887,N_13836);
nand UO_0 (O_0,N_14595,N_14498);
or UO_1 (O_1,N_14793,N_14963);
nor UO_2 (O_2,N_14489,N_14400);
xor UO_3 (O_3,N_14887,N_14845);
xnor UO_4 (O_4,N_14404,N_14384);
nor UO_5 (O_5,N_14602,N_14657);
nand UO_6 (O_6,N_14648,N_14539);
nand UO_7 (O_7,N_14905,N_14477);
and UO_8 (O_8,N_14521,N_14062);
and UO_9 (O_9,N_14307,N_14399);
nor UO_10 (O_10,N_14204,N_14779);
nor UO_11 (O_11,N_14169,N_14168);
nand UO_12 (O_12,N_14997,N_14805);
nor UO_13 (O_13,N_14527,N_14067);
or UO_14 (O_14,N_14170,N_14330);
nor UO_15 (O_15,N_14876,N_14323);
or UO_16 (O_16,N_14809,N_14255);
and UO_17 (O_17,N_14747,N_14233);
nand UO_18 (O_18,N_14059,N_14299);
nor UO_19 (O_19,N_14916,N_14829);
xnor UO_20 (O_20,N_14538,N_14254);
xor UO_21 (O_21,N_14003,N_14136);
nand UO_22 (O_22,N_14275,N_14720);
xor UO_23 (O_23,N_14245,N_14519);
or UO_24 (O_24,N_14155,N_14135);
nor UO_25 (O_25,N_14686,N_14695);
or UO_26 (O_26,N_14199,N_14162);
xor UO_27 (O_27,N_14556,N_14069);
nor UO_28 (O_28,N_14201,N_14085);
nor UO_29 (O_29,N_14397,N_14572);
xor UO_30 (O_30,N_14732,N_14965);
xnor UO_31 (O_31,N_14510,N_14919);
nor UO_32 (O_32,N_14278,N_14023);
nand UO_33 (O_33,N_14601,N_14774);
xnor UO_34 (O_34,N_14978,N_14923);
and UO_35 (O_35,N_14093,N_14993);
and UO_36 (O_36,N_14957,N_14277);
nand UO_37 (O_37,N_14269,N_14493);
nand UO_38 (O_38,N_14403,N_14821);
and UO_39 (O_39,N_14529,N_14703);
nand UO_40 (O_40,N_14195,N_14799);
and UO_41 (O_41,N_14267,N_14303);
nor UO_42 (O_42,N_14710,N_14457);
and UO_43 (O_43,N_14760,N_14421);
and UO_44 (O_44,N_14584,N_14224);
xor UO_45 (O_45,N_14724,N_14347);
nand UO_46 (O_46,N_14262,N_14927);
nand UO_47 (O_47,N_14435,N_14209);
nor UO_48 (O_48,N_14836,N_14105);
xnor UO_49 (O_49,N_14746,N_14202);
xnor UO_50 (O_50,N_14315,N_14882);
nor UO_51 (O_51,N_14653,N_14164);
and UO_52 (O_52,N_14322,N_14427);
xor UO_53 (O_53,N_14637,N_14026);
nand UO_54 (O_54,N_14551,N_14979);
or UO_55 (O_55,N_14659,N_14042);
nor UO_56 (O_56,N_14718,N_14412);
xnor UO_57 (O_57,N_14175,N_14426);
nor UO_58 (O_58,N_14128,N_14509);
and UO_59 (O_59,N_14674,N_14054);
nor UO_60 (O_60,N_14989,N_14460);
nand UO_61 (O_61,N_14088,N_14032);
and UO_62 (O_62,N_14331,N_14487);
xor UO_63 (O_63,N_14068,N_14604);
nand UO_64 (O_64,N_14897,N_14665);
and UO_65 (O_65,N_14043,N_14543);
nor UO_66 (O_66,N_14050,N_14259);
nor UO_67 (O_67,N_14574,N_14818);
and UO_68 (O_68,N_14146,N_14995);
nor UO_69 (O_69,N_14933,N_14292);
xor UO_70 (O_70,N_14681,N_14367);
nand UO_71 (O_71,N_14906,N_14496);
nor UO_72 (O_72,N_14723,N_14279);
and UO_73 (O_73,N_14512,N_14375);
and UO_74 (O_74,N_14180,N_14148);
or UO_75 (O_75,N_14008,N_14038);
nand UO_76 (O_76,N_14865,N_14896);
or UO_77 (O_77,N_14630,N_14097);
xnor UO_78 (O_78,N_14900,N_14691);
nor UO_79 (O_79,N_14358,N_14327);
xnor UO_80 (O_80,N_14232,N_14930);
xnor UO_81 (O_81,N_14939,N_14791);
nor UO_82 (O_82,N_14757,N_14454);
or UO_83 (O_83,N_14482,N_14272);
or UO_84 (O_84,N_14260,N_14242);
xnor UO_85 (O_85,N_14123,N_14725);
or UO_86 (O_86,N_14861,N_14531);
xnor UO_87 (O_87,N_14632,N_14899);
nor UO_88 (O_88,N_14176,N_14355);
nor UO_89 (O_89,N_14607,N_14109);
nor UO_90 (O_90,N_14309,N_14745);
and UO_91 (O_91,N_14895,N_14541);
nand UO_92 (O_92,N_14571,N_14415);
nor UO_93 (O_93,N_14219,N_14444);
nor UO_94 (O_94,N_14785,N_14321);
nand UO_95 (O_95,N_14915,N_14391);
and UO_96 (O_96,N_14727,N_14768);
nor UO_97 (O_97,N_14949,N_14300);
nor UO_98 (O_98,N_14436,N_14328);
xor UO_99 (O_99,N_14382,N_14127);
xnor UO_100 (O_100,N_14177,N_14667);
xor UO_101 (O_101,N_14077,N_14223);
and UO_102 (O_102,N_14302,N_14185);
xnor UO_103 (O_103,N_14153,N_14040);
nand UO_104 (O_104,N_14117,N_14335);
or UO_105 (O_105,N_14886,N_14449);
nor UO_106 (O_106,N_14563,N_14020);
and UO_107 (O_107,N_14439,N_14516);
xnor UO_108 (O_108,N_14474,N_14893);
nor UO_109 (O_109,N_14075,N_14430);
or UO_110 (O_110,N_14542,N_14221);
nor UO_111 (O_111,N_14470,N_14557);
or UO_112 (O_112,N_14783,N_14972);
or UO_113 (O_113,N_14287,N_14904);
xnor UO_114 (O_114,N_14668,N_14264);
nand UO_115 (O_115,N_14431,N_14152);
or UO_116 (O_116,N_14110,N_14612);
nor UO_117 (O_117,N_14787,N_14958);
nand UO_118 (O_118,N_14121,N_14765);
and UO_119 (O_119,N_14012,N_14837);
and UO_120 (O_120,N_14986,N_14846);
xor UO_121 (O_121,N_14789,N_14802);
or UO_122 (O_122,N_14405,N_14049);
nor UO_123 (O_123,N_14140,N_14348);
nand UO_124 (O_124,N_14285,N_14687);
and UO_125 (O_125,N_14658,N_14592);
nand UO_126 (O_126,N_14810,N_14084);
and UO_127 (O_127,N_14633,N_14337);
xnor UO_128 (O_128,N_14617,N_14453);
nand UO_129 (O_129,N_14597,N_14850);
nor UO_130 (O_130,N_14812,N_14840);
nor UO_131 (O_131,N_14317,N_14740);
xnor UO_132 (O_132,N_14418,N_14621);
nand UO_133 (O_133,N_14875,N_14877);
or UO_134 (O_134,N_14420,N_14540);
nor UO_135 (O_135,N_14490,N_14590);
nor UO_136 (O_136,N_14273,N_14644);
or UO_137 (O_137,N_14971,N_14263);
nor UO_138 (O_138,N_14374,N_14800);
nand UO_139 (O_139,N_14499,N_14781);
and UO_140 (O_140,N_14606,N_14094);
nor UO_141 (O_141,N_14000,N_14005);
nor UO_142 (O_142,N_14932,N_14294);
xor UO_143 (O_143,N_14425,N_14599);
and UO_144 (O_144,N_14652,N_14343);
xor UO_145 (O_145,N_14329,N_14610);
nor UO_146 (O_146,N_14742,N_14194);
or UO_147 (O_147,N_14848,N_14238);
xnor UO_148 (O_148,N_14346,N_14773);
or UO_149 (O_149,N_14689,N_14605);
xnor UO_150 (O_150,N_14318,N_14464);
or UO_151 (O_151,N_14838,N_14060);
xor UO_152 (O_152,N_14553,N_14118);
nand UO_153 (O_153,N_14145,N_14467);
or UO_154 (O_154,N_14371,N_14623);
and UO_155 (O_155,N_14664,N_14650);
nor UO_156 (O_156,N_14853,N_14296);
xor UO_157 (O_157,N_14562,N_14138);
xnor UO_158 (O_158,N_14844,N_14713);
nand UO_159 (O_159,N_14929,N_14295);
nand UO_160 (O_160,N_14226,N_14596);
or UO_161 (O_161,N_14922,N_14924);
and UO_162 (O_162,N_14181,N_14053);
nor UO_163 (O_163,N_14361,N_14173);
nor UO_164 (O_164,N_14547,N_14210);
xnor UO_165 (O_165,N_14411,N_14268);
nor UO_166 (O_166,N_14847,N_14549);
xnor UO_167 (O_167,N_14640,N_14578);
xor UO_168 (O_168,N_14763,N_14398);
nor UO_169 (O_169,N_14353,N_14390);
and UO_170 (O_170,N_14860,N_14332);
xnor UO_171 (O_171,N_14910,N_14207);
and UO_172 (O_172,N_14830,N_14786);
and UO_173 (O_173,N_14828,N_14651);
and UO_174 (O_174,N_14506,N_14702);
or UO_175 (O_175,N_14734,N_14743);
and UO_176 (O_176,N_14526,N_14305);
nand UO_177 (O_177,N_14434,N_14834);
nor UO_178 (O_178,N_14282,N_14873);
xor UO_179 (O_179,N_14554,N_14767);
xor UO_180 (O_180,N_14437,N_14912);
or UO_181 (O_181,N_14780,N_14911);
and UO_182 (O_182,N_14172,N_14517);
xor UO_183 (O_183,N_14407,N_14946);
and UO_184 (O_184,N_14593,N_14715);
nand UO_185 (O_185,N_14334,N_14647);
nand UO_186 (O_186,N_14045,N_14485);
nor UO_187 (O_187,N_14120,N_14566);
or UO_188 (O_188,N_14766,N_14937);
xnor UO_189 (O_189,N_14947,N_14338);
nand UO_190 (O_190,N_14885,N_14313);
and UO_191 (O_191,N_14580,N_14814);
or UO_192 (O_192,N_14133,N_14306);
nor UO_193 (O_193,N_14953,N_14684);
or UO_194 (O_194,N_14641,N_14649);
or UO_195 (O_195,N_14792,N_14680);
and UO_196 (O_196,N_14729,N_14615);
nor UO_197 (O_197,N_14141,N_14225);
and UO_198 (O_198,N_14033,N_14483);
xnor UO_199 (O_199,N_14211,N_14007);
xnor UO_200 (O_200,N_14627,N_14197);
nor UO_201 (O_201,N_14356,N_14868);
nor UO_202 (O_202,N_14274,N_14316);
or UO_203 (O_203,N_14469,N_14761);
nor UO_204 (O_204,N_14662,N_14835);
and UO_205 (O_205,N_14102,N_14611);
nand UO_206 (O_206,N_14585,N_14183);
or UO_207 (O_207,N_14749,N_14721);
nor UO_208 (O_208,N_14991,N_14236);
or UO_209 (O_209,N_14530,N_14826);
xnor UO_210 (O_210,N_14212,N_14402);
or UO_211 (O_211,N_14270,N_14824);
and UO_212 (O_212,N_14770,N_14708);
nor UO_213 (O_213,N_14620,N_14345);
nand UO_214 (O_214,N_14645,N_14283);
and UO_215 (O_215,N_14975,N_14258);
or UO_216 (O_216,N_14643,N_14119);
nor UO_217 (O_217,N_14017,N_14737);
nor UO_218 (O_218,N_14064,N_14942);
nand UO_219 (O_219,N_14235,N_14862);
or UO_220 (O_220,N_14728,N_14962);
or UO_221 (O_221,N_14872,N_14031);
and UO_222 (O_222,N_14669,N_14090);
nand UO_223 (O_223,N_14815,N_14735);
xnor UO_224 (O_224,N_14406,N_14699);
xor UO_225 (O_225,N_14992,N_14220);
nor UO_226 (O_226,N_14717,N_14881);
xnor UO_227 (O_227,N_14944,N_14030);
or UO_228 (O_228,N_14558,N_14304);
xnor UO_229 (O_229,N_14484,N_14750);
and UO_230 (O_230,N_14945,N_14581);
or UO_231 (O_231,N_14214,N_14925);
nand UO_232 (O_232,N_14513,N_14446);
xor UO_233 (O_233,N_14113,N_14480);
or UO_234 (O_234,N_14871,N_14794);
xor UO_235 (O_235,N_14998,N_14174);
nand UO_236 (O_236,N_14336,N_14672);
or UO_237 (O_237,N_14660,N_14798);
nand UO_238 (O_238,N_14290,N_14970);
or UO_239 (O_239,N_14753,N_14276);
xnor UO_240 (O_240,N_14381,N_14352);
or UO_241 (O_241,N_14368,N_14186);
nor UO_242 (O_242,N_14363,N_14739);
nor UO_243 (O_243,N_14086,N_14428);
xor UO_244 (O_244,N_14982,N_14806);
and UO_245 (O_245,N_14072,N_14114);
xnor UO_246 (O_246,N_14491,N_14308);
or UO_247 (O_247,N_14822,N_14618);
or UO_248 (O_248,N_14429,N_14079);
and UO_249 (O_249,N_14104,N_14246);
and UO_250 (O_250,N_14994,N_14624);
or UO_251 (O_251,N_14646,N_14070);
xnor UO_252 (O_252,N_14366,N_14159);
or UO_253 (O_253,N_14522,N_14414);
nand UO_254 (O_254,N_14560,N_14216);
and UO_255 (O_255,N_14073,N_14936);
nor UO_256 (O_256,N_14021,N_14001);
nand UO_257 (O_257,N_14171,N_14187);
nand UO_258 (O_258,N_14445,N_14150);
or UO_259 (O_259,N_14011,N_14416);
xor UO_260 (O_260,N_14379,N_14333);
nand UO_261 (O_261,N_14964,N_14364);
xnor UO_262 (O_262,N_14843,N_14310);
xnor UO_263 (O_263,N_14298,N_14143);
xnor UO_264 (O_264,N_14555,N_14100);
and UO_265 (O_265,N_14854,N_14369);
nand UO_266 (O_266,N_14413,N_14663);
and UO_267 (O_267,N_14111,N_14249);
and UO_268 (O_268,N_14476,N_14980);
nand UO_269 (O_269,N_14320,N_14576);
and UO_270 (O_270,N_14999,N_14771);
and UO_271 (O_271,N_14507,N_14488);
nand UO_272 (O_272,N_14443,N_14864);
or UO_273 (O_273,N_14676,N_14813);
and UO_274 (O_274,N_14018,N_14544);
nand UO_275 (O_275,N_14524,N_14206);
nor UO_276 (O_276,N_14515,N_14811);
or UO_277 (O_277,N_14514,N_14564);
and UO_278 (O_278,N_14670,N_14548);
xor UO_279 (O_279,N_14473,N_14888);
nor UO_280 (O_280,N_14990,N_14178);
nor UO_281 (O_281,N_14777,N_14055);
nor UO_282 (O_282,N_14248,N_14132);
nor UO_283 (O_283,N_14587,N_14433);
nand UO_284 (O_284,N_14025,N_14378);
and UO_285 (O_285,N_14827,N_14909);
xor UO_286 (O_286,N_14376,N_14231);
nand UO_287 (O_287,N_14227,N_14711);
nand UO_288 (O_288,N_14362,N_14208);
nor UO_289 (O_289,N_14385,N_14856);
and UO_290 (O_290,N_14442,N_14311);
and UO_291 (O_291,N_14738,N_14149);
xor UO_292 (O_292,N_14511,N_14908);
and UO_293 (O_293,N_14807,N_14688);
xor UO_294 (O_294,N_14189,N_14901);
nor UO_295 (O_295,N_14503,N_14839);
nor UO_296 (O_296,N_14230,N_14631);
nor UO_297 (O_297,N_14692,N_14913);
xor UO_298 (O_298,N_14504,N_14481);
nor UO_299 (O_299,N_14969,N_14797);
xnor UO_300 (O_300,N_14619,N_14126);
xnor UO_301 (O_301,N_14301,N_14389);
or UO_302 (O_302,N_14525,N_14694);
or UO_303 (O_303,N_14182,N_14098);
nor UO_304 (O_304,N_14016,N_14714);
or UO_305 (O_305,N_14387,N_14215);
and UO_306 (O_306,N_14479,N_14092);
nand UO_307 (O_307,N_14907,N_14679);
and UO_308 (O_308,N_14319,N_14066);
nand UO_309 (O_309,N_14061,N_14696);
or UO_310 (O_310,N_14239,N_14466);
xnor UO_311 (O_311,N_14459,N_14833);
or UO_312 (O_312,N_14096,N_14058);
xnor UO_313 (O_313,N_14409,N_14029);
nand UO_314 (O_314,N_14565,N_14591);
xnor UO_315 (O_315,N_14920,N_14154);
or UO_316 (O_316,N_14167,N_14698);
nand UO_317 (O_317,N_14165,N_14577);
nand UO_318 (O_318,N_14796,N_14447);
nor UO_319 (O_319,N_14324,N_14472);
or UO_320 (O_320,N_14700,N_14056);
xnor UO_321 (O_321,N_14626,N_14987);
xnor UO_322 (O_322,N_14934,N_14751);
or UO_323 (O_323,N_14921,N_14917);
and UO_324 (O_324,N_14758,N_14816);
and UO_325 (O_325,N_14004,N_14754);
and UO_326 (O_326,N_14065,N_14655);
nand UO_327 (O_327,N_14790,N_14423);
nor UO_328 (O_328,N_14465,N_14393);
or UO_329 (O_329,N_14122,N_14261);
and UO_330 (O_330,N_14396,N_14716);
nand UO_331 (O_331,N_14424,N_14157);
nand UO_332 (O_332,N_14508,N_14603);
and UO_333 (O_333,N_14325,N_14961);
xnor UO_334 (O_334,N_14938,N_14891);
xnor UO_335 (O_335,N_14951,N_14191);
nand UO_336 (O_336,N_14196,N_14981);
and UO_337 (O_337,N_14625,N_14218);
xnor UO_338 (O_338,N_14408,N_14450);
nor UO_339 (O_339,N_14952,N_14831);
xnor UO_340 (O_340,N_14440,N_14756);
and UO_341 (O_341,N_14213,N_14253);
or UO_342 (O_342,N_14222,N_14083);
or UO_343 (O_343,N_14350,N_14037);
and UO_344 (O_344,N_14410,N_14520);
nand UO_345 (O_345,N_14190,N_14588);
nor UO_346 (O_346,N_14297,N_14028);
or UO_347 (O_347,N_14985,N_14432);
and UO_348 (O_348,N_14567,N_14266);
and UO_349 (O_349,N_14795,N_14200);
nor UO_350 (O_350,N_14629,N_14741);
nand UO_351 (O_351,N_14392,N_14046);
or UO_352 (O_352,N_14163,N_14501);
or UO_353 (O_353,N_14825,N_14874);
or UO_354 (O_354,N_14523,N_14036);
nand UO_355 (O_355,N_14257,N_14842);
nor UO_356 (O_356,N_14351,N_14788);
and UO_357 (O_357,N_14044,N_14528);
nand UO_358 (O_358,N_14247,N_14022);
nor UO_359 (O_359,N_14339,N_14976);
nand UO_360 (O_360,N_14286,N_14636);
nand UO_361 (O_361,N_14707,N_14251);
or UO_362 (O_362,N_14468,N_14583);
nor UO_363 (O_363,N_14748,N_14203);
xnor UO_364 (O_364,N_14139,N_14395);
and UO_365 (O_365,N_14948,N_14284);
xnor UO_366 (O_366,N_14857,N_14115);
or UO_367 (O_367,N_14455,N_14288);
nand UO_368 (O_368,N_14451,N_14863);
nand UO_369 (O_369,N_14074,N_14866);
or UO_370 (O_370,N_14492,N_14142);
nand UO_371 (O_371,N_14616,N_14372);
and UO_372 (O_372,N_14561,N_14701);
and UO_373 (O_373,N_14820,N_14456);
nor UO_374 (O_374,N_14956,N_14063);
nand UO_375 (O_375,N_14582,N_14107);
and UO_376 (O_376,N_14841,N_14678);
and UO_377 (O_377,N_14095,N_14638);
nand UO_378 (O_378,N_14984,N_14486);
nand UO_379 (O_379,N_14144,N_14733);
nand UO_380 (O_380,N_14589,N_14744);
nand UO_381 (O_381,N_14575,N_14101);
nand UO_382 (O_382,N_14996,N_14081);
and UO_383 (O_383,N_14719,N_14495);
nor UO_384 (O_384,N_14250,N_14441);
and UO_385 (O_385,N_14883,N_14609);
or UO_386 (O_386,N_14326,N_14778);
xor UO_387 (O_387,N_14931,N_14918);
nand UO_388 (O_388,N_14394,N_14198);
xnor UO_389 (O_389,N_14188,N_14752);
or UO_390 (O_390,N_14052,N_14808);
nor UO_391 (O_391,N_14417,N_14106);
or UO_392 (O_392,N_14704,N_14009);
xor UO_393 (O_393,N_14764,N_14902);
nand UO_394 (O_394,N_14158,N_14772);
and UO_395 (O_395,N_14628,N_14463);
and UO_396 (O_396,N_14505,N_14401);
and UO_397 (O_397,N_14131,N_14341);
and UO_398 (O_398,N_14685,N_14817);
and UO_399 (O_399,N_14419,N_14769);
or UO_400 (O_400,N_14988,N_14047);
or UO_401 (O_401,N_14697,N_14977);
nand UO_402 (O_402,N_14775,N_14705);
and UO_403 (O_403,N_14823,N_14130);
nor UO_404 (O_404,N_14010,N_14293);
nor UO_405 (O_405,N_14002,N_14974);
xor UO_406 (O_406,N_14314,N_14013);
and UO_407 (O_407,N_14832,N_14265);
xnor UO_408 (O_408,N_14879,N_14359);
nor UO_409 (O_409,N_14365,N_14935);
and UO_410 (O_410,N_14535,N_14386);
and UO_411 (O_411,N_14654,N_14869);
nand UO_412 (O_412,N_14855,N_14613);
nor UO_413 (O_413,N_14950,N_14099);
nand UO_414 (O_414,N_14661,N_14966);
xnor UO_415 (O_415,N_14289,N_14642);
and UO_416 (O_416,N_14237,N_14438);
nand UO_417 (O_417,N_14666,N_14878);
nand UO_418 (O_418,N_14914,N_14851);
xor UO_419 (O_419,N_14884,N_14500);
xor UO_420 (O_420,N_14955,N_14041);
and UO_421 (O_421,N_14867,N_14967);
or UO_422 (O_422,N_14370,N_14048);
xnor UO_423 (O_423,N_14518,N_14388);
nor UO_424 (O_424,N_14690,N_14377);
nand UO_425 (O_425,N_14570,N_14546);
and UO_426 (O_426,N_14722,N_14373);
and UO_427 (O_427,N_14147,N_14234);
or UO_428 (O_428,N_14677,N_14903);
and UO_429 (O_429,N_14252,N_14545);
nand UO_430 (O_430,N_14103,N_14635);
nand UO_431 (O_431,N_14634,N_14536);
and UO_432 (O_432,N_14349,N_14360);
nor UO_433 (O_433,N_14755,N_14859);
or UO_434 (O_434,N_14229,N_14091);
nor UO_435 (O_435,N_14870,N_14383);
xnor UO_436 (O_436,N_14452,N_14532);
or UO_437 (O_437,N_14586,N_14550);
nand UO_438 (O_438,N_14458,N_14940);
and UO_439 (O_439,N_14344,N_14478);
or UO_440 (O_440,N_14594,N_14240);
or UO_441 (O_441,N_14600,N_14819);
nand UO_442 (O_442,N_14494,N_14983);
nor UO_443 (O_443,N_14803,N_14709);
nand UO_444 (O_444,N_14502,N_14759);
nand UO_445 (O_445,N_14614,N_14080);
nor UO_446 (O_446,N_14166,N_14954);
nand UO_447 (O_447,N_14726,N_14804);
or UO_448 (O_448,N_14639,N_14014);
and UO_449 (O_449,N_14244,N_14968);
or UO_450 (O_450,N_14608,N_14858);
nor UO_451 (O_451,N_14736,N_14656);
and UO_452 (O_452,N_14568,N_14019);
xnor UO_453 (O_453,N_14475,N_14024);
and UO_454 (O_454,N_14280,N_14354);
or UO_455 (O_455,N_14683,N_14682);
nand UO_456 (O_456,N_14462,N_14161);
xnor UO_457 (O_457,N_14027,N_14497);
nand UO_458 (O_458,N_14534,N_14960);
xor UO_459 (O_459,N_14849,N_14552);
or UO_460 (O_460,N_14730,N_14559);
nor UO_461 (O_461,N_14693,N_14137);
xnor UO_462 (O_462,N_14928,N_14422);
nor UO_463 (O_463,N_14057,N_14731);
nand UO_464 (O_464,N_14160,N_14112);
xor UO_465 (O_465,N_14134,N_14448);
nor UO_466 (O_466,N_14089,N_14712);
and UO_467 (O_467,N_14898,N_14471);
xor UO_468 (O_468,N_14342,N_14039);
or UO_469 (O_469,N_14241,N_14087);
or UO_470 (O_470,N_14129,N_14894);
or UO_471 (O_471,N_14579,N_14943);
or UO_472 (O_472,N_14281,N_14179);
nand UO_473 (O_473,N_14184,N_14291);
or UO_474 (O_474,N_14271,N_14380);
and UO_475 (O_475,N_14959,N_14573);
nor UO_476 (O_476,N_14941,N_14973);
nand UO_477 (O_477,N_14193,N_14034);
nand UO_478 (O_478,N_14706,N_14784);
or UO_479 (O_479,N_14801,N_14890);
xor UO_480 (O_480,N_14569,N_14762);
or UO_481 (O_481,N_14051,N_14006);
nand UO_482 (O_482,N_14852,N_14782);
and UO_483 (O_483,N_14108,N_14312);
nor UO_484 (O_484,N_14078,N_14892);
nor UO_485 (O_485,N_14675,N_14125);
and UO_486 (O_486,N_14340,N_14124);
xnor UO_487 (O_487,N_14076,N_14015);
nor UO_488 (O_488,N_14622,N_14192);
xor UO_489 (O_489,N_14461,N_14035);
or UO_490 (O_490,N_14156,N_14926);
xnor UO_491 (O_491,N_14889,N_14533);
or UO_492 (O_492,N_14598,N_14673);
xnor UO_493 (O_493,N_14228,N_14205);
nand UO_494 (O_494,N_14357,N_14537);
or UO_495 (O_495,N_14776,N_14082);
and UO_496 (O_496,N_14256,N_14217);
or UO_497 (O_497,N_14151,N_14243);
nand UO_498 (O_498,N_14671,N_14880);
or UO_499 (O_499,N_14071,N_14116);
xnor UO_500 (O_500,N_14129,N_14251);
nand UO_501 (O_501,N_14737,N_14246);
nor UO_502 (O_502,N_14780,N_14518);
xor UO_503 (O_503,N_14802,N_14945);
nand UO_504 (O_504,N_14776,N_14745);
and UO_505 (O_505,N_14636,N_14775);
or UO_506 (O_506,N_14020,N_14864);
xor UO_507 (O_507,N_14110,N_14114);
nand UO_508 (O_508,N_14340,N_14581);
nor UO_509 (O_509,N_14191,N_14528);
or UO_510 (O_510,N_14662,N_14135);
or UO_511 (O_511,N_14359,N_14728);
and UO_512 (O_512,N_14540,N_14194);
or UO_513 (O_513,N_14821,N_14874);
nand UO_514 (O_514,N_14500,N_14609);
and UO_515 (O_515,N_14705,N_14148);
and UO_516 (O_516,N_14194,N_14518);
nor UO_517 (O_517,N_14561,N_14223);
nor UO_518 (O_518,N_14439,N_14181);
or UO_519 (O_519,N_14238,N_14737);
nor UO_520 (O_520,N_14392,N_14617);
nand UO_521 (O_521,N_14327,N_14417);
xor UO_522 (O_522,N_14908,N_14485);
or UO_523 (O_523,N_14799,N_14053);
nand UO_524 (O_524,N_14633,N_14312);
and UO_525 (O_525,N_14371,N_14655);
xnor UO_526 (O_526,N_14315,N_14187);
nand UO_527 (O_527,N_14146,N_14447);
or UO_528 (O_528,N_14775,N_14344);
nand UO_529 (O_529,N_14611,N_14636);
nor UO_530 (O_530,N_14886,N_14844);
xnor UO_531 (O_531,N_14089,N_14241);
xor UO_532 (O_532,N_14767,N_14440);
and UO_533 (O_533,N_14227,N_14526);
nor UO_534 (O_534,N_14934,N_14128);
xnor UO_535 (O_535,N_14570,N_14843);
and UO_536 (O_536,N_14428,N_14654);
or UO_537 (O_537,N_14752,N_14684);
nand UO_538 (O_538,N_14621,N_14378);
or UO_539 (O_539,N_14325,N_14900);
nand UO_540 (O_540,N_14843,N_14883);
or UO_541 (O_541,N_14961,N_14602);
nor UO_542 (O_542,N_14776,N_14154);
nor UO_543 (O_543,N_14416,N_14972);
xnor UO_544 (O_544,N_14399,N_14669);
nand UO_545 (O_545,N_14029,N_14956);
nand UO_546 (O_546,N_14824,N_14559);
xnor UO_547 (O_547,N_14851,N_14930);
or UO_548 (O_548,N_14706,N_14186);
nand UO_549 (O_549,N_14915,N_14305);
nor UO_550 (O_550,N_14347,N_14336);
and UO_551 (O_551,N_14215,N_14384);
xnor UO_552 (O_552,N_14275,N_14886);
xnor UO_553 (O_553,N_14378,N_14518);
nor UO_554 (O_554,N_14163,N_14091);
and UO_555 (O_555,N_14266,N_14663);
nor UO_556 (O_556,N_14236,N_14964);
or UO_557 (O_557,N_14354,N_14620);
nand UO_558 (O_558,N_14206,N_14732);
nor UO_559 (O_559,N_14801,N_14389);
nor UO_560 (O_560,N_14081,N_14700);
nor UO_561 (O_561,N_14624,N_14348);
nand UO_562 (O_562,N_14356,N_14957);
xnor UO_563 (O_563,N_14546,N_14505);
or UO_564 (O_564,N_14107,N_14360);
nor UO_565 (O_565,N_14967,N_14987);
and UO_566 (O_566,N_14956,N_14363);
nand UO_567 (O_567,N_14061,N_14259);
xnor UO_568 (O_568,N_14714,N_14565);
nor UO_569 (O_569,N_14080,N_14603);
nand UO_570 (O_570,N_14429,N_14256);
nand UO_571 (O_571,N_14237,N_14358);
xnor UO_572 (O_572,N_14459,N_14815);
nor UO_573 (O_573,N_14391,N_14659);
xor UO_574 (O_574,N_14267,N_14050);
xnor UO_575 (O_575,N_14110,N_14868);
xor UO_576 (O_576,N_14491,N_14380);
and UO_577 (O_577,N_14271,N_14908);
nand UO_578 (O_578,N_14013,N_14531);
or UO_579 (O_579,N_14599,N_14780);
xor UO_580 (O_580,N_14359,N_14090);
nor UO_581 (O_581,N_14684,N_14281);
nor UO_582 (O_582,N_14658,N_14504);
xor UO_583 (O_583,N_14274,N_14353);
nor UO_584 (O_584,N_14600,N_14842);
nor UO_585 (O_585,N_14820,N_14911);
xor UO_586 (O_586,N_14426,N_14333);
xnor UO_587 (O_587,N_14852,N_14506);
and UO_588 (O_588,N_14786,N_14052);
nand UO_589 (O_589,N_14998,N_14421);
nand UO_590 (O_590,N_14611,N_14078);
or UO_591 (O_591,N_14401,N_14821);
nand UO_592 (O_592,N_14030,N_14352);
xnor UO_593 (O_593,N_14080,N_14121);
nor UO_594 (O_594,N_14676,N_14207);
and UO_595 (O_595,N_14605,N_14042);
nand UO_596 (O_596,N_14884,N_14869);
nor UO_597 (O_597,N_14710,N_14993);
xor UO_598 (O_598,N_14474,N_14999);
nor UO_599 (O_599,N_14836,N_14216);
nor UO_600 (O_600,N_14487,N_14387);
xnor UO_601 (O_601,N_14091,N_14124);
nand UO_602 (O_602,N_14955,N_14199);
xor UO_603 (O_603,N_14041,N_14032);
xnor UO_604 (O_604,N_14682,N_14854);
nor UO_605 (O_605,N_14678,N_14065);
and UO_606 (O_606,N_14424,N_14847);
and UO_607 (O_607,N_14211,N_14428);
xnor UO_608 (O_608,N_14061,N_14676);
nor UO_609 (O_609,N_14348,N_14948);
nor UO_610 (O_610,N_14943,N_14468);
xor UO_611 (O_611,N_14906,N_14864);
nor UO_612 (O_612,N_14508,N_14284);
or UO_613 (O_613,N_14665,N_14143);
nor UO_614 (O_614,N_14331,N_14554);
nor UO_615 (O_615,N_14096,N_14611);
nand UO_616 (O_616,N_14341,N_14072);
xor UO_617 (O_617,N_14228,N_14719);
or UO_618 (O_618,N_14780,N_14500);
nor UO_619 (O_619,N_14198,N_14643);
and UO_620 (O_620,N_14010,N_14515);
and UO_621 (O_621,N_14253,N_14942);
xor UO_622 (O_622,N_14467,N_14696);
xnor UO_623 (O_623,N_14603,N_14546);
or UO_624 (O_624,N_14394,N_14134);
or UO_625 (O_625,N_14360,N_14781);
nor UO_626 (O_626,N_14636,N_14815);
xnor UO_627 (O_627,N_14844,N_14001);
and UO_628 (O_628,N_14209,N_14676);
nand UO_629 (O_629,N_14640,N_14519);
nor UO_630 (O_630,N_14640,N_14701);
or UO_631 (O_631,N_14693,N_14266);
and UO_632 (O_632,N_14592,N_14528);
nand UO_633 (O_633,N_14679,N_14921);
nor UO_634 (O_634,N_14857,N_14935);
nor UO_635 (O_635,N_14180,N_14121);
nand UO_636 (O_636,N_14254,N_14165);
or UO_637 (O_637,N_14238,N_14254);
or UO_638 (O_638,N_14639,N_14363);
and UO_639 (O_639,N_14914,N_14104);
and UO_640 (O_640,N_14239,N_14283);
xor UO_641 (O_641,N_14127,N_14476);
nand UO_642 (O_642,N_14276,N_14361);
nand UO_643 (O_643,N_14062,N_14400);
nand UO_644 (O_644,N_14413,N_14184);
xnor UO_645 (O_645,N_14117,N_14128);
or UO_646 (O_646,N_14962,N_14434);
nand UO_647 (O_647,N_14821,N_14174);
and UO_648 (O_648,N_14644,N_14589);
and UO_649 (O_649,N_14328,N_14180);
nor UO_650 (O_650,N_14601,N_14638);
and UO_651 (O_651,N_14473,N_14592);
and UO_652 (O_652,N_14471,N_14468);
nor UO_653 (O_653,N_14617,N_14739);
nand UO_654 (O_654,N_14211,N_14129);
nor UO_655 (O_655,N_14087,N_14171);
xnor UO_656 (O_656,N_14110,N_14542);
and UO_657 (O_657,N_14786,N_14023);
or UO_658 (O_658,N_14610,N_14258);
nand UO_659 (O_659,N_14435,N_14144);
nor UO_660 (O_660,N_14530,N_14231);
nor UO_661 (O_661,N_14602,N_14858);
xnor UO_662 (O_662,N_14328,N_14017);
and UO_663 (O_663,N_14182,N_14653);
and UO_664 (O_664,N_14958,N_14078);
or UO_665 (O_665,N_14266,N_14741);
or UO_666 (O_666,N_14739,N_14355);
xor UO_667 (O_667,N_14707,N_14618);
or UO_668 (O_668,N_14140,N_14585);
nand UO_669 (O_669,N_14335,N_14196);
nor UO_670 (O_670,N_14677,N_14703);
nand UO_671 (O_671,N_14340,N_14121);
and UO_672 (O_672,N_14424,N_14965);
xnor UO_673 (O_673,N_14064,N_14655);
or UO_674 (O_674,N_14032,N_14528);
nand UO_675 (O_675,N_14998,N_14592);
nand UO_676 (O_676,N_14886,N_14442);
nor UO_677 (O_677,N_14701,N_14229);
and UO_678 (O_678,N_14252,N_14762);
and UO_679 (O_679,N_14867,N_14489);
xor UO_680 (O_680,N_14392,N_14093);
nor UO_681 (O_681,N_14368,N_14675);
or UO_682 (O_682,N_14633,N_14674);
nor UO_683 (O_683,N_14265,N_14583);
or UO_684 (O_684,N_14928,N_14352);
and UO_685 (O_685,N_14488,N_14926);
or UO_686 (O_686,N_14446,N_14322);
or UO_687 (O_687,N_14920,N_14356);
or UO_688 (O_688,N_14541,N_14019);
nand UO_689 (O_689,N_14004,N_14982);
nand UO_690 (O_690,N_14099,N_14796);
or UO_691 (O_691,N_14652,N_14853);
nor UO_692 (O_692,N_14670,N_14533);
nor UO_693 (O_693,N_14926,N_14593);
or UO_694 (O_694,N_14072,N_14707);
and UO_695 (O_695,N_14025,N_14939);
or UO_696 (O_696,N_14230,N_14601);
and UO_697 (O_697,N_14830,N_14799);
nor UO_698 (O_698,N_14396,N_14454);
and UO_699 (O_699,N_14121,N_14133);
or UO_700 (O_700,N_14955,N_14643);
and UO_701 (O_701,N_14597,N_14869);
or UO_702 (O_702,N_14647,N_14938);
and UO_703 (O_703,N_14972,N_14848);
xnor UO_704 (O_704,N_14771,N_14638);
nand UO_705 (O_705,N_14726,N_14910);
nand UO_706 (O_706,N_14867,N_14092);
nand UO_707 (O_707,N_14310,N_14215);
nand UO_708 (O_708,N_14104,N_14849);
or UO_709 (O_709,N_14208,N_14798);
xor UO_710 (O_710,N_14988,N_14793);
xor UO_711 (O_711,N_14097,N_14705);
and UO_712 (O_712,N_14957,N_14494);
or UO_713 (O_713,N_14304,N_14809);
xor UO_714 (O_714,N_14867,N_14974);
and UO_715 (O_715,N_14743,N_14125);
or UO_716 (O_716,N_14383,N_14215);
or UO_717 (O_717,N_14084,N_14791);
nor UO_718 (O_718,N_14793,N_14283);
nor UO_719 (O_719,N_14276,N_14736);
nor UO_720 (O_720,N_14364,N_14818);
or UO_721 (O_721,N_14899,N_14635);
and UO_722 (O_722,N_14818,N_14621);
xor UO_723 (O_723,N_14777,N_14087);
xor UO_724 (O_724,N_14884,N_14611);
or UO_725 (O_725,N_14106,N_14651);
or UO_726 (O_726,N_14574,N_14757);
and UO_727 (O_727,N_14380,N_14207);
nor UO_728 (O_728,N_14099,N_14393);
or UO_729 (O_729,N_14306,N_14391);
nand UO_730 (O_730,N_14807,N_14088);
or UO_731 (O_731,N_14042,N_14347);
nor UO_732 (O_732,N_14378,N_14435);
nand UO_733 (O_733,N_14753,N_14162);
nand UO_734 (O_734,N_14677,N_14284);
nor UO_735 (O_735,N_14619,N_14856);
or UO_736 (O_736,N_14088,N_14030);
and UO_737 (O_737,N_14481,N_14055);
nand UO_738 (O_738,N_14762,N_14390);
and UO_739 (O_739,N_14005,N_14661);
nand UO_740 (O_740,N_14935,N_14094);
nor UO_741 (O_741,N_14826,N_14446);
nor UO_742 (O_742,N_14791,N_14513);
nand UO_743 (O_743,N_14126,N_14800);
or UO_744 (O_744,N_14804,N_14802);
nor UO_745 (O_745,N_14659,N_14507);
nand UO_746 (O_746,N_14088,N_14031);
or UO_747 (O_747,N_14984,N_14556);
or UO_748 (O_748,N_14510,N_14519);
and UO_749 (O_749,N_14984,N_14913);
nor UO_750 (O_750,N_14503,N_14376);
and UO_751 (O_751,N_14095,N_14477);
or UO_752 (O_752,N_14087,N_14492);
xor UO_753 (O_753,N_14296,N_14526);
nor UO_754 (O_754,N_14918,N_14396);
xor UO_755 (O_755,N_14251,N_14715);
xor UO_756 (O_756,N_14822,N_14433);
nor UO_757 (O_757,N_14023,N_14831);
or UO_758 (O_758,N_14733,N_14303);
or UO_759 (O_759,N_14617,N_14450);
nor UO_760 (O_760,N_14316,N_14069);
xor UO_761 (O_761,N_14136,N_14041);
or UO_762 (O_762,N_14496,N_14992);
and UO_763 (O_763,N_14508,N_14920);
xor UO_764 (O_764,N_14276,N_14351);
xor UO_765 (O_765,N_14506,N_14041);
nor UO_766 (O_766,N_14336,N_14075);
and UO_767 (O_767,N_14901,N_14847);
and UO_768 (O_768,N_14941,N_14002);
nand UO_769 (O_769,N_14977,N_14766);
and UO_770 (O_770,N_14509,N_14975);
xor UO_771 (O_771,N_14961,N_14098);
and UO_772 (O_772,N_14344,N_14543);
or UO_773 (O_773,N_14138,N_14396);
and UO_774 (O_774,N_14091,N_14386);
nand UO_775 (O_775,N_14112,N_14113);
xor UO_776 (O_776,N_14494,N_14617);
xor UO_777 (O_777,N_14911,N_14824);
xor UO_778 (O_778,N_14112,N_14750);
xnor UO_779 (O_779,N_14362,N_14434);
nor UO_780 (O_780,N_14131,N_14384);
or UO_781 (O_781,N_14698,N_14894);
nand UO_782 (O_782,N_14962,N_14694);
nor UO_783 (O_783,N_14965,N_14280);
or UO_784 (O_784,N_14927,N_14274);
xor UO_785 (O_785,N_14936,N_14411);
or UO_786 (O_786,N_14214,N_14679);
nor UO_787 (O_787,N_14884,N_14085);
or UO_788 (O_788,N_14364,N_14359);
or UO_789 (O_789,N_14299,N_14435);
and UO_790 (O_790,N_14252,N_14076);
xnor UO_791 (O_791,N_14653,N_14127);
nand UO_792 (O_792,N_14628,N_14943);
or UO_793 (O_793,N_14227,N_14032);
and UO_794 (O_794,N_14757,N_14898);
xor UO_795 (O_795,N_14287,N_14391);
nor UO_796 (O_796,N_14547,N_14845);
and UO_797 (O_797,N_14994,N_14400);
and UO_798 (O_798,N_14035,N_14658);
or UO_799 (O_799,N_14688,N_14109);
nor UO_800 (O_800,N_14107,N_14250);
nand UO_801 (O_801,N_14466,N_14150);
and UO_802 (O_802,N_14651,N_14344);
xor UO_803 (O_803,N_14153,N_14246);
nor UO_804 (O_804,N_14966,N_14184);
xnor UO_805 (O_805,N_14855,N_14732);
nand UO_806 (O_806,N_14995,N_14889);
nor UO_807 (O_807,N_14180,N_14381);
and UO_808 (O_808,N_14986,N_14570);
xor UO_809 (O_809,N_14163,N_14631);
nand UO_810 (O_810,N_14594,N_14691);
xor UO_811 (O_811,N_14085,N_14982);
nor UO_812 (O_812,N_14652,N_14873);
nor UO_813 (O_813,N_14101,N_14135);
nor UO_814 (O_814,N_14751,N_14891);
nor UO_815 (O_815,N_14781,N_14193);
or UO_816 (O_816,N_14678,N_14408);
nand UO_817 (O_817,N_14917,N_14616);
or UO_818 (O_818,N_14397,N_14305);
and UO_819 (O_819,N_14938,N_14628);
nor UO_820 (O_820,N_14862,N_14818);
or UO_821 (O_821,N_14430,N_14986);
nand UO_822 (O_822,N_14909,N_14292);
and UO_823 (O_823,N_14658,N_14686);
nand UO_824 (O_824,N_14667,N_14941);
and UO_825 (O_825,N_14146,N_14340);
and UO_826 (O_826,N_14449,N_14987);
nand UO_827 (O_827,N_14008,N_14578);
nor UO_828 (O_828,N_14022,N_14117);
and UO_829 (O_829,N_14970,N_14386);
or UO_830 (O_830,N_14135,N_14625);
nor UO_831 (O_831,N_14963,N_14139);
or UO_832 (O_832,N_14358,N_14896);
or UO_833 (O_833,N_14575,N_14841);
nand UO_834 (O_834,N_14540,N_14314);
nand UO_835 (O_835,N_14735,N_14133);
and UO_836 (O_836,N_14802,N_14480);
and UO_837 (O_837,N_14686,N_14970);
xnor UO_838 (O_838,N_14361,N_14574);
or UO_839 (O_839,N_14728,N_14729);
and UO_840 (O_840,N_14837,N_14477);
nand UO_841 (O_841,N_14189,N_14753);
or UO_842 (O_842,N_14202,N_14404);
nand UO_843 (O_843,N_14402,N_14779);
or UO_844 (O_844,N_14689,N_14881);
or UO_845 (O_845,N_14068,N_14693);
and UO_846 (O_846,N_14411,N_14904);
nand UO_847 (O_847,N_14606,N_14911);
and UO_848 (O_848,N_14678,N_14236);
nor UO_849 (O_849,N_14051,N_14743);
nor UO_850 (O_850,N_14801,N_14257);
or UO_851 (O_851,N_14636,N_14496);
or UO_852 (O_852,N_14990,N_14499);
nor UO_853 (O_853,N_14801,N_14545);
or UO_854 (O_854,N_14844,N_14670);
nand UO_855 (O_855,N_14982,N_14321);
and UO_856 (O_856,N_14547,N_14404);
and UO_857 (O_857,N_14657,N_14146);
or UO_858 (O_858,N_14237,N_14031);
xor UO_859 (O_859,N_14146,N_14761);
nor UO_860 (O_860,N_14169,N_14348);
and UO_861 (O_861,N_14727,N_14392);
nor UO_862 (O_862,N_14471,N_14938);
xnor UO_863 (O_863,N_14607,N_14709);
xnor UO_864 (O_864,N_14256,N_14845);
or UO_865 (O_865,N_14641,N_14702);
and UO_866 (O_866,N_14064,N_14755);
xor UO_867 (O_867,N_14008,N_14372);
and UO_868 (O_868,N_14635,N_14002);
xor UO_869 (O_869,N_14946,N_14236);
or UO_870 (O_870,N_14426,N_14458);
xnor UO_871 (O_871,N_14772,N_14025);
and UO_872 (O_872,N_14089,N_14142);
or UO_873 (O_873,N_14349,N_14314);
nand UO_874 (O_874,N_14716,N_14793);
nor UO_875 (O_875,N_14321,N_14837);
or UO_876 (O_876,N_14013,N_14651);
nand UO_877 (O_877,N_14653,N_14534);
or UO_878 (O_878,N_14832,N_14549);
or UO_879 (O_879,N_14471,N_14585);
xnor UO_880 (O_880,N_14898,N_14109);
and UO_881 (O_881,N_14344,N_14999);
xnor UO_882 (O_882,N_14092,N_14021);
nand UO_883 (O_883,N_14695,N_14279);
and UO_884 (O_884,N_14044,N_14103);
xnor UO_885 (O_885,N_14427,N_14577);
xnor UO_886 (O_886,N_14825,N_14067);
nand UO_887 (O_887,N_14164,N_14773);
or UO_888 (O_888,N_14711,N_14080);
xor UO_889 (O_889,N_14528,N_14786);
nor UO_890 (O_890,N_14362,N_14198);
or UO_891 (O_891,N_14322,N_14480);
nand UO_892 (O_892,N_14257,N_14991);
and UO_893 (O_893,N_14781,N_14796);
nand UO_894 (O_894,N_14363,N_14555);
and UO_895 (O_895,N_14144,N_14999);
nand UO_896 (O_896,N_14232,N_14220);
and UO_897 (O_897,N_14619,N_14604);
xor UO_898 (O_898,N_14848,N_14760);
or UO_899 (O_899,N_14506,N_14562);
nor UO_900 (O_900,N_14385,N_14149);
nand UO_901 (O_901,N_14895,N_14585);
nand UO_902 (O_902,N_14838,N_14441);
xnor UO_903 (O_903,N_14570,N_14699);
and UO_904 (O_904,N_14433,N_14676);
nor UO_905 (O_905,N_14508,N_14562);
xor UO_906 (O_906,N_14501,N_14211);
or UO_907 (O_907,N_14083,N_14494);
nor UO_908 (O_908,N_14969,N_14780);
nand UO_909 (O_909,N_14543,N_14471);
nand UO_910 (O_910,N_14397,N_14932);
nand UO_911 (O_911,N_14728,N_14784);
and UO_912 (O_912,N_14707,N_14823);
and UO_913 (O_913,N_14377,N_14187);
nor UO_914 (O_914,N_14400,N_14984);
and UO_915 (O_915,N_14693,N_14735);
and UO_916 (O_916,N_14361,N_14495);
nand UO_917 (O_917,N_14122,N_14255);
xor UO_918 (O_918,N_14298,N_14983);
nand UO_919 (O_919,N_14909,N_14993);
or UO_920 (O_920,N_14509,N_14241);
and UO_921 (O_921,N_14117,N_14383);
nor UO_922 (O_922,N_14563,N_14127);
and UO_923 (O_923,N_14340,N_14553);
nand UO_924 (O_924,N_14100,N_14895);
or UO_925 (O_925,N_14472,N_14376);
xor UO_926 (O_926,N_14088,N_14738);
or UO_927 (O_927,N_14594,N_14042);
nor UO_928 (O_928,N_14850,N_14322);
nand UO_929 (O_929,N_14582,N_14391);
nor UO_930 (O_930,N_14089,N_14069);
nor UO_931 (O_931,N_14721,N_14147);
nand UO_932 (O_932,N_14994,N_14992);
nand UO_933 (O_933,N_14084,N_14703);
and UO_934 (O_934,N_14009,N_14859);
nand UO_935 (O_935,N_14523,N_14003);
nand UO_936 (O_936,N_14361,N_14721);
nand UO_937 (O_937,N_14901,N_14382);
or UO_938 (O_938,N_14811,N_14634);
and UO_939 (O_939,N_14282,N_14735);
or UO_940 (O_940,N_14561,N_14723);
nand UO_941 (O_941,N_14017,N_14151);
and UO_942 (O_942,N_14687,N_14427);
or UO_943 (O_943,N_14552,N_14345);
and UO_944 (O_944,N_14542,N_14799);
and UO_945 (O_945,N_14769,N_14199);
or UO_946 (O_946,N_14590,N_14122);
xor UO_947 (O_947,N_14966,N_14667);
nand UO_948 (O_948,N_14616,N_14452);
or UO_949 (O_949,N_14734,N_14370);
nor UO_950 (O_950,N_14967,N_14671);
nor UO_951 (O_951,N_14985,N_14511);
nand UO_952 (O_952,N_14511,N_14200);
nor UO_953 (O_953,N_14012,N_14296);
or UO_954 (O_954,N_14153,N_14863);
and UO_955 (O_955,N_14814,N_14322);
and UO_956 (O_956,N_14744,N_14055);
or UO_957 (O_957,N_14429,N_14884);
and UO_958 (O_958,N_14730,N_14911);
xor UO_959 (O_959,N_14419,N_14206);
and UO_960 (O_960,N_14032,N_14293);
or UO_961 (O_961,N_14956,N_14468);
xnor UO_962 (O_962,N_14095,N_14848);
nor UO_963 (O_963,N_14623,N_14763);
or UO_964 (O_964,N_14854,N_14218);
nand UO_965 (O_965,N_14074,N_14589);
xnor UO_966 (O_966,N_14856,N_14445);
and UO_967 (O_967,N_14474,N_14271);
xnor UO_968 (O_968,N_14437,N_14406);
or UO_969 (O_969,N_14714,N_14020);
xnor UO_970 (O_970,N_14148,N_14241);
and UO_971 (O_971,N_14078,N_14724);
or UO_972 (O_972,N_14937,N_14236);
nor UO_973 (O_973,N_14608,N_14573);
or UO_974 (O_974,N_14935,N_14900);
or UO_975 (O_975,N_14913,N_14654);
nand UO_976 (O_976,N_14085,N_14322);
or UO_977 (O_977,N_14778,N_14538);
xor UO_978 (O_978,N_14047,N_14524);
nand UO_979 (O_979,N_14569,N_14379);
and UO_980 (O_980,N_14660,N_14050);
or UO_981 (O_981,N_14432,N_14092);
xor UO_982 (O_982,N_14393,N_14265);
nand UO_983 (O_983,N_14646,N_14285);
nor UO_984 (O_984,N_14398,N_14098);
xor UO_985 (O_985,N_14566,N_14535);
and UO_986 (O_986,N_14889,N_14725);
and UO_987 (O_987,N_14991,N_14724);
xnor UO_988 (O_988,N_14550,N_14176);
and UO_989 (O_989,N_14185,N_14187);
and UO_990 (O_990,N_14488,N_14967);
nand UO_991 (O_991,N_14356,N_14608);
and UO_992 (O_992,N_14634,N_14379);
nand UO_993 (O_993,N_14738,N_14191);
nand UO_994 (O_994,N_14493,N_14722);
nand UO_995 (O_995,N_14795,N_14959);
nor UO_996 (O_996,N_14274,N_14411);
nor UO_997 (O_997,N_14962,N_14718);
or UO_998 (O_998,N_14450,N_14967);
or UO_999 (O_999,N_14541,N_14388);
nor UO_1000 (O_1000,N_14312,N_14744);
nand UO_1001 (O_1001,N_14564,N_14611);
xor UO_1002 (O_1002,N_14638,N_14272);
and UO_1003 (O_1003,N_14604,N_14419);
or UO_1004 (O_1004,N_14069,N_14948);
xnor UO_1005 (O_1005,N_14147,N_14572);
nor UO_1006 (O_1006,N_14038,N_14840);
nor UO_1007 (O_1007,N_14015,N_14960);
or UO_1008 (O_1008,N_14095,N_14523);
nor UO_1009 (O_1009,N_14528,N_14487);
xor UO_1010 (O_1010,N_14525,N_14126);
or UO_1011 (O_1011,N_14862,N_14711);
xor UO_1012 (O_1012,N_14368,N_14102);
nor UO_1013 (O_1013,N_14917,N_14964);
nand UO_1014 (O_1014,N_14249,N_14004);
and UO_1015 (O_1015,N_14238,N_14301);
and UO_1016 (O_1016,N_14565,N_14093);
nand UO_1017 (O_1017,N_14329,N_14159);
nor UO_1018 (O_1018,N_14047,N_14544);
and UO_1019 (O_1019,N_14422,N_14903);
xor UO_1020 (O_1020,N_14833,N_14391);
nor UO_1021 (O_1021,N_14363,N_14768);
and UO_1022 (O_1022,N_14157,N_14135);
nor UO_1023 (O_1023,N_14523,N_14375);
or UO_1024 (O_1024,N_14131,N_14088);
nor UO_1025 (O_1025,N_14892,N_14739);
and UO_1026 (O_1026,N_14790,N_14414);
or UO_1027 (O_1027,N_14571,N_14675);
xor UO_1028 (O_1028,N_14586,N_14483);
xor UO_1029 (O_1029,N_14786,N_14679);
or UO_1030 (O_1030,N_14645,N_14520);
and UO_1031 (O_1031,N_14209,N_14222);
xor UO_1032 (O_1032,N_14180,N_14205);
nand UO_1033 (O_1033,N_14813,N_14810);
and UO_1034 (O_1034,N_14957,N_14501);
nand UO_1035 (O_1035,N_14278,N_14925);
or UO_1036 (O_1036,N_14959,N_14308);
nor UO_1037 (O_1037,N_14950,N_14074);
and UO_1038 (O_1038,N_14412,N_14619);
or UO_1039 (O_1039,N_14458,N_14143);
xor UO_1040 (O_1040,N_14182,N_14492);
xnor UO_1041 (O_1041,N_14887,N_14434);
nand UO_1042 (O_1042,N_14938,N_14488);
or UO_1043 (O_1043,N_14476,N_14274);
or UO_1044 (O_1044,N_14433,N_14064);
or UO_1045 (O_1045,N_14217,N_14668);
xnor UO_1046 (O_1046,N_14035,N_14610);
nand UO_1047 (O_1047,N_14972,N_14076);
nand UO_1048 (O_1048,N_14167,N_14501);
xnor UO_1049 (O_1049,N_14043,N_14166);
or UO_1050 (O_1050,N_14693,N_14945);
nor UO_1051 (O_1051,N_14584,N_14268);
nor UO_1052 (O_1052,N_14952,N_14446);
and UO_1053 (O_1053,N_14102,N_14159);
nand UO_1054 (O_1054,N_14355,N_14675);
nor UO_1055 (O_1055,N_14780,N_14470);
nand UO_1056 (O_1056,N_14908,N_14279);
nand UO_1057 (O_1057,N_14808,N_14673);
nor UO_1058 (O_1058,N_14142,N_14863);
nand UO_1059 (O_1059,N_14227,N_14079);
or UO_1060 (O_1060,N_14389,N_14478);
nor UO_1061 (O_1061,N_14830,N_14630);
nand UO_1062 (O_1062,N_14312,N_14532);
and UO_1063 (O_1063,N_14726,N_14925);
nand UO_1064 (O_1064,N_14873,N_14168);
nand UO_1065 (O_1065,N_14425,N_14303);
nor UO_1066 (O_1066,N_14541,N_14194);
nand UO_1067 (O_1067,N_14160,N_14940);
xor UO_1068 (O_1068,N_14676,N_14751);
nand UO_1069 (O_1069,N_14151,N_14649);
or UO_1070 (O_1070,N_14427,N_14887);
and UO_1071 (O_1071,N_14855,N_14164);
nor UO_1072 (O_1072,N_14980,N_14401);
nor UO_1073 (O_1073,N_14408,N_14643);
nand UO_1074 (O_1074,N_14899,N_14245);
nand UO_1075 (O_1075,N_14724,N_14344);
and UO_1076 (O_1076,N_14172,N_14800);
nand UO_1077 (O_1077,N_14978,N_14779);
nor UO_1078 (O_1078,N_14025,N_14872);
and UO_1079 (O_1079,N_14283,N_14868);
nor UO_1080 (O_1080,N_14769,N_14953);
or UO_1081 (O_1081,N_14125,N_14732);
xnor UO_1082 (O_1082,N_14976,N_14954);
and UO_1083 (O_1083,N_14348,N_14922);
xor UO_1084 (O_1084,N_14435,N_14776);
xor UO_1085 (O_1085,N_14618,N_14336);
nor UO_1086 (O_1086,N_14483,N_14609);
and UO_1087 (O_1087,N_14436,N_14607);
or UO_1088 (O_1088,N_14343,N_14071);
nor UO_1089 (O_1089,N_14478,N_14617);
xnor UO_1090 (O_1090,N_14599,N_14196);
xnor UO_1091 (O_1091,N_14198,N_14887);
nor UO_1092 (O_1092,N_14980,N_14038);
nor UO_1093 (O_1093,N_14244,N_14150);
xnor UO_1094 (O_1094,N_14357,N_14970);
and UO_1095 (O_1095,N_14872,N_14019);
and UO_1096 (O_1096,N_14962,N_14088);
nor UO_1097 (O_1097,N_14246,N_14711);
nand UO_1098 (O_1098,N_14638,N_14795);
or UO_1099 (O_1099,N_14852,N_14774);
nand UO_1100 (O_1100,N_14291,N_14197);
xnor UO_1101 (O_1101,N_14561,N_14391);
or UO_1102 (O_1102,N_14508,N_14429);
or UO_1103 (O_1103,N_14427,N_14745);
xor UO_1104 (O_1104,N_14569,N_14511);
and UO_1105 (O_1105,N_14047,N_14697);
nand UO_1106 (O_1106,N_14767,N_14915);
nand UO_1107 (O_1107,N_14094,N_14905);
and UO_1108 (O_1108,N_14217,N_14889);
nor UO_1109 (O_1109,N_14993,N_14154);
or UO_1110 (O_1110,N_14694,N_14237);
nor UO_1111 (O_1111,N_14281,N_14603);
and UO_1112 (O_1112,N_14426,N_14018);
and UO_1113 (O_1113,N_14350,N_14090);
xnor UO_1114 (O_1114,N_14041,N_14548);
or UO_1115 (O_1115,N_14111,N_14405);
or UO_1116 (O_1116,N_14439,N_14451);
nor UO_1117 (O_1117,N_14603,N_14556);
and UO_1118 (O_1118,N_14113,N_14366);
nand UO_1119 (O_1119,N_14605,N_14010);
nand UO_1120 (O_1120,N_14690,N_14584);
xnor UO_1121 (O_1121,N_14999,N_14266);
or UO_1122 (O_1122,N_14915,N_14588);
xor UO_1123 (O_1123,N_14349,N_14199);
nor UO_1124 (O_1124,N_14900,N_14572);
nor UO_1125 (O_1125,N_14453,N_14677);
or UO_1126 (O_1126,N_14542,N_14528);
nor UO_1127 (O_1127,N_14838,N_14591);
nand UO_1128 (O_1128,N_14926,N_14277);
nor UO_1129 (O_1129,N_14389,N_14929);
and UO_1130 (O_1130,N_14630,N_14925);
nor UO_1131 (O_1131,N_14838,N_14806);
xor UO_1132 (O_1132,N_14757,N_14217);
nand UO_1133 (O_1133,N_14088,N_14670);
nand UO_1134 (O_1134,N_14251,N_14660);
xor UO_1135 (O_1135,N_14853,N_14220);
nor UO_1136 (O_1136,N_14361,N_14352);
nand UO_1137 (O_1137,N_14565,N_14097);
or UO_1138 (O_1138,N_14702,N_14034);
xor UO_1139 (O_1139,N_14033,N_14133);
nand UO_1140 (O_1140,N_14480,N_14761);
xnor UO_1141 (O_1141,N_14568,N_14747);
xnor UO_1142 (O_1142,N_14272,N_14831);
nor UO_1143 (O_1143,N_14681,N_14661);
and UO_1144 (O_1144,N_14914,N_14467);
and UO_1145 (O_1145,N_14956,N_14711);
nor UO_1146 (O_1146,N_14646,N_14219);
and UO_1147 (O_1147,N_14269,N_14734);
and UO_1148 (O_1148,N_14016,N_14694);
nand UO_1149 (O_1149,N_14370,N_14419);
xor UO_1150 (O_1150,N_14083,N_14135);
xnor UO_1151 (O_1151,N_14878,N_14251);
xnor UO_1152 (O_1152,N_14966,N_14954);
nand UO_1153 (O_1153,N_14368,N_14570);
nand UO_1154 (O_1154,N_14004,N_14984);
nand UO_1155 (O_1155,N_14112,N_14636);
xnor UO_1156 (O_1156,N_14589,N_14154);
and UO_1157 (O_1157,N_14530,N_14145);
and UO_1158 (O_1158,N_14516,N_14419);
and UO_1159 (O_1159,N_14232,N_14730);
nand UO_1160 (O_1160,N_14474,N_14084);
or UO_1161 (O_1161,N_14213,N_14032);
and UO_1162 (O_1162,N_14943,N_14517);
nand UO_1163 (O_1163,N_14044,N_14547);
xnor UO_1164 (O_1164,N_14281,N_14192);
and UO_1165 (O_1165,N_14078,N_14615);
xor UO_1166 (O_1166,N_14002,N_14856);
nor UO_1167 (O_1167,N_14120,N_14943);
or UO_1168 (O_1168,N_14523,N_14218);
and UO_1169 (O_1169,N_14010,N_14475);
nor UO_1170 (O_1170,N_14654,N_14540);
xnor UO_1171 (O_1171,N_14246,N_14129);
nand UO_1172 (O_1172,N_14455,N_14452);
nand UO_1173 (O_1173,N_14500,N_14865);
and UO_1174 (O_1174,N_14413,N_14774);
and UO_1175 (O_1175,N_14547,N_14792);
nand UO_1176 (O_1176,N_14924,N_14672);
or UO_1177 (O_1177,N_14245,N_14592);
and UO_1178 (O_1178,N_14735,N_14164);
xnor UO_1179 (O_1179,N_14315,N_14419);
nor UO_1180 (O_1180,N_14723,N_14948);
and UO_1181 (O_1181,N_14405,N_14662);
and UO_1182 (O_1182,N_14901,N_14306);
xor UO_1183 (O_1183,N_14155,N_14781);
nor UO_1184 (O_1184,N_14358,N_14176);
xor UO_1185 (O_1185,N_14112,N_14673);
xnor UO_1186 (O_1186,N_14312,N_14491);
nor UO_1187 (O_1187,N_14888,N_14445);
and UO_1188 (O_1188,N_14706,N_14997);
xnor UO_1189 (O_1189,N_14158,N_14356);
nor UO_1190 (O_1190,N_14762,N_14698);
xor UO_1191 (O_1191,N_14554,N_14560);
nand UO_1192 (O_1192,N_14441,N_14897);
or UO_1193 (O_1193,N_14701,N_14566);
or UO_1194 (O_1194,N_14005,N_14932);
or UO_1195 (O_1195,N_14905,N_14703);
nand UO_1196 (O_1196,N_14884,N_14256);
and UO_1197 (O_1197,N_14537,N_14943);
nand UO_1198 (O_1198,N_14093,N_14460);
nand UO_1199 (O_1199,N_14321,N_14057);
xnor UO_1200 (O_1200,N_14654,N_14455);
and UO_1201 (O_1201,N_14769,N_14492);
xor UO_1202 (O_1202,N_14581,N_14084);
xnor UO_1203 (O_1203,N_14850,N_14778);
nor UO_1204 (O_1204,N_14301,N_14433);
nor UO_1205 (O_1205,N_14686,N_14123);
nand UO_1206 (O_1206,N_14145,N_14852);
and UO_1207 (O_1207,N_14089,N_14845);
nand UO_1208 (O_1208,N_14659,N_14593);
nor UO_1209 (O_1209,N_14618,N_14278);
and UO_1210 (O_1210,N_14667,N_14973);
or UO_1211 (O_1211,N_14030,N_14907);
or UO_1212 (O_1212,N_14830,N_14590);
or UO_1213 (O_1213,N_14860,N_14612);
nand UO_1214 (O_1214,N_14558,N_14454);
nor UO_1215 (O_1215,N_14041,N_14699);
nor UO_1216 (O_1216,N_14823,N_14141);
xnor UO_1217 (O_1217,N_14596,N_14305);
nor UO_1218 (O_1218,N_14456,N_14226);
nor UO_1219 (O_1219,N_14110,N_14458);
and UO_1220 (O_1220,N_14272,N_14182);
or UO_1221 (O_1221,N_14628,N_14428);
or UO_1222 (O_1222,N_14893,N_14131);
nand UO_1223 (O_1223,N_14670,N_14772);
nor UO_1224 (O_1224,N_14288,N_14967);
xor UO_1225 (O_1225,N_14436,N_14434);
or UO_1226 (O_1226,N_14942,N_14361);
nand UO_1227 (O_1227,N_14663,N_14904);
nor UO_1228 (O_1228,N_14371,N_14414);
or UO_1229 (O_1229,N_14035,N_14573);
xnor UO_1230 (O_1230,N_14396,N_14700);
xor UO_1231 (O_1231,N_14841,N_14754);
nand UO_1232 (O_1232,N_14911,N_14077);
and UO_1233 (O_1233,N_14394,N_14732);
or UO_1234 (O_1234,N_14445,N_14211);
and UO_1235 (O_1235,N_14357,N_14360);
or UO_1236 (O_1236,N_14932,N_14888);
or UO_1237 (O_1237,N_14501,N_14880);
and UO_1238 (O_1238,N_14103,N_14085);
xor UO_1239 (O_1239,N_14092,N_14520);
nand UO_1240 (O_1240,N_14921,N_14982);
and UO_1241 (O_1241,N_14939,N_14266);
and UO_1242 (O_1242,N_14401,N_14679);
nor UO_1243 (O_1243,N_14418,N_14692);
and UO_1244 (O_1244,N_14899,N_14131);
and UO_1245 (O_1245,N_14121,N_14061);
nand UO_1246 (O_1246,N_14989,N_14967);
nor UO_1247 (O_1247,N_14960,N_14545);
and UO_1248 (O_1248,N_14069,N_14606);
nand UO_1249 (O_1249,N_14120,N_14333);
or UO_1250 (O_1250,N_14408,N_14965);
nor UO_1251 (O_1251,N_14173,N_14640);
nor UO_1252 (O_1252,N_14560,N_14824);
xnor UO_1253 (O_1253,N_14991,N_14285);
xor UO_1254 (O_1254,N_14466,N_14270);
xor UO_1255 (O_1255,N_14653,N_14704);
and UO_1256 (O_1256,N_14326,N_14963);
or UO_1257 (O_1257,N_14563,N_14841);
and UO_1258 (O_1258,N_14643,N_14748);
and UO_1259 (O_1259,N_14966,N_14417);
and UO_1260 (O_1260,N_14020,N_14584);
or UO_1261 (O_1261,N_14326,N_14962);
xor UO_1262 (O_1262,N_14420,N_14903);
nand UO_1263 (O_1263,N_14431,N_14703);
or UO_1264 (O_1264,N_14461,N_14489);
nor UO_1265 (O_1265,N_14475,N_14215);
and UO_1266 (O_1266,N_14784,N_14528);
nor UO_1267 (O_1267,N_14410,N_14711);
xnor UO_1268 (O_1268,N_14596,N_14030);
xor UO_1269 (O_1269,N_14404,N_14496);
nand UO_1270 (O_1270,N_14223,N_14648);
nand UO_1271 (O_1271,N_14278,N_14734);
xnor UO_1272 (O_1272,N_14194,N_14590);
or UO_1273 (O_1273,N_14240,N_14011);
and UO_1274 (O_1274,N_14581,N_14089);
nand UO_1275 (O_1275,N_14043,N_14021);
and UO_1276 (O_1276,N_14243,N_14315);
xnor UO_1277 (O_1277,N_14479,N_14037);
nand UO_1278 (O_1278,N_14082,N_14839);
xnor UO_1279 (O_1279,N_14814,N_14653);
and UO_1280 (O_1280,N_14843,N_14440);
or UO_1281 (O_1281,N_14654,N_14080);
or UO_1282 (O_1282,N_14008,N_14282);
xor UO_1283 (O_1283,N_14594,N_14533);
nor UO_1284 (O_1284,N_14370,N_14936);
nor UO_1285 (O_1285,N_14311,N_14016);
nand UO_1286 (O_1286,N_14682,N_14608);
nand UO_1287 (O_1287,N_14465,N_14876);
nor UO_1288 (O_1288,N_14219,N_14856);
xor UO_1289 (O_1289,N_14557,N_14404);
nor UO_1290 (O_1290,N_14688,N_14465);
nor UO_1291 (O_1291,N_14605,N_14243);
nor UO_1292 (O_1292,N_14011,N_14905);
nand UO_1293 (O_1293,N_14063,N_14897);
xor UO_1294 (O_1294,N_14190,N_14209);
nor UO_1295 (O_1295,N_14257,N_14648);
and UO_1296 (O_1296,N_14080,N_14489);
nor UO_1297 (O_1297,N_14697,N_14100);
nor UO_1298 (O_1298,N_14056,N_14395);
nor UO_1299 (O_1299,N_14251,N_14953);
xor UO_1300 (O_1300,N_14604,N_14486);
xor UO_1301 (O_1301,N_14752,N_14947);
xnor UO_1302 (O_1302,N_14547,N_14791);
xor UO_1303 (O_1303,N_14244,N_14596);
nand UO_1304 (O_1304,N_14469,N_14369);
and UO_1305 (O_1305,N_14920,N_14755);
and UO_1306 (O_1306,N_14118,N_14297);
nor UO_1307 (O_1307,N_14801,N_14724);
xnor UO_1308 (O_1308,N_14273,N_14555);
nand UO_1309 (O_1309,N_14654,N_14569);
or UO_1310 (O_1310,N_14708,N_14170);
xor UO_1311 (O_1311,N_14168,N_14610);
nand UO_1312 (O_1312,N_14732,N_14781);
and UO_1313 (O_1313,N_14362,N_14294);
or UO_1314 (O_1314,N_14325,N_14497);
nand UO_1315 (O_1315,N_14888,N_14069);
or UO_1316 (O_1316,N_14558,N_14402);
and UO_1317 (O_1317,N_14814,N_14043);
and UO_1318 (O_1318,N_14939,N_14223);
or UO_1319 (O_1319,N_14822,N_14535);
nand UO_1320 (O_1320,N_14659,N_14535);
nand UO_1321 (O_1321,N_14815,N_14148);
nand UO_1322 (O_1322,N_14948,N_14457);
or UO_1323 (O_1323,N_14540,N_14779);
nor UO_1324 (O_1324,N_14021,N_14414);
nand UO_1325 (O_1325,N_14135,N_14667);
nor UO_1326 (O_1326,N_14033,N_14189);
xor UO_1327 (O_1327,N_14351,N_14909);
xor UO_1328 (O_1328,N_14612,N_14888);
or UO_1329 (O_1329,N_14879,N_14915);
or UO_1330 (O_1330,N_14836,N_14589);
or UO_1331 (O_1331,N_14069,N_14262);
xor UO_1332 (O_1332,N_14219,N_14529);
xnor UO_1333 (O_1333,N_14397,N_14390);
nor UO_1334 (O_1334,N_14786,N_14418);
or UO_1335 (O_1335,N_14974,N_14949);
nor UO_1336 (O_1336,N_14039,N_14905);
nor UO_1337 (O_1337,N_14415,N_14114);
and UO_1338 (O_1338,N_14719,N_14636);
nand UO_1339 (O_1339,N_14712,N_14818);
nor UO_1340 (O_1340,N_14645,N_14138);
xnor UO_1341 (O_1341,N_14096,N_14065);
or UO_1342 (O_1342,N_14561,N_14901);
nand UO_1343 (O_1343,N_14844,N_14740);
and UO_1344 (O_1344,N_14344,N_14687);
and UO_1345 (O_1345,N_14098,N_14684);
nor UO_1346 (O_1346,N_14400,N_14011);
nand UO_1347 (O_1347,N_14689,N_14892);
nand UO_1348 (O_1348,N_14286,N_14351);
nand UO_1349 (O_1349,N_14092,N_14041);
xnor UO_1350 (O_1350,N_14354,N_14403);
xnor UO_1351 (O_1351,N_14860,N_14893);
nor UO_1352 (O_1352,N_14216,N_14014);
and UO_1353 (O_1353,N_14784,N_14952);
nand UO_1354 (O_1354,N_14055,N_14803);
or UO_1355 (O_1355,N_14625,N_14681);
nor UO_1356 (O_1356,N_14310,N_14881);
nor UO_1357 (O_1357,N_14408,N_14236);
xor UO_1358 (O_1358,N_14087,N_14939);
and UO_1359 (O_1359,N_14116,N_14568);
nand UO_1360 (O_1360,N_14074,N_14426);
nor UO_1361 (O_1361,N_14452,N_14054);
nor UO_1362 (O_1362,N_14745,N_14659);
xor UO_1363 (O_1363,N_14640,N_14454);
nor UO_1364 (O_1364,N_14670,N_14034);
and UO_1365 (O_1365,N_14547,N_14675);
nor UO_1366 (O_1366,N_14125,N_14439);
nor UO_1367 (O_1367,N_14711,N_14477);
or UO_1368 (O_1368,N_14079,N_14485);
xor UO_1369 (O_1369,N_14465,N_14512);
or UO_1370 (O_1370,N_14111,N_14620);
xor UO_1371 (O_1371,N_14497,N_14247);
xnor UO_1372 (O_1372,N_14273,N_14938);
and UO_1373 (O_1373,N_14672,N_14387);
and UO_1374 (O_1374,N_14346,N_14364);
and UO_1375 (O_1375,N_14360,N_14093);
nand UO_1376 (O_1376,N_14417,N_14550);
and UO_1377 (O_1377,N_14190,N_14356);
nand UO_1378 (O_1378,N_14116,N_14574);
and UO_1379 (O_1379,N_14179,N_14567);
nand UO_1380 (O_1380,N_14723,N_14350);
or UO_1381 (O_1381,N_14318,N_14958);
xnor UO_1382 (O_1382,N_14847,N_14773);
xor UO_1383 (O_1383,N_14009,N_14265);
xnor UO_1384 (O_1384,N_14510,N_14040);
nor UO_1385 (O_1385,N_14336,N_14997);
or UO_1386 (O_1386,N_14263,N_14131);
nand UO_1387 (O_1387,N_14183,N_14070);
xnor UO_1388 (O_1388,N_14384,N_14603);
and UO_1389 (O_1389,N_14885,N_14251);
or UO_1390 (O_1390,N_14091,N_14945);
or UO_1391 (O_1391,N_14066,N_14115);
xor UO_1392 (O_1392,N_14150,N_14890);
and UO_1393 (O_1393,N_14156,N_14328);
and UO_1394 (O_1394,N_14484,N_14695);
nand UO_1395 (O_1395,N_14470,N_14513);
nand UO_1396 (O_1396,N_14963,N_14930);
or UO_1397 (O_1397,N_14954,N_14513);
or UO_1398 (O_1398,N_14435,N_14237);
and UO_1399 (O_1399,N_14413,N_14251);
nand UO_1400 (O_1400,N_14504,N_14494);
nand UO_1401 (O_1401,N_14949,N_14164);
nand UO_1402 (O_1402,N_14639,N_14927);
and UO_1403 (O_1403,N_14568,N_14006);
nor UO_1404 (O_1404,N_14241,N_14721);
and UO_1405 (O_1405,N_14449,N_14160);
xor UO_1406 (O_1406,N_14097,N_14660);
xor UO_1407 (O_1407,N_14839,N_14764);
xnor UO_1408 (O_1408,N_14565,N_14288);
nand UO_1409 (O_1409,N_14362,N_14535);
nand UO_1410 (O_1410,N_14822,N_14108);
nor UO_1411 (O_1411,N_14301,N_14645);
xnor UO_1412 (O_1412,N_14447,N_14952);
nand UO_1413 (O_1413,N_14130,N_14013);
and UO_1414 (O_1414,N_14852,N_14970);
xor UO_1415 (O_1415,N_14675,N_14589);
xor UO_1416 (O_1416,N_14263,N_14084);
and UO_1417 (O_1417,N_14500,N_14796);
and UO_1418 (O_1418,N_14393,N_14754);
nand UO_1419 (O_1419,N_14881,N_14228);
xor UO_1420 (O_1420,N_14445,N_14179);
xnor UO_1421 (O_1421,N_14017,N_14423);
nand UO_1422 (O_1422,N_14205,N_14444);
xnor UO_1423 (O_1423,N_14266,N_14755);
or UO_1424 (O_1424,N_14366,N_14761);
nand UO_1425 (O_1425,N_14279,N_14498);
and UO_1426 (O_1426,N_14863,N_14316);
nand UO_1427 (O_1427,N_14080,N_14439);
and UO_1428 (O_1428,N_14765,N_14535);
or UO_1429 (O_1429,N_14902,N_14547);
and UO_1430 (O_1430,N_14196,N_14537);
nand UO_1431 (O_1431,N_14045,N_14729);
nand UO_1432 (O_1432,N_14801,N_14853);
xnor UO_1433 (O_1433,N_14875,N_14186);
nand UO_1434 (O_1434,N_14766,N_14941);
nor UO_1435 (O_1435,N_14772,N_14606);
xnor UO_1436 (O_1436,N_14921,N_14195);
nand UO_1437 (O_1437,N_14043,N_14016);
or UO_1438 (O_1438,N_14788,N_14252);
nand UO_1439 (O_1439,N_14489,N_14331);
xnor UO_1440 (O_1440,N_14638,N_14219);
and UO_1441 (O_1441,N_14032,N_14351);
nor UO_1442 (O_1442,N_14887,N_14248);
and UO_1443 (O_1443,N_14208,N_14489);
xor UO_1444 (O_1444,N_14373,N_14802);
nand UO_1445 (O_1445,N_14583,N_14837);
nand UO_1446 (O_1446,N_14586,N_14522);
and UO_1447 (O_1447,N_14916,N_14838);
nand UO_1448 (O_1448,N_14774,N_14202);
nor UO_1449 (O_1449,N_14540,N_14874);
or UO_1450 (O_1450,N_14044,N_14640);
and UO_1451 (O_1451,N_14627,N_14866);
or UO_1452 (O_1452,N_14080,N_14279);
and UO_1453 (O_1453,N_14086,N_14722);
and UO_1454 (O_1454,N_14565,N_14752);
or UO_1455 (O_1455,N_14738,N_14900);
nand UO_1456 (O_1456,N_14626,N_14910);
nor UO_1457 (O_1457,N_14096,N_14748);
and UO_1458 (O_1458,N_14826,N_14879);
or UO_1459 (O_1459,N_14632,N_14427);
nand UO_1460 (O_1460,N_14171,N_14567);
xor UO_1461 (O_1461,N_14289,N_14377);
or UO_1462 (O_1462,N_14813,N_14011);
xnor UO_1463 (O_1463,N_14574,N_14522);
nand UO_1464 (O_1464,N_14649,N_14075);
nand UO_1465 (O_1465,N_14280,N_14196);
nor UO_1466 (O_1466,N_14113,N_14716);
xnor UO_1467 (O_1467,N_14958,N_14289);
nor UO_1468 (O_1468,N_14063,N_14207);
and UO_1469 (O_1469,N_14264,N_14341);
nor UO_1470 (O_1470,N_14496,N_14060);
nor UO_1471 (O_1471,N_14074,N_14827);
and UO_1472 (O_1472,N_14457,N_14817);
and UO_1473 (O_1473,N_14857,N_14388);
and UO_1474 (O_1474,N_14421,N_14549);
or UO_1475 (O_1475,N_14843,N_14058);
nor UO_1476 (O_1476,N_14173,N_14527);
or UO_1477 (O_1477,N_14474,N_14403);
xnor UO_1478 (O_1478,N_14020,N_14185);
xor UO_1479 (O_1479,N_14319,N_14906);
nor UO_1480 (O_1480,N_14582,N_14603);
nand UO_1481 (O_1481,N_14547,N_14623);
or UO_1482 (O_1482,N_14516,N_14769);
or UO_1483 (O_1483,N_14942,N_14070);
or UO_1484 (O_1484,N_14165,N_14622);
nor UO_1485 (O_1485,N_14352,N_14279);
nor UO_1486 (O_1486,N_14525,N_14866);
nor UO_1487 (O_1487,N_14154,N_14106);
or UO_1488 (O_1488,N_14947,N_14954);
or UO_1489 (O_1489,N_14089,N_14578);
nor UO_1490 (O_1490,N_14059,N_14874);
xnor UO_1491 (O_1491,N_14743,N_14032);
nor UO_1492 (O_1492,N_14457,N_14326);
xor UO_1493 (O_1493,N_14017,N_14137);
nor UO_1494 (O_1494,N_14175,N_14081);
xnor UO_1495 (O_1495,N_14219,N_14841);
and UO_1496 (O_1496,N_14922,N_14783);
nand UO_1497 (O_1497,N_14872,N_14981);
xnor UO_1498 (O_1498,N_14088,N_14523);
nor UO_1499 (O_1499,N_14701,N_14963);
xnor UO_1500 (O_1500,N_14228,N_14243);
nor UO_1501 (O_1501,N_14053,N_14577);
nor UO_1502 (O_1502,N_14561,N_14769);
nand UO_1503 (O_1503,N_14798,N_14964);
nand UO_1504 (O_1504,N_14511,N_14267);
nor UO_1505 (O_1505,N_14834,N_14425);
nand UO_1506 (O_1506,N_14866,N_14228);
xor UO_1507 (O_1507,N_14594,N_14639);
and UO_1508 (O_1508,N_14630,N_14551);
xnor UO_1509 (O_1509,N_14073,N_14771);
and UO_1510 (O_1510,N_14753,N_14644);
or UO_1511 (O_1511,N_14265,N_14860);
or UO_1512 (O_1512,N_14331,N_14777);
nor UO_1513 (O_1513,N_14536,N_14232);
nor UO_1514 (O_1514,N_14873,N_14099);
xor UO_1515 (O_1515,N_14294,N_14016);
and UO_1516 (O_1516,N_14252,N_14036);
and UO_1517 (O_1517,N_14322,N_14384);
nand UO_1518 (O_1518,N_14495,N_14582);
nor UO_1519 (O_1519,N_14523,N_14719);
or UO_1520 (O_1520,N_14364,N_14474);
or UO_1521 (O_1521,N_14336,N_14125);
and UO_1522 (O_1522,N_14618,N_14662);
nor UO_1523 (O_1523,N_14429,N_14844);
xnor UO_1524 (O_1524,N_14019,N_14572);
and UO_1525 (O_1525,N_14370,N_14622);
nor UO_1526 (O_1526,N_14778,N_14129);
nand UO_1527 (O_1527,N_14413,N_14762);
xor UO_1528 (O_1528,N_14497,N_14722);
xor UO_1529 (O_1529,N_14566,N_14992);
nand UO_1530 (O_1530,N_14961,N_14119);
nor UO_1531 (O_1531,N_14391,N_14587);
xnor UO_1532 (O_1532,N_14785,N_14567);
xor UO_1533 (O_1533,N_14181,N_14802);
or UO_1534 (O_1534,N_14425,N_14913);
nand UO_1535 (O_1535,N_14383,N_14559);
or UO_1536 (O_1536,N_14133,N_14348);
nor UO_1537 (O_1537,N_14827,N_14913);
nor UO_1538 (O_1538,N_14348,N_14249);
nor UO_1539 (O_1539,N_14979,N_14244);
xnor UO_1540 (O_1540,N_14062,N_14436);
nand UO_1541 (O_1541,N_14266,N_14696);
nor UO_1542 (O_1542,N_14492,N_14764);
xor UO_1543 (O_1543,N_14497,N_14061);
or UO_1544 (O_1544,N_14395,N_14432);
and UO_1545 (O_1545,N_14191,N_14868);
or UO_1546 (O_1546,N_14396,N_14574);
nand UO_1547 (O_1547,N_14705,N_14672);
nand UO_1548 (O_1548,N_14787,N_14485);
nand UO_1549 (O_1549,N_14933,N_14619);
nor UO_1550 (O_1550,N_14882,N_14877);
nor UO_1551 (O_1551,N_14457,N_14177);
nand UO_1552 (O_1552,N_14059,N_14001);
nand UO_1553 (O_1553,N_14233,N_14517);
nor UO_1554 (O_1554,N_14903,N_14328);
nand UO_1555 (O_1555,N_14515,N_14899);
and UO_1556 (O_1556,N_14452,N_14703);
or UO_1557 (O_1557,N_14787,N_14258);
nand UO_1558 (O_1558,N_14047,N_14869);
xnor UO_1559 (O_1559,N_14588,N_14549);
or UO_1560 (O_1560,N_14789,N_14627);
or UO_1561 (O_1561,N_14197,N_14840);
and UO_1562 (O_1562,N_14466,N_14339);
or UO_1563 (O_1563,N_14901,N_14952);
nand UO_1564 (O_1564,N_14034,N_14127);
or UO_1565 (O_1565,N_14458,N_14062);
xor UO_1566 (O_1566,N_14746,N_14264);
nand UO_1567 (O_1567,N_14146,N_14822);
or UO_1568 (O_1568,N_14593,N_14778);
and UO_1569 (O_1569,N_14215,N_14573);
xor UO_1570 (O_1570,N_14782,N_14664);
xnor UO_1571 (O_1571,N_14031,N_14043);
nor UO_1572 (O_1572,N_14494,N_14732);
nand UO_1573 (O_1573,N_14451,N_14745);
nand UO_1574 (O_1574,N_14039,N_14434);
nand UO_1575 (O_1575,N_14778,N_14459);
or UO_1576 (O_1576,N_14125,N_14222);
xnor UO_1577 (O_1577,N_14252,N_14872);
nor UO_1578 (O_1578,N_14087,N_14342);
or UO_1579 (O_1579,N_14510,N_14525);
nor UO_1580 (O_1580,N_14202,N_14380);
and UO_1581 (O_1581,N_14847,N_14985);
nand UO_1582 (O_1582,N_14283,N_14949);
nor UO_1583 (O_1583,N_14438,N_14549);
nand UO_1584 (O_1584,N_14184,N_14353);
and UO_1585 (O_1585,N_14430,N_14575);
and UO_1586 (O_1586,N_14747,N_14580);
nand UO_1587 (O_1587,N_14946,N_14331);
nand UO_1588 (O_1588,N_14387,N_14893);
xor UO_1589 (O_1589,N_14297,N_14496);
and UO_1590 (O_1590,N_14586,N_14682);
xor UO_1591 (O_1591,N_14719,N_14815);
nor UO_1592 (O_1592,N_14552,N_14261);
nor UO_1593 (O_1593,N_14930,N_14840);
or UO_1594 (O_1594,N_14273,N_14034);
or UO_1595 (O_1595,N_14265,N_14089);
nor UO_1596 (O_1596,N_14352,N_14357);
nand UO_1597 (O_1597,N_14535,N_14484);
nor UO_1598 (O_1598,N_14539,N_14329);
xor UO_1599 (O_1599,N_14346,N_14278);
nand UO_1600 (O_1600,N_14515,N_14821);
nand UO_1601 (O_1601,N_14077,N_14378);
nand UO_1602 (O_1602,N_14842,N_14899);
nor UO_1603 (O_1603,N_14732,N_14489);
xnor UO_1604 (O_1604,N_14623,N_14863);
nor UO_1605 (O_1605,N_14682,N_14775);
or UO_1606 (O_1606,N_14787,N_14779);
or UO_1607 (O_1607,N_14675,N_14889);
xor UO_1608 (O_1608,N_14750,N_14404);
and UO_1609 (O_1609,N_14433,N_14808);
nand UO_1610 (O_1610,N_14285,N_14868);
and UO_1611 (O_1611,N_14320,N_14256);
xor UO_1612 (O_1612,N_14569,N_14000);
nor UO_1613 (O_1613,N_14705,N_14313);
xor UO_1614 (O_1614,N_14005,N_14834);
nand UO_1615 (O_1615,N_14284,N_14036);
xnor UO_1616 (O_1616,N_14203,N_14652);
and UO_1617 (O_1617,N_14560,N_14357);
nor UO_1618 (O_1618,N_14519,N_14645);
nand UO_1619 (O_1619,N_14005,N_14615);
and UO_1620 (O_1620,N_14382,N_14352);
or UO_1621 (O_1621,N_14944,N_14938);
and UO_1622 (O_1622,N_14226,N_14937);
and UO_1623 (O_1623,N_14203,N_14278);
or UO_1624 (O_1624,N_14309,N_14487);
nand UO_1625 (O_1625,N_14765,N_14367);
nand UO_1626 (O_1626,N_14045,N_14278);
or UO_1627 (O_1627,N_14905,N_14124);
and UO_1628 (O_1628,N_14532,N_14793);
nor UO_1629 (O_1629,N_14788,N_14569);
or UO_1630 (O_1630,N_14548,N_14329);
xor UO_1631 (O_1631,N_14997,N_14283);
nand UO_1632 (O_1632,N_14466,N_14235);
nand UO_1633 (O_1633,N_14486,N_14156);
nand UO_1634 (O_1634,N_14307,N_14522);
xor UO_1635 (O_1635,N_14240,N_14138);
xnor UO_1636 (O_1636,N_14021,N_14640);
and UO_1637 (O_1637,N_14422,N_14125);
xnor UO_1638 (O_1638,N_14571,N_14406);
nor UO_1639 (O_1639,N_14813,N_14354);
and UO_1640 (O_1640,N_14702,N_14232);
xor UO_1641 (O_1641,N_14883,N_14680);
nor UO_1642 (O_1642,N_14851,N_14023);
or UO_1643 (O_1643,N_14970,N_14060);
or UO_1644 (O_1644,N_14635,N_14513);
nor UO_1645 (O_1645,N_14514,N_14511);
xor UO_1646 (O_1646,N_14969,N_14883);
or UO_1647 (O_1647,N_14484,N_14566);
nor UO_1648 (O_1648,N_14774,N_14659);
xor UO_1649 (O_1649,N_14983,N_14893);
nand UO_1650 (O_1650,N_14362,N_14018);
nand UO_1651 (O_1651,N_14738,N_14167);
nor UO_1652 (O_1652,N_14685,N_14988);
xnor UO_1653 (O_1653,N_14344,N_14571);
or UO_1654 (O_1654,N_14061,N_14282);
nand UO_1655 (O_1655,N_14495,N_14722);
and UO_1656 (O_1656,N_14605,N_14357);
nand UO_1657 (O_1657,N_14207,N_14920);
and UO_1658 (O_1658,N_14643,N_14872);
xor UO_1659 (O_1659,N_14540,N_14295);
xnor UO_1660 (O_1660,N_14982,N_14160);
nand UO_1661 (O_1661,N_14386,N_14276);
nand UO_1662 (O_1662,N_14705,N_14494);
xor UO_1663 (O_1663,N_14317,N_14147);
nor UO_1664 (O_1664,N_14090,N_14391);
xnor UO_1665 (O_1665,N_14185,N_14749);
xor UO_1666 (O_1666,N_14418,N_14552);
and UO_1667 (O_1667,N_14321,N_14893);
xnor UO_1668 (O_1668,N_14600,N_14141);
nor UO_1669 (O_1669,N_14838,N_14647);
nor UO_1670 (O_1670,N_14170,N_14015);
or UO_1671 (O_1671,N_14786,N_14455);
and UO_1672 (O_1672,N_14248,N_14391);
and UO_1673 (O_1673,N_14587,N_14611);
xnor UO_1674 (O_1674,N_14986,N_14128);
xor UO_1675 (O_1675,N_14651,N_14088);
nor UO_1676 (O_1676,N_14012,N_14265);
and UO_1677 (O_1677,N_14306,N_14055);
nor UO_1678 (O_1678,N_14196,N_14259);
xnor UO_1679 (O_1679,N_14186,N_14979);
xnor UO_1680 (O_1680,N_14268,N_14031);
and UO_1681 (O_1681,N_14104,N_14192);
and UO_1682 (O_1682,N_14031,N_14795);
nor UO_1683 (O_1683,N_14095,N_14061);
nand UO_1684 (O_1684,N_14661,N_14397);
xor UO_1685 (O_1685,N_14251,N_14420);
or UO_1686 (O_1686,N_14082,N_14342);
nor UO_1687 (O_1687,N_14420,N_14679);
and UO_1688 (O_1688,N_14025,N_14521);
nand UO_1689 (O_1689,N_14886,N_14990);
xor UO_1690 (O_1690,N_14673,N_14381);
and UO_1691 (O_1691,N_14172,N_14868);
nor UO_1692 (O_1692,N_14046,N_14260);
xnor UO_1693 (O_1693,N_14850,N_14458);
xnor UO_1694 (O_1694,N_14368,N_14957);
or UO_1695 (O_1695,N_14267,N_14859);
or UO_1696 (O_1696,N_14877,N_14571);
nand UO_1697 (O_1697,N_14326,N_14664);
nor UO_1698 (O_1698,N_14783,N_14195);
nor UO_1699 (O_1699,N_14147,N_14171);
nand UO_1700 (O_1700,N_14579,N_14108);
and UO_1701 (O_1701,N_14818,N_14136);
and UO_1702 (O_1702,N_14988,N_14783);
and UO_1703 (O_1703,N_14534,N_14415);
xor UO_1704 (O_1704,N_14672,N_14182);
nor UO_1705 (O_1705,N_14914,N_14735);
or UO_1706 (O_1706,N_14210,N_14317);
or UO_1707 (O_1707,N_14802,N_14926);
xnor UO_1708 (O_1708,N_14452,N_14485);
and UO_1709 (O_1709,N_14332,N_14221);
or UO_1710 (O_1710,N_14776,N_14953);
and UO_1711 (O_1711,N_14142,N_14245);
xnor UO_1712 (O_1712,N_14328,N_14002);
nor UO_1713 (O_1713,N_14310,N_14792);
and UO_1714 (O_1714,N_14778,N_14269);
nor UO_1715 (O_1715,N_14782,N_14586);
xor UO_1716 (O_1716,N_14261,N_14541);
or UO_1717 (O_1717,N_14562,N_14718);
or UO_1718 (O_1718,N_14846,N_14124);
xor UO_1719 (O_1719,N_14576,N_14520);
nand UO_1720 (O_1720,N_14775,N_14406);
nand UO_1721 (O_1721,N_14952,N_14430);
nor UO_1722 (O_1722,N_14682,N_14626);
and UO_1723 (O_1723,N_14229,N_14467);
nand UO_1724 (O_1724,N_14021,N_14510);
xor UO_1725 (O_1725,N_14398,N_14772);
xor UO_1726 (O_1726,N_14912,N_14293);
and UO_1727 (O_1727,N_14165,N_14087);
and UO_1728 (O_1728,N_14902,N_14113);
or UO_1729 (O_1729,N_14209,N_14725);
and UO_1730 (O_1730,N_14396,N_14634);
nand UO_1731 (O_1731,N_14159,N_14336);
or UO_1732 (O_1732,N_14127,N_14151);
nor UO_1733 (O_1733,N_14561,N_14228);
nand UO_1734 (O_1734,N_14883,N_14627);
nor UO_1735 (O_1735,N_14802,N_14567);
nor UO_1736 (O_1736,N_14503,N_14897);
nand UO_1737 (O_1737,N_14369,N_14947);
nand UO_1738 (O_1738,N_14356,N_14015);
nand UO_1739 (O_1739,N_14362,N_14122);
xnor UO_1740 (O_1740,N_14205,N_14459);
or UO_1741 (O_1741,N_14392,N_14175);
and UO_1742 (O_1742,N_14677,N_14951);
and UO_1743 (O_1743,N_14396,N_14349);
xnor UO_1744 (O_1744,N_14496,N_14104);
nand UO_1745 (O_1745,N_14786,N_14058);
nand UO_1746 (O_1746,N_14628,N_14118);
xor UO_1747 (O_1747,N_14427,N_14416);
or UO_1748 (O_1748,N_14987,N_14727);
and UO_1749 (O_1749,N_14340,N_14842);
nand UO_1750 (O_1750,N_14684,N_14139);
or UO_1751 (O_1751,N_14023,N_14181);
or UO_1752 (O_1752,N_14904,N_14671);
nand UO_1753 (O_1753,N_14349,N_14347);
nand UO_1754 (O_1754,N_14284,N_14255);
nand UO_1755 (O_1755,N_14178,N_14094);
xnor UO_1756 (O_1756,N_14835,N_14065);
and UO_1757 (O_1757,N_14958,N_14167);
nor UO_1758 (O_1758,N_14656,N_14615);
xnor UO_1759 (O_1759,N_14738,N_14185);
nor UO_1760 (O_1760,N_14794,N_14901);
and UO_1761 (O_1761,N_14662,N_14569);
xnor UO_1762 (O_1762,N_14509,N_14979);
nand UO_1763 (O_1763,N_14488,N_14180);
nand UO_1764 (O_1764,N_14886,N_14995);
nor UO_1765 (O_1765,N_14516,N_14046);
nand UO_1766 (O_1766,N_14224,N_14034);
xor UO_1767 (O_1767,N_14397,N_14416);
xnor UO_1768 (O_1768,N_14005,N_14948);
and UO_1769 (O_1769,N_14935,N_14168);
or UO_1770 (O_1770,N_14244,N_14819);
or UO_1771 (O_1771,N_14235,N_14707);
xor UO_1772 (O_1772,N_14013,N_14084);
nand UO_1773 (O_1773,N_14679,N_14678);
nand UO_1774 (O_1774,N_14984,N_14447);
nand UO_1775 (O_1775,N_14842,N_14594);
xor UO_1776 (O_1776,N_14075,N_14301);
xor UO_1777 (O_1777,N_14359,N_14384);
and UO_1778 (O_1778,N_14582,N_14381);
or UO_1779 (O_1779,N_14783,N_14880);
nor UO_1780 (O_1780,N_14117,N_14990);
and UO_1781 (O_1781,N_14594,N_14839);
or UO_1782 (O_1782,N_14095,N_14186);
xor UO_1783 (O_1783,N_14801,N_14641);
or UO_1784 (O_1784,N_14205,N_14016);
nor UO_1785 (O_1785,N_14188,N_14548);
and UO_1786 (O_1786,N_14111,N_14134);
xor UO_1787 (O_1787,N_14265,N_14701);
or UO_1788 (O_1788,N_14294,N_14196);
nor UO_1789 (O_1789,N_14080,N_14402);
or UO_1790 (O_1790,N_14240,N_14453);
or UO_1791 (O_1791,N_14986,N_14150);
nand UO_1792 (O_1792,N_14328,N_14923);
and UO_1793 (O_1793,N_14697,N_14039);
xor UO_1794 (O_1794,N_14118,N_14697);
nor UO_1795 (O_1795,N_14474,N_14750);
nand UO_1796 (O_1796,N_14671,N_14606);
or UO_1797 (O_1797,N_14234,N_14892);
xnor UO_1798 (O_1798,N_14969,N_14656);
nand UO_1799 (O_1799,N_14788,N_14835);
and UO_1800 (O_1800,N_14445,N_14444);
and UO_1801 (O_1801,N_14798,N_14062);
nand UO_1802 (O_1802,N_14464,N_14378);
xor UO_1803 (O_1803,N_14373,N_14515);
or UO_1804 (O_1804,N_14113,N_14807);
and UO_1805 (O_1805,N_14567,N_14879);
and UO_1806 (O_1806,N_14831,N_14656);
and UO_1807 (O_1807,N_14925,N_14273);
xnor UO_1808 (O_1808,N_14668,N_14269);
and UO_1809 (O_1809,N_14082,N_14784);
nand UO_1810 (O_1810,N_14333,N_14354);
nand UO_1811 (O_1811,N_14432,N_14038);
nor UO_1812 (O_1812,N_14151,N_14890);
xor UO_1813 (O_1813,N_14134,N_14537);
xnor UO_1814 (O_1814,N_14616,N_14004);
nand UO_1815 (O_1815,N_14270,N_14266);
xor UO_1816 (O_1816,N_14829,N_14630);
xor UO_1817 (O_1817,N_14894,N_14354);
or UO_1818 (O_1818,N_14086,N_14941);
or UO_1819 (O_1819,N_14208,N_14157);
or UO_1820 (O_1820,N_14581,N_14442);
xnor UO_1821 (O_1821,N_14498,N_14817);
nor UO_1822 (O_1822,N_14824,N_14135);
nor UO_1823 (O_1823,N_14039,N_14734);
nand UO_1824 (O_1824,N_14378,N_14371);
and UO_1825 (O_1825,N_14307,N_14406);
or UO_1826 (O_1826,N_14045,N_14634);
or UO_1827 (O_1827,N_14560,N_14011);
or UO_1828 (O_1828,N_14566,N_14841);
nand UO_1829 (O_1829,N_14571,N_14659);
nor UO_1830 (O_1830,N_14279,N_14754);
or UO_1831 (O_1831,N_14838,N_14083);
nand UO_1832 (O_1832,N_14499,N_14801);
nor UO_1833 (O_1833,N_14955,N_14884);
nand UO_1834 (O_1834,N_14053,N_14809);
nand UO_1835 (O_1835,N_14157,N_14320);
nand UO_1836 (O_1836,N_14348,N_14469);
and UO_1837 (O_1837,N_14832,N_14514);
or UO_1838 (O_1838,N_14184,N_14802);
nand UO_1839 (O_1839,N_14911,N_14235);
nor UO_1840 (O_1840,N_14882,N_14434);
and UO_1841 (O_1841,N_14013,N_14775);
nor UO_1842 (O_1842,N_14554,N_14206);
nor UO_1843 (O_1843,N_14565,N_14687);
and UO_1844 (O_1844,N_14710,N_14844);
xor UO_1845 (O_1845,N_14750,N_14629);
xor UO_1846 (O_1846,N_14152,N_14322);
and UO_1847 (O_1847,N_14064,N_14773);
or UO_1848 (O_1848,N_14421,N_14139);
and UO_1849 (O_1849,N_14942,N_14943);
and UO_1850 (O_1850,N_14420,N_14022);
nor UO_1851 (O_1851,N_14118,N_14337);
nor UO_1852 (O_1852,N_14153,N_14072);
nand UO_1853 (O_1853,N_14703,N_14215);
nand UO_1854 (O_1854,N_14215,N_14870);
or UO_1855 (O_1855,N_14360,N_14862);
or UO_1856 (O_1856,N_14523,N_14354);
xnor UO_1857 (O_1857,N_14931,N_14526);
xnor UO_1858 (O_1858,N_14380,N_14348);
and UO_1859 (O_1859,N_14515,N_14922);
nand UO_1860 (O_1860,N_14122,N_14078);
or UO_1861 (O_1861,N_14935,N_14774);
xor UO_1862 (O_1862,N_14242,N_14126);
nand UO_1863 (O_1863,N_14952,N_14139);
or UO_1864 (O_1864,N_14811,N_14130);
nor UO_1865 (O_1865,N_14440,N_14165);
and UO_1866 (O_1866,N_14053,N_14980);
and UO_1867 (O_1867,N_14580,N_14366);
nand UO_1868 (O_1868,N_14425,N_14321);
or UO_1869 (O_1869,N_14243,N_14263);
or UO_1870 (O_1870,N_14724,N_14642);
nand UO_1871 (O_1871,N_14570,N_14411);
xor UO_1872 (O_1872,N_14909,N_14539);
or UO_1873 (O_1873,N_14021,N_14914);
nor UO_1874 (O_1874,N_14030,N_14382);
xnor UO_1875 (O_1875,N_14023,N_14559);
and UO_1876 (O_1876,N_14907,N_14680);
and UO_1877 (O_1877,N_14609,N_14242);
and UO_1878 (O_1878,N_14461,N_14915);
or UO_1879 (O_1879,N_14717,N_14229);
xnor UO_1880 (O_1880,N_14629,N_14180);
nand UO_1881 (O_1881,N_14470,N_14481);
and UO_1882 (O_1882,N_14996,N_14552);
xnor UO_1883 (O_1883,N_14382,N_14610);
xnor UO_1884 (O_1884,N_14531,N_14712);
or UO_1885 (O_1885,N_14277,N_14136);
and UO_1886 (O_1886,N_14093,N_14002);
or UO_1887 (O_1887,N_14286,N_14659);
xnor UO_1888 (O_1888,N_14063,N_14713);
nor UO_1889 (O_1889,N_14565,N_14974);
or UO_1890 (O_1890,N_14484,N_14977);
or UO_1891 (O_1891,N_14190,N_14327);
or UO_1892 (O_1892,N_14128,N_14030);
and UO_1893 (O_1893,N_14101,N_14036);
xnor UO_1894 (O_1894,N_14939,N_14633);
and UO_1895 (O_1895,N_14183,N_14243);
or UO_1896 (O_1896,N_14433,N_14191);
and UO_1897 (O_1897,N_14318,N_14733);
nand UO_1898 (O_1898,N_14620,N_14163);
nand UO_1899 (O_1899,N_14084,N_14362);
nor UO_1900 (O_1900,N_14918,N_14731);
xor UO_1901 (O_1901,N_14581,N_14736);
nand UO_1902 (O_1902,N_14944,N_14159);
xor UO_1903 (O_1903,N_14010,N_14113);
nor UO_1904 (O_1904,N_14784,N_14643);
and UO_1905 (O_1905,N_14108,N_14923);
nand UO_1906 (O_1906,N_14604,N_14628);
nor UO_1907 (O_1907,N_14091,N_14799);
nor UO_1908 (O_1908,N_14976,N_14582);
or UO_1909 (O_1909,N_14062,N_14673);
and UO_1910 (O_1910,N_14287,N_14998);
nand UO_1911 (O_1911,N_14615,N_14022);
nand UO_1912 (O_1912,N_14297,N_14108);
xnor UO_1913 (O_1913,N_14649,N_14228);
and UO_1914 (O_1914,N_14194,N_14736);
nor UO_1915 (O_1915,N_14290,N_14619);
and UO_1916 (O_1916,N_14607,N_14604);
nor UO_1917 (O_1917,N_14086,N_14408);
nand UO_1918 (O_1918,N_14384,N_14447);
and UO_1919 (O_1919,N_14315,N_14085);
or UO_1920 (O_1920,N_14061,N_14337);
nor UO_1921 (O_1921,N_14856,N_14524);
or UO_1922 (O_1922,N_14158,N_14790);
and UO_1923 (O_1923,N_14177,N_14951);
xnor UO_1924 (O_1924,N_14739,N_14628);
xor UO_1925 (O_1925,N_14130,N_14771);
nor UO_1926 (O_1926,N_14117,N_14562);
nor UO_1927 (O_1927,N_14768,N_14489);
nor UO_1928 (O_1928,N_14574,N_14278);
or UO_1929 (O_1929,N_14226,N_14815);
nand UO_1930 (O_1930,N_14935,N_14165);
nand UO_1931 (O_1931,N_14672,N_14700);
nor UO_1932 (O_1932,N_14435,N_14786);
and UO_1933 (O_1933,N_14316,N_14448);
or UO_1934 (O_1934,N_14857,N_14845);
nand UO_1935 (O_1935,N_14378,N_14140);
nand UO_1936 (O_1936,N_14509,N_14494);
xnor UO_1937 (O_1937,N_14003,N_14298);
xor UO_1938 (O_1938,N_14360,N_14602);
xnor UO_1939 (O_1939,N_14931,N_14085);
and UO_1940 (O_1940,N_14790,N_14952);
nor UO_1941 (O_1941,N_14858,N_14399);
or UO_1942 (O_1942,N_14563,N_14001);
xnor UO_1943 (O_1943,N_14875,N_14892);
xnor UO_1944 (O_1944,N_14723,N_14898);
and UO_1945 (O_1945,N_14849,N_14069);
or UO_1946 (O_1946,N_14219,N_14874);
and UO_1947 (O_1947,N_14735,N_14211);
nand UO_1948 (O_1948,N_14744,N_14125);
nor UO_1949 (O_1949,N_14140,N_14334);
nor UO_1950 (O_1950,N_14177,N_14468);
and UO_1951 (O_1951,N_14681,N_14735);
xor UO_1952 (O_1952,N_14678,N_14509);
nand UO_1953 (O_1953,N_14800,N_14599);
xor UO_1954 (O_1954,N_14760,N_14268);
or UO_1955 (O_1955,N_14054,N_14414);
or UO_1956 (O_1956,N_14933,N_14608);
or UO_1957 (O_1957,N_14517,N_14355);
nand UO_1958 (O_1958,N_14419,N_14030);
or UO_1959 (O_1959,N_14680,N_14338);
xnor UO_1960 (O_1960,N_14898,N_14651);
nor UO_1961 (O_1961,N_14421,N_14854);
xor UO_1962 (O_1962,N_14356,N_14969);
nor UO_1963 (O_1963,N_14390,N_14532);
nor UO_1964 (O_1964,N_14321,N_14148);
nor UO_1965 (O_1965,N_14468,N_14636);
and UO_1966 (O_1966,N_14947,N_14832);
nor UO_1967 (O_1967,N_14952,N_14504);
nand UO_1968 (O_1968,N_14516,N_14138);
xor UO_1969 (O_1969,N_14557,N_14230);
and UO_1970 (O_1970,N_14073,N_14907);
nand UO_1971 (O_1971,N_14293,N_14348);
or UO_1972 (O_1972,N_14850,N_14219);
xor UO_1973 (O_1973,N_14467,N_14225);
nand UO_1974 (O_1974,N_14572,N_14269);
and UO_1975 (O_1975,N_14979,N_14720);
nor UO_1976 (O_1976,N_14625,N_14064);
xor UO_1977 (O_1977,N_14247,N_14903);
and UO_1978 (O_1978,N_14604,N_14335);
or UO_1979 (O_1979,N_14563,N_14828);
nor UO_1980 (O_1980,N_14762,N_14775);
xnor UO_1981 (O_1981,N_14785,N_14105);
nor UO_1982 (O_1982,N_14045,N_14736);
nand UO_1983 (O_1983,N_14702,N_14513);
or UO_1984 (O_1984,N_14585,N_14258);
or UO_1985 (O_1985,N_14125,N_14803);
nor UO_1986 (O_1986,N_14673,N_14326);
nor UO_1987 (O_1987,N_14774,N_14082);
nor UO_1988 (O_1988,N_14898,N_14790);
and UO_1989 (O_1989,N_14991,N_14793);
or UO_1990 (O_1990,N_14598,N_14181);
or UO_1991 (O_1991,N_14100,N_14231);
xnor UO_1992 (O_1992,N_14766,N_14732);
nor UO_1993 (O_1993,N_14824,N_14704);
and UO_1994 (O_1994,N_14743,N_14582);
nor UO_1995 (O_1995,N_14962,N_14233);
and UO_1996 (O_1996,N_14317,N_14742);
or UO_1997 (O_1997,N_14310,N_14551);
or UO_1998 (O_1998,N_14717,N_14027);
xnor UO_1999 (O_1999,N_14973,N_14923);
endmodule