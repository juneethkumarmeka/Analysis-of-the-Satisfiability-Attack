module basic_1000_10000_1500_100_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_417,In_599);
nor U1 (N_1,In_57,In_37);
or U2 (N_2,In_825,In_921);
nor U3 (N_3,In_384,In_59);
nand U4 (N_4,In_873,In_756);
nand U5 (N_5,In_304,In_966);
xor U6 (N_6,In_475,In_908);
nor U7 (N_7,In_725,In_31);
xnor U8 (N_8,In_227,In_918);
xor U9 (N_9,In_977,In_915);
nor U10 (N_10,In_834,In_487);
nor U11 (N_11,In_865,In_525);
nand U12 (N_12,In_814,In_416);
nand U13 (N_13,In_269,In_617);
nand U14 (N_14,In_690,In_598);
and U15 (N_15,In_137,In_892);
and U16 (N_16,In_249,In_243);
nand U17 (N_17,In_512,In_491);
nor U18 (N_18,In_537,In_857);
or U19 (N_19,In_15,In_801);
and U20 (N_20,In_765,In_419);
nand U21 (N_21,In_202,In_608);
nand U22 (N_22,In_478,In_531);
and U23 (N_23,In_767,In_300);
nand U24 (N_24,In_647,In_997);
nand U25 (N_25,In_119,In_861);
xor U26 (N_26,In_118,In_917);
and U27 (N_27,In_46,In_664);
or U28 (N_28,In_792,In_841);
nor U29 (N_29,In_611,In_586);
or U30 (N_30,In_728,In_541);
nor U31 (N_31,In_935,In_649);
nor U32 (N_32,In_214,In_708);
nor U33 (N_33,In_9,In_99);
or U34 (N_34,In_499,In_235);
nor U35 (N_35,In_442,In_833);
or U36 (N_36,In_200,In_631);
nand U37 (N_37,In_518,In_602);
nor U38 (N_38,In_674,In_652);
nand U39 (N_39,In_775,In_239);
or U40 (N_40,In_964,In_153);
nand U41 (N_41,In_629,In_845);
and U42 (N_42,In_558,In_69);
and U43 (N_43,In_48,In_712);
and U44 (N_44,In_275,In_511);
or U45 (N_45,In_687,In_314);
nor U46 (N_46,In_796,In_392);
nor U47 (N_47,In_658,In_711);
or U48 (N_48,In_783,In_643);
nor U49 (N_49,In_62,In_359);
and U50 (N_50,In_853,In_123);
xor U51 (N_51,In_571,In_36);
nor U52 (N_52,In_467,In_879);
nor U53 (N_53,In_484,In_578);
nor U54 (N_54,In_999,In_898);
or U55 (N_55,In_75,In_887);
or U56 (N_56,In_672,In_747);
and U57 (N_57,In_313,In_919);
nor U58 (N_58,In_221,In_950);
nand U59 (N_59,In_585,In_798);
nor U60 (N_60,In_899,In_931);
or U61 (N_61,In_544,In_210);
or U62 (N_62,In_581,In_78);
or U63 (N_63,In_398,In_191);
and U64 (N_64,In_576,In_922);
xnor U65 (N_65,In_949,In_545);
or U66 (N_66,In_588,In_688);
or U67 (N_67,In_878,In_969);
and U68 (N_68,In_670,In_987);
and U69 (N_69,In_691,In_567);
and U70 (N_70,In_379,In_973);
nand U71 (N_71,In_257,In_373);
xor U72 (N_72,In_109,In_583);
nand U73 (N_73,In_874,In_176);
or U74 (N_74,In_340,In_749);
and U75 (N_75,In_136,In_183);
nand U76 (N_76,In_569,In_284);
nor U77 (N_77,In_242,In_911);
nand U78 (N_78,In_315,In_897);
and U79 (N_79,In_293,In_718);
xnor U80 (N_80,In_420,In_816);
nor U81 (N_81,In_286,In_152);
or U82 (N_82,In_77,In_208);
nor U83 (N_83,In_944,In_372);
nand U84 (N_84,In_240,In_199);
and U85 (N_85,In_422,In_470);
or U86 (N_86,In_822,In_258);
or U87 (N_87,In_233,In_364);
nor U88 (N_88,In_490,In_761);
or U89 (N_89,In_157,In_510);
xnor U90 (N_90,In_913,In_509);
or U91 (N_91,In_529,In_967);
and U92 (N_92,In_716,In_958);
nand U93 (N_93,In_939,In_843);
nor U94 (N_94,In_645,In_669);
and U95 (N_95,In_14,In_338);
and U96 (N_96,In_523,In_804);
nor U97 (N_97,In_87,In_805);
nand U98 (N_98,In_7,In_410);
nor U99 (N_99,In_836,In_425);
or U100 (N_100,In_391,N_45);
nor U101 (N_101,In_353,In_327);
nand U102 (N_102,In_3,In_395);
nand U103 (N_103,In_970,In_633);
nand U104 (N_104,In_319,In_22);
nor U105 (N_105,In_554,In_591);
nand U106 (N_106,In_984,In_341);
and U107 (N_107,In_682,In_339);
nand U108 (N_108,In_53,N_78);
nand U109 (N_109,In_308,In_961);
nand U110 (N_110,In_130,In_55);
nor U111 (N_111,In_486,In_234);
or U112 (N_112,In_182,In_306);
nor U113 (N_113,In_852,In_637);
nand U114 (N_114,In_705,In_122);
and U115 (N_115,In_360,In_132);
and U116 (N_116,In_330,In_255);
nand U117 (N_117,In_642,In_365);
nor U118 (N_118,In_847,In_806);
nor U119 (N_119,In_24,In_505);
xnor U120 (N_120,In_253,In_877);
nand U121 (N_121,In_582,N_29);
nor U122 (N_122,In_292,In_981);
xnor U123 (N_123,In_495,In_216);
nand U124 (N_124,In_536,In_423);
or U125 (N_125,In_324,In_433);
or U126 (N_126,In_809,In_923);
or U127 (N_127,In_476,In_207);
or U128 (N_128,N_37,In_303);
nand U129 (N_129,In_826,In_477);
nor U130 (N_130,In_768,N_51);
nor U131 (N_131,In_107,In_177);
or U132 (N_132,In_851,In_100);
nor U133 (N_133,In_550,In_80);
and U134 (N_134,In_979,In_355);
nand U135 (N_135,In_776,In_600);
or U136 (N_136,In_203,In_400);
and U137 (N_137,In_817,In_219);
xnor U138 (N_138,In_677,In_882);
or U139 (N_139,In_12,N_86);
or U140 (N_140,In_829,In_368);
or U141 (N_141,In_875,In_19);
and U142 (N_142,In_13,In_524);
nand U143 (N_143,In_409,In_727);
or U144 (N_144,In_115,In_593);
and U145 (N_145,N_70,In_165);
nor U146 (N_146,In_223,In_555);
xnor U147 (N_147,In_318,In_18);
nand U148 (N_148,In_884,In_789);
nand U149 (N_149,In_66,In_974);
or U150 (N_150,In_68,In_194);
or U151 (N_151,In_256,In_634);
xor U152 (N_152,In_406,In_627);
xor U153 (N_153,In_613,N_49);
or U154 (N_154,In_127,In_685);
nor U155 (N_155,In_86,In_457);
or U156 (N_156,N_74,In_720);
or U157 (N_157,In_596,In_704);
nor U158 (N_158,In_237,In_0);
nor U159 (N_159,In_676,In_699);
nand U160 (N_160,In_232,In_247);
and U161 (N_161,In_197,In_595);
and U162 (N_162,In_660,In_111);
nor U163 (N_163,In_496,In_837);
or U164 (N_164,In_781,In_560);
xnor U165 (N_165,In_871,In_421);
nor U166 (N_166,In_213,In_782);
nor U167 (N_167,In_838,In_606);
or U168 (N_168,In_262,In_320);
or U169 (N_169,N_76,In_696);
and U170 (N_170,In_519,N_95);
nor U171 (N_171,In_626,In_515);
xor U172 (N_172,In_146,In_797);
and U173 (N_173,N_6,In_357);
xor U174 (N_174,In_920,In_787);
or U175 (N_175,In_793,In_4);
or U176 (N_176,N_71,In_35);
xnor U177 (N_177,In_501,In_85);
nor U178 (N_178,In_835,N_65);
nor U179 (N_179,In_312,In_568);
nor U180 (N_180,In_868,In_988);
and U181 (N_181,In_955,In_745);
or U182 (N_182,In_686,N_9);
nor U183 (N_183,In_962,In_252);
or U184 (N_184,In_51,In_26);
and U185 (N_185,In_448,In_196);
xor U186 (N_186,In_985,N_43);
nor U187 (N_187,In_678,In_800);
nor U188 (N_188,In_276,In_881);
nand U189 (N_189,In_362,In_790);
nor U190 (N_190,In_700,In_785);
nand U191 (N_191,N_16,In_251);
and U192 (N_192,In_231,In_818);
and U193 (N_193,In_497,In_823);
and U194 (N_194,In_810,In_311);
and U195 (N_195,In_807,In_367);
and U196 (N_196,In_722,In_415);
nand U197 (N_197,N_93,In_780);
nor U198 (N_198,In_166,N_34);
and U199 (N_199,In_883,In_366);
or U200 (N_200,N_157,In_862);
or U201 (N_201,In_748,In_492);
nand U202 (N_202,In_620,In_820);
and U203 (N_203,In_169,In_103);
xnor U204 (N_204,In_894,In_706);
nor U205 (N_205,In_819,In_996);
xnor U206 (N_206,In_474,In_993);
and U207 (N_207,In_155,N_189);
nor U208 (N_208,In_795,In_886);
nand U209 (N_209,In_436,In_336);
or U210 (N_210,In_186,In_942);
xor U211 (N_211,In_390,N_54);
xnor U212 (N_212,In_241,In_738);
nand U213 (N_213,In_580,In_23);
nor U214 (N_214,N_82,In_564);
and U215 (N_215,In_173,In_735);
and U216 (N_216,In_297,In_291);
nor U217 (N_217,In_383,In_855);
or U218 (N_218,N_15,In_799);
and U219 (N_219,In_743,In_171);
xor U220 (N_220,N_61,In_450);
and U221 (N_221,In_454,In_407);
or U222 (N_222,In_813,In_557);
nand U223 (N_223,In_552,In_498);
and U224 (N_224,In_105,In_959);
nand U225 (N_225,In_896,In_803);
and U226 (N_226,N_105,In_762);
or U227 (N_227,In_84,N_87);
xor U228 (N_228,N_136,In_666);
nand U229 (N_229,In_925,N_115);
nor U230 (N_230,In_134,In_278);
nand U231 (N_231,N_27,In_302);
nand U232 (N_232,N_118,In_47);
xnor U233 (N_233,In_615,In_158);
and U234 (N_234,In_370,In_547);
and U235 (N_235,In_697,In_609);
nand U236 (N_236,In_172,In_983);
nor U237 (N_237,In_244,In_363);
nor U238 (N_238,In_25,N_119);
and U239 (N_239,In_126,In_263);
or U240 (N_240,In_97,In_681);
nand U241 (N_241,In_565,In_140);
nor U242 (N_242,N_102,In_434);
nor U243 (N_243,N_146,In_72);
nor U244 (N_244,In_856,In_211);
xor U245 (N_245,In_926,In_755);
xor U246 (N_246,N_179,In_542);
nor U247 (N_247,N_110,In_880);
nor U248 (N_248,In_671,In_456);
or U249 (N_249,N_73,In_16);
xnor U250 (N_250,N_8,In_724);
nor U251 (N_251,N_84,In_27);
xor U252 (N_252,In_483,In_358);
and U253 (N_253,In_352,N_81);
or U254 (N_254,In_228,N_199);
xor U255 (N_255,In_522,N_97);
nand U256 (N_256,In_195,In_759);
xnor U257 (N_257,In_389,In_839);
nor U258 (N_258,N_25,In_689);
nor U259 (N_259,In_131,In_732);
nand U260 (N_260,In_774,In_701);
or U261 (N_261,In_890,In_288);
nand U262 (N_262,In_412,In_938);
nor U263 (N_263,In_551,In_205);
nand U264 (N_264,In_117,N_154);
or U265 (N_265,N_131,In_471);
or U266 (N_266,N_153,In_414);
and U267 (N_267,N_85,In_411);
nand U268 (N_268,In_936,N_94);
xor U269 (N_269,N_137,N_123);
nand U270 (N_270,In_342,N_163);
or U271 (N_271,In_181,In_50);
or U272 (N_272,N_69,In_968);
or U273 (N_273,N_18,In_264);
xor U274 (N_274,In_750,In_610);
or U275 (N_275,In_430,N_140);
or U276 (N_276,In_254,In_374);
or U277 (N_277,In_112,N_59);
and U278 (N_278,In_125,N_127);
or U279 (N_279,In_133,In_193);
and U280 (N_280,In_513,In_124);
nor U281 (N_281,N_135,In_659);
xnor U282 (N_282,N_33,N_196);
and U283 (N_283,In_95,In_636);
and U284 (N_284,In_106,In_891);
nor U285 (N_285,In_82,In_770);
nand U286 (N_286,In_371,In_488);
nor U287 (N_287,In_348,In_440);
or U288 (N_288,N_106,In_198);
and U289 (N_289,N_162,In_579);
nor U290 (N_290,N_28,In_914);
or U291 (N_291,In_628,N_22);
nor U292 (N_292,In_404,N_174);
xor U293 (N_293,In_549,In_904);
nand U294 (N_294,In_94,In_533);
or U295 (N_295,In_698,In_451);
xor U296 (N_296,N_96,In_64);
xor U297 (N_297,In_587,In_405);
nor U298 (N_298,In_945,N_31);
and U299 (N_299,In_566,In_889);
nor U300 (N_300,In_535,In_88);
nand U301 (N_301,In_577,In_885);
xor U302 (N_302,In_184,In_361);
and U303 (N_303,In_58,In_559);
and U304 (N_304,In_432,In_40);
nor U305 (N_305,In_449,In_329);
nor U306 (N_306,N_42,In_39);
and U307 (N_307,In_464,N_58);
or U308 (N_308,In_438,In_89);
nor U309 (N_309,In_399,N_231);
nor U310 (N_310,In_54,N_241);
xnor U311 (N_311,In_299,N_291);
or U312 (N_312,N_60,N_248);
nand U313 (N_313,N_276,In_614);
nand U314 (N_314,In_872,In_731);
xor U315 (N_315,In_744,In_347);
nor U316 (N_316,In_849,N_19);
and U317 (N_317,In_334,In_447);
xor U318 (N_318,In_840,In_466);
and U319 (N_319,In_733,In_639);
nor U320 (N_320,In_846,In_343);
xnor U321 (N_321,N_206,N_120);
nor U322 (N_322,In_651,In_250);
and U323 (N_323,In_713,N_177);
nor U324 (N_324,In_656,In_493);
nor U325 (N_325,In_382,N_138);
and U326 (N_326,In_638,In_38);
or U327 (N_327,In_842,In_139);
and U328 (N_328,N_68,In_957);
nor U329 (N_329,In_532,In_956);
and U330 (N_330,In_683,N_5);
nand U331 (N_331,In_589,In_52);
nor U332 (N_332,N_281,In_236);
xor U333 (N_333,In_472,N_11);
or U334 (N_334,In_325,N_250);
or U335 (N_335,In_933,In_468);
nor U336 (N_336,In_70,In_93);
nor U337 (N_337,N_10,N_262);
nand U338 (N_338,N_139,N_21);
nand U339 (N_339,N_183,In_60);
and U340 (N_340,In_574,In_943);
and U341 (N_341,N_12,In_396);
xor U342 (N_342,In_646,N_224);
and U343 (N_343,In_502,N_173);
or U344 (N_344,N_284,In_741);
or U345 (N_345,In_90,In_632);
nor U346 (N_346,In_215,N_292);
xnor U347 (N_347,N_235,In_61);
nor U348 (N_348,In_96,N_133);
or U349 (N_349,In_429,In_91);
nand U350 (N_350,In_684,In_204);
nor U351 (N_351,In_528,In_590);
xnor U352 (N_352,N_212,In_317);
xnor U353 (N_353,In_65,N_229);
and U354 (N_354,N_62,In_42);
nand U355 (N_355,N_155,In_693);
nor U356 (N_356,In_831,In_378);
and U357 (N_357,N_186,In_665);
nor U358 (N_358,In_272,N_14);
nor U359 (N_359,In_323,N_52);
or U360 (N_360,N_207,In_791);
or U361 (N_361,In_516,N_265);
xnor U362 (N_362,In_248,In_960);
nand U363 (N_363,In_773,N_104);
or U364 (N_364,N_79,In_481);
and U365 (N_365,In_946,In_377);
or U366 (N_366,N_147,In_346);
nand U367 (N_367,In_539,N_228);
nand U368 (N_368,N_285,In_266);
or U369 (N_369,In_900,N_158);
and U370 (N_370,In_444,In_159);
and U371 (N_371,In_2,In_730);
xor U372 (N_372,In_556,In_296);
nand U373 (N_373,In_888,N_144);
or U374 (N_374,In_952,In_723);
nor U375 (N_375,N_90,N_63);
or U376 (N_376,N_113,N_190);
and U377 (N_377,In_408,In_463);
nor U378 (N_378,N_116,N_176);
nand U379 (N_379,N_252,In_503);
or U380 (N_380,In_459,In_349);
nand U381 (N_381,In_514,In_764);
and U382 (N_382,In_827,N_129);
nand U383 (N_383,In_28,In_703);
and U384 (N_384,N_187,In_648);
or U385 (N_385,In_980,In_494);
nor U386 (N_386,In_369,In_56);
or U387 (N_387,In_641,In_772);
xor U388 (N_388,In_116,In_212);
and U389 (N_389,In_44,In_734);
xnor U390 (N_390,N_299,In_445);
and U391 (N_391,N_171,In_867);
or U392 (N_392,In_848,In_859);
nor U393 (N_393,In_114,In_736);
or U394 (N_394,N_277,In_356);
and U395 (N_395,In_605,In_473);
or U396 (N_396,In_937,N_184);
xnor U397 (N_397,N_208,In_758);
or U398 (N_398,In_462,In_508);
or U399 (N_399,N_67,N_209);
or U400 (N_400,N_294,N_261);
nor U401 (N_401,N_121,N_275);
nand U402 (N_402,In_129,N_237);
and U403 (N_403,In_766,In_553);
or U404 (N_404,In_187,N_216);
nand U405 (N_405,N_46,In_778);
nor U406 (N_406,N_395,In_635);
or U407 (N_407,In_209,In_850);
or U408 (N_408,In_351,N_333);
or U409 (N_409,In_273,In_828);
nor U410 (N_410,In_680,In_621);
nor U411 (N_411,In_930,In_261);
xnor U412 (N_412,In_655,In_443);
or U413 (N_413,N_364,In_121);
or U414 (N_414,N_278,In_333);
or U415 (N_415,In_802,N_343);
nor U416 (N_416,In_461,N_166);
or U417 (N_417,N_373,N_101);
or U418 (N_418,N_357,In_188);
xnor U419 (N_419,In_866,N_204);
nor U420 (N_420,N_256,In_387);
or U421 (N_421,In_189,N_341);
xnor U422 (N_422,N_236,In_623);
nor U423 (N_423,In_268,In_175);
and U424 (N_424,N_347,N_376);
nor U425 (N_425,N_198,N_254);
or U426 (N_426,N_111,In_386);
nor U427 (N_427,In_245,N_214);
nor U428 (N_428,N_362,In_141);
nor U429 (N_429,N_234,N_23);
or U430 (N_430,N_48,N_342);
or U431 (N_431,In_328,In_954);
nand U432 (N_432,N_322,N_338);
or U433 (N_433,In_815,In_540);
and U434 (N_434,In_603,N_103);
xnor U435 (N_435,In_707,In_285);
nor U436 (N_436,In_179,N_142);
nor U437 (N_437,In_870,N_319);
and U438 (N_438,In_739,In_517);
nor U439 (N_439,In_538,In_79);
and U440 (N_440,In_570,N_356);
or U441 (N_441,N_100,In_201);
or U442 (N_442,N_371,In_489);
nor U443 (N_443,N_353,In_283);
and U444 (N_444,N_389,N_287);
or U445 (N_445,In_910,In_8);
nand U446 (N_446,In_113,In_821);
nand U447 (N_447,In_281,N_107);
nand U448 (N_448,In_34,In_108);
nand U449 (N_449,In_563,In_963);
nand U450 (N_450,N_50,In_128);
and U451 (N_451,N_351,N_75);
xnor U452 (N_452,N_239,In_893);
or U453 (N_453,N_367,N_361);
and U454 (N_454,N_197,In_76);
or U455 (N_455,In_662,N_167);
and U456 (N_456,N_246,In_757);
nor U457 (N_457,In_479,N_225);
nand U458 (N_458,In_667,In_630);
nor U459 (N_459,In_418,In_310);
and U460 (N_460,N_26,N_263);
nor U461 (N_461,N_38,N_374);
nor U462 (N_462,In_616,N_245);
or U463 (N_463,N_308,In_354);
or U464 (N_464,In_534,N_217);
or U465 (N_465,In_863,In_994);
or U466 (N_466,In_344,N_243);
and U467 (N_467,In_143,In_927);
or U468 (N_468,N_365,N_390);
or U469 (N_469,N_298,N_230);
xnor U470 (N_470,In_709,In_206);
xnor U471 (N_471,N_80,In_694);
nand U472 (N_472,N_39,In_480);
nand U473 (N_473,In_279,N_349);
nand U474 (N_474,In_982,N_314);
nand U475 (N_475,In_226,In_185);
nor U476 (N_476,In_504,N_297);
or U477 (N_477,N_112,In_71);
nor U478 (N_478,In_572,N_91);
nor U479 (N_479,N_344,N_172);
nor U480 (N_480,In_45,In_975);
xnor U481 (N_481,In_224,In_661);
and U482 (N_482,In_751,N_378);
nor U483 (N_483,In_719,N_363);
and U484 (N_484,In_452,In_168);
or U485 (N_485,In_104,N_92);
and U486 (N_486,N_145,N_273);
or U487 (N_487,In_895,In_811);
nand U488 (N_488,In_527,N_170);
nor U489 (N_489,In_149,In_294);
nor U490 (N_490,In_679,In_729);
nand U491 (N_491,N_150,In_287);
or U492 (N_492,In_238,In_692);
or U493 (N_493,N_255,N_310);
or U494 (N_494,N_337,N_384);
xor U495 (N_495,N_394,In_506);
nand U496 (N_496,N_117,In_520);
or U497 (N_497,In_932,N_244);
nor U498 (N_498,In_947,N_181);
or U499 (N_499,N_320,In_458);
nand U500 (N_500,N_331,N_178);
nor U501 (N_501,N_413,N_431);
xor U502 (N_502,N_288,N_488);
nor U503 (N_503,In_469,N_290);
nor U504 (N_504,N_98,In_844);
or U505 (N_505,N_192,N_175);
or U506 (N_506,N_414,In_32);
and U507 (N_507,N_156,N_1);
nand U508 (N_508,N_412,In_657);
and U509 (N_509,N_203,In_161);
and U510 (N_510,In_190,In_485);
nor U511 (N_511,N_56,N_211);
xnor U512 (N_512,In_67,In_151);
or U513 (N_513,In_695,In_167);
or U514 (N_514,N_114,In_869);
nand U515 (N_515,N_202,In_543);
xnor U516 (N_516,N_169,N_370);
nand U517 (N_517,In_332,In_426);
and U518 (N_518,N_326,In_854);
or U519 (N_519,N_180,In_902);
nor U520 (N_520,In_49,N_403);
nand U521 (N_521,N_435,In_500);
nand U522 (N_522,N_77,N_423);
or U523 (N_523,N_340,In_101);
xor U524 (N_524,N_7,In_280);
or U525 (N_525,N_327,N_477);
nand U526 (N_526,N_332,N_482);
nand U527 (N_527,In_217,N_474);
nor U528 (N_528,N_484,In_380);
nand U529 (N_529,N_383,N_450);
xor U530 (N_530,N_160,In_309);
nor U531 (N_531,In_305,N_311);
or U532 (N_532,In_1,N_44);
xnor U533 (N_533,N_433,In_909);
and U534 (N_534,N_329,In_375);
nand U535 (N_535,N_257,In_530);
nand U536 (N_536,In_948,In_858);
nand U537 (N_537,In_110,N_258);
or U538 (N_538,N_397,In_170);
and U539 (N_539,In_431,N_195);
nand U540 (N_540,N_312,In_246);
xnor U541 (N_541,In_991,N_432);
and U542 (N_542,N_53,In_573);
nor U543 (N_543,N_41,N_483);
and U544 (N_544,N_24,N_440);
xor U545 (N_545,In_784,N_321);
or U546 (N_546,In_618,In_376);
and U547 (N_547,In_742,N_148);
or U548 (N_548,In_976,In_345);
nand U549 (N_549,N_289,N_221);
nor U550 (N_550,In_941,In_597);
or U551 (N_551,N_463,N_99);
nor U552 (N_552,N_305,In_710);
nor U553 (N_553,N_478,In_120);
nand U554 (N_554,In_607,In_928);
and U555 (N_555,N_200,N_443);
or U556 (N_556,N_191,N_266);
and U557 (N_557,In_274,In_714);
or U558 (N_558,In_277,In_575);
nand U559 (N_559,In_331,N_421);
nor U560 (N_560,N_411,In_322);
nor U561 (N_561,In_737,In_41);
or U562 (N_562,In_546,In_63);
xor U563 (N_563,N_451,In_978);
and U564 (N_564,N_232,N_132);
nand U565 (N_565,In_990,In_92);
nand U566 (N_566,In_995,N_419);
and U567 (N_567,In_282,N_122);
nand U568 (N_568,In_465,N_323);
nand U569 (N_569,In_316,In_427);
and U570 (N_570,N_410,In_220);
nor U571 (N_571,In_754,N_466);
nor U572 (N_572,In_526,In_594);
nor U573 (N_573,N_487,N_369);
and U574 (N_574,N_447,N_489);
or U575 (N_575,N_213,In_752);
nor U576 (N_576,N_247,N_406);
and U577 (N_577,N_300,N_380);
nand U578 (N_578,In_164,N_220);
nand U579 (N_579,N_108,N_3);
and U580 (N_580,In_779,N_40);
nor U581 (N_581,In_321,N_89);
and U582 (N_582,In_622,N_194);
and U583 (N_583,In_763,N_475);
or U584 (N_584,In_860,In_397);
and U585 (N_585,N_126,N_182);
and U586 (N_586,N_476,N_377);
xnor U587 (N_587,In_903,N_32);
and U588 (N_588,In_147,In_43);
xor U589 (N_589,In_788,In_403);
or U590 (N_590,In_740,N_185);
and U591 (N_591,In_148,N_30);
nor U592 (N_592,In_653,In_394);
or U593 (N_593,N_215,N_164);
and U594 (N_594,N_469,In_289);
nor U595 (N_595,N_223,In_640);
nand U596 (N_596,N_497,N_405);
nand U597 (N_597,In_326,N_251);
nand U598 (N_598,N_442,N_339);
and U599 (N_599,N_457,N_490);
nand U600 (N_600,N_424,N_159);
nand U601 (N_601,In_906,In_265);
nand U602 (N_602,In_953,N_417);
and U603 (N_603,In_222,N_149);
nand U604 (N_604,In_259,N_388);
and U605 (N_605,N_72,N_165);
xnor U606 (N_606,N_492,In_548);
xnor U607 (N_607,In_604,N_521);
xor U608 (N_608,In_726,N_309);
and U609 (N_609,N_566,N_188);
or U610 (N_610,N_592,N_471);
or U611 (N_611,In_808,In_350);
nand U612 (N_612,In_663,In_402);
nor U613 (N_613,In_428,N_533);
or U614 (N_614,In_11,N_372);
nand U615 (N_615,N_346,N_218);
nand U616 (N_616,In_753,In_5);
or U617 (N_617,N_560,In_295);
and U618 (N_618,In_624,N_539);
or U619 (N_619,N_532,N_461);
or U620 (N_620,N_13,N_379);
or U621 (N_621,In_298,In_437);
and U622 (N_622,N_523,N_502);
or U623 (N_623,In_385,N_124);
nor U624 (N_624,N_400,N_448);
nor U625 (N_625,In_156,In_992);
or U626 (N_626,N_472,In_715);
or U627 (N_627,N_561,In_584);
or U628 (N_628,N_535,N_399);
nor U629 (N_629,N_35,In_145);
nand U630 (N_630,In_507,N_582);
and U631 (N_631,In_794,In_812);
nor U632 (N_632,N_425,In_21);
xor U633 (N_633,N_280,N_317);
nor U634 (N_634,N_529,N_408);
nor U635 (N_635,N_480,N_355);
xor U636 (N_636,N_473,N_452);
nand U637 (N_637,N_467,N_485);
nand U638 (N_638,N_438,N_501);
and U639 (N_639,N_543,In_832);
nor U640 (N_640,N_563,In_455);
and U641 (N_641,In_225,N_496);
nor U642 (N_642,N_345,N_143);
nor U643 (N_643,N_546,N_161);
or U644 (N_644,N_510,N_227);
nand U645 (N_645,N_503,N_446);
nor U646 (N_646,N_286,N_306);
and U647 (N_647,N_307,N_325);
nor U648 (N_648,N_520,In_644);
nor U649 (N_649,N_499,In_924);
and U650 (N_650,N_386,N_303);
and U651 (N_651,In_435,N_576);
nor U652 (N_652,N_454,N_552);
or U653 (N_653,In_138,N_282);
or U654 (N_654,N_570,N_494);
nand U655 (N_655,N_549,N_575);
xnor U656 (N_656,In_73,N_456);
and U657 (N_657,In_98,In_381);
and U658 (N_658,N_437,In_989);
and U659 (N_659,In_769,N_427);
nor U660 (N_660,N_572,In_601);
nor U661 (N_661,N_550,N_420);
nand U662 (N_662,N_283,N_522);
nand U663 (N_663,N_268,In_393);
nand U664 (N_664,N_556,In_102);
xnor U665 (N_665,N_577,N_459);
or U666 (N_666,In_592,N_589);
xor U667 (N_667,In_824,In_230);
nand U668 (N_668,In_986,N_436);
or U669 (N_669,N_493,In_150);
xnor U670 (N_670,N_530,N_519);
xnor U671 (N_671,N_313,N_555);
nand U672 (N_672,N_587,In_401);
nand U673 (N_673,N_449,In_951);
or U674 (N_674,N_381,In_30);
and U675 (N_675,In_998,N_542);
or U676 (N_676,N_409,N_269);
nor U677 (N_677,N_64,In_760);
xnor U678 (N_678,N_508,N_36);
nand U679 (N_679,N_415,N_260);
nor U680 (N_680,In_625,In_307);
nand U681 (N_681,In_17,N_210);
nor U682 (N_682,N_596,N_55);
and U683 (N_683,In_290,In_174);
xor U684 (N_684,In_675,N_525);
and U685 (N_685,In_650,N_516);
nor U686 (N_686,N_441,N_350);
xnor U687 (N_687,N_554,N_528);
or U688 (N_688,N_540,In_721);
xnor U689 (N_689,In_482,N_481);
and U690 (N_690,N_4,N_491);
or U691 (N_691,N_242,N_272);
or U692 (N_692,N_418,In_912);
or U693 (N_693,In_424,N_498);
or U694 (N_694,In_441,In_335);
nand U695 (N_695,N_548,N_201);
nor U696 (N_696,N_428,N_295);
xor U697 (N_697,N_302,In_20);
or U698 (N_698,N_512,In_271);
or U699 (N_699,N_393,N_293);
nand U700 (N_700,N_640,In_180);
and U701 (N_701,N_628,N_430);
nor U702 (N_702,N_564,N_652);
or U703 (N_703,N_88,N_657);
and U704 (N_704,N_604,N_109);
and U705 (N_705,N_270,N_661);
or U706 (N_706,N_680,N_407);
or U707 (N_707,N_274,N_382);
nor U708 (N_708,N_581,N_264);
xnor U709 (N_709,In_154,N_271);
and U710 (N_710,N_699,N_694);
nor U711 (N_711,N_392,N_585);
nor U712 (N_712,N_462,N_591);
or U713 (N_713,N_324,N_655);
and U714 (N_714,N_368,N_651);
nor U715 (N_715,N_599,In_135);
and U716 (N_716,N_559,N_396);
nand U717 (N_717,N_676,N_553);
and U718 (N_718,N_562,N_193);
or U719 (N_719,N_617,N_697);
nand U720 (N_720,N_656,In_267);
nand U721 (N_721,N_219,N_679);
or U722 (N_722,N_568,N_622);
xor U723 (N_723,N_578,N_690);
and U724 (N_724,N_504,N_439);
nor U725 (N_725,N_375,In_702);
nor U726 (N_726,In_301,N_515);
nor U727 (N_727,N_593,N_642);
nor U728 (N_728,In_771,In_446);
or U729 (N_729,N_465,N_238);
xnor U730 (N_730,In_144,N_434);
nand U731 (N_731,In_905,In_521);
nor U732 (N_732,In_163,N_253);
and U733 (N_733,N_444,N_233);
nor U734 (N_734,N_621,N_460);
nand U735 (N_735,N_531,N_641);
nor U736 (N_736,N_620,N_598);
and U737 (N_737,N_387,N_17);
or U738 (N_738,N_588,In_460);
or U739 (N_739,N_315,N_416);
or U740 (N_740,N_486,N_625);
and U741 (N_741,In_916,N_663);
nand U742 (N_742,N_334,N_354);
nand U743 (N_743,N_573,N_569);
and U744 (N_744,N_0,N_685);
nor U745 (N_745,In_830,N_316);
and U746 (N_746,N_616,N_259);
xnor U747 (N_747,N_675,N_691);
and U748 (N_748,N_20,N_506);
or U749 (N_749,N_335,N_630);
and U750 (N_750,N_571,N_686);
and U751 (N_751,N_688,In_777);
and U752 (N_752,N_662,N_429);
nand U753 (N_753,N_594,N_629);
and U754 (N_754,N_611,N_301);
or U755 (N_755,N_360,In_746);
and U756 (N_756,N_518,N_385);
or U757 (N_757,N_401,N_619);
and U758 (N_758,N_304,N_606);
nor U759 (N_759,N_682,In_717);
xnor U760 (N_760,In_439,In_229);
nand U761 (N_761,N_668,N_398);
nor U762 (N_762,N_318,In_965);
nand U763 (N_763,In_10,N_692);
nor U764 (N_764,N_647,N_66);
nor U765 (N_765,N_479,N_128);
xor U766 (N_766,N_57,In_971);
nand U767 (N_767,N_673,N_538);
nor U768 (N_768,N_565,N_267);
nand U769 (N_769,In_160,N_404);
nor U770 (N_770,N_511,N_495);
nand U771 (N_771,N_627,In_218);
and U772 (N_772,N_600,N_152);
nand U773 (N_773,In_33,In_934);
and U774 (N_774,N_83,In_83);
xor U775 (N_775,N_659,In_562);
nand U776 (N_776,N_633,N_687);
and U777 (N_777,N_130,N_650);
or U778 (N_778,N_358,N_537);
nor U779 (N_779,N_649,N_500);
nand U780 (N_780,N_222,N_453);
nor U781 (N_781,N_683,N_644);
or U782 (N_782,N_47,N_597);
or U783 (N_783,In_786,N_534);
and U784 (N_784,N_671,N_674);
nand U785 (N_785,N_125,N_464);
and U786 (N_786,N_551,N_653);
and U787 (N_787,N_141,N_359);
or U788 (N_788,N_517,In_142);
or U789 (N_789,In_972,N_2);
nand U790 (N_790,N_580,N_470);
nor U791 (N_791,N_590,In_619);
nand U792 (N_792,N_643,In_668);
nand U793 (N_793,N_669,N_296);
nor U794 (N_794,In_29,In_81);
nor U795 (N_795,N_426,N_605);
and U796 (N_796,N_696,In_74);
nand U797 (N_797,In_654,N_402);
and U798 (N_798,N_583,N_279);
or U799 (N_799,N_678,N_509);
nor U800 (N_800,N_782,N_613);
and U801 (N_801,N_623,N_557);
nor U802 (N_802,N_706,N_787);
or U803 (N_803,N_710,N_741);
nor U804 (N_804,N_793,N_586);
or U805 (N_805,N_742,N_527);
nor U806 (N_806,N_739,In_876);
nand U807 (N_807,N_711,N_777);
nand U808 (N_808,N_788,N_601);
nand U809 (N_809,N_660,N_713);
nand U810 (N_810,N_794,N_541);
or U811 (N_811,N_746,N_749);
and U812 (N_812,N_615,N_752);
nor U813 (N_813,N_775,N_645);
xnor U814 (N_814,N_757,N_134);
and U815 (N_815,N_703,In_178);
or U816 (N_816,N_748,N_328);
and U817 (N_817,N_689,In_270);
or U818 (N_818,In_388,N_781);
or U819 (N_819,N_765,N_545);
or U820 (N_820,N_603,N_779);
nand U821 (N_821,N_731,N_718);
nand U822 (N_822,N_733,In_337);
nand U823 (N_823,N_524,N_772);
nor U824 (N_824,N_579,N_745);
or U825 (N_825,N_709,N_634);
nor U826 (N_826,N_744,N_612);
and U827 (N_827,N_799,N_730);
and U828 (N_828,N_736,N_584);
nor U829 (N_829,N_768,N_769);
nor U830 (N_830,N_762,N_226);
xor U831 (N_831,N_786,N_670);
nand U832 (N_832,N_778,N_755);
or U833 (N_833,N_507,N_205);
nand U834 (N_834,N_614,N_737);
nor U835 (N_835,N_505,In_162);
or U836 (N_836,N_151,N_352);
and U837 (N_837,N_797,N_658);
xor U838 (N_838,N_608,N_526);
nor U839 (N_839,N_723,N_547);
or U840 (N_840,N_672,N_240);
or U841 (N_841,N_455,N_609);
nand U842 (N_842,N_727,In_929);
nand U843 (N_843,N_664,N_761);
or U844 (N_844,N_695,N_758);
xor U845 (N_845,N_714,In_413);
and U846 (N_846,N_789,N_725);
nand U847 (N_847,In_6,N_631);
and U848 (N_848,N_795,N_767);
xnor U849 (N_849,N_638,N_602);
nor U850 (N_850,N_722,In_940);
and U851 (N_851,N_784,N_780);
nand U852 (N_852,N_665,N_763);
nor U853 (N_853,N_756,N_618);
nor U854 (N_854,N_708,N_636);
nor U855 (N_855,N_783,In_561);
nor U856 (N_856,N_724,N_760);
and U857 (N_857,In_612,N_468);
nand U858 (N_858,N_719,N_698);
xnor U859 (N_859,N_707,N_677);
or U860 (N_860,N_750,N_798);
nand U861 (N_861,N_422,N_595);
nand U862 (N_862,N_716,N_705);
nor U863 (N_863,N_624,N_646);
or U864 (N_864,In_453,N_536);
nand U865 (N_865,N_544,N_770);
and U866 (N_866,In_192,N_348);
and U867 (N_867,N_759,N_693);
or U868 (N_868,N_771,N_632);
nor U869 (N_869,N_702,N_754);
nand U870 (N_870,N_610,N_704);
nand U871 (N_871,N_785,N_567);
nor U872 (N_872,N_445,N_667);
and U873 (N_873,N_735,In_260);
or U874 (N_874,N_639,N_607);
xnor U875 (N_875,N_330,N_684);
nor U876 (N_876,N_654,N_513);
nand U877 (N_877,N_729,N_720);
nand U878 (N_878,N_336,N_791);
and U879 (N_879,N_635,N_681);
nor U880 (N_880,N_701,N_514);
or U881 (N_881,In_901,N_743);
and U882 (N_882,N_458,In_673);
or U883 (N_883,N_712,N_666);
nand U884 (N_884,N_715,N_700);
and U885 (N_885,N_792,N_776);
xnor U886 (N_886,N_773,N_747);
and U887 (N_887,N_391,N_558);
xor U888 (N_888,N_574,N_753);
nor U889 (N_889,N_648,N_249);
nor U890 (N_890,N_366,N_717);
nor U891 (N_891,N_732,N_796);
and U892 (N_892,N_721,N_751);
nor U893 (N_893,N_637,N_726);
and U894 (N_894,N_766,In_907);
nand U895 (N_895,N_738,N_764);
or U896 (N_896,N_626,N_790);
or U897 (N_897,N_740,N_774);
and U898 (N_898,N_734,N_168);
nor U899 (N_899,In_864,N_728);
nor U900 (N_900,N_865,N_885);
xor U901 (N_901,N_820,N_812);
nand U902 (N_902,N_821,N_841);
or U903 (N_903,N_894,N_818);
and U904 (N_904,N_853,N_825);
or U905 (N_905,N_870,N_886);
and U906 (N_906,N_801,N_891);
nor U907 (N_907,N_855,N_840);
nand U908 (N_908,N_842,N_830);
and U909 (N_909,N_811,N_857);
or U910 (N_910,N_806,N_882);
nand U911 (N_911,N_858,N_892);
and U912 (N_912,N_815,N_829);
or U913 (N_913,N_863,N_844);
and U914 (N_914,N_896,N_826);
nor U915 (N_915,N_890,N_834);
or U916 (N_916,N_872,N_819);
or U917 (N_917,N_805,N_835);
nand U918 (N_918,N_846,N_897);
nand U919 (N_919,N_809,N_836);
xor U920 (N_920,N_850,N_889);
and U921 (N_921,N_864,N_831);
nand U922 (N_922,N_851,N_800);
nand U923 (N_923,N_848,N_843);
or U924 (N_924,N_832,N_883);
or U925 (N_925,N_827,N_875);
nor U926 (N_926,N_899,N_822);
and U927 (N_927,N_849,N_868);
or U928 (N_928,N_880,N_845);
and U929 (N_929,N_871,N_808);
nor U930 (N_930,N_881,N_833);
nand U931 (N_931,N_803,N_823);
and U932 (N_932,N_895,N_867);
nor U933 (N_933,N_802,N_866);
xnor U934 (N_934,N_876,N_877);
nor U935 (N_935,N_807,N_887);
and U936 (N_936,N_837,N_856);
nor U937 (N_937,N_884,N_893);
nand U938 (N_938,N_860,N_859);
nand U939 (N_939,N_898,N_879);
xnor U940 (N_940,N_852,N_869);
and U941 (N_941,N_862,N_828);
nor U942 (N_942,N_847,N_816);
xnor U943 (N_943,N_817,N_814);
nor U944 (N_944,N_804,N_824);
xnor U945 (N_945,N_838,N_813);
nand U946 (N_946,N_839,N_873);
nor U947 (N_947,N_874,N_854);
and U948 (N_948,N_888,N_878);
xor U949 (N_949,N_861,N_810);
xor U950 (N_950,N_856,N_839);
nand U951 (N_951,N_860,N_879);
xor U952 (N_952,N_846,N_817);
nor U953 (N_953,N_888,N_851);
nor U954 (N_954,N_809,N_878);
nand U955 (N_955,N_821,N_809);
xor U956 (N_956,N_863,N_899);
and U957 (N_957,N_868,N_850);
or U958 (N_958,N_894,N_811);
and U959 (N_959,N_863,N_894);
or U960 (N_960,N_826,N_872);
nand U961 (N_961,N_878,N_894);
nand U962 (N_962,N_837,N_812);
nor U963 (N_963,N_808,N_881);
and U964 (N_964,N_813,N_884);
and U965 (N_965,N_841,N_850);
nor U966 (N_966,N_808,N_883);
nand U967 (N_967,N_827,N_864);
or U968 (N_968,N_895,N_893);
and U969 (N_969,N_800,N_841);
or U970 (N_970,N_898,N_855);
nand U971 (N_971,N_823,N_843);
and U972 (N_972,N_871,N_879);
and U973 (N_973,N_847,N_835);
xnor U974 (N_974,N_819,N_840);
or U975 (N_975,N_805,N_859);
or U976 (N_976,N_865,N_835);
or U977 (N_977,N_830,N_871);
and U978 (N_978,N_891,N_874);
and U979 (N_979,N_835,N_867);
nand U980 (N_980,N_800,N_852);
and U981 (N_981,N_817,N_873);
nand U982 (N_982,N_837,N_888);
nand U983 (N_983,N_870,N_856);
or U984 (N_984,N_827,N_851);
and U985 (N_985,N_891,N_892);
nand U986 (N_986,N_891,N_864);
or U987 (N_987,N_829,N_855);
and U988 (N_988,N_840,N_843);
nor U989 (N_989,N_820,N_824);
nand U990 (N_990,N_807,N_896);
nor U991 (N_991,N_838,N_827);
nor U992 (N_992,N_861,N_889);
nand U993 (N_993,N_855,N_883);
and U994 (N_994,N_827,N_815);
or U995 (N_995,N_817,N_887);
nand U996 (N_996,N_802,N_829);
nor U997 (N_997,N_894,N_859);
nor U998 (N_998,N_835,N_862);
xnor U999 (N_999,N_820,N_894);
nand U1000 (N_1000,N_953,N_959);
or U1001 (N_1001,N_969,N_962);
nor U1002 (N_1002,N_997,N_927);
and U1003 (N_1003,N_972,N_910);
nor U1004 (N_1004,N_929,N_915);
nand U1005 (N_1005,N_983,N_943);
or U1006 (N_1006,N_996,N_973);
and U1007 (N_1007,N_919,N_950);
nand U1008 (N_1008,N_930,N_964);
nor U1009 (N_1009,N_914,N_986);
nor U1010 (N_1010,N_981,N_912);
or U1011 (N_1011,N_957,N_989);
nand U1012 (N_1012,N_988,N_935);
xor U1013 (N_1013,N_967,N_918);
nand U1014 (N_1014,N_960,N_991);
or U1015 (N_1015,N_965,N_951);
or U1016 (N_1016,N_924,N_907);
and U1017 (N_1017,N_976,N_999);
nor U1018 (N_1018,N_944,N_926);
or U1019 (N_1019,N_990,N_977);
or U1020 (N_1020,N_921,N_925);
nand U1021 (N_1021,N_928,N_987);
or U1022 (N_1022,N_932,N_931);
xor U1023 (N_1023,N_971,N_985);
and U1024 (N_1024,N_994,N_992);
nand U1025 (N_1025,N_945,N_948);
or U1026 (N_1026,N_966,N_934);
xor U1027 (N_1027,N_938,N_940);
nor U1028 (N_1028,N_949,N_908);
and U1029 (N_1029,N_903,N_958);
xor U1030 (N_1030,N_946,N_970);
or U1031 (N_1031,N_942,N_980);
nand U1032 (N_1032,N_954,N_933);
nor U1033 (N_1033,N_916,N_979);
nand U1034 (N_1034,N_920,N_998);
and U1035 (N_1035,N_913,N_917);
and U1036 (N_1036,N_936,N_905);
nor U1037 (N_1037,N_961,N_923);
nor U1038 (N_1038,N_911,N_922);
nand U1039 (N_1039,N_974,N_955);
nor U1040 (N_1040,N_984,N_909);
or U1041 (N_1041,N_975,N_937);
or U1042 (N_1042,N_978,N_906);
or U1043 (N_1043,N_902,N_900);
or U1044 (N_1044,N_963,N_995);
or U1045 (N_1045,N_901,N_952);
xor U1046 (N_1046,N_993,N_956);
nor U1047 (N_1047,N_947,N_968);
nand U1048 (N_1048,N_939,N_982);
nand U1049 (N_1049,N_941,N_904);
nor U1050 (N_1050,N_950,N_912);
nand U1051 (N_1051,N_947,N_983);
or U1052 (N_1052,N_929,N_905);
or U1053 (N_1053,N_921,N_988);
and U1054 (N_1054,N_919,N_995);
and U1055 (N_1055,N_925,N_919);
or U1056 (N_1056,N_918,N_981);
nand U1057 (N_1057,N_909,N_957);
nand U1058 (N_1058,N_983,N_991);
or U1059 (N_1059,N_992,N_920);
or U1060 (N_1060,N_999,N_962);
nor U1061 (N_1061,N_934,N_919);
nor U1062 (N_1062,N_904,N_998);
nand U1063 (N_1063,N_963,N_938);
nand U1064 (N_1064,N_943,N_996);
and U1065 (N_1065,N_987,N_943);
and U1066 (N_1066,N_988,N_924);
or U1067 (N_1067,N_946,N_971);
nand U1068 (N_1068,N_950,N_967);
nand U1069 (N_1069,N_994,N_941);
and U1070 (N_1070,N_991,N_927);
and U1071 (N_1071,N_956,N_977);
nor U1072 (N_1072,N_968,N_951);
or U1073 (N_1073,N_972,N_932);
nor U1074 (N_1074,N_959,N_967);
xnor U1075 (N_1075,N_907,N_991);
xnor U1076 (N_1076,N_940,N_992);
nand U1077 (N_1077,N_957,N_928);
and U1078 (N_1078,N_900,N_970);
xnor U1079 (N_1079,N_954,N_900);
and U1080 (N_1080,N_999,N_914);
nor U1081 (N_1081,N_923,N_978);
xor U1082 (N_1082,N_916,N_923);
nor U1083 (N_1083,N_983,N_935);
nand U1084 (N_1084,N_946,N_975);
nor U1085 (N_1085,N_905,N_968);
or U1086 (N_1086,N_987,N_977);
nand U1087 (N_1087,N_923,N_944);
and U1088 (N_1088,N_988,N_930);
nand U1089 (N_1089,N_962,N_903);
and U1090 (N_1090,N_992,N_946);
or U1091 (N_1091,N_981,N_933);
xor U1092 (N_1092,N_924,N_926);
nor U1093 (N_1093,N_904,N_972);
and U1094 (N_1094,N_945,N_930);
and U1095 (N_1095,N_941,N_971);
xnor U1096 (N_1096,N_958,N_983);
or U1097 (N_1097,N_989,N_928);
or U1098 (N_1098,N_987,N_960);
nor U1099 (N_1099,N_943,N_907);
and U1100 (N_1100,N_1037,N_1026);
and U1101 (N_1101,N_1016,N_1080);
nand U1102 (N_1102,N_1014,N_1095);
and U1103 (N_1103,N_1041,N_1059);
or U1104 (N_1104,N_1058,N_1086);
or U1105 (N_1105,N_1042,N_1072);
or U1106 (N_1106,N_1035,N_1065);
nor U1107 (N_1107,N_1084,N_1028);
nand U1108 (N_1108,N_1009,N_1075);
and U1109 (N_1109,N_1052,N_1082);
and U1110 (N_1110,N_1060,N_1043);
and U1111 (N_1111,N_1044,N_1064);
or U1112 (N_1112,N_1068,N_1013);
and U1113 (N_1113,N_1021,N_1054);
or U1114 (N_1114,N_1077,N_1098);
or U1115 (N_1115,N_1020,N_1039);
nand U1116 (N_1116,N_1004,N_1074);
nor U1117 (N_1117,N_1025,N_1003);
and U1118 (N_1118,N_1081,N_1007);
and U1119 (N_1119,N_1079,N_1036);
nand U1120 (N_1120,N_1018,N_1034);
nand U1121 (N_1121,N_1033,N_1023);
xnor U1122 (N_1122,N_1071,N_1076);
or U1123 (N_1123,N_1002,N_1019);
nor U1124 (N_1124,N_1083,N_1047);
or U1125 (N_1125,N_1073,N_1012);
or U1126 (N_1126,N_1040,N_1001);
nand U1127 (N_1127,N_1069,N_1048);
nand U1128 (N_1128,N_1045,N_1057);
nand U1129 (N_1129,N_1062,N_1032);
and U1130 (N_1130,N_1091,N_1099);
nand U1131 (N_1131,N_1031,N_1017);
xor U1132 (N_1132,N_1046,N_1066);
xnor U1133 (N_1133,N_1063,N_1049);
nor U1134 (N_1134,N_1096,N_1030);
and U1135 (N_1135,N_1056,N_1006);
nor U1136 (N_1136,N_1093,N_1094);
nand U1137 (N_1137,N_1038,N_1088);
or U1138 (N_1138,N_1011,N_1029);
and U1139 (N_1139,N_1097,N_1067);
or U1140 (N_1140,N_1027,N_1089);
nand U1141 (N_1141,N_1055,N_1000);
nor U1142 (N_1142,N_1070,N_1090);
and U1143 (N_1143,N_1005,N_1022);
and U1144 (N_1144,N_1015,N_1010);
or U1145 (N_1145,N_1053,N_1092);
nor U1146 (N_1146,N_1061,N_1087);
or U1147 (N_1147,N_1078,N_1024);
or U1148 (N_1148,N_1008,N_1051);
xnor U1149 (N_1149,N_1050,N_1085);
nand U1150 (N_1150,N_1039,N_1022);
and U1151 (N_1151,N_1038,N_1077);
and U1152 (N_1152,N_1051,N_1062);
and U1153 (N_1153,N_1099,N_1067);
or U1154 (N_1154,N_1026,N_1094);
and U1155 (N_1155,N_1047,N_1092);
nand U1156 (N_1156,N_1036,N_1017);
nand U1157 (N_1157,N_1021,N_1027);
or U1158 (N_1158,N_1056,N_1066);
or U1159 (N_1159,N_1014,N_1088);
and U1160 (N_1160,N_1081,N_1087);
nor U1161 (N_1161,N_1062,N_1043);
nand U1162 (N_1162,N_1065,N_1077);
nor U1163 (N_1163,N_1055,N_1002);
and U1164 (N_1164,N_1081,N_1008);
and U1165 (N_1165,N_1057,N_1085);
or U1166 (N_1166,N_1084,N_1058);
nand U1167 (N_1167,N_1048,N_1036);
and U1168 (N_1168,N_1083,N_1040);
and U1169 (N_1169,N_1010,N_1048);
nor U1170 (N_1170,N_1002,N_1044);
or U1171 (N_1171,N_1020,N_1041);
or U1172 (N_1172,N_1077,N_1032);
or U1173 (N_1173,N_1046,N_1021);
nand U1174 (N_1174,N_1022,N_1047);
or U1175 (N_1175,N_1061,N_1082);
or U1176 (N_1176,N_1024,N_1043);
nor U1177 (N_1177,N_1058,N_1021);
or U1178 (N_1178,N_1037,N_1018);
or U1179 (N_1179,N_1018,N_1073);
or U1180 (N_1180,N_1018,N_1065);
and U1181 (N_1181,N_1012,N_1050);
or U1182 (N_1182,N_1055,N_1037);
and U1183 (N_1183,N_1061,N_1044);
nor U1184 (N_1184,N_1088,N_1062);
nand U1185 (N_1185,N_1056,N_1020);
nand U1186 (N_1186,N_1098,N_1023);
nand U1187 (N_1187,N_1058,N_1088);
nor U1188 (N_1188,N_1021,N_1014);
or U1189 (N_1189,N_1088,N_1018);
nand U1190 (N_1190,N_1012,N_1064);
and U1191 (N_1191,N_1041,N_1095);
and U1192 (N_1192,N_1046,N_1047);
nand U1193 (N_1193,N_1011,N_1040);
and U1194 (N_1194,N_1090,N_1069);
nand U1195 (N_1195,N_1053,N_1031);
nor U1196 (N_1196,N_1037,N_1020);
xor U1197 (N_1197,N_1004,N_1053);
or U1198 (N_1198,N_1064,N_1031);
or U1199 (N_1199,N_1058,N_1032);
and U1200 (N_1200,N_1127,N_1107);
and U1201 (N_1201,N_1168,N_1134);
xor U1202 (N_1202,N_1105,N_1102);
nand U1203 (N_1203,N_1131,N_1137);
or U1204 (N_1204,N_1124,N_1192);
nand U1205 (N_1205,N_1184,N_1186);
nor U1206 (N_1206,N_1103,N_1143);
or U1207 (N_1207,N_1125,N_1163);
nor U1208 (N_1208,N_1179,N_1159);
xor U1209 (N_1209,N_1120,N_1130);
or U1210 (N_1210,N_1144,N_1135);
and U1211 (N_1211,N_1140,N_1198);
and U1212 (N_1212,N_1191,N_1149);
xor U1213 (N_1213,N_1172,N_1101);
nor U1214 (N_1214,N_1132,N_1142);
and U1215 (N_1215,N_1171,N_1187);
or U1216 (N_1216,N_1161,N_1166);
or U1217 (N_1217,N_1146,N_1164);
or U1218 (N_1218,N_1177,N_1100);
and U1219 (N_1219,N_1139,N_1126);
and U1220 (N_1220,N_1196,N_1112);
nor U1221 (N_1221,N_1173,N_1128);
nand U1222 (N_1222,N_1188,N_1118);
nor U1223 (N_1223,N_1147,N_1169);
and U1224 (N_1224,N_1162,N_1133);
nor U1225 (N_1225,N_1197,N_1190);
nand U1226 (N_1226,N_1167,N_1178);
nor U1227 (N_1227,N_1180,N_1115);
or U1228 (N_1228,N_1106,N_1151);
or U1229 (N_1229,N_1138,N_1189);
nand U1230 (N_1230,N_1104,N_1183);
and U1231 (N_1231,N_1170,N_1160);
nor U1232 (N_1232,N_1150,N_1185);
nor U1233 (N_1233,N_1108,N_1155);
or U1234 (N_1234,N_1195,N_1182);
or U1235 (N_1235,N_1123,N_1114);
nor U1236 (N_1236,N_1157,N_1199);
nor U1237 (N_1237,N_1117,N_1141);
xor U1238 (N_1238,N_1194,N_1113);
xnor U1239 (N_1239,N_1110,N_1148);
and U1240 (N_1240,N_1111,N_1174);
nand U1241 (N_1241,N_1156,N_1129);
xnor U1242 (N_1242,N_1109,N_1165);
xnor U1243 (N_1243,N_1175,N_1121);
or U1244 (N_1244,N_1158,N_1153);
nor U1245 (N_1245,N_1154,N_1116);
xnor U1246 (N_1246,N_1136,N_1176);
and U1247 (N_1247,N_1152,N_1119);
nand U1248 (N_1248,N_1122,N_1145);
and U1249 (N_1249,N_1193,N_1181);
and U1250 (N_1250,N_1178,N_1117);
and U1251 (N_1251,N_1133,N_1164);
nand U1252 (N_1252,N_1183,N_1161);
nor U1253 (N_1253,N_1115,N_1156);
nor U1254 (N_1254,N_1169,N_1178);
or U1255 (N_1255,N_1186,N_1107);
or U1256 (N_1256,N_1181,N_1177);
or U1257 (N_1257,N_1125,N_1194);
and U1258 (N_1258,N_1120,N_1181);
or U1259 (N_1259,N_1167,N_1118);
and U1260 (N_1260,N_1133,N_1134);
and U1261 (N_1261,N_1170,N_1127);
and U1262 (N_1262,N_1192,N_1102);
nor U1263 (N_1263,N_1126,N_1116);
or U1264 (N_1264,N_1180,N_1197);
xor U1265 (N_1265,N_1122,N_1112);
nor U1266 (N_1266,N_1157,N_1172);
nor U1267 (N_1267,N_1170,N_1132);
and U1268 (N_1268,N_1131,N_1194);
nand U1269 (N_1269,N_1128,N_1107);
or U1270 (N_1270,N_1140,N_1167);
nand U1271 (N_1271,N_1132,N_1126);
xor U1272 (N_1272,N_1193,N_1186);
or U1273 (N_1273,N_1139,N_1156);
nand U1274 (N_1274,N_1177,N_1109);
or U1275 (N_1275,N_1100,N_1181);
nand U1276 (N_1276,N_1171,N_1191);
and U1277 (N_1277,N_1125,N_1178);
and U1278 (N_1278,N_1186,N_1179);
or U1279 (N_1279,N_1147,N_1142);
nand U1280 (N_1280,N_1119,N_1182);
or U1281 (N_1281,N_1103,N_1100);
nand U1282 (N_1282,N_1167,N_1101);
and U1283 (N_1283,N_1179,N_1136);
and U1284 (N_1284,N_1141,N_1142);
or U1285 (N_1285,N_1140,N_1184);
xor U1286 (N_1286,N_1179,N_1197);
and U1287 (N_1287,N_1135,N_1145);
nand U1288 (N_1288,N_1198,N_1129);
or U1289 (N_1289,N_1171,N_1197);
or U1290 (N_1290,N_1181,N_1159);
nor U1291 (N_1291,N_1119,N_1199);
xor U1292 (N_1292,N_1113,N_1134);
or U1293 (N_1293,N_1186,N_1135);
nand U1294 (N_1294,N_1175,N_1157);
and U1295 (N_1295,N_1133,N_1167);
nand U1296 (N_1296,N_1127,N_1192);
nand U1297 (N_1297,N_1132,N_1152);
nand U1298 (N_1298,N_1182,N_1113);
xnor U1299 (N_1299,N_1154,N_1195);
nor U1300 (N_1300,N_1297,N_1223);
and U1301 (N_1301,N_1285,N_1278);
nand U1302 (N_1302,N_1243,N_1286);
xnor U1303 (N_1303,N_1260,N_1221);
and U1304 (N_1304,N_1235,N_1263);
or U1305 (N_1305,N_1245,N_1284);
or U1306 (N_1306,N_1292,N_1236);
nand U1307 (N_1307,N_1222,N_1290);
xor U1308 (N_1308,N_1206,N_1287);
nor U1309 (N_1309,N_1214,N_1282);
nor U1310 (N_1310,N_1209,N_1280);
nor U1311 (N_1311,N_1211,N_1269);
and U1312 (N_1312,N_1213,N_1219);
and U1313 (N_1313,N_1264,N_1216);
or U1314 (N_1314,N_1289,N_1298);
or U1315 (N_1315,N_1239,N_1225);
nand U1316 (N_1316,N_1217,N_1205);
xnor U1317 (N_1317,N_1266,N_1279);
or U1318 (N_1318,N_1210,N_1224);
nand U1319 (N_1319,N_1227,N_1267);
and U1320 (N_1320,N_1248,N_1262);
and U1321 (N_1321,N_1207,N_1247);
nand U1322 (N_1322,N_1231,N_1203);
or U1323 (N_1323,N_1230,N_1277);
or U1324 (N_1324,N_1252,N_1253);
and U1325 (N_1325,N_1275,N_1291);
xnor U1326 (N_1326,N_1258,N_1240);
nor U1327 (N_1327,N_1215,N_1273);
nor U1328 (N_1328,N_1272,N_1265);
nor U1329 (N_1329,N_1274,N_1233);
and U1330 (N_1330,N_1228,N_1212);
nor U1331 (N_1331,N_1208,N_1256);
or U1332 (N_1332,N_1259,N_1255);
and U1333 (N_1333,N_1261,N_1246);
or U1334 (N_1334,N_1270,N_1232);
nor U1335 (N_1335,N_1201,N_1281);
and U1336 (N_1336,N_1276,N_1200);
xor U1337 (N_1337,N_1234,N_1294);
nor U1338 (N_1338,N_1241,N_1202);
or U1339 (N_1339,N_1218,N_1238);
and U1340 (N_1340,N_1249,N_1254);
nor U1341 (N_1341,N_1251,N_1244);
nor U1342 (N_1342,N_1242,N_1257);
nand U1343 (N_1343,N_1296,N_1283);
xor U1344 (N_1344,N_1220,N_1293);
or U1345 (N_1345,N_1295,N_1268);
or U1346 (N_1346,N_1250,N_1229);
or U1347 (N_1347,N_1271,N_1226);
nor U1348 (N_1348,N_1204,N_1237);
or U1349 (N_1349,N_1288,N_1299);
and U1350 (N_1350,N_1249,N_1286);
nand U1351 (N_1351,N_1265,N_1211);
and U1352 (N_1352,N_1287,N_1237);
nor U1353 (N_1353,N_1288,N_1242);
nor U1354 (N_1354,N_1221,N_1288);
nand U1355 (N_1355,N_1277,N_1286);
xor U1356 (N_1356,N_1206,N_1293);
nand U1357 (N_1357,N_1290,N_1237);
and U1358 (N_1358,N_1252,N_1251);
nor U1359 (N_1359,N_1290,N_1213);
xnor U1360 (N_1360,N_1244,N_1242);
or U1361 (N_1361,N_1246,N_1208);
or U1362 (N_1362,N_1234,N_1276);
nand U1363 (N_1363,N_1286,N_1273);
and U1364 (N_1364,N_1293,N_1277);
and U1365 (N_1365,N_1216,N_1219);
and U1366 (N_1366,N_1247,N_1273);
and U1367 (N_1367,N_1203,N_1220);
and U1368 (N_1368,N_1295,N_1269);
nor U1369 (N_1369,N_1272,N_1237);
nor U1370 (N_1370,N_1294,N_1274);
nor U1371 (N_1371,N_1208,N_1235);
xor U1372 (N_1372,N_1246,N_1294);
nand U1373 (N_1373,N_1214,N_1292);
nand U1374 (N_1374,N_1280,N_1272);
nor U1375 (N_1375,N_1201,N_1238);
and U1376 (N_1376,N_1275,N_1242);
or U1377 (N_1377,N_1222,N_1225);
nand U1378 (N_1378,N_1216,N_1286);
and U1379 (N_1379,N_1233,N_1200);
xnor U1380 (N_1380,N_1256,N_1219);
xor U1381 (N_1381,N_1237,N_1278);
and U1382 (N_1382,N_1225,N_1200);
nand U1383 (N_1383,N_1272,N_1292);
and U1384 (N_1384,N_1278,N_1290);
or U1385 (N_1385,N_1265,N_1229);
or U1386 (N_1386,N_1272,N_1261);
nand U1387 (N_1387,N_1211,N_1292);
and U1388 (N_1388,N_1204,N_1229);
nand U1389 (N_1389,N_1279,N_1252);
or U1390 (N_1390,N_1217,N_1209);
and U1391 (N_1391,N_1283,N_1214);
and U1392 (N_1392,N_1235,N_1285);
or U1393 (N_1393,N_1244,N_1240);
or U1394 (N_1394,N_1237,N_1277);
and U1395 (N_1395,N_1209,N_1247);
and U1396 (N_1396,N_1241,N_1243);
nand U1397 (N_1397,N_1296,N_1256);
and U1398 (N_1398,N_1267,N_1294);
or U1399 (N_1399,N_1245,N_1246);
nand U1400 (N_1400,N_1322,N_1301);
nand U1401 (N_1401,N_1336,N_1342);
nand U1402 (N_1402,N_1339,N_1318);
nand U1403 (N_1403,N_1350,N_1381);
nor U1404 (N_1404,N_1356,N_1377);
and U1405 (N_1405,N_1370,N_1354);
nor U1406 (N_1406,N_1366,N_1363);
xnor U1407 (N_1407,N_1379,N_1305);
and U1408 (N_1408,N_1308,N_1303);
and U1409 (N_1409,N_1395,N_1384);
or U1410 (N_1410,N_1357,N_1347);
or U1411 (N_1411,N_1398,N_1394);
or U1412 (N_1412,N_1364,N_1331);
nand U1413 (N_1413,N_1326,N_1399);
or U1414 (N_1414,N_1324,N_1343);
nand U1415 (N_1415,N_1375,N_1351);
or U1416 (N_1416,N_1320,N_1321);
or U1417 (N_1417,N_1365,N_1374);
nand U1418 (N_1418,N_1376,N_1349);
nor U1419 (N_1419,N_1313,N_1360);
or U1420 (N_1420,N_1341,N_1361);
or U1421 (N_1421,N_1330,N_1314);
nand U1422 (N_1422,N_1345,N_1355);
nor U1423 (N_1423,N_1389,N_1329);
or U1424 (N_1424,N_1380,N_1302);
xor U1425 (N_1425,N_1387,N_1306);
xnor U1426 (N_1426,N_1319,N_1332);
and U1427 (N_1427,N_1352,N_1369);
or U1428 (N_1428,N_1388,N_1396);
nand U1429 (N_1429,N_1304,N_1335);
and U1430 (N_1430,N_1386,N_1373);
nor U1431 (N_1431,N_1311,N_1358);
nand U1432 (N_1432,N_1315,N_1372);
nor U1433 (N_1433,N_1367,N_1378);
or U1434 (N_1434,N_1393,N_1323);
nor U1435 (N_1435,N_1397,N_1338);
nand U1436 (N_1436,N_1317,N_1348);
nor U1437 (N_1437,N_1337,N_1383);
nor U1438 (N_1438,N_1371,N_1385);
nand U1439 (N_1439,N_1310,N_1334);
xor U1440 (N_1440,N_1344,N_1327);
nand U1441 (N_1441,N_1325,N_1362);
and U1442 (N_1442,N_1328,N_1346);
and U1443 (N_1443,N_1307,N_1391);
nor U1444 (N_1444,N_1300,N_1333);
nand U1445 (N_1445,N_1382,N_1312);
and U1446 (N_1446,N_1309,N_1316);
nand U1447 (N_1447,N_1340,N_1353);
nand U1448 (N_1448,N_1359,N_1390);
nand U1449 (N_1449,N_1392,N_1368);
and U1450 (N_1450,N_1333,N_1338);
and U1451 (N_1451,N_1378,N_1329);
nor U1452 (N_1452,N_1301,N_1348);
nand U1453 (N_1453,N_1308,N_1300);
nand U1454 (N_1454,N_1322,N_1369);
and U1455 (N_1455,N_1339,N_1325);
or U1456 (N_1456,N_1301,N_1305);
nor U1457 (N_1457,N_1333,N_1382);
and U1458 (N_1458,N_1365,N_1335);
nand U1459 (N_1459,N_1386,N_1316);
nand U1460 (N_1460,N_1305,N_1340);
nor U1461 (N_1461,N_1394,N_1388);
or U1462 (N_1462,N_1333,N_1334);
nand U1463 (N_1463,N_1390,N_1357);
or U1464 (N_1464,N_1396,N_1346);
and U1465 (N_1465,N_1389,N_1320);
and U1466 (N_1466,N_1385,N_1357);
nand U1467 (N_1467,N_1348,N_1392);
nand U1468 (N_1468,N_1303,N_1304);
and U1469 (N_1469,N_1350,N_1341);
xor U1470 (N_1470,N_1301,N_1354);
nor U1471 (N_1471,N_1351,N_1377);
and U1472 (N_1472,N_1382,N_1364);
and U1473 (N_1473,N_1310,N_1337);
and U1474 (N_1474,N_1302,N_1351);
nand U1475 (N_1475,N_1361,N_1344);
nor U1476 (N_1476,N_1377,N_1337);
nand U1477 (N_1477,N_1305,N_1346);
nor U1478 (N_1478,N_1316,N_1344);
nor U1479 (N_1479,N_1393,N_1303);
or U1480 (N_1480,N_1345,N_1320);
or U1481 (N_1481,N_1339,N_1306);
or U1482 (N_1482,N_1325,N_1309);
nand U1483 (N_1483,N_1324,N_1317);
nand U1484 (N_1484,N_1347,N_1389);
and U1485 (N_1485,N_1377,N_1374);
nor U1486 (N_1486,N_1312,N_1384);
nand U1487 (N_1487,N_1396,N_1354);
and U1488 (N_1488,N_1353,N_1369);
xnor U1489 (N_1489,N_1305,N_1330);
nand U1490 (N_1490,N_1351,N_1331);
nand U1491 (N_1491,N_1313,N_1348);
nor U1492 (N_1492,N_1324,N_1308);
nand U1493 (N_1493,N_1380,N_1315);
nor U1494 (N_1494,N_1337,N_1351);
nor U1495 (N_1495,N_1340,N_1311);
and U1496 (N_1496,N_1300,N_1356);
nand U1497 (N_1497,N_1395,N_1397);
nor U1498 (N_1498,N_1364,N_1352);
nor U1499 (N_1499,N_1398,N_1364);
and U1500 (N_1500,N_1431,N_1427);
nand U1501 (N_1501,N_1487,N_1439);
or U1502 (N_1502,N_1495,N_1408);
nand U1503 (N_1503,N_1492,N_1489);
or U1504 (N_1504,N_1464,N_1404);
xnor U1505 (N_1505,N_1474,N_1433);
or U1506 (N_1506,N_1402,N_1463);
nand U1507 (N_1507,N_1472,N_1453);
nand U1508 (N_1508,N_1468,N_1441);
and U1509 (N_1509,N_1443,N_1432);
or U1510 (N_1510,N_1419,N_1455);
or U1511 (N_1511,N_1410,N_1490);
nor U1512 (N_1512,N_1478,N_1493);
nor U1513 (N_1513,N_1449,N_1494);
nand U1514 (N_1514,N_1460,N_1421);
nor U1515 (N_1515,N_1413,N_1436);
and U1516 (N_1516,N_1451,N_1459);
nand U1517 (N_1517,N_1496,N_1454);
or U1518 (N_1518,N_1497,N_1471);
nand U1519 (N_1519,N_1477,N_1424);
nand U1520 (N_1520,N_1405,N_1444);
or U1521 (N_1521,N_1461,N_1442);
and U1522 (N_1522,N_1425,N_1417);
xor U1523 (N_1523,N_1452,N_1475);
or U1524 (N_1524,N_1437,N_1446);
nor U1525 (N_1525,N_1418,N_1476);
and U1526 (N_1526,N_1457,N_1447);
nand U1527 (N_1527,N_1440,N_1435);
nand U1528 (N_1528,N_1467,N_1434);
nand U1529 (N_1529,N_1466,N_1479);
or U1530 (N_1530,N_1486,N_1416);
or U1531 (N_1531,N_1426,N_1450);
nand U1532 (N_1532,N_1438,N_1462);
or U1533 (N_1533,N_1403,N_1473);
or U1534 (N_1534,N_1485,N_1412);
nor U1535 (N_1535,N_1420,N_1458);
nor U1536 (N_1536,N_1411,N_1480);
nand U1537 (N_1537,N_1445,N_1481);
or U1538 (N_1538,N_1428,N_1401);
nand U1539 (N_1539,N_1499,N_1400);
and U1540 (N_1540,N_1488,N_1484);
nand U1541 (N_1541,N_1470,N_1448);
nor U1542 (N_1542,N_1415,N_1456);
or U1543 (N_1543,N_1414,N_1491);
or U1544 (N_1544,N_1483,N_1422);
nor U1545 (N_1545,N_1407,N_1482);
nand U1546 (N_1546,N_1465,N_1429);
and U1547 (N_1547,N_1409,N_1406);
or U1548 (N_1548,N_1423,N_1430);
or U1549 (N_1549,N_1469,N_1498);
nor U1550 (N_1550,N_1404,N_1479);
and U1551 (N_1551,N_1439,N_1457);
or U1552 (N_1552,N_1474,N_1493);
or U1553 (N_1553,N_1499,N_1447);
or U1554 (N_1554,N_1402,N_1413);
and U1555 (N_1555,N_1495,N_1489);
nor U1556 (N_1556,N_1472,N_1414);
nand U1557 (N_1557,N_1424,N_1400);
and U1558 (N_1558,N_1450,N_1453);
and U1559 (N_1559,N_1493,N_1486);
and U1560 (N_1560,N_1411,N_1420);
or U1561 (N_1561,N_1486,N_1497);
nor U1562 (N_1562,N_1471,N_1472);
and U1563 (N_1563,N_1485,N_1419);
nor U1564 (N_1564,N_1434,N_1423);
nand U1565 (N_1565,N_1481,N_1452);
or U1566 (N_1566,N_1493,N_1441);
nor U1567 (N_1567,N_1420,N_1495);
or U1568 (N_1568,N_1417,N_1432);
nor U1569 (N_1569,N_1459,N_1484);
and U1570 (N_1570,N_1429,N_1445);
and U1571 (N_1571,N_1467,N_1495);
or U1572 (N_1572,N_1482,N_1493);
nor U1573 (N_1573,N_1423,N_1444);
or U1574 (N_1574,N_1446,N_1474);
and U1575 (N_1575,N_1493,N_1460);
nand U1576 (N_1576,N_1414,N_1454);
xor U1577 (N_1577,N_1417,N_1442);
and U1578 (N_1578,N_1468,N_1406);
and U1579 (N_1579,N_1408,N_1407);
nand U1580 (N_1580,N_1445,N_1457);
and U1581 (N_1581,N_1404,N_1423);
and U1582 (N_1582,N_1456,N_1419);
nor U1583 (N_1583,N_1436,N_1449);
xnor U1584 (N_1584,N_1456,N_1431);
xor U1585 (N_1585,N_1489,N_1497);
or U1586 (N_1586,N_1457,N_1415);
nor U1587 (N_1587,N_1458,N_1492);
or U1588 (N_1588,N_1442,N_1423);
xor U1589 (N_1589,N_1433,N_1465);
xnor U1590 (N_1590,N_1494,N_1417);
or U1591 (N_1591,N_1456,N_1428);
nand U1592 (N_1592,N_1403,N_1427);
nand U1593 (N_1593,N_1457,N_1400);
or U1594 (N_1594,N_1428,N_1458);
and U1595 (N_1595,N_1460,N_1479);
and U1596 (N_1596,N_1457,N_1499);
and U1597 (N_1597,N_1473,N_1488);
nand U1598 (N_1598,N_1480,N_1495);
and U1599 (N_1599,N_1433,N_1405);
nor U1600 (N_1600,N_1504,N_1500);
and U1601 (N_1601,N_1528,N_1559);
and U1602 (N_1602,N_1580,N_1545);
nand U1603 (N_1603,N_1587,N_1519);
and U1604 (N_1604,N_1551,N_1574);
or U1605 (N_1605,N_1588,N_1595);
nor U1606 (N_1606,N_1563,N_1526);
nor U1607 (N_1607,N_1584,N_1564);
xor U1608 (N_1608,N_1536,N_1514);
xor U1609 (N_1609,N_1581,N_1593);
nand U1610 (N_1610,N_1531,N_1555);
or U1611 (N_1611,N_1511,N_1599);
or U1612 (N_1612,N_1538,N_1512);
or U1613 (N_1613,N_1523,N_1592);
and U1614 (N_1614,N_1565,N_1549);
or U1615 (N_1615,N_1594,N_1527);
nor U1616 (N_1616,N_1515,N_1517);
and U1617 (N_1617,N_1502,N_1522);
nor U1618 (N_1618,N_1510,N_1572);
nor U1619 (N_1619,N_1579,N_1586);
or U1620 (N_1620,N_1547,N_1590);
xnor U1621 (N_1621,N_1550,N_1524);
and U1622 (N_1622,N_1567,N_1552);
or U1623 (N_1623,N_1521,N_1597);
nand U1624 (N_1624,N_1503,N_1591);
xor U1625 (N_1625,N_1577,N_1509);
or U1626 (N_1626,N_1582,N_1562);
and U1627 (N_1627,N_1561,N_1553);
nand U1628 (N_1628,N_1530,N_1507);
or U1629 (N_1629,N_1573,N_1557);
nor U1630 (N_1630,N_1505,N_1529);
nor U1631 (N_1631,N_1516,N_1558);
nor U1632 (N_1632,N_1598,N_1506);
and U1633 (N_1633,N_1540,N_1543);
xnor U1634 (N_1634,N_1542,N_1560);
nor U1635 (N_1635,N_1501,N_1589);
or U1636 (N_1636,N_1535,N_1532);
or U1637 (N_1637,N_1546,N_1568);
or U1638 (N_1638,N_1534,N_1508);
or U1639 (N_1639,N_1570,N_1533);
nor U1640 (N_1640,N_1539,N_1566);
and U1641 (N_1641,N_1554,N_1518);
nor U1642 (N_1642,N_1571,N_1537);
nor U1643 (N_1643,N_1548,N_1541);
nor U1644 (N_1644,N_1556,N_1544);
nor U1645 (N_1645,N_1583,N_1585);
and U1646 (N_1646,N_1569,N_1576);
nand U1647 (N_1647,N_1520,N_1596);
nand U1648 (N_1648,N_1525,N_1513);
xnor U1649 (N_1649,N_1578,N_1575);
and U1650 (N_1650,N_1563,N_1509);
nor U1651 (N_1651,N_1591,N_1519);
or U1652 (N_1652,N_1593,N_1546);
xor U1653 (N_1653,N_1583,N_1575);
nand U1654 (N_1654,N_1538,N_1584);
nand U1655 (N_1655,N_1541,N_1559);
and U1656 (N_1656,N_1597,N_1513);
or U1657 (N_1657,N_1568,N_1528);
nand U1658 (N_1658,N_1545,N_1533);
nor U1659 (N_1659,N_1592,N_1585);
or U1660 (N_1660,N_1515,N_1535);
nand U1661 (N_1661,N_1533,N_1527);
nor U1662 (N_1662,N_1547,N_1506);
or U1663 (N_1663,N_1572,N_1592);
nor U1664 (N_1664,N_1575,N_1540);
xnor U1665 (N_1665,N_1558,N_1543);
xnor U1666 (N_1666,N_1542,N_1548);
nand U1667 (N_1667,N_1516,N_1565);
or U1668 (N_1668,N_1562,N_1537);
or U1669 (N_1669,N_1523,N_1536);
xor U1670 (N_1670,N_1575,N_1512);
nand U1671 (N_1671,N_1556,N_1568);
or U1672 (N_1672,N_1502,N_1578);
nor U1673 (N_1673,N_1545,N_1569);
and U1674 (N_1674,N_1591,N_1508);
or U1675 (N_1675,N_1591,N_1576);
nand U1676 (N_1676,N_1597,N_1591);
nand U1677 (N_1677,N_1560,N_1510);
nor U1678 (N_1678,N_1550,N_1580);
nor U1679 (N_1679,N_1514,N_1551);
nor U1680 (N_1680,N_1545,N_1576);
nor U1681 (N_1681,N_1559,N_1581);
nand U1682 (N_1682,N_1501,N_1579);
nand U1683 (N_1683,N_1507,N_1590);
nor U1684 (N_1684,N_1554,N_1591);
nor U1685 (N_1685,N_1525,N_1595);
and U1686 (N_1686,N_1545,N_1549);
nor U1687 (N_1687,N_1529,N_1532);
nor U1688 (N_1688,N_1566,N_1579);
nor U1689 (N_1689,N_1571,N_1565);
or U1690 (N_1690,N_1567,N_1539);
nand U1691 (N_1691,N_1578,N_1588);
nor U1692 (N_1692,N_1547,N_1544);
xnor U1693 (N_1693,N_1594,N_1540);
and U1694 (N_1694,N_1530,N_1512);
nand U1695 (N_1695,N_1555,N_1561);
and U1696 (N_1696,N_1584,N_1583);
or U1697 (N_1697,N_1550,N_1567);
nor U1698 (N_1698,N_1521,N_1582);
xnor U1699 (N_1699,N_1575,N_1542);
and U1700 (N_1700,N_1643,N_1685);
or U1701 (N_1701,N_1689,N_1694);
nand U1702 (N_1702,N_1606,N_1691);
nand U1703 (N_1703,N_1642,N_1627);
nor U1704 (N_1704,N_1692,N_1610);
nand U1705 (N_1705,N_1673,N_1626);
nor U1706 (N_1706,N_1618,N_1663);
nor U1707 (N_1707,N_1630,N_1658);
nand U1708 (N_1708,N_1639,N_1678);
or U1709 (N_1709,N_1657,N_1615);
and U1710 (N_1710,N_1687,N_1697);
and U1711 (N_1711,N_1611,N_1617);
nand U1712 (N_1712,N_1662,N_1631);
nand U1713 (N_1713,N_1634,N_1651);
xor U1714 (N_1714,N_1655,N_1601);
nor U1715 (N_1715,N_1613,N_1609);
or U1716 (N_1716,N_1652,N_1688);
and U1717 (N_1717,N_1637,N_1644);
nand U1718 (N_1718,N_1649,N_1620);
nor U1719 (N_1719,N_1602,N_1698);
nand U1720 (N_1720,N_1612,N_1614);
or U1721 (N_1721,N_1603,N_1635);
nand U1722 (N_1722,N_1660,N_1674);
nor U1723 (N_1723,N_1661,N_1619);
nand U1724 (N_1724,N_1675,N_1669);
or U1725 (N_1725,N_1621,N_1682);
xnor U1726 (N_1726,N_1671,N_1654);
nor U1727 (N_1727,N_1665,N_1667);
nand U1728 (N_1728,N_1676,N_1664);
nor U1729 (N_1729,N_1629,N_1625);
xor U1730 (N_1730,N_1672,N_1693);
nor U1731 (N_1731,N_1670,N_1648);
nor U1732 (N_1732,N_1636,N_1690);
and U1733 (N_1733,N_1645,N_1607);
and U1734 (N_1734,N_1600,N_1647);
nor U1735 (N_1735,N_1659,N_1624);
nor U1736 (N_1736,N_1638,N_1668);
or U1737 (N_1737,N_1623,N_1666);
nand U1738 (N_1738,N_1684,N_1699);
nand U1739 (N_1739,N_1616,N_1683);
nand U1740 (N_1740,N_1604,N_1633);
nand U1741 (N_1741,N_1656,N_1641);
or U1742 (N_1742,N_1622,N_1646);
and U1743 (N_1743,N_1650,N_1608);
nand U1744 (N_1744,N_1628,N_1680);
or U1745 (N_1745,N_1677,N_1605);
and U1746 (N_1746,N_1695,N_1640);
nand U1747 (N_1747,N_1632,N_1679);
and U1748 (N_1748,N_1686,N_1696);
xnor U1749 (N_1749,N_1653,N_1681);
and U1750 (N_1750,N_1600,N_1678);
nand U1751 (N_1751,N_1623,N_1677);
nand U1752 (N_1752,N_1695,N_1604);
and U1753 (N_1753,N_1637,N_1672);
or U1754 (N_1754,N_1689,N_1632);
nor U1755 (N_1755,N_1658,N_1613);
nand U1756 (N_1756,N_1636,N_1692);
and U1757 (N_1757,N_1645,N_1665);
nand U1758 (N_1758,N_1653,N_1638);
nor U1759 (N_1759,N_1665,N_1616);
xor U1760 (N_1760,N_1685,N_1645);
nand U1761 (N_1761,N_1655,N_1691);
nand U1762 (N_1762,N_1696,N_1610);
and U1763 (N_1763,N_1663,N_1624);
nand U1764 (N_1764,N_1694,N_1683);
xnor U1765 (N_1765,N_1613,N_1603);
or U1766 (N_1766,N_1697,N_1676);
nor U1767 (N_1767,N_1625,N_1670);
or U1768 (N_1768,N_1630,N_1664);
and U1769 (N_1769,N_1690,N_1666);
xnor U1770 (N_1770,N_1690,N_1693);
nand U1771 (N_1771,N_1645,N_1641);
nand U1772 (N_1772,N_1647,N_1609);
and U1773 (N_1773,N_1653,N_1650);
or U1774 (N_1774,N_1679,N_1628);
or U1775 (N_1775,N_1695,N_1692);
and U1776 (N_1776,N_1654,N_1666);
nand U1777 (N_1777,N_1659,N_1682);
and U1778 (N_1778,N_1601,N_1648);
xor U1779 (N_1779,N_1663,N_1638);
nor U1780 (N_1780,N_1628,N_1653);
or U1781 (N_1781,N_1653,N_1611);
xnor U1782 (N_1782,N_1630,N_1651);
and U1783 (N_1783,N_1624,N_1689);
nand U1784 (N_1784,N_1645,N_1667);
nor U1785 (N_1785,N_1624,N_1685);
nand U1786 (N_1786,N_1639,N_1638);
nand U1787 (N_1787,N_1669,N_1612);
nand U1788 (N_1788,N_1621,N_1648);
nand U1789 (N_1789,N_1644,N_1605);
and U1790 (N_1790,N_1626,N_1676);
xor U1791 (N_1791,N_1693,N_1625);
xnor U1792 (N_1792,N_1630,N_1618);
or U1793 (N_1793,N_1693,N_1623);
nand U1794 (N_1794,N_1628,N_1659);
and U1795 (N_1795,N_1628,N_1609);
nand U1796 (N_1796,N_1699,N_1640);
xnor U1797 (N_1797,N_1664,N_1610);
xnor U1798 (N_1798,N_1615,N_1651);
and U1799 (N_1799,N_1637,N_1665);
nand U1800 (N_1800,N_1798,N_1725);
nor U1801 (N_1801,N_1726,N_1773);
and U1802 (N_1802,N_1786,N_1799);
and U1803 (N_1803,N_1724,N_1771);
or U1804 (N_1804,N_1791,N_1733);
nor U1805 (N_1805,N_1760,N_1743);
and U1806 (N_1806,N_1759,N_1779);
or U1807 (N_1807,N_1736,N_1778);
or U1808 (N_1808,N_1731,N_1762);
or U1809 (N_1809,N_1764,N_1742);
nor U1810 (N_1810,N_1752,N_1765);
and U1811 (N_1811,N_1777,N_1706);
or U1812 (N_1812,N_1701,N_1793);
or U1813 (N_1813,N_1792,N_1775);
nand U1814 (N_1814,N_1723,N_1789);
or U1815 (N_1815,N_1715,N_1711);
and U1816 (N_1816,N_1780,N_1721);
or U1817 (N_1817,N_1737,N_1730);
nor U1818 (N_1818,N_1782,N_1710);
or U1819 (N_1819,N_1785,N_1763);
xnor U1820 (N_1820,N_1797,N_1716);
nand U1821 (N_1821,N_1748,N_1790);
or U1822 (N_1822,N_1722,N_1795);
nand U1823 (N_1823,N_1702,N_1761);
nand U1824 (N_1824,N_1741,N_1705);
nand U1825 (N_1825,N_1707,N_1734);
and U1826 (N_1826,N_1787,N_1770);
nor U1827 (N_1827,N_1745,N_1758);
or U1828 (N_1828,N_1796,N_1750);
or U1829 (N_1829,N_1766,N_1703);
nor U1830 (N_1830,N_1749,N_1776);
and U1831 (N_1831,N_1794,N_1754);
nand U1832 (N_1832,N_1738,N_1727);
or U1833 (N_1833,N_1718,N_1744);
and U1834 (N_1834,N_1747,N_1714);
and U1835 (N_1835,N_1788,N_1772);
nor U1836 (N_1836,N_1729,N_1755);
nor U1837 (N_1837,N_1719,N_1712);
or U1838 (N_1838,N_1700,N_1751);
nand U1839 (N_1839,N_1783,N_1739);
or U1840 (N_1840,N_1768,N_1746);
nor U1841 (N_1841,N_1735,N_1769);
or U1842 (N_1842,N_1781,N_1784);
nand U1843 (N_1843,N_1708,N_1757);
and U1844 (N_1844,N_1713,N_1756);
xnor U1845 (N_1845,N_1732,N_1740);
nand U1846 (N_1846,N_1704,N_1774);
nand U1847 (N_1847,N_1709,N_1728);
and U1848 (N_1848,N_1717,N_1753);
nor U1849 (N_1849,N_1720,N_1767);
nor U1850 (N_1850,N_1712,N_1774);
nand U1851 (N_1851,N_1746,N_1710);
xnor U1852 (N_1852,N_1726,N_1721);
and U1853 (N_1853,N_1767,N_1790);
nor U1854 (N_1854,N_1718,N_1747);
nor U1855 (N_1855,N_1761,N_1790);
nand U1856 (N_1856,N_1762,N_1787);
or U1857 (N_1857,N_1763,N_1769);
or U1858 (N_1858,N_1798,N_1736);
nor U1859 (N_1859,N_1798,N_1757);
xnor U1860 (N_1860,N_1729,N_1727);
nand U1861 (N_1861,N_1791,N_1788);
nor U1862 (N_1862,N_1720,N_1765);
nor U1863 (N_1863,N_1787,N_1799);
nand U1864 (N_1864,N_1724,N_1759);
or U1865 (N_1865,N_1759,N_1723);
and U1866 (N_1866,N_1773,N_1744);
and U1867 (N_1867,N_1764,N_1766);
nor U1868 (N_1868,N_1763,N_1793);
and U1869 (N_1869,N_1702,N_1778);
nand U1870 (N_1870,N_1769,N_1736);
and U1871 (N_1871,N_1769,N_1730);
nor U1872 (N_1872,N_1741,N_1754);
xnor U1873 (N_1873,N_1757,N_1782);
and U1874 (N_1874,N_1720,N_1751);
xor U1875 (N_1875,N_1754,N_1705);
nor U1876 (N_1876,N_1713,N_1712);
and U1877 (N_1877,N_1794,N_1728);
xnor U1878 (N_1878,N_1727,N_1799);
xor U1879 (N_1879,N_1708,N_1754);
or U1880 (N_1880,N_1797,N_1727);
nor U1881 (N_1881,N_1709,N_1768);
nor U1882 (N_1882,N_1742,N_1762);
nor U1883 (N_1883,N_1776,N_1729);
nand U1884 (N_1884,N_1746,N_1715);
or U1885 (N_1885,N_1747,N_1745);
nand U1886 (N_1886,N_1717,N_1755);
and U1887 (N_1887,N_1708,N_1799);
or U1888 (N_1888,N_1700,N_1757);
or U1889 (N_1889,N_1772,N_1738);
nor U1890 (N_1890,N_1791,N_1703);
and U1891 (N_1891,N_1702,N_1710);
xor U1892 (N_1892,N_1711,N_1747);
xor U1893 (N_1893,N_1764,N_1775);
or U1894 (N_1894,N_1799,N_1703);
nand U1895 (N_1895,N_1749,N_1708);
and U1896 (N_1896,N_1735,N_1728);
or U1897 (N_1897,N_1792,N_1758);
and U1898 (N_1898,N_1766,N_1740);
nand U1899 (N_1899,N_1756,N_1718);
or U1900 (N_1900,N_1873,N_1809);
and U1901 (N_1901,N_1898,N_1816);
xor U1902 (N_1902,N_1842,N_1843);
nand U1903 (N_1903,N_1896,N_1806);
or U1904 (N_1904,N_1859,N_1862);
or U1905 (N_1905,N_1846,N_1833);
xor U1906 (N_1906,N_1866,N_1865);
xnor U1907 (N_1907,N_1849,N_1861);
and U1908 (N_1908,N_1805,N_1814);
nor U1909 (N_1909,N_1844,N_1808);
nor U1910 (N_1910,N_1800,N_1830);
nor U1911 (N_1911,N_1860,N_1883);
nand U1912 (N_1912,N_1819,N_1855);
nor U1913 (N_1913,N_1858,N_1825);
and U1914 (N_1914,N_1810,N_1812);
or U1915 (N_1915,N_1890,N_1889);
nand U1916 (N_1916,N_1869,N_1894);
or U1917 (N_1917,N_1831,N_1881);
nand U1918 (N_1918,N_1836,N_1815);
and U1919 (N_1919,N_1879,N_1804);
and U1920 (N_1920,N_1875,N_1828);
nor U1921 (N_1921,N_1897,N_1884);
nor U1922 (N_1922,N_1895,N_1863);
nor U1923 (N_1923,N_1886,N_1803);
nor U1924 (N_1924,N_1877,N_1848);
nor U1925 (N_1925,N_1823,N_1829);
and U1926 (N_1926,N_1834,N_1892);
xor U1927 (N_1927,N_1839,N_1847);
nor U1928 (N_1928,N_1824,N_1871);
and U1929 (N_1929,N_1872,N_1838);
and U1930 (N_1930,N_1885,N_1888);
nor U1931 (N_1931,N_1841,N_1826);
or U1932 (N_1932,N_1801,N_1802);
nand U1933 (N_1933,N_1853,N_1856);
xor U1934 (N_1934,N_1882,N_1891);
nand U1935 (N_1935,N_1832,N_1887);
nand U1936 (N_1936,N_1807,N_1850);
nor U1937 (N_1937,N_1837,N_1817);
or U1938 (N_1938,N_1854,N_1852);
and U1939 (N_1939,N_1870,N_1857);
xnor U1940 (N_1940,N_1820,N_1864);
or U1941 (N_1941,N_1822,N_1851);
xnor U1942 (N_1942,N_1867,N_1878);
nor U1943 (N_1943,N_1845,N_1811);
nand U1944 (N_1944,N_1880,N_1868);
nor U1945 (N_1945,N_1821,N_1835);
and U1946 (N_1946,N_1840,N_1874);
nor U1947 (N_1947,N_1818,N_1893);
or U1948 (N_1948,N_1813,N_1899);
or U1949 (N_1949,N_1827,N_1876);
nand U1950 (N_1950,N_1880,N_1890);
and U1951 (N_1951,N_1819,N_1883);
nor U1952 (N_1952,N_1814,N_1857);
nand U1953 (N_1953,N_1882,N_1850);
nand U1954 (N_1954,N_1822,N_1898);
nor U1955 (N_1955,N_1882,N_1834);
or U1956 (N_1956,N_1892,N_1800);
nand U1957 (N_1957,N_1830,N_1816);
nand U1958 (N_1958,N_1870,N_1859);
xor U1959 (N_1959,N_1841,N_1860);
or U1960 (N_1960,N_1812,N_1861);
or U1961 (N_1961,N_1847,N_1817);
and U1962 (N_1962,N_1896,N_1843);
and U1963 (N_1963,N_1866,N_1806);
or U1964 (N_1964,N_1846,N_1881);
or U1965 (N_1965,N_1820,N_1894);
nor U1966 (N_1966,N_1897,N_1808);
xnor U1967 (N_1967,N_1817,N_1812);
nor U1968 (N_1968,N_1898,N_1888);
or U1969 (N_1969,N_1834,N_1873);
or U1970 (N_1970,N_1830,N_1820);
and U1971 (N_1971,N_1837,N_1811);
nand U1972 (N_1972,N_1824,N_1872);
nor U1973 (N_1973,N_1834,N_1869);
nand U1974 (N_1974,N_1821,N_1877);
or U1975 (N_1975,N_1837,N_1849);
nand U1976 (N_1976,N_1808,N_1813);
nor U1977 (N_1977,N_1866,N_1856);
and U1978 (N_1978,N_1858,N_1865);
or U1979 (N_1979,N_1842,N_1808);
nor U1980 (N_1980,N_1853,N_1831);
xnor U1981 (N_1981,N_1866,N_1820);
nor U1982 (N_1982,N_1832,N_1803);
xnor U1983 (N_1983,N_1804,N_1890);
nor U1984 (N_1984,N_1875,N_1801);
nand U1985 (N_1985,N_1893,N_1842);
nor U1986 (N_1986,N_1873,N_1850);
nor U1987 (N_1987,N_1831,N_1816);
or U1988 (N_1988,N_1850,N_1831);
or U1989 (N_1989,N_1850,N_1877);
nand U1990 (N_1990,N_1803,N_1869);
nand U1991 (N_1991,N_1857,N_1884);
or U1992 (N_1992,N_1892,N_1888);
nand U1993 (N_1993,N_1808,N_1880);
xnor U1994 (N_1994,N_1890,N_1841);
and U1995 (N_1995,N_1891,N_1884);
or U1996 (N_1996,N_1865,N_1892);
and U1997 (N_1997,N_1857,N_1862);
or U1998 (N_1998,N_1867,N_1881);
or U1999 (N_1999,N_1852,N_1872);
nand U2000 (N_2000,N_1979,N_1927);
and U2001 (N_2001,N_1900,N_1914);
nand U2002 (N_2002,N_1972,N_1947);
nand U2003 (N_2003,N_1970,N_1988);
xor U2004 (N_2004,N_1958,N_1986);
xnor U2005 (N_2005,N_1995,N_1930);
and U2006 (N_2006,N_1918,N_1937);
xnor U2007 (N_2007,N_1998,N_1977);
nor U2008 (N_2008,N_1917,N_1993);
nand U2009 (N_2009,N_1905,N_1926);
nand U2010 (N_2010,N_1908,N_1954);
or U2011 (N_2011,N_1941,N_1973);
xor U2012 (N_2012,N_1922,N_1902);
or U2013 (N_2013,N_1971,N_1967);
or U2014 (N_2014,N_1983,N_1975);
nor U2015 (N_2015,N_1932,N_1963);
nand U2016 (N_2016,N_1911,N_1981);
xnor U2017 (N_2017,N_1934,N_1940);
or U2018 (N_2018,N_1945,N_1968);
and U2019 (N_2019,N_1969,N_1985);
or U2020 (N_2020,N_1912,N_1938);
xnor U2021 (N_2021,N_1987,N_1915);
and U2022 (N_2022,N_1956,N_1957);
nor U2023 (N_2023,N_1939,N_1976);
or U2024 (N_2024,N_1997,N_1966);
or U2025 (N_2025,N_1955,N_1929);
and U2026 (N_2026,N_1959,N_1953);
or U2027 (N_2027,N_1907,N_1903);
and U2028 (N_2028,N_1990,N_1933);
nand U2029 (N_2029,N_1980,N_1962);
nor U2030 (N_2030,N_1943,N_1961);
xor U2031 (N_2031,N_1991,N_1910);
xnor U2032 (N_2032,N_1951,N_1906);
nor U2033 (N_2033,N_1923,N_1950);
or U2034 (N_2034,N_1996,N_1982);
nor U2035 (N_2035,N_1960,N_1919);
or U2036 (N_2036,N_1909,N_1925);
nor U2037 (N_2037,N_1935,N_1946);
nand U2038 (N_2038,N_1901,N_1992);
or U2039 (N_2039,N_1952,N_1989);
or U2040 (N_2040,N_1928,N_1949);
and U2041 (N_2041,N_1913,N_1944);
nand U2042 (N_2042,N_1984,N_1999);
nand U2043 (N_2043,N_1916,N_1965);
or U2044 (N_2044,N_1936,N_1920);
xnor U2045 (N_2045,N_1921,N_1974);
and U2046 (N_2046,N_1994,N_1904);
and U2047 (N_2047,N_1931,N_1948);
and U2048 (N_2048,N_1924,N_1978);
nor U2049 (N_2049,N_1942,N_1964);
xor U2050 (N_2050,N_1954,N_1919);
nor U2051 (N_2051,N_1987,N_1975);
or U2052 (N_2052,N_1949,N_1960);
nand U2053 (N_2053,N_1981,N_1909);
and U2054 (N_2054,N_1952,N_1961);
or U2055 (N_2055,N_1916,N_1913);
nor U2056 (N_2056,N_1908,N_1974);
and U2057 (N_2057,N_1978,N_1975);
and U2058 (N_2058,N_1908,N_1964);
or U2059 (N_2059,N_1965,N_1947);
and U2060 (N_2060,N_1903,N_1958);
nor U2061 (N_2061,N_1985,N_1948);
or U2062 (N_2062,N_1905,N_1915);
nor U2063 (N_2063,N_1959,N_1970);
xnor U2064 (N_2064,N_1970,N_1917);
nor U2065 (N_2065,N_1979,N_1917);
or U2066 (N_2066,N_1942,N_1973);
nand U2067 (N_2067,N_1983,N_1927);
nor U2068 (N_2068,N_1914,N_1912);
nand U2069 (N_2069,N_1946,N_1936);
nand U2070 (N_2070,N_1934,N_1900);
or U2071 (N_2071,N_1984,N_1928);
nand U2072 (N_2072,N_1940,N_1949);
nor U2073 (N_2073,N_1971,N_1910);
nor U2074 (N_2074,N_1917,N_1925);
nor U2075 (N_2075,N_1909,N_1905);
xor U2076 (N_2076,N_1993,N_1928);
xor U2077 (N_2077,N_1922,N_1956);
and U2078 (N_2078,N_1973,N_1974);
nor U2079 (N_2079,N_1953,N_1900);
and U2080 (N_2080,N_1989,N_1972);
and U2081 (N_2081,N_1930,N_1915);
xor U2082 (N_2082,N_1953,N_1988);
nand U2083 (N_2083,N_1980,N_1928);
nand U2084 (N_2084,N_1983,N_1954);
xor U2085 (N_2085,N_1927,N_1955);
and U2086 (N_2086,N_1976,N_1978);
and U2087 (N_2087,N_1957,N_1978);
nand U2088 (N_2088,N_1954,N_1973);
and U2089 (N_2089,N_1943,N_1915);
and U2090 (N_2090,N_1956,N_1988);
nand U2091 (N_2091,N_1998,N_1914);
nor U2092 (N_2092,N_1908,N_1901);
nand U2093 (N_2093,N_1962,N_1946);
xor U2094 (N_2094,N_1985,N_1991);
and U2095 (N_2095,N_1930,N_1906);
nor U2096 (N_2096,N_1956,N_1900);
and U2097 (N_2097,N_1992,N_1990);
and U2098 (N_2098,N_1980,N_1933);
xnor U2099 (N_2099,N_1918,N_1903);
and U2100 (N_2100,N_2041,N_2092);
and U2101 (N_2101,N_2002,N_2010);
and U2102 (N_2102,N_2077,N_2031);
xnor U2103 (N_2103,N_2011,N_2063);
nand U2104 (N_2104,N_2037,N_2085);
and U2105 (N_2105,N_2027,N_2097);
or U2106 (N_2106,N_2042,N_2022);
or U2107 (N_2107,N_2080,N_2009);
and U2108 (N_2108,N_2008,N_2075);
or U2109 (N_2109,N_2015,N_2083);
and U2110 (N_2110,N_2053,N_2049);
nand U2111 (N_2111,N_2045,N_2003);
nor U2112 (N_2112,N_2098,N_2014);
nand U2113 (N_2113,N_2034,N_2068);
or U2114 (N_2114,N_2035,N_2094);
or U2115 (N_2115,N_2067,N_2069);
and U2116 (N_2116,N_2001,N_2084);
or U2117 (N_2117,N_2023,N_2090);
or U2118 (N_2118,N_2005,N_2047);
nand U2119 (N_2119,N_2028,N_2051);
or U2120 (N_2120,N_2089,N_2024);
nor U2121 (N_2121,N_2012,N_2029);
nand U2122 (N_2122,N_2036,N_2086);
nand U2123 (N_2123,N_2060,N_2070);
xnor U2124 (N_2124,N_2006,N_2026);
xnor U2125 (N_2125,N_2032,N_2081);
or U2126 (N_2126,N_2046,N_2062);
xor U2127 (N_2127,N_2043,N_2044);
xnor U2128 (N_2128,N_2019,N_2071);
xnor U2129 (N_2129,N_2065,N_2064);
and U2130 (N_2130,N_2033,N_2048);
nand U2131 (N_2131,N_2030,N_2000);
and U2132 (N_2132,N_2096,N_2038);
nand U2133 (N_2133,N_2007,N_2078);
xor U2134 (N_2134,N_2016,N_2066);
nor U2135 (N_2135,N_2061,N_2091);
nor U2136 (N_2136,N_2054,N_2087);
nor U2137 (N_2137,N_2099,N_2021);
and U2138 (N_2138,N_2076,N_2004);
and U2139 (N_2139,N_2082,N_2025);
nand U2140 (N_2140,N_2052,N_2058);
and U2141 (N_2141,N_2018,N_2073);
and U2142 (N_2142,N_2095,N_2079);
or U2143 (N_2143,N_2056,N_2040);
nand U2144 (N_2144,N_2074,N_2020);
and U2145 (N_2145,N_2057,N_2039);
nand U2146 (N_2146,N_2017,N_2072);
nor U2147 (N_2147,N_2093,N_2050);
or U2148 (N_2148,N_2088,N_2013);
or U2149 (N_2149,N_2059,N_2055);
nand U2150 (N_2150,N_2077,N_2022);
or U2151 (N_2151,N_2002,N_2075);
and U2152 (N_2152,N_2093,N_2001);
or U2153 (N_2153,N_2050,N_2083);
and U2154 (N_2154,N_2093,N_2070);
or U2155 (N_2155,N_2047,N_2072);
nor U2156 (N_2156,N_2049,N_2082);
or U2157 (N_2157,N_2029,N_2013);
or U2158 (N_2158,N_2071,N_2069);
nor U2159 (N_2159,N_2041,N_2014);
nand U2160 (N_2160,N_2064,N_2050);
and U2161 (N_2161,N_2052,N_2071);
and U2162 (N_2162,N_2009,N_2092);
or U2163 (N_2163,N_2017,N_2091);
nor U2164 (N_2164,N_2096,N_2032);
and U2165 (N_2165,N_2063,N_2003);
nand U2166 (N_2166,N_2040,N_2066);
and U2167 (N_2167,N_2023,N_2092);
nor U2168 (N_2168,N_2055,N_2013);
nand U2169 (N_2169,N_2063,N_2075);
or U2170 (N_2170,N_2081,N_2021);
and U2171 (N_2171,N_2068,N_2078);
nor U2172 (N_2172,N_2021,N_2093);
xnor U2173 (N_2173,N_2095,N_2002);
and U2174 (N_2174,N_2030,N_2001);
nand U2175 (N_2175,N_2083,N_2041);
nor U2176 (N_2176,N_2090,N_2096);
or U2177 (N_2177,N_2004,N_2098);
or U2178 (N_2178,N_2058,N_2027);
xnor U2179 (N_2179,N_2001,N_2064);
nor U2180 (N_2180,N_2062,N_2071);
and U2181 (N_2181,N_2069,N_2076);
and U2182 (N_2182,N_2041,N_2064);
and U2183 (N_2183,N_2032,N_2024);
xnor U2184 (N_2184,N_2015,N_2039);
nand U2185 (N_2185,N_2002,N_2079);
nor U2186 (N_2186,N_2046,N_2060);
nor U2187 (N_2187,N_2039,N_2006);
nand U2188 (N_2188,N_2067,N_2042);
or U2189 (N_2189,N_2097,N_2072);
or U2190 (N_2190,N_2086,N_2085);
nor U2191 (N_2191,N_2074,N_2033);
and U2192 (N_2192,N_2075,N_2022);
nand U2193 (N_2193,N_2013,N_2052);
nand U2194 (N_2194,N_2090,N_2016);
xnor U2195 (N_2195,N_2000,N_2051);
or U2196 (N_2196,N_2040,N_2057);
nor U2197 (N_2197,N_2002,N_2052);
nor U2198 (N_2198,N_2049,N_2069);
and U2199 (N_2199,N_2017,N_2047);
nand U2200 (N_2200,N_2196,N_2122);
nor U2201 (N_2201,N_2130,N_2125);
nor U2202 (N_2202,N_2188,N_2180);
or U2203 (N_2203,N_2116,N_2134);
nor U2204 (N_2204,N_2106,N_2166);
nor U2205 (N_2205,N_2189,N_2157);
or U2206 (N_2206,N_2186,N_2154);
nand U2207 (N_2207,N_2113,N_2162);
nand U2208 (N_2208,N_2149,N_2129);
or U2209 (N_2209,N_2194,N_2120);
nor U2210 (N_2210,N_2185,N_2139);
and U2211 (N_2211,N_2173,N_2158);
and U2212 (N_2212,N_2163,N_2124);
or U2213 (N_2213,N_2132,N_2136);
nand U2214 (N_2214,N_2114,N_2121);
or U2215 (N_2215,N_2170,N_2126);
nand U2216 (N_2216,N_2156,N_2169);
and U2217 (N_2217,N_2128,N_2153);
and U2218 (N_2218,N_2109,N_2164);
and U2219 (N_2219,N_2102,N_2195);
nor U2220 (N_2220,N_2111,N_2100);
nand U2221 (N_2221,N_2107,N_2197);
and U2222 (N_2222,N_2112,N_2198);
nor U2223 (N_2223,N_2131,N_2167);
nand U2224 (N_2224,N_2160,N_2191);
nor U2225 (N_2225,N_2155,N_2177);
or U2226 (N_2226,N_2135,N_2184);
xnor U2227 (N_2227,N_2144,N_2104);
and U2228 (N_2228,N_2183,N_2165);
and U2229 (N_2229,N_2187,N_2176);
nor U2230 (N_2230,N_2138,N_2115);
or U2231 (N_2231,N_2174,N_2127);
or U2232 (N_2232,N_2148,N_2123);
nor U2233 (N_2233,N_2152,N_2171);
xor U2234 (N_2234,N_2151,N_2108);
and U2235 (N_2235,N_2147,N_2137);
nand U2236 (N_2236,N_2179,N_2150);
xor U2237 (N_2237,N_2175,N_2181);
or U2238 (N_2238,N_2168,N_2199);
or U2239 (N_2239,N_2119,N_2117);
nand U2240 (N_2240,N_2103,N_2143);
or U2241 (N_2241,N_2161,N_2146);
and U2242 (N_2242,N_2118,N_2141);
or U2243 (N_2243,N_2105,N_2192);
and U2244 (N_2244,N_2190,N_2159);
nor U2245 (N_2245,N_2172,N_2140);
nand U2246 (N_2246,N_2178,N_2110);
or U2247 (N_2247,N_2133,N_2145);
and U2248 (N_2248,N_2182,N_2142);
nor U2249 (N_2249,N_2101,N_2193);
xnor U2250 (N_2250,N_2155,N_2183);
nor U2251 (N_2251,N_2179,N_2117);
or U2252 (N_2252,N_2184,N_2101);
nor U2253 (N_2253,N_2138,N_2178);
nor U2254 (N_2254,N_2143,N_2118);
nor U2255 (N_2255,N_2130,N_2104);
nand U2256 (N_2256,N_2128,N_2112);
nor U2257 (N_2257,N_2103,N_2180);
nand U2258 (N_2258,N_2184,N_2157);
or U2259 (N_2259,N_2162,N_2153);
nand U2260 (N_2260,N_2185,N_2190);
and U2261 (N_2261,N_2132,N_2191);
and U2262 (N_2262,N_2102,N_2130);
nand U2263 (N_2263,N_2139,N_2147);
or U2264 (N_2264,N_2185,N_2183);
and U2265 (N_2265,N_2134,N_2174);
and U2266 (N_2266,N_2127,N_2194);
nor U2267 (N_2267,N_2100,N_2108);
and U2268 (N_2268,N_2180,N_2111);
nand U2269 (N_2269,N_2177,N_2140);
or U2270 (N_2270,N_2124,N_2189);
and U2271 (N_2271,N_2171,N_2126);
and U2272 (N_2272,N_2167,N_2112);
nand U2273 (N_2273,N_2183,N_2116);
xnor U2274 (N_2274,N_2162,N_2155);
xor U2275 (N_2275,N_2123,N_2198);
xor U2276 (N_2276,N_2171,N_2180);
nand U2277 (N_2277,N_2162,N_2103);
nand U2278 (N_2278,N_2109,N_2153);
nand U2279 (N_2279,N_2122,N_2125);
or U2280 (N_2280,N_2106,N_2193);
or U2281 (N_2281,N_2111,N_2138);
or U2282 (N_2282,N_2141,N_2161);
nand U2283 (N_2283,N_2141,N_2121);
and U2284 (N_2284,N_2198,N_2109);
or U2285 (N_2285,N_2195,N_2162);
nor U2286 (N_2286,N_2130,N_2174);
nand U2287 (N_2287,N_2145,N_2155);
or U2288 (N_2288,N_2128,N_2133);
or U2289 (N_2289,N_2170,N_2166);
nand U2290 (N_2290,N_2129,N_2126);
or U2291 (N_2291,N_2125,N_2135);
and U2292 (N_2292,N_2107,N_2187);
and U2293 (N_2293,N_2173,N_2199);
nor U2294 (N_2294,N_2140,N_2166);
nor U2295 (N_2295,N_2109,N_2116);
nor U2296 (N_2296,N_2129,N_2107);
xnor U2297 (N_2297,N_2124,N_2178);
or U2298 (N_2298,N_2104,N_2132);
and U2299 (N_2299,N_2134,N_2140);
nand U2300 (N_2300,N_2201,N_2265);
xnor U2301 (N_2301,N_2223,N_2263);
and U2302 (N_2302,N_2207,N_2229);
nor U2303 (N_2303,N_2225,N_2296);
or U2304 (N_2304,N_2295,N_2210);
nand U2305 (N_2305,N_2213,N_2259);
xnor U2306 (N_2306,N_2278,N_2242);
or U2307 (N_2307,N_2299,N_2232);
xor U2308 (N_2308,N_2240,N_2234);
nand U2309 (N_2309,N_2251,N_2206);
nor U2310 (N_2310,N_2224,N_2264);
nor U2311 (N_2311,N_2291,N_2260);
and U2312 (N_2312,N_2287,N_2244);
nand U2313 (N_2313,N_2288,N_2238);
and U2314 (N_2314,N_2211,N_2246);
and U2315 (N_2315,N_2237,N_2255);
nand U2316 (N_2316,N_2272,N_2256);
nor U2317 (N_2317,N_2205,N_2273);
nor U2318 (N_2318,N_2239,N_2290);
nor U2319 (N_2319,N_2292,N_2297);
nor U2320 (N_2320,N_2218,N_2261);
nor U2321 (N_2321,N_2217,N_2243);
and U2322 (N_2322,N_2233,N_2227);
nor U2323 (N_2323,N_2216,N_2279);
or U2324 (N_2324,N_2268,N_2289);
nor U2325 (N_2325,N_2274,N_2285);
nor U2326 (N_2326,N_2267,N_2258);
xor U2327 (N_2327,N_2235,N_2269);
nor U2328 (N_2328,N_2271,N_2298);
nor U2329 (N_2329,N_2286,N_2294);
xnor U2330 (N_2330,N_2280,N_2204);
xor U2331 (N_2331,N_2247,N_2277);
xor U2332 (N_2332,N_2254,N_2209);
nand U2333 (N_2333,N_2249,N_2208);
xor U2334 (N_2334,N_2252,N_2276);
nor U2335 (N_2335,N_2226,N_2270);
xnor U2336 (N_2336,N_2214,N_2283);
nand U2337 (N_2337,N_2284,N_2222);
and U2338 (N_2338,N_2281,N_2212);
xor U2339 (N_2339,N_2202,N_2220);
nor U2340 (N_2340,N_2282,N_2275);
nor U2341 (N_2341,N_2230,N_2215);
and U2342 (N_2342,N_2228,N_2231);
or U2343 (N_2343,N_2262,N_2219);
or U2344 (N_2344,N_2293,N_2248);
or U2345 (N_2345,N_2253,N_2257);
nand U2346 (N_2346,N_2236,N_2241);
nor U2347 (N_2347,N_2203,N_2250);
or U2348 (N_2348,N_2245,N_2200);
nand U2349 (N_2349,N_2266,N_2221);
nor U2350 (N_2350,N_2294,N_2251);
or U2351 (N_2351,N_2289,N_2242);
nor U2352 (N_2352,N_2238,N_2249);
nor U2353 (N_2353,N_2260,N_2299);
nor U2354 (N_2354,N_2255,N_2299);
nor U2355 (N_2355,N_2274,N_2267);
and U2356 (N_2356,N_2238,N_2278);
and U2357 (N_2357,N_2207,N_2240);
and U2358 (N_2358,N_2203,N_2273);
nand U2359 (N_2359,N_2239,N_2229);
nor U2360 (N_2360,N_2244,N_2271);
xnor U2361 (N_2361,N_2218,N_2272);
nand U2362 (N_2362,N_2204,N_2286);
nand U2363 (N_2363,N_2285,N_2290);
and U2364 (N_2364,N_2277,N_2265);
and U2365 (N_2365,N_2252,N_2201);
xor U2366 (N_2366,N_2288,N_2247);
and U2367 (N_2367,N_2259,N_2229);
or U2368 (N_2368,N_2291,N_2282);
nand U2369 (N_2369,N_2296,N_2289);
and U2370 (N_2370,N_2216,N_2209);
or U2371 (N_2371,N_2261,N_2200);
nor U2372 (N_2372,N_2239,N_2243);
or U2373 (N_2373,N_2280,N_2298);
nand U2374 (N_2374,N_2266,N_2219);
nor U2375 (N_2375,N_2269,N_2297);
nand U2376 (N_2376,N_2273,N_2204);
nor U2377 (N_2377,N_2203,N_2263);
or U2378 (N_2378,N_2229,N_2242);
nor U2379 (N_2379,N_2270,N_2219);
or U2380 (N_2380,N_2212,N_2244);
xor U2381 (N_2381,N_2238,N_2209);
and U2382 (N_2382,N_2222,N_2281);
and U2383 (N_2383,N_2252,N_2260);
or U2384 (N_2384,N_2283,N_2230);
and U2385 (N_2385,N_2232,N_2227);
nand U2386 (N_2386,N_2223,N_2233);
nand U2387 (N_2387,N_2247,N_2221);
nor U2388 (N_2388,N_2286,N_2220);
nor U2389 (N_2389,N_2242,N_2285);
nor U2390 (N_2390,N_2200,N_2277);
nand U2391 (N_2391,N_2210,N_2249);
nand U2392 (N_2392,N_2244,N_2258);
nand U2393 (N_2393,N_2248,N_2250);
nor U2394 (N_2394,N_2205,N_2230);
nand U2395 (N_2395,N_2287,N_2202);
or U2396 (N_2396,N_2284,N_2209);
and U2397 (N_2397,N_2220,N_2242);
or U2398 (N_2398,N_2285,N_2284);
and U2399 (N_2399,N_2207,N_2203);
or U2400 (N_2400,N_2385,N_2310);
and U2401 (N_2401,N_2316,N_2378);
and U2402 (N_2402,N_2339,N_2374);
nand U2403 (N_2403,N_2341,N_2358);
nor U2404 (N_2404,N_2312,N_2338);
nor U2405 (N_2405,N_2307,N_2364);
and U2406 (N_2406,N_2354,N_2396);
and U2407 (N_2407,N_2365,N_2332);
nor U2408 (N_2408,N_2387,N_2397);
and U2409 (N_2409,N_2327,N_2389);
nor U2410 (N_2410,N_2323,N_2321);
nor U2411 (N_2411,N_2383,N_2359);
nand U2412 (N_2412,N_2353,N_2388);
nor U2413 (N_2413,N_2320,N_2352);
nor U2414 (N_2414,N_2382,N_2308);
or U2415 (N_2415,N_2319,N_2399);
nor U2416 (N_2416,N_2363,N_2326);
and U2417 (N_2417,N_2330,N_2313);
nor U2418 (N_2418,N_2336,N_2318);
nor U2419 (N_2419,N_2340,N_2305);
and U2420 (N_2420,N_2377,N_2350);
nand U2421 (N_2421,N_2306,N_2315);
nor U2422 (N_2422,N_2394,N_2391);
or U2423 (N_2423,N_2311,N_2301);
nand U2424 (N_2424,N_2333,N_2347);
nor U2425 (N_2425,N_2368,N_2325);
nor U2426 (N_2426,N_2334,N_2349);
nor U2427 (N_2427,N_2371,N_2348);
nand U2428 (N_2428,N_2366,N_2376);
nand U2429 (N_2429,N_2369,N_2380);
nor U2430 (N_2430,N_2373,N_2302);
and U2431 (N_2431,N_2335,N_2355);
or U2432 (N_2432,N_2324,N_2390);
xor U2433 (N_2433,N_2375,N_2343);
and U2434 (N_2434,N_2346,N_2342);
nand U2435 (N_2435,N_2303,N_2393);
and U2436 (N_2436,N_2381,N_2367);
nor U2437 (N_2437,N_2344,N_2351);
and U2438 (N_2438,N_2395,N_2379);
or U2439 (N_2439,N_2331,N_2356);
nand U2440 (N_2440,N_2398,N_2357);
and U2441 (N_2441,N_2361,N_2314);
xor U2442 (N_2442,N_2300,N_2372);
nor U2443 (N_2443,N_2328,N_2345);
nor U2444 (N_2444,N_2329,N_2304);
or U2445 (N_2445,N_2370,N_2317);
nand U2446 (N_2446,N_2337,N_2362);
and U2447 (N_2447,N_2384,N_2392);
or U2448 (N_2448,N_2322,N_2360);
and U2449 (N_2449,N_2309,N_2386);
nor U2450 (N_2450,N_2374,N_2359);
nand U2451 (N_2451,N_2398,N_2388);
nor U2452 (N_2452,N_2398,N_2392);
nor U2453 (N_2453,N_2333,N_2385);
nand U2454 (N_2454,N_2307,N_2390);
or U2455 (N_2455,N_2389,N_2357);
or U2456 (N_2456,N_2352,N_2306);
or U2457 (N_2457,N_2374,N_2378);
or U2458 (N_2458,N_2348,N_2338);
and U2459 (N_2459,N_2377,N_2313);
and U2460 (N_2460,N_2340,N_2335);
or U2461 (N_2461,N_2330,N_2374);
xor U2462 (N_2462,N_2374,N_2317);
or U2463 (N_2463,N_2306,N_2393);
or U2464 (N_2464,N_2349,N_2394);
nand U2465 (N_2465,N_2300,N_2322);
nor U2466 (N_2466,N_2329,N_2358);
nand U2467 (N_2467,N_2353,N_2348);
or U2468 (N_2468,N_2311,N_2307);
xnor U2469 (N_2469,N_2398,N_2374);
or U2470 (N_2470,N_2381,N_2399);
xnor U2471 (N_2471,N_2313,N_2393);
and U2472 (N_2472,N_2358,N_2300);
or U2473 (N_2473,N_2375,N_2308);
nor U2474 (N_2474,N_2324,N_2388);
xnor U2475 (N_2475,N_2386,N_2363);
nor U2476 (N_2476,N_2397,N_2301);
xnor U2477 (N_2477,N_2399,N_2325);
or U2478 (N_2478,N_2361,N_2392);
or U2479 (N_2479,N_2345,N_2394);
xor U2480 (N_2480,N_2333,N_2341);
or U2481 (N_2481,N_2320,N_2316);
nand U2482 (N_2482,N_2347,N_2394);
xnor U2483 (N_2483,N_2341,N_2300);
nor U2484 (N_2484,N_2311,N_2336);
or U2485 (N_2485,N_2312,N_2336);
nand U2486 (N_2486,N_2359,N_2358);
nand U2487 (N_2487,N_2375,N_2367);
xnor U2488 (N_2488,N_2365,N_2375);
xor U2489 (N_2489,N_2347,N_2318);
nand U2490 (N_2490,N_2311,N_2396);
or U2491 (N_2491,N_2335,N_2348);
nor U2492 (N_2492,N_2331,N_2372);
and U2493 (N_2493,N_2378,N_2348);
nor U2494 (N_2494,N_2305,N_2394);
and U2495 (N_2495,N_2314,N_2396);
and U2496 (N_2496,N_2365,N_2354);
xor U2497 (N_2497,N_2398,N_2360);
or U2498 (N_2498,N_2363,N_2366);
and U2499 (N_2499,N_2393,N_2341);
nor U2500 (N_2500,N_2442,N_2469);
xor U2501 (N_2501,N_2408,N_2468);
nand U2502 (N_2502,N_2453,N_2406);
or U2503 (N_2503,N_2438,N_2467);
and U2504 (N_2504,N_2458,N_2459);
nand U2505 (N_2505,N_2462,N_2483);
nand U2506 (N_2506,N_2414,N_2487);
and U2507 (N_2507,N_2429,N_2444);
or U2508 (N_2508,N_2417,N_2427);
or U2509 (N_2509,N_2477,N_2426);
or U2510 (N_2510,N_2412,N_2454);
nand U2511 (N_2511,N_2488,N_2432);
or U2512 (N_2512,N_2484,N_2430);
nand U2513 (N_2513,N_2478,N_2496);
and U2514 (N_2514,N_2470,N_2413);
or U2515 (N_2515,N_2441,N_2425);
and U2516 (N_2516,N_2420,N_2464);
and U2517 (N_2517,N_2410,N_2482);
or U2518 (N_2518,N_2466,N_2465);
or U2519 (N_2519,N_2440,N_2434);
nor U2520 (N_2520,N_2492,N_2452);
nand U2521 (N_2521,N_2421,N_2472);
nand U2522 (N_2522,N_2435,N_2486);
nor U2523 (N_2523,N_2471,N_2445);
and U2524 (N_2524,N_2409,N_2455);
and U2525 (N_2525,N_2415,N_2423);
and U2526 (N_2526,N_2495,N_2463);
or U2527 (N_2527,N_2456,N_2491);
xnor U2528 (N_2528,N_2402,N_2479);
nand U2529 (N_2529,N_2473,N_2447);
nand U2530 (N_2530,N_2480,N_2476);
nor U2531 (N_2531,N_2433,N_2405);
nor U2532 (N_2532,N_2439,N_2407);
nor U2533 (N_2533,N_2461,N_2449);
and U2534 (N_2534,N_2411,N_2443);
or U2535 (N_2535,N_2494,N_2424);
and U2536 (N_2536,N_2400,N_2450);
nor U2537 (N_2537,N_2403,N_2418);
xnor U2538 (N_2538,N_2436,N_2497);
and U2539 (N_2539,N_2448,N_2460);
and U2540 (N_2540,N_2489,N_2431);
and U2541 (N_2541,N_2416,N_2485);
nor U2542 (N_2542,N_2446,N_2437);
nor U2543 (N_2543,N_2499,N_2474);
or U2544 (N_2544,N_2457,N_2428);
and U2545 (N_2545,N_2498,N_2419);
nand U2546 (N_2546,N_2404,N_2451);
nand U2547 (N_2547,N_2401,N_2475);
and U2548 (N_2548,N_2493,N_2490);
nor U2549 (N_2549,N_2481,N_2422);
and U2550 (N_2550,N_2485,N_2450);
or U2551 (N_2551,N_2452,N_2407);
or U2552 (N_2552,N_2437,N_2441);
xnor U2553 (N_2553,N_2412,N_2450);
or U2554 (N_2554,N_2412,N_2417);
or U2555 (N_2555,N_2461,N_2499);
or U2556 (N_2556,N_2468,N_2486);
and U2557 (N_2557,N_2494,N_2437);
nor U2558 (N_2558,N_2442,N_2492);
nand U2559 (N_2559,N_2469,N_2491);
and U2560 (N_2560,N_2464,N_2452);
nand U2561 (N_2561,N_2451,N_2435);
or U2562 (N_2562,N_2436,N_2429);
and U2563 (N_2563,N_2400,N_2435);
and U2564 (N_2564,N_2474,N_2466);
xor U2565 (N_2565,N_2443,N_2469);
nand U2566 (N_2566,N_2471,N_2441);
nor U2567 (N_2567,N_2412,N_2480);
nor U2568 (N_2568,N_2497,N_2451);
or U2569 (N_2569,N_2412,N_2496);
nor U2570 (N_2570,N_2403,N_2438);
and U2571 (N_2571,N_2439,N_2463);
or U2572 (N_2572,N_2477,N_2456);
or U2573 (N_2573,N_2442,N_2455);
nor U2574 (N_2574,N_2423,N_2461);
or U2575 (N_2575,N_2401,N_2420);
or U2576 (N_2576,N_2486,N_2464);
xor U2577 (N_2577,N_2402,N_2404);
and U2578 (N_2578,N_2413,N_2441);
and U2579 (N_2579,N_2467,N_2458);
or U2580 (N_2580,N_2484,N_2413);
xnor U2581 (N_2581,N_2478,N_2469);
or U2582 (N_2582,N_2425,N_2471);
nand U2583 (N_2583,N_2472,N_2451);
xnor U2584 (N_2584,N_2467,N_2443);
and U2585 (N_2585,N_2481,N_2433);
nor U2586 (N_2586,N_2466,N_2400);
nand U2587 (N_2587,N_2447,N_2423);
nand U2588 (N_2588,N_2480,N_2437);
nor U2589 (N_2589,N_2452,N_2430);
nor U2590 (N_2590,N_2450,N_2464);
nand U2591 (N_2591,N_2409,N_2444);
and U2592 (N_2592,N_2476,N_2466);
nor U2593 (N_2593,N_2439,N_2470);
nor U2594 (N_2594,N_2433,N_2463);
nand U2595 (N_2595,N_2491,N_2487);
or U2596 (N_2596,N_2460,N_2452);
and U2597 (N_2597,N_2420,N_2462);
xnor U2598 (N_2598,N_2446,N_2442);
and U2599 (N_2599,N_2457,N_2420);
or U2600 (N_2600,N_2552,N_2553);
and U2601 (N_2601,N_2567,N_2561);
xnor U2602 (N_2602,N_2536,N_2572);
nor U2603 (N_2603,N_2509,N_2559);
nor U2604 (N_2604,N_2542,N_2598);
or U2605 (N_2605,N_2505,N_2594);
and U2606 (N_2606,N_2517,N_2550);
nand U2607 (N_2607,N_2581,N_2500);
nand U2608 (N_2608,N_2587,N_2525);
nor U2609 (N_2609,N_2514,N_2590);
nor U2610 (N_2610,N_2560,N_2522);
nor U2611 (N_2611,N_2555,N_2596);
or U2612 (N_2612,N_2586,N_2564);
nand U2613 (N_2613,N_2518,N_2510);
xnor U2614 (N_2614,N_2541,N_2511);
or U2615 (N_2615,N_2575,N_2589);
nand U2616 (N_2616,N_2568,N_2591);
and U2617 (N_2617,N_2570,N_2515);
nand U2618 (N_2618,N_2537,N_2529);
nor U2619 (N_2619,N_2538,N_2562);
nor U2620 (N_2620,N_2593,N_2502);
nand U2621 (N_2621,N_2521,N_2588);
nor U2622 (N_2622,N_2584,N_2571);
and U2623 (N_2623,N_2513,N_2543);
xor U2624 (N_2624,N_2595,N_2506);
nand U2625 (N_2625,N_2577,N_2566);
nor U2626 (N_2626,N_2534,N_2539);
xnor U2627 (N_2627,N_2527,N_2523);
or U2628 (N_2628,N_2530,N_2546);
and U2629 (N_2629,N_2599,N_2574);
nand U2630 (N_2630,N_2516,N_2533);
or U2631 (N_2631,N_2547,N_2551);
nand U2632 (N_2632,N_2512,N_2544);
nand U2633 (N_2633,N_2526,N_2558);
nor U2634 (N_2634,N_2540,N_2528);
or U2635 (N_2635,N_2520,N_2548);
nor U2636 (N_2636,N_2578,N_2532);
nand U2637 (N_2637,N_2583,N_2503);
or U2638 (N_2638,N_2545,N_2582);
nor U2639 (N_2639,N_2579,N_2524);
xnor U2640 (N_2640,N_2508,N_2576);
and U2641 (N_2641,N_2556,N_2563);
nor U2642 (N_2642,N_2531,N_2585);
nor U2643 (N_2643,N_2519,N_2501);
or U2644 (N_2644,N_2597,N_2507);
nor U2645 (N_2645,N_2569,N_2573);
or U2646 (N_2646,N_2580,N_2535);
nor U2647 (N_2647,N_2554,N_2557);
nand U2648 (N_2648,N_2592,N_2549);
nor U2649 (N_2649,N_2565,N_2504);
nor U2650 (N_2650,N_2529,N_2571);
nor U2651 (N_2651,N_2515,N_2519);
nor U2652 (N_2652,N_2523,N_2541);
or U2653 (N_2653,N_2554,N_2582);
or U2654 (N_2654,N_2551,N_2585);
or U2655 (N_2655,N_2520,N_2524);
nand U2656 (N_2656,N_2557,N_2550);
nand U2657 (N_2657,N_2533,N_2545);
nand U2658 (N_2658,N_2529,N_2595);
or U2659 (N_2659,N_2526,N_2587);
and U2660 (N_2660,N_2595,N_2593);
and U2661 (N_2661,N_2565,N_2567);
and U2662 (N_2662,N_2523,N_2545);
nor U2663 (N_2663,N_2513,N_2529);
and U2664 (N_2664,N_2529,N_2552);
nand U2665 (N_2665,N_2504,N_2587);
nor U2666 (N_2666,N_2598,N_2584);
and U2667 (N_2667,N_2568,N_2582);
nor U2668 (N_2668,N_2551,N_2533);
and U2669 (N_2669,N_2578,N_2548);
nor U2670 (N_2670,N_2537,N_2548);
nor U2671 (N_2671,N_2524,N_2542);
xnor U2672 (N_2672,N_2574,N_2560);
nand U2673 (N_2673,N_2518,N_2561);
or U2674 (N_2674,N_2560,N_2597);
or U2675 (N_2675,N_2599,N_2533);
and U2676 (N_2676,N_2597,N_2585);
or U2677 (N_2677,N_2569,N_2541);
and U2678 (N_2678,N_2599,N_2517);
or U2679 (N_2679,N_2598,N_2544);
nand U2680 (N_2680,N_2578,N_2549);
nor U2681 (N_2681,N_2599,N_2563);
nor U2682 (N_2682,N_2564,N_2523);
and U2683 (N_2683,N_2516,N_2572);
or U2684 (N_2684,N_2507,N_2580);
xnor U2685 (N_2685,N_2586,N_2584);
or U2686 (N_2686,N_2533,N_2547);
xor U2687 (N_2687,N_2531,N_2568);
nand U2688 (N_2688,N_2586,N_2542);
and U2689 (N_2689,N_2523,N_2540);
nand U2690 (N_2690,N_2506,N_2513);
nor U2691 (N_2691,N_2539,N_2511);
xor U2692 (N_2692,N_2580,N_2556);
nand U2693 (N_2693,N_2591,N_2589);
and U2694 (N_2694,N_2551,N_2529);
nor U2695 (N_2695,N_2506,N_2586);
nand U2696 (N_2696,N_2557,N_2536);
or U2697 (N_2697,N_2519,N_2549);
and U2698 (N_2698,N_2564,N_2546);
nand U2699 (N_2699,N_2568,N_2556);
or U2700 (N_2700,N_2678,N_2692);
nand U2701 (N_2701,N_2613,N_2610);
nand U2702 (N_2702,N_2620,N_2645);
and U2703 (N_2703,N_2656,N_2695);
xnor U2704 (N_2704,N_2666,N_2607);
and U2705 (N_2705,N_2627,N_2616);
nor U2706 (N_2706,N_2693,N_2604);
or U2707 (N_2707,N_2651,N_2662);
and U2708 (N_2708,N_2630,N_2623);
and U2709 (N_2709,N_2679,N_2684);
and U2710 (N_2710,N_2622,N_2697);
and U2711 (N_2711,N_2661,N_2672);
and U2712 (N_2712,N_2650,N_2639);
nand U2713 (N_2713,N_2624,N_2600);
nor U2714 (N_2714,N_2690,N_2626);
nor U2715 (N_2715,N_2605,N_2649);
nand U2716 (N_2716,N_2634,N_2667);
or U2717 (N_2717,N_2655,N_2643);
and U2718 (N_2718,N_2625,N_2682);
or U2719 (N_2719,N_2674,N_2698);
or U2720 (N_2720,N_2631,N_2676);
nor U2721 (N_2721,N_2621,N_2646);
and U2722 (N_2722,N_2603,N_2669);
nor U2723 (N_2723,N_2632,N_2602);
or U2724 (N_2724,N_2658,N_2647);
nand U2725 (N_2725,N_2691,N_2664);
and U2726 (N_2726,N_2671,N_2611);
or U2727 (N_2727,N_2694,N_2619);
nand U2728 (N_2728,N_2677,N_2644);
and U2729 (N_2729,N_2635,N_2685);
nor U2730 (N_2730,N_2601,N_2657);
nand U2731 (N_2731,N_2615,N_2628);
nor U2732 (N_2732,N_2606,N_2608);
and U2733 (N_2733,N_2688,N_2681);
nor U2734 (N_2734,N_2637,N_2668);
nor U2735 (N_2735,N_2652,N_2696);
nor U2736 (N_2736,N_2648,N_2680);
and U2737 (N_2737,N_2683,N_2614);
and U2738 (N_2738,N_2699,N_2638);
and U2739 (N_2739,N_2633,N_2653);
nand U2740 (N_2740,N_2654,N_2618);
and U2741 (N_2741,N_2687,N_2640);
nor U2742 (N_2742,N_2617,N_2665);
and U2743 (N_2743,N_2686,N_2673);
xnor U2744 (N_2744,N_2659,N_2670);
nand U2745 (N_2745,N_2629,N_2641);
and U2746 (N_2746,N_2636,N_2689);
or U2747 (N_2747,N_2675,N_2663);
nor U2748 (N_2748,N_2612,N_2642);
or U2749 (N_2749,N_2609,N_2660);
and U2750 (N_2750,N_2657,N_2614);
nand U2751 (N_2751,N_2621,N_2652);
xnor U2752 (N_2752,N_2651,N_2619);
nor U2753 (N_2753,N_2601,N_2668);
xnor U2754 (N_2754,N_2649,N_2620);
or U2755 (N_2755,N_2610,N_2675);
or U2756 (N_2756,N_2641,N_2654);
nand U2757 (N_2757,N_2639,N_2658);
or U2758 (N_2758,N_2649,N_2610);
nor U2759 (N_2759,N_2637,N_2647);
xor U2760 (N_2760,N_2660,N_2693);
nor U2761 (N_2761,N_2604,N_2655);
or U2762 (N_2762,N_2690,N_2638);
nand U2763 (N_2763,N_2625,N_2684);
and U2764 (N_2764,N_2655,N_2674);
and U2765 (N_2765,N_2613,N_2653);
xor U2766 (N_2766,N_2615,N_2650);
or U2767 (N_2767,N_2645,N_2697);
xor U2768 (N_2768,N_2693,N_2608);
xor U2769 (N_2769,N_2633,N_2603);
nand U2770 (N_2770,N_2692,N_2646);
xnor U2771 (N_2771,N_2665,N_2626);
and U2772 (N_2772,N_2686,N_2605);
nand U2773 (N_2773,N_2665,N_2601);
and U2774 (N_2774,N_2650,N_2614);
nand U2775 (N_2775,N_2654,N_2628);
or U2776 (N_2776,N_2672,N_2616);
nand U2777 (N_2777,N_2646,N_2605);
nor U2778 (N_2778,N_2601,N_2675);
nand U2779 (N_2779,N_2645,N_2623);
nand U2780 (N_2780,N_2604,N_2665);
and U2781 (N_2781,N_2608,N_2662);
nor U2782 (N_2782,N_2663,N_2667);
nand U2783 (N_2783,N_2665,N_2699);
and U2784 (N_2784,N_2697,N_2636);
xor U2785 (N_2785,N_2689,N_2625);
nor U2786 (N_2786,N_2617,N_2679);
nor U2787 (N_2787,N_2650,N_2600);
nand U2788 (N_2788,N_2628,N_2612);
and U2789 (N_2789,N_2675,N_2656);
nor U2790 (N_2790,N_2603,N_2674);
nand U2791 (N_2791,N_2643,N_2684);
or U2792 (N_2792,N_2653,N_2649);
or U2793 (N_2793,N_2670,N_2635);
or U2794 (N_2794,N_2616,N_2601);
xnor U2795 (N_2795,N_2619,N_2641);
or U2796 (N_2796,N_2614,N_2652);
and U2797 (N_2797,N_2667,N_2645);
nor U2798 (N_2798,N_2600,N_2664);
or U2799 (N_2799,N_2622,N_2664);
nor U2800 (N_2800,N_2700,N_2781);
nor U2801 (N_2801,N_2782,N_2711);
and U2802 (N_2802,N_2775,N_2744);
or U2803 (N_2803,N_2783,N_2704);
nor U2804 (N_2804,N_2789,N_2753);
nor U2805 (N_2805,N_2766,N_2702);
or U2806 (N_2806,N_2799,N_2726);
nand U2807 (N_2807,N_2715,N_2752);
or U2808 (N_2808,N_2735,N_2798);
xnor U2809 (N_2809,N_2756,N_2733);
and U2810 (N_2810,N_2746,N_2768);
nor U2811 (N_2811,N_2763,N_2788);
or U2812 (N_2812,N_2739,N_2703);
nand U2813 (N_2813,N_2732,N_2708);
or U2814 (N_2814,N_2751,N_2705);
nor U2815 (N_2815,N_2759,N_2776);
xor U2816 (N_2816,N_2794,N_2757);
nand U2817 (N_2817,N_2710,N_2765);
and U2818 (N_2818,N_2730,N_2796);
or U2819 (N_2819,N_2707,N_2755);
or U2820 (N_2820,N_2709,N_2792);
or U2821 (N_2821,N_2721,N_2731);
nand U2822 (N_2822,N_2769,N_2738);
and U2823 (N_2823,N_2712,N_2724);
and U2824 (N_2824,N_2719,N_2740);
and U2825 (N_2825,N_2761,N_2787);
or U2826 (N_2826,N_2734,N_2743);
nand U2827 (N_2827,N_2771,N_2748);
and U2828 (N_2828,N_2736,N_2785);
nand U2829 (N_2829,N_2773,N_2701);
nor U2830 (N_2830,N_2713,N_2780);
or U2831 (N_2831,N_2716,N_2714);
and U2832 (N_2832,N_2790,N_2764);
and U2833 (N_2833,N_2784,N_2728);
nor U2834 (N_2834,N_2718,N_2777);
and U2835 (N_2835,N_2779,N_2772);
nand U2836 (N_2836,N_2745,N_2737);
nor U2837 (N_2837,N_2717,N_2791);
nand U2838 (N_2838,N_2720,N_2706);
nand U2839 (N_2839,N_2786,N_2778);
or U2840 (N_2840,N_2754,N_2793);
nand U2841 (N_2841,N_2727,N_2722);
nor U2842 (N_2842,N_2774,N_2770);
or U2843 (N_2843,N_2725,N_2758);
nand U2844 (N_2844,N_2767,N_2742);
and U2845 (N_2845,N_2750,N_2760);
or U2846 (N_2846,N_2797,N_2747);
and U2847 (N_2847,N_2795,N_2741);
or U2848 (N_2848,N_2729,N_2723);
and U2849 (N_2849,N_2749,N_2762);
or U2850 (N_2850,N_2713,N_2790);
nor U2851 (N_2851,N_2742,N_2774);
nand U2852 (N_2852,N_2771,N_2792);
nand U2853 (N_2853,N_2701,N_2798);
and U2854 (N_2854,N_2780,N_2706);
or U2855 (N_2855,N_2734,N_2726);
nor U2856 (N_2856,N_2785,N_2755);
xor U2857 (N_2857,N_2720,N_2703);
or U2858 (N_2858,N_2703,N_2785);
or U2859 (N_2859,N_2789,N_2757);
and U2860 (N_2860,N_2748,N_2733);
and U2861 (N_2861,N_2734,N_2741);
nand U2862 (N_2862,N_2724,N_2741);
nor U2863 (N_2863,N_2743,N_2771);
or U2864 (N_2864,N_2700,N_2729);
xor U2865 (N_2865,N_2777,N_2716);
xor U2866 (N_2866,N_2728,N_2750);
and U2867 (N_2867,N_2770,N_2760);
nor U2868 (N_2868,N_2739,N_2765);
nand U2869 (N_2869,N_2760,N_2748);
nand U2870 (N_2870,N_2706,N_2769);
or U2871 (N_2871,N_2774,N_2717);
and U2872 (N_2872,N_2702,N_2779);
nand U2873 (N_2873,N_2732,N_2738);
nand U2874 (N_2874,N_2710,N_2751);
and U2875 (N_2875,N_2730,N_2793);
nand U2876 (N_2876,N_2747,N_2744);
or U2877 (N_2877,N_2711,N_2704);
or U2878 (N_2878,N_2724,N_2732);
and U2879 (N_2879,N_2794,N_2775);
nand U2880 (N_2880,N_2716,N_2723);
or U2881 (N_2881,N_2715,N_2722);
nor U2882 (N_2882,N_2752,N_2747);
nor U2883 (N_2883,N_2710,N_2790);
xor U2884 (N_2884,N_2796,N_2795);
or U2885 (N_2885,N_2774,N_2746);
nand U2886 (N_2886,N_2791,N_2716);
nand U2887 (N_2887,N_2734,N_2737);
nor U2888 (N_2888,N_2722,N_2798);
xor U2889 (N_2889,N_2712,N_2792);
nor U2890 (N_2890,N_2763,N_2752);
nand U2891 (N_2891,N_2775,N_2710);
nand U2892 (N_2892,N_2759,N_2738);
and U2893 (N_2893,N_2720,N_2723);
or U2894 (N_2894,N_2788,N_2748);
or U2895 (N_2895,N_2730,N_2733);
or U2896 (N_2896,N_2797,N_2749);
or U2897 (N_2897,N_2789,N_2717);
or U2898 (N_2898,N_2730,N_2720);
xor U2899 (N_2899,N_2701,N_2751);
and U2900 (N_2900,N_2821,N_2899);
or U2901 (N_2901,N_2857,N_2839);
nand U2902 (N_2902,N_2875,N_2881);
nand U2903 (N_2903,N_2824,N_2813);
or U2904 (N_2904,N_2818,N_2878);
or U2905 (N_2905,N_2887,N_2853);
nand U2906 (N_2906,N_2866,N_2849);
nor U2907 (N_2907,N_2890,N_2804);
and U2908 (N_2908,N_2838,N_2852);
nor U2909 (N_2909,N_2802,N_2819);
nor U2910 (N_2910,N_2871,N_2889);
or U2911 (N_2911,N_2808,N_2843);
nand U2912 (N_2912,N_2830,N_2873);
or U2913 (N_2913,N_2833,N_2879);
xor U2914 (N_2914,N_2891,N_2847);
nor U2915 (N_2915,N_2888,N_2895);
nand U2916 (N_2916,N_2874,N_2844);
or U2917 (N_2917,N_2841,N_2867);
and U2918 (N_2918,N_2805,N_2886);
xor U2919 (N_2919,N_2893,N_2883);
nand U2920 (N_2920,N_2816,N_2861);
nor U2921 (N_2921,N_2825,N_2820);
and U2922 (N_2922,N_2864,N_2806);
and U2923 (N_2923,N_2801,N_2845);
nor U2924 (N_2924,N_2860,N_2803);
and U2925 (N_2925,N_2836,N_2846);
nor U2926 (N_2926,N_2800,N_2826);
nand U2927 (N_2927,N_2898,N_2856);
nor U2928 (N_2928,N_2823,N_2834);
or U2929 (N_2929,N_2854,N_2872);
nor U2930 (N_2930,N_2885,N_2832);
or U2931 (N_2931,N_2815,N_2884);
or U2932 (N_2932,N_2863,N_2892);
or U2933 (N_2933,N_2870,N_2850);
nor U2934 (N_2934,N_2862,N_2848);
nor U2935 (N_2935,N_2828,N_2817);
nand U2936 (N_2936,N_2877,N_2896);
and U2937 (N_2937,N_2835,N_2876);
nor U2938 (N_2938,N_2842,N_2882);
nand U2939 (N_2939,N_2858,N_2807);
and U2940 (N_2940,N_2810,N_2831);
or U2941 (N_2941,N_2840,N_2865);
or U2942 (N_2942,N_2809,N_2814);
or U2943 (N_2943,N_2851,N_2859);
nor U2944 (N_2944,N_2894,N_2868);
or U2945 (N_2945,N_2837,N_2880);
and U2946 (N_2946,N_2869,N_2855);
and U2947 (N_2947,N_2811,N_2822);
nand U2948 (N_2948,N_2827,N_2829);
or U2949 (N_2949,N_2812,N_2897);
xor U2950 (N_2950,N_2829,N_2845);
nor U2951 (N_2951,N_2821,N_2844);
or U2952 (N_2952,N_2899,N_2842);
or U2953 (N_2953,N_2867,N_2802);
nand U2954 (N_2954,N_2832,N_2827);
nand U2955 (N_2955,N_2810,N_2806);
or U2956 (N_2956,N_2838,N_2803);
nor U2957 (N_2957,N_2857,N_2869);
and U2958 (N_2958,N_2870,N_2815);
nand U2959 (N_2959,N_2854,N_2891);
or U2960 (N_2960,N_2846,N_2859);
or U2961 (N_2961,N_2801,N_2811);
nor U2962 (N_2962,N_2866,N_2816);
nand U2963 (N_2963,N_2800,N_2848);
or U2964 (N_2964,N_2875,N_2868);
xnor U2965 (N_2965,N_2813,N_2809);
nand U2966 (N_2966,N_2816,N_2846);
or U2967 (N_2967,N_2811,N_2863);
and U2968 (N_2968,N_2899,N_2819);
nor U2969 (N_2969,N_2871,N_2840);
nor U2970 (N_2970,N_2851,N_2848);
nand U2971 (N_2971,N_2896,N_2866);
nand U2972 (N_2972,N_2816,N_2808);
nand U2973 (N_2973,N_2818,N_2868);
nand U2974 (N_2974,N_2854,N_2866);
nor U2975 (N_2975,N_2882,N_2838);
and U2976 (N_2976,N_2822,N_2885);
nor U2977 (N_2977,N_2879,N_2885);
xor U2978 (N_2978,N_2824,N_2812);
or U2979 (N_2979,N_2870,N_2840);
and U2980 (N_2980,N_2880,N_2834);
nor U2981 (N_2981,N_2803,N_2807);
or U2982 (N_2982,N_2882,N_2866);
and U2983 (N_2983,N_2823,N_2898);
nor U2984 (N_2984,N_2882,N_2861);
nand U2985 (N_2985,N_2821,N_2857);
nor U2986 (N_2986,N_2853,N_2885);
or U2987 (N_2987,N_2841,N_2895);
or U2988 (N_2988,N_2803,N_2893);
nand U2989 (N_2989,N_2806,N_2891);
or U2990 (N_2990,N_2880,N_2829);
nand U2991 (N_2991,N_2853,N_2832);
nand U2992 (N_2992,N_2830,N_2835);
xnor U2993 (N_2993,N_2862,N_2889);
nor U2994 (N_2994,N_2810,N_2892);
nand U2995 (N_2995,N_2887,N_2892);
or U2996 (N_2996,N_2894,N_2800);
xnor U2997 (N_2997,N_2857,N_2897);
nor U2998 (N_2998,N_2854,N_2831);
nand U2999 (N_2999,N_2887,N_2874);
or U3000 (N_3000,N_2991,N_2945);
and U3001 (N_3001,N_2943,N_2971);
and U3002 (N_3002,N_2970,N_2996);
nor U3003 (N_3003,N_2935,N_2930);
nand U3004 (N_3004,N_2908,N_2963);
nor U3005 (N_3005,N_2967,N_2920);
or U3006 (N_3006,N_2909,N_2907);
and U3007 (N_3007,N_2954,N_2923);
nand U3008 (N_3008,N_2999,N_2982);
nor U3009 (N_3009,N_2992,N_2917);
and U3010 (N_3010,N_2926,N_2903);
nand U3011 (N_3011,N_2912,N_2989);
and U3012 (N_3012,N_2902,N_2948);
xor U3013 (N_3013,N_2952,N_2906);
or U3014 (N_3014,N_2984,N_2977);
nor U3015 (N_3015,N_2990,N_2998);
nor U3016 (N_3016,N_2965,N_2934);
nor U3017 (N_3017,N_2981,N_2947);
nor U3018 (N_3018,N_2939,N_2933);
or U3019 (N_3019,N_2946,N_2913);
or U3020 (N_3020,N_2927,N_2951);
nand U3021 (N_3021,N_2941,N_2938);
and U3022 (N_3022,N_2916,N_2932);
nor U3023 (N_3023,N_2957,N_2980);
xor U3024 (N_3024,N_2944,N_2964);
xor U3025 (N_3025,N_2949,N_2914);
and U3026 (N_3026,N_2962,N_2973);
or U3027 (N_3027,N_2928,N_2911);
and U3028 (N_3028,N_2995,N_2950);
nand U3029 (N_3029,N_2931,N_2961);
and U3030 (N_3030,N_2924,N_2922);
or U3031 (N_3031,N_2905,N_2919);
nor U3032 (N_3032,N_2985,N_2986);
and U3033 (N_3033,N_2929,N_2936);
or U3034 (N_3034,N_2918,N_2955);
xor U3035 (N_3035,N_2937,N_2983);
nor U3036 (N_3036,N_2988,N_2993);
nand U3037 (N_3037,N_2900,N_2910);
nand U3038 (N_3038,N_2969,N_2958);
or U3039 (N_3039,N_2966,N_2953);
nor U3040 (N_3040,N_2975,N_2979);
nand U3041 (N_3041,N_2978,N_2942);
and U3042 (N_3042,N_2921,N_2994);
and U3043 (N_3043,N_2959,N_2968);
nand U3044 (N_3044,N_2976,N_2956);
or U3045 (N_3045,N_2987,N_2972);
or U3046 (N_3046,N_2940,N_2915);
or U3047 (N_3047,N_2901,N_2960);
and U3048 (N_3048,N_2904,N_2997);
or U3049 (N_3049,N_2974,N_2925);
and U3050 (N_3050,N_2947,N_2986);
and U3051 (N_3051,N_2956,N_2965);
nand U3052 (N_3052,N_2923,N_2905);
and U3053 (N_3053,N_2969,N_2991);
and U3054 (N_3054,N_2926,N_2998);
nand U3055 (N_3055,N_2963,N_2968);
and U3056 (N_3056,N_2942,N_2998);
or U3057 (N_3057,N_2949,N_2953);
nand U3058 (N_3058,N_2974,N_2958);
and U3059 (N_3059,N_2908,N_2920);
nor U3060 (N_3060,N_2903,N_2947);
nand U3061 (N_3061,N_2943,N_2958);
and U3062 (N_3062,N_2915,N_2966);
and U3063 (N_3063,N_2962,N_2933);
nand U3064 (N_3064,N_2984,N_2907);
and U3065 (N_3065,N_2961,N_2979);
and U3066 (N_3066,N_2913,N_2933);
nand U3067 (N_3067,N_2939,N_2937);
and U3068 (N_3068,N_2976,N_2939);
nor U3069 (N_3069,N_2944,N_2973);
nand U3070 (N_3070,N_2979,N_2934);
xor U3071 (N_3071,N_2947,N_2962);
nor U3072 (N_3072,N_2991,N_2947);
xnor U3073 (N_3073,N_2909,N_2977);
nor U3074 (N_3074,N_2977,N_2924);
nand U3075 (N_3075,N_2983,N_2988);
nand U3076 (N_3076,N_2952,N_2958);
xnor U3077 (N_3077,N_2901,N_2977);
nand U3078 (N_3078,N_2967,N_2925);
nand U3079 (N_3079,N_2987,N_2991);
nand U3080 (N_3080,N_2902,N_2976);
nor U3081 (N_3081,N_2985,N_2979);
or U3082 (N_3082,N_2989,N_2986);
nor U3083 (N_3083,N_2952,N_2962);
and U3084 (N_3084,N_2979,N_2994);
or U3085 (N_3085,N_2914,N_2953);
or U3086 (N_3086,N_2971,N_2932);
or U3087 (N_3087,N_2968,N_2951);
and U3088 (N_3088,N_2951,N_2963);
or U3089 (N_3089,N_2940,N_2917);
nand U3090 (N_3090,N_2908,N_2910);
nor U3091 (N_3091,N_2913,N_2996);
xor U3092 (N_3092,N_2915,N_2907);
xnor U3093 (N_3093,N_2955,N_2904);
xor U3094 (N_3094,N_2983,N_2910);
xor U3095 (N_3095,N_2916,N_2967);
xor U3096 (N_3096,N_2957,N_2913);
or U3097 (N_3097,N_2948,N_2967);
nand U3098 (N_3098,N_2933,N_2937);
nand U3099 (N_3099,N_2947,N_2954);
nor U3100 (N_3100,N_3095,N_3092);
or U3101 (N_3101,N_3067,N_3057);
nor U3102 (N_3102,N_3063,N_3098);
or U3103 (N_3103,N_3079,N_3049);
or U3104 (N_3104,N_3077,N_3082);
nor U3105 (N_3105,N_3054,N_3010);
and U3106 (N_3106,N_3004,N_3091);
or U3107 (N_3107,N_3056,N_3089);
nor U3108 (N_3108,N_3068,N_3002);
or U3109 (N_3109,N_3043,N_3024);
xnor U3110 (N_3110,N_3058,N_3061);
nand U3111 (N_3111,N_3086,N_3062);
or U3112 (N_3112,N_3020,N_3066);
or U3113 (N_3113,N_3069,N_3084);
nor U3114 (N_3114,N_3023,N_3074);
or U3115 (N_3115,N_3064,N_3022);
xor U3116 (N_3116,N_3031,N_3036);
nor U3117 (N_3117,N_3080,N_3039);
nand U3118 (N_3118,N_3011,N_3017);
nor U3119 (N_3119,N_3019,N_3038);
and U3120 (N_3120,N_3033,N_3044);
or U3121 (N_3121,N_3050,N_3087);
or U3122 (N_3122,N_3045,N_3037);
or U3123 (N_3123,N_3083,N_3001);
or U3124 (N_3124,N_3042,N_3096);
nand U3125 (N_3125,N_3055,N_3081);
nand U3126 (N_3126,N_3073,N_3070);
and U3127 (N_3127,N_3097,N_3000);
xor U3128 (N_3128,N_3026,N_3003);
or U3129 (N_3129,N_3005,N_3072);
nor U3130 (N_3130,N_3099,N_3046);
nor U3131 (N_3131,N_3012,N_3093);
nand U3132 (N_3132,N_3014,N_3040);
and U3133 (N_3133,N_3048,N_3016);
or U3134 (N_3134,N_3025,N_3094);
nand U3135 (N_3135,N_3009,N_3034);
nor U3136 (N_3136,N_3015,N_3088);
nand U3137 (N_3137,N_3059,N_3076);
and U3138 (N_3138,N_3085,N_3071);
nor U3139 (N_3139,N_3027,N_3021);
or U3140 (N_3140,N_3008,N_3030);
nor U3141 (N_3141,N_3047,N_3035);
nor U3142 (N_3142,N_3052,N_3013);
or U3143 (N_3143,N_3028,N_3053);
and U3144 (N_3144,N_3032,N_3075);
xor U3145 (N_3145,N_3041,N_3060);
xor U3146 (N_3146,N_3065,N_3006);
nor U3147 (N_3147,N_3018,N_3090);
nor U3148 (N_3148,N_3078,N_3029);
nand U3149 (N_3149,N_3051,N_3007);
nor U3150 (N_3150,N_3054,N_3023);
and U3151 (N_3151,N_3080,N_3044);
and U3152 (N_3152,N_3061,N_3040);
or U3153 (N_3153,N_3043,N_3037);
and U3154 (N_3154,N_3005,N_3018);
nor U3155 (N_3155,N_3072,N_3065);
nor U3156 (N_3156,N_3084,N_3008);
and U3157 (N_3157,N_3001,N_3066);
and U3158 (N_3158,N_3066,N_3006);
and U3159 (N_3159,N_3018,N_3000);
and U3160 (N_3160,N_3052,N_3074);
nand U3161 (N_3161,N_3082,N_3053);
or U3162 (N_3162,N_3077,N_3013);
and U3163 (N_3163,N_3028,N_3035);
nand U3164 (N_3164,N_3072,N_3068);
xnor U3165 (N_3165,N_3007,N_3080);
nor U3166 (N_3166,N_3077,N_3067);
nand U3167 (N_3167,N_3005,N_3001);
and U3168 (N_3168,N_3050,N_3032);
xnor U3169 (N_3169,N_3097,N_3088);
and U3170 (N_3170,N_3042,N_3029);
xnor U3171 (N_3171,N_3073,N_3015);
and U3172 (N_3172,N_3046,N_3053);
xor U3173 (N_3173,N_3046,N_3058);
nand U3174 (N_3174,N_3061,N_3026);
or U3175 (N_3175,N_3055,N_3036);
and U3176 (N_3176,N_3074,N_3022);
nor U3177 (N_3177,N_3065,N_3093);
or U3178 (N_3178,N_3018,N_3073);
and U3179 (N_3179,N_3001,N_3011);
or U3180 (N_3180,N_3022,N_3014);
xnor U3181 (N_3181,N_3099,N_3012);
xnor U3182 (N_3182,N_3067,N_3086);
and U3183 (N_3183,N_3044,N_3006);
or U3184 (N_3184,N_3012,N_3022);
nor U3185 (N_3185,N_3057,N_3007);
nand U3186 (N_3186,N_3098,N_3051);
nor U3187 (N_3187,N_3019,N_3034);
xor U3188 (N_3188,N_3058,N_3030);
nor U3189 (N_3189,N_3036,N_3073);
nand U3190 (N_3190,N_3022,N_3006);
and U3191 (N_3191,N_3043,N_3023);
nor U3192 (N_3192,N_3011,N_3006);
nand U3193 (N_3193,N_3090,N_3047);
nor U3194 (N_3194,N_3017,N_3000);
or U3195 (N_3195,N_3076,N_3051);
nand U3196 (N_3196,N_3067,N_3069);
nand U3197 (N_3197,N_3017,N_3047);
nand U3198 (N_3198,N_3055,N_3031);
or U3199 (N_3199,N_3022,N_3077);
xor U3200 (N_3200,N_3153,N_3199);
nand U3201 (N_3201,N_3192,N_3157);
nand U3202 (N_3202,N_3102,N_3143);
nor U3203 (N_3203,N_3128,N_3168);
xor U3204 (N_3204,N_3105,N_3152);
or U3205 (N_3205,N_3137,N_3124);
nor U3206 (N_3206,N_3136,N_3138);
and U3207 (N_3207,N_3181,N_3195);
and U3208 (N_3208,N_3183,N_3161);
and U3209 (N_3209,N_3185,N_3174);
nand U3210 (N_3210,N_3176,N_3180);
and U3211 (N_3211,N_3141,N_3177);
and U3212 (N_3212,N_3133,N_3155);
nand U3213 (N_3213,N_3134,N_3147);
or U3214 (N_3214,N_3198,N_3164);
nor U3215 (N_3215,N_3126,N_3166);
or U3216 (N_3216,N_3165,N_3100);
or U3217 (N_3217,N_3197,N_3112);
nor U3218 (N_3218,N_3169,N_3117);
nor U3219 (N_3219,N_3130,N_3160);
and U3220 (N_3220,N_3162,N_3150);
nor U3221 (N_3221,N_3163,N_3116);
or U3222 (N_3222,N_3107,N_3175);
and U3223 (N_3223,N_3148,N_3122);
and U3224 (N_3224,N_3156,N_3104);
nor U3225 (N_3225,N_3142,N_3159);
nor U3226 (N_3226,N_3193,N_3190);
or U3227 (N_3227,N_3140,N_3101);
or U3228 (N_3228,N_3187,N_3196);
or U3229 (N_3229,N_3145,N_3131);
or U3230 (N_3230,N_3139,N_3149);
xnor U3231 (N_3231,N_3172,N_3121);
nand U3232 (N_3232,N_3127,N_3110);
nor U3233 (N_3233,N_3167,N_3171);
and U3234 (N_3234,N_3184,N_3103);
nor U3235 (N_3235,N_3158,N_3178);
xnor U3236 (N_3236,N_3115,N_3114);
nand U3237 (N_3237,N_3151,N_3144);
or U3238 (N_3238,N_3154,N_3182);
nor U3239 (N_3239,N_3106,N_3119);
nand U3240 (N_3240,N_3111,N_3189);
nand U3241 (N_3241,N_3109,N_3135);
nand U3242 (N_3242,N_3125,N_3146);
or U3243 (N_3243,N_3120,N_3170);
nor U3244 (N_3244,N_3179,N_3188);
nand U3245 (N_3245,N_3132,N_3129);
xnor U3246 (N_3246,N_3173,N_3123);
and U3247 (N_3247,N_3118,N_3191);
and U3248 (N_3248,N_3186,N_3108);
and U3249 (N_3249,N_3113,N_3194);
nor U3250 (N_3250,N_3143,N_3193);
nor U3251 (N_3251,N_3182,N_3139);
xor U3252 (N_3252,N_3178,N_3163);
nand U3253 (N_3253,N_3141,N_3123);
or U3254 (N_3254,N_3162,N_3179);
nand U3255 (N_3255,N_3132,N_3189);
or U3256 (N_3256,N_3196,N_3188);
or U3257 (N_3257,N_3170,N_3179);
nand U3258 (N_3258,N_3170,N_3151);
nand U3259 (N_3259,N_3182,N_3141);
nor U3260 (N_3260,N_3177,N_3112);
and U3261 (N_3261,N_3176,N_3192);
or U3262 (N_3262,N_3164,N_3122);
and U3263 (N_3263,N_3162,N_3126);
xnor U3264 (N_3264,N_3188,N_3172);
and U3265 (N_3265,N_3173,N_3165);
and U3266 (N_3266,N_3130,N_3123);
nor U3267 (N_3267,N_3135,N_3198);
nand U3268 (N_3268,N_3157,N_3199);
xor U3269 (N_3269,N_3101,N_3131);
nand U3270 (N_3270,N_3143,N_3116);
nor U3271 (N_3271,N_3102,N_3140);
and U3272 (N_3272,N_3158,N_3115);
nand U3273 (N_3273,N_3134,N_3132);
nor U3274 (N_3274,N_3193,N_3170);
nor U3275 (N_3275,N_3199,N_3118);
nand U3276 (N_3276,N_3169,N_3131);
or U3277 (N_3277,N_3149,N_3155);
nor U3278 (N_3278,N_3116,N_3111);
nand U3279 (N_3279,N_3103,N_3196);
and U3280 (N_3280,N_3170,N_3146);
and U3281 (N_3281,N_3189,N_3147);
xnor U3282 (N_3282,N_3186,N_3147);
and U3283 (N_3283,N_3128,N_3177);
and U3284 (N_3284,N_3194,N_3173);
nor U3285 (N_3285,N_3169,N_3191);
or U3286 (N_3286,N_3158,N_3124);
nor U3287 (N_3287,N_3128,N_3152);
or U3288 (N_3288,N_3161,N_3137);
nand U3289 (N_3289,N_3133,N_3136);
nand U3290 (N_3290,N_3138,N_3122);
nand U3291 (N_3291,N_3135,N_3197);
nand U3292 (N_3292,N_3142,N_3165);
or U3293 (N_3293,N_3103,N_3189);
nand U3294 (N_3294,N_3163,N_3148);
and U3295 (N_3295,N_3199,N_3188);
nand U3296 (N_3296,N_3196,N_3191);
nor U3297 (N_3297,N_3127,N_3142);
or U3298 (N_3298,N_3176,N_3150);
or U3299 (N_3299,N_3112,N_3129);
nor U3300 (N_3300,N_3298,N_3266);
nand U3301 (N_3301,N_3293,N_3245);
or U3302 (N_3302,N_3216,N_3228);
and U3303 (N_3303,N_3270,N_3213);
and U3304 (N_3304,N_3272,N_3277);
nor U3305 (N_3305,N_3225,N_3279);
nor U3306 (N_3306,N_3233,N_3235);
nand U3307 (N_3307,N_3258,N_3290);
nand U3308 (N_3308,N_3241,N_3267);
nor U3309 (N_3309,N_3202,N_3240);
nand U3310 (N_3310,N_3204,N_3250);
xor U3311 (N_3311,N_3207,N_3208);
nor U3312 (N_3312,N_3227,N_3221);
nand U3313 (N_3313,N_3271,N_3275);
or U3314 (N_3314,N_3291,N_3237);
and U3315 (N_3315,N_3222,N_3249);
or U3316 (N_3316,N_3214,N_3259);
and U3317 (N_3317,N_3283,N_3210);
nand U3318 (N_3318,N_3253,N_3285);
and U3319 (N_3319,N_3223,N_3206);
nand U3320 (N_3320,N_3244,N_3242);
nand U3321 (N_3321,N_3281,N_3280);
and U3322 (N_3322,N_3247,N_3200);
nand U3323 (N_3323,N_3218,N_3287);
nor U3324 (N_3324,N_3203,N_3292);
nand U3325 (N_3325,N_3297,N_3274);
and U3326 (N_3326,N_3231,N_3251);
nor U3327 (N_3327,N_3209,N_3246);
xnor U3328 (N_3328,N_3226,N_3295);
nor U3329 (N_3329,N_3289,N_3238);
nor U3330 (N_3330,N_3265,N_3269);
nand U3331 (N_3331,N_3299,N_3286);
nand U3332 (N_3332,N_3268,N_3219);
nor U3333 (N_3333,N_3232,N_3224);
xor U3334 (N_3334,N_3239,N_3217);
or U3335 (N_3335,N_3255,N_3211);
nor U3336 (N_3336,N_3212,N_3229);
xor U3337 (N_3337,N_3201,N_3261);
nor U3338 (N_3338,N_3273,N_3243);
and U3339 (N_3339,N_3220,N_3236);
and U3340 (N_3340,N_3276,N_3215);
nor U3341 (N_3341,N_3288,N_3256);
nor U3342 (N_3342,N_3262,N_3294);
nand U3343 (N_3343,N_3205,N_3234);
nand U3344 (N_3344,N_3260,N_3254);
nor U3345 (N_3345,N_3284,N_3252);
or U3346 (N_3346,N_3248,N_3264);
nand U3347 (N_3347,N_3278,N_3230);
nand U3348 (N_3348,N_3263,N_3282);
nor U3349 (N_3349,N_3296,N_3257);
xor U3350 (N_3350,N_3252,N_3276);
nor U3351 (N_3351,N_3283,N_3230);
nor U3352 (N_3352,N_3263,N_3244);
nor U3353 (N_3353,N_3296,N_3218);
nand U3354 (N_3354,N_3224,N_3211);
xnor U3355 (N_3355,N_3285,N_3296);
or U3356 (N_3356,N_3216,N_3245);
and U3357 (N_3357,N_3254,N_3267);
nand U3358 (N_3358,N_3220,N_3287);
nand U3359 (N_3359,N_3277,N_3211);
or U3360 (N_3360,N_3222,N_3285);
nand U3361 (N_3361,N_3279,N_3274);
nand U3362 (N_3362,N_3283,N_3206);
nand U3363 (N_3363,N_3205,N_3261);
nor U3364 (N_3364,N_3242,N_3263);
or U3365 (N_3365,N_3254,N_3253);
and U3366 (N_3366,N_3273,N_3200);
or U3367 (N_3367,N_3277,N_3293);
xnor U3368 (N_3368,N_3287,N_3270);
xnor U3369 (N_3369,N_3271,N_3239);
or U3370 (N_3370,N_3226,N_3265);
or U3371 (N_3371,N_3266,N_3227);
nor U3372 (N_3372,N_3287,N_3285);
nand U3373 (N_3373,N_3243,N_3298);
or U3374 (N_3374,N_3254,N_3276);
nor U3375 (N_3375,N_3212,N_3241);
nand U3376 (N_3376,N_3227,N_3243);
and U3377 (N_3377,N_3202,N_3252);
nor U3378 (N_3378,N_3239,N_3218);
nand U3379 (N_3379,N_3243,N_3286);
or U3380 (N_3380,N_3248,N_3220);
or U3381 (N_3381,N_3254,N_3242);
nor U3382 (N_3382,N_3279,N_3265);
nand U3383 (N_3383,N_3263,N_3228);
xnor U3384 (N_3384,N_3236,N_3248);
and U3385 (N_3385,N_3249,N_3279);
nand U3386 (N_3386,N_3227,N_3232);
nand U3387 (N_3387,N_3275,N_3214);
and U3388 (N_3388,N_3276,N_3248);
or U3389 (N_3389,N_3293,N_3239);
xnor U3390 (N_3390,N_3213,N_3252);
nand U3391 (N_3391,N_3219,N_3280);
nor U3392 (N_3392,N_3277,N_3290);
and U3393 (N_3393,N_3205,N_3250);
and U3394 (N_3394,N_3238,N_3230);
nand U3395 (N_3395,N_3248,N_3222);
nor U3396 (N_3396,N_3221,N_3226);
nor U3397 (N_3397,N_3241,N_3210);
nor U3398 (N_3398,N_3280,N_3215);
nand U3399 (N_3399,N_3267,N_3216);
or U3400 (N_3400,N_3326,N_3372);
or U3401 (N_3401,N_3373,N_3303);
nand U3402 (N_3402,N_3301,N_3369);
nor U3403 (N_3403,N_3300,N_3358);
and U3404 (N_3404,N_3390,N_3386);
and U3405 (N_3405,N_3309,N_3376);
or U3406 (N_3406,N_3322,N_3387);
xor U3407 (N_3407,N_3361,N_3347);
nand U3408 (N_3408,N_3351,N_3362);
and U3409 (N_3409,N_3344,N_3350);
nor U3410 (N_3410,N_3320,N_3341);
and U3411 (N_3411,N_3364,N_3308);
and U3412 (N_3412,N_3332,N_3330);
nand U3413 (N_3413,N_3323,N_3315);
or U3414 (N_3414,N_3336,N_3342);
or U3415 (N_3415,N_3359,N_3375);
nand U3416 (N_3416,N_3324,N_3382);
nor U3417 (N_3417,N_3345,N_3377);
nor U3418 (N_3418,N_3321,N_3381);
nand U3419 (N_3419,N_3370,N_3319);
nor U3420 (N_3420,N_3395,N_3317);
or U3421 (N_3421,N_3318,N_3346);
or U3422 (N_3422,N_3339,N_3312);
or U3423 (N_3423,N_3393,N_3316);
nand U3424 (N_3424,N_3325,N_3337);
nor U3425 (N_3425,N_3366,N_3310);
or U3426 (N_3426,N_3307,N_3343);
or U3427 (N_3427,N_3314,N_3397);
or U3428 (N_3428,N_3380,N_3333);
and U3429 (N_3429,N_3334,N_3371);
and U3430 (N_3430,N_3335,N_3313);
nand U3431 (N_3431,N_3354,N_3391);
or U3432 (N_3432,N_3384,N_3349);
nand U3433 (N_3433,N_3360,N_3340);
nand U3434 (N_3434,N_3355,N_3363);
nand U3435 (N_3435,N_3353,N_3394);
or U3436 (N_3436,N_3383,N_3367);
xor U3437 (N_3437,N_3329,N_3328);
or U3438 (N_3438,N_3398,N_3389);
xor U3439 (N_3439,N_3338,N_3356);
nor U3440 (N_3440,N_3352,N_3379);
and U3441 (N_3441,N_3368,N_3327);
nor U3442 (N_3442,N_3396,N_3348);
or U3443 (N_3443,N_3311,N_3331);
and U3444 (N_3444,N_3305,N_3392);
or U3445 (N_3445,N_3302,N_3374);
nand U3446 (N_3446,N_3399,N_3306);
nand U3447 (N_3447,N_3357,N_3378);
nand U3448 (N_3448,N_3388,N_3365);
and U3449 (N_3449,N_3304,N_3385);
or U3450 (N_3450,N_3366,N_3378);
or U3451 (N_3451,N_3316,N_3358);
nand U3452 (N_3452,N_3326,N_3355);
and U3453 (N_3453,N_3367,N_3318);
nor U3454 (N_3454,N_3340,N_3366);
nor U3455 (N_3455,N_3304,N_3365);
and U3456 (N_3456,N_3379,N_3348);
nand U3457 (N_3457,N_3331,N_3327);
nand U3458 (N_3458,N_3359,N_3314);
or U3459 (N_3459,N_3326,N_3316);
and U3460 (N_3460,N_3374,N_3315);
nor U3461 (N_3461,N_3321,N_3332);
nor U3462 (N_3462,N_3309,N_3363);
xor U3463 (N_3463,N_3344,N_3378);
and U3464 (N_3464,N_3328,N_3316);
nand U3465 (N_3465,N_3368,N_3359);
nand U3466 (N_3466,N_3324,N_3372);
nor U3467 (N_3467,N_3322,N_3360);
xnor U3468 (N_3468,N_3330,N_3300);
xnor U3469 (N_3469,N_3331,N_3321);
and U3470 (N_3470,N_3352,N_3306);
nor U3471 (N_3471,N_3357,N_3367);
and U3472 (N_3472,N_3341,N_3314);
nor U3473 (N_3473,N_3368,N_3329);
nor U3474 (N_3474,N_3364,N_3332);
and U3475 (N_3475,N_3353,N_3382);
nand U3476 (N_3476,N_3336,N_3300);
nor U3477 (N_3477,N_3381,N_3303);
nand U3478 (N_3478,N_3374,N_3319);
nor U3479 (N_3479,N_3348,N_3306);
nand U3480 (N_3480,N_3384,N_3320);
nor U3481 (N_3481,N_3336,N_3393);
nand U3482 (N_3482,N_3378,N_3390);
nor U3483 (N_3483,N_3328,N_3310);
xnor U3484 (N_3484,N_3386,N_3392);
xnor U3485 (N_3485,N_3359,N_3330);
and U3486 (N_3486,N_3387,N_3373);
or U3487 (N_3487,N_3386,N_3383);
nand U3488 (N_3488,N_3325,N_3359);
nor U3489 (N_3489,N_3377,N_3394);
nor U3490 (N_3490,N_3303,N_3318);
xor U3491 (N_3491,N_3362,N_3382);
or U3492 (N_3492,N_3359,N_3354);
and U3493 (N_3493,N_3344,N_3387);
nand U3494 (N_3494,N_3390,N_3321);
nand U3495 (N_3495,N_3302,N_3349);
and U3496 (N_3496,N_3317,N_3396);
or U3497 (N_3497,N_3309,N_3354);
nand U3498 (N_3498,N_3395,N_3396);
nor U3499 (N_3499,N_3397,N_3333);
or U3500 (N_3500,N_3446,N_3438);
or U3501 (N_3501,N_3422,N_3432);
xnor U3502 (N_3502,N_3489,N_3488);
nor U3503 (N_3503,N_3463,N_3459);
or U3504 (N_3504,N_3475,N_3419);
nor U3505 (N_3505,N_3495,N_3445);
nor U3506 (N_3506,N_3498,N_3487);
nor U3507 (N_3507,N_3484,N_3409);
xor U3508 (N_3508,N_3454,N_3449);
or U3509 (N_3509,N_3442,N_3464);
nand U3510 (N_3510,N_3428,N_3465);
xor U3511 (N_3511,N_3444,N_3435);
nor U3512 (N_3512,N_3408,N_3482);
xnor U3513 (N_3513,N_3405,N_3407);
or U3514 (N_3514,N_3470,N_3424);
or U3515 (N_3515,N_3461,N_3417);
nand U3516 (N_3516,N_3425,N_3418);
nor U3517 (N_3517,N_3416,N_3473);
or U3518 (N_3518,N_3452,N_3443);
or U3519 (N_3519,N_3496,N_3455);
nand U3520 (N_3520,N_3457,N_3441);
or U3521 (N_3521,N_3490,N_3404);
nand U3522 (N_3522,N_3493,N_3494);
and U3523 (N_3523,N_3471,N_3402);
and U3524 (N_3524,N_3448,N_3476);
nor U3525 (N_3525,N_3400,N_3410);
nand U3526 (N_3526,N_3492,N_3421);
or U3527 (N_3527,N_3413,N_3433);
or U3528 (N_3528,N_3453,N_3477);
nor U3529 (N_3529,N_3403,N_3460);
and U3530 (N_3530,N_3486,N_3472);
and U3531 (N_3531,N_3479,N_3458);
and U3532 (N_3532,N_3415,N_3467);
nor U3533 (N_3533,N_3406,N_3431);
or U3534 (N_3534,N_3497,N_3483);
xnor U3535 (N_3535,N_3469,N_3478);
or U3536 (N_3536,N_3468,N_3480);
nor U3537 (N_3537,N_3412,N_3420);
xnor U3538 (N_3538,N_3485,N_3401);
or U3539 (N_3539,N_3440,N_3414);
and U3540 (N_3540,N_3426,N_3456);
and U3541 (N_3541,N_3447,N_3430);
or U3542 (N_3542,N_3499,N_3434);
or U3543 (N_3543,N_3474,N_3429);
and U3544 (N_3544,N_3423,N_3491);
nor U3545 (N_3545,N_3450,N_3411);
or U3546 (N_3546,N_3437,N_3427);
nand U3547 (N_3547,N_3436,N_3451);
and U3548 (N_3548,N_3462,N_3481);
and U3549 (N_3549,N_3439,N_3466);
or U3550 (N_3550,N_3437,N_3480);
or U3551 (N_3551,N_3421,N_3428);
and U3552 (N_3552,N_3485,N_3481);
nor U3553 (N_3553,N_3469,N_3467);
and U3554 (N_3554,N_3444,N_3469);
nand U3555 (N_3555,N_3426,N_3431);
nor U3556 (N_3556,N_3492,N_3425);
nand U3557 (N_3557,N_3469,N_3454);
or U3558 (N_3558,N_3420,N_3474);
nor U3559 (N_3559,N_3483,N_3442);
xnor U3560 (N_3560,N_3452,N_3467);
and U3561 (N_3561,N_3411,N_3414);
nand U3562 (N_3562,N_3484,N_3481);
nor U3563 (N_3563,N_3430,N_3444);
nor U3564 (N_3564,N_3414,N_3402);
xnor U3565 (N_3565,N_3473,N_3462);
or U3566 (N_3566,N_3457,N_3448);
nor U3567 (N_3567,N_3440,N_3490);
nand U3568 (N_3568,N_3451,N_3418);
and U3569 (N_3569,N_3422,N_3489);
nand U3570 (N_3570,N_3455,N_3446);
and U3571 (N_3571,N_3439,N_3443);
xor U3572 (N_3572,N_3490,N_3429);
nand U3573 (N_3573,N_3422,N_3455);
and U3574 (N_3574,N_3406,N_3484);
and U3575 (N_3575,N_3420,N_3451);
nor U3576 (N_3576,N_3440,N_3403);
and U3577 (N_3577,N_3409,N_3498);
or U3578 (N_3578,N_3405,N_3490);
nor U3579 (N_3579,N_3465,N_3403);
xor U3580 (N_3580,N_3470,N_3499);
nor U3581 (N_3581,N_3438,N_3488);
nor U3582 (N_3582,N_3449,N_3402);
nand U3583 (N_3583,N_3489,N_3496);
or U3584 (N_3584,N_3487,N_3401);
nand U3585 (N_3585,N_3466,N_3489);
xor U3586 (N_3586,N_3435,N_3464);
nor U3587 (N_3587,N_3425,N_3436);
nor U3588 (N_3588,N_3452,N_3456);
nor U3589 (N_3589,N_3499,N_3461);
nor U3590 (N_3590,N_3486,N_3488);
xor U3591 (N_3591,N_3477,N_3467);
nand U3592 (N_3592,N_3429,N_3424);
nor U3593 (N_3593,N_3434,N_3408);
nor U3594 (N_3594,N_3480,N_3417);
xor U3595 (N_3595,N_3496,N_3443);
xor U3596 (N_3596,N_3448,N_3432);
nand U3597 (N_3597,N_3470,N_3494);
xnor U3598 (N_3598,N_3408,N_3471);
and U3599 (N_3599,N_3414,N_3474);
and U3600 (N_3600,N_3567,N_3595);
or U3601 (N_3601,N_3569,N_3546);
or U3602 (N_3602,N_3549,N_3599);
nor U3603 (N_3603,N_3550,N_3570);
or U3604 (N_3604,N_3572,N_3517);
or U3605 (N_3605,N_3508,N_3539);
nand U3606 (N_3606,N_3574,N_3582);
or U3607 (N_3607,N_3533,N_3536);
and U3608 (N_3608,N_3575,N_3505);
and U3609 (N_3609,N_3556,N_3591);
and U3610 (N_3610,N_3548,N_3581);
nor U3611 (N_3611,N_3514,N_3525);
or U3612 (N_3612,N_3585,N_3588);
and U3613 (N_3613,N_3590,N_3502);
nor U3614 (N_3614,N_3560,N_3520);
and U3615 (N_3615,N_3530,N_3566);
or U3616 (N_3616,N_3542,N_3532);
nor U3617 (N_3617,N_3512,N_3522);
nand U3618 (N_3618,N_3503,N_3562);
nand U3619 (N_3619,N_3579,N_3552);
nand U3620 (N_3620,N_3564,N_3557);
or U3621 (N_3621,N_3565,N_3523);
nand U3622 (N_3622,N_3535,N_3541);
or U3623 (N_3623,N_3596,N_3510);
and U3624 (N_3624,N_3513,N_3584);
nand U3625 (N_3625,N_3504,N_3515);
or U3626 (N_3626,N_3547,N_3559);
and U3627 (N_3627,N_3555,N_3534);
and U3628 (N_3628,N_3568,N_3563);
nand U3629 (N_3629,N_3586,N_3580);
and U3630 (N_3630,N_3551,N_3501);
nor U3631 (N_3631,N_3524,N_3558);
nor U3632 (N_3632,N_3545,N_3516);
nor U3633 (N_3633,N_3561,N_3507);
nand U3634 (N_3634,N_3500,N_3594);
nor U3635 (N_3635,N_3598,N_3529);
nor U3636 (N_3636,N_3592,N_3554);
nor U3637 (N_3637,N_3537,N_3571);
or U3638 (N_3638,N_3519,N_3589);
and U3639 (N_3639,N_3511,N_3597);
xnor U3640 (N_3640,N_3583,N_3538);
or U3641 (N_3641,N_3528,N_3593);
nor U3642 (N_3642,N_3544,N_3543);
xor U3643 (N_3643,N_3518,N_3531);
and U3644 (N_3644,N_3509,N_3553);
nand U3645 (N_3645,N_3521,N_3527);
nand U3646 (N_3646,N_3577,N_3573);
nor U3647 (N_3647,N_3526,N_3578);
nor U3648 (N_3648,N_3576,N_3506);
or U3649 (N_3649,N_3540,N_3587);
nor U3650 (N_3650,N_3501,N_3517);
and U3651 (N_3651,N_3507,N_3538);
and U3652 (N_3652,N_3518,N_3521);
or U3653 (N_3653,N_3507,N_3579);
nor U3654 (N_3654,N_3579,N_3595);
nor U3655 (N_3655,N_3560,N_3510);
or U3656 (N_3656,N_3584,N_3525);
nor U3657 (N_3657,N_3575,N_3510);
or U3658 (N_3658,N_3562,N_3597);
or U3659 (N_3659,N_3579,N_3560);
xor U3660 (N_3660,N_3558,N_3513);
and U3661 (N_3661,N_3515,N_3503);
and U3662 (N_3662,N_3588,N_3515);
or U3663 (N_3663,N_3575,N_3521);
xnor U3664 (N_3664,N_3540,N_3584);
or U3665 (N_3665,N_3518,N_3572);
or U3666 (N_3666,N_3586,N_3562);
or U3667 (N_3667,N_3521,N_3547);
nor U3668 (N_3668,N_3516,N_3554);
and U3669 (N_3669,N_3575,N_3586);
nand U3670 (N_3670,N_3540,N_3570);
nor U3671 (N_3671,N_3592,N_3506);
and U3672 (N_3672,N_3540,N_3589);
nand U3673 (N_3673,N_3579,N_3589);
xnor U3674 (N_3674,N_3520,N_3535);
or U3675 (N_3675,N_3570,N_3562);
or U3676 (N_3676,N_3570,N_3524);
and U3677 (N_3677,N_3534,N_3577);
nor U3678 (N_3678,N_3545,N_3587);
or U3679 (N_3679,N_3551,N_3583);
nand U3680 (N_3680,N_3595,N_3546);
or U3681 (N_3681,N_3576,N_3512);
nand U3682 (N_3682,N_3544,N_3538);
and U3683 (N_3683,N_3551,N_3544);
nor U3684 (N_3684,N_3569,N_3532);
nand U3685 (N_3685,N_3580,N_3525);
and U3686 (N_3686,N_3506,N_3572);
nand U3687 (N_3687,N_3533,N_3508);
xnor U3688 (N_3688,N_3527,N_3572);
nand U3689 (N_3689,N_3515,N_3520);
nor U3690 (N_3690,N_3567,N_3547);
or U3691 (N_3691,N_3523,N_3534);
or U3692 (N_3692,N_3509,N_3565);
nor U3693 (N_3693,N_3588,N_3580);
or U3694 (N_3694,N_3563,N_3597);
nor U3695 (N_3695,N_3531,N_3563);
or U3696 (N_3696,N_3515,N_3586);
or U3697 (N_3697,N_3584,N_3511);
or U3698 (N_3698,N_3504,N_3507);
or U3699 (N_3699,N_3527,N_3505);
and U3700 (N_3700,N_3629,N_3635);
or U3701 (N_3701,N_3628,N_3672);
or U3702 (N_3702,N_3691,N_3699);
xnor U3703 (N_3703,N_3606,N_3654);
nor U3704 (N_3704,N_3631,N_3682);
nand U3705 (N_3705,N_3621,N_3617);
and U3706 (N_3706,N_3668,N_3626);
and U3707 (N_3707,N_3605,N_3680);
nand U3708 (N_3708,N_3664,N_3646);
and U3709 (N_3709,N_3641,N_3647);
nand U3710 (N_3710,N_3639,N_3645);
nor U3711 (N_3711,N_3665,N_3658);
nor U3712 (N_3712,N_3677,N_3640);
nand U3713 (N_3713,N_3697,N_3600);
nand U3714 (N_3714,N_3627,N_3657);
nand U3715 (N_3715,N_3688,N_3663);
and U3716 (N_3716,N_3624,N_3684);
or U3717 (N_3717,N_3695,N_3620);
and U3718 (N_3718,N_3634,N_3681);
and U3719 (N_3719,N_3690,N_3610);
nand U3720 (N_3720,N_3696,N_3643);
nand U3721 (N_3721,N_3604,N_3651);
or U3722 (N_3722,N_3611,N_3659);
nor U3723 (N_3723,N_3666,N_3667);
and U3724 (N_3724,N_3674,N_3670);
or U3725 (N_3725,N_3687,N_3622);
nand U3726 (N_3726,N_3648,N_3686);
and U3727 (N_3727,N_3673,N_3694);
nor U3728 (N_3728,N_3618,N_3669);
and U3729 (N_3729,N_3671,N_3607);
or U3730 (N_3730,N_3661,N_3601);
nor U3731 (N_3731,N_3655,N_3683);
nor U3732 (N_3732,N_3649,N_3698);
and U3733 (N_3733,N_3679,N_3614);
or U3734 (N_3734,N_3662,N_3632);
and U3735 (N_3735,N_3619,N_3676);
and U3736 (N_3736,N_3638,N_3608);
xor U3737 (N_3737,N_3637,N_3615);
xnor U3738 (N_3738,N_3644,N_3660);
or U3739 (N_3739,N_3616,N_3685);
xor U3740 (N_3740,N_3630,N_3612);
nand U3741 (N_3741,N_3675,N_3650);
and U3742 (N_3742,N_3653,N_3603);
nor U3743 (N_3743,N_3636,N_3609);
nand U3744 (N_3744,N_3693,N_3692);
or U3745 (N_3745,N_3642,N_3689);
nand U3746 (N_3746,N_3613,N_3633);
nor U3747 (N_3747,N_3678,N_3652);
nand U3748 (N_3748,N_3602,N_3625);
and U3749 (N_3749,N_3656,N_3623);
or U3750 (N_3750,N_3658,N_3666);
xor U3751 (N_3751,N_3695,N_3671);
and U3752 (N_3752,N_3626,N_3687);
or U3753 (N_3753,N_3609,N_3660);
xor U3754 (N_3754,N_3667,N_3673);
nand U3755 (N_3755,N_3621,N_3686);
or U3756 (N_3756,N_3619,N_3698);
xnor U3757 (N_3757,N_3693,N_3645);
nand U3758 (N_3758,N_3661,N_3671);
or U3759 (N_3759,N_3620,N_3651);
or U3760 (N_3760,N_3604,N_3680);
and U3761 (N_3761,N_3660,N_3617);
and U3762 (N_3762,N_3674,N_3692);
nor U3763 (N_3763,N_3601,N_3648);
nand U3764 (N_3764,N_3620,N_3691);
nor U3765 (N_3765,N_3672,N_3629);
xnor U3766 (N_3766,N_3682,N_3657);
and U3767 (N_3767,N_3695,N_3689);
xor U3768 (N_3768,N_3651,N_3602);
nand U3769 (N_3769,N_3642,N_3602);
nand U3770 (N_3770,N_3605,N_3637);
or U3771 (N_3771,N_3654,N_3628);
or U3772 (N_3772,N_3608,N_3669);
or U3773 (N_3773,N_3658,N_3640);
or U3774 (N_3774,N_3629,N_3675);
nor U3775 (N_3775,N_3637,N_3608);
nor U3776 (N_3776,N_3625,N_3671);
and U3777 (N_3777,N_3665,N_3695);
nor U3778 (N_3778,N_3682,N_3656);
and U3779 (N_3779,N_3665,N_3636);
nor U3780 (N_3780,N_3603,N_3617);
and U3781 (N_3781,N_3662,N_3601);
or U3782 (N_3782,N_3674,N_3655);
and U3783 (N_3783,N_3601,N_3630);
nand U3784 (N_3784,N_3689,N_3680);
or U3785 (N_3785,N_3657,N_3634);
or U3786 (N_3786,N_3657,N_3602);
and U3787 (N_3787,N_3660,N_3671);
nor U3788 (N_3788,N_3663,N_3641);
and U3789 (N_3789,N_3626,N_3605);
nor U3790 (N_3790,N_3643,N_3642);
nor U3791 (N_3791,N_3654,N_3649);
nand U3792 (N_3792,N_3617,N_3679);
nor U3793 (N_3793,N_3618,N_3651);
nor U3794 (N_3794,N_3679,N_3618);
and U3795 (N_3795,N_3613,N_3690);
or U3796 (N_3796,N_3661,N_3634);
or U3797 (N_3797,N_3608,N_3604);
nor U3798 (N_3798,N_3608,N_3652);
nor U3799 (N_3799,N_3663,N_3622);
xnor U3800 (N_3800,N_3720,N_3710);
or U3801 (N_3801,N_3725,N_3779);
or U3802 (N_3802,N_3756,N_3732);
xnor U3803 (N_3803,N_3711,N_3727);
nor U3804 (N_3804,N_3762,N_3731);
nor U3805 (N_3805,N_3778,N_3791);
nand U3806 (N_3806,N_3703,N_3726);
nor U3807 (N_3807,N_3713,N_3790);
nor U3808 (N_3808,N_3760,N_3772);
or U3809 (N_3809,N_3787,N_3723);
and U3810 (N_3810,N_3753,N_3741);
nor U3811 (N_3811,N_3748,N_3707);
nand U3812 (N_3812,N_3769,N_3767);
nor U3813 (N_3813,N_3724,N_3746);
nor U3814 (N_3814,N_3734,N_3783);
or U3815 (N_3815,N_3782,N_3708);
and U3816 (N_3816,N_3722,N_3754);
nor U3817 (N_3817,N_3792,N_3771);
or U3818 (N_3818,N_3757,N_3750);
or U3819 (N_3819,N_3752,N_3737);
or U3820 (N_3820,N_3793,N_3716);
nor U3821 (N_3821,N_3763,N_3788);
nor U3822 (N_3822,N_3701,N_3796);
nand U3823 (N_3823,N_3781,N_3758);
or U3824 (N_3824,N_3755,N_3797);
nand U3825 (N_3825,N_3728,N_3798);
nand U3826 (N_3826,N_3789,N_3706);
or U3827 (N_3827,N_3736,N_3774);
nor U3828 (N_3828,N_3744,N_3773);
and U3829 (N_3829,N_3738,N_3785);
xnor U3830 (N_3830,N_3761,N_3751);
xor U3831 (N_3831,N_3714,N_3733);
nand U3832 (N_3832,N_3730,N_3718);
xnor U3833 (N_3833,N_3799,N_3794);
and U3834 (N_3834,N_3780,N_3766);
or U3835 (N_3835,N_3759,N_3776);
or U3836 (N_3836,N_3775,N_3739);
nor U3837 (N_3837,N_3729,N_3719);
and U3838 (N_3838,N_3721,N_3704);
or U3839 (N_3839,N_3709,N_3735);
or U3840 (N_3840,N_3712,N_3743);
nor U3841 (N_3841,N_3777,N_3705);
and U3842 (N_3842,N_3740,N_3768);
nor U3843 (N_3843,N_3770,N_3749);
or U3844 (N_3844,N_3786,N_3784);
or U3845 (N_3845,N_3745,N_3702);
or U3846 (N_3846,N_3717,N_3715);
or U3847 (N_3847,N_3700,N_3742);
xnor U3848 (N_3848,N_3795,N_3747);
and U3849 (N_3849,N_3764,N_3765);
or U3850 (N_3850,N_3790,N_3740);
or U3851 (N_3851,N_3706,N_3785);
xnor U3852 (N_3852,N_3797,N_3779);
nand U3853 (N_3853,N_3726,N_3788);
nor U3854 (N_3854,N_3765,N_3753);
or U3855 (N_3855,N_3758,N_3796);
and U3856 (N_3856,N_3741,N_3750);
nand U3857 (N_3857,N_3752,N_3743);
or U3858 (N_3858,N_3778,N_3720);
nor U3859 (N_3859,N_3765,N_3715);
and U3860 (N_3860,N_3761,N_3748);
nor U3861 (N_3861,N_3726,N_3708);
and U3862 (N_3862,N_3711,N_3766);
nand U3863 (N_3863,N_3726,N_3798);
nand U3864 (N_3864,N_3778,N_3710);
and U3865 (N_3865,N_3776,N_3725);
or U3866 (N_3866,N_3778,N_3746);
nand U3867 (N_3867,N_3732,N_3779);
xor U3868 (N_3868,N_3760,N_3747);
and U3869 (N_3869,N_3734,N_3709);
and U3870 (N_3870,N_3788,N_3724);
nand U3871 (N_3871,N_3776,N_3737);
nand U3872 (N_3872,N_3770,N_3771);
and U3873 (N_3873,N_3731,N_3733);
nor U3874 (N_3874,N_3739,N_3710);
nor U3875 (N_3875,N_3743,N_3751);
and U3876 (N_3876,N_3719,N_3733);
nand U3877 (N_3877,N_3789,N_3781);
xnor U3878 (N_3878,N_3794,N_3792);
nor U3879 (N_3879,N_3766,N_3770);
xnor U3880 (N_3880,N_3723,N_3755);
nand U3881 (N_3881,N_3721,N_3712);
or U3882 (N_3882,N_3744,N_3722);
or U3883 (N_3883,N_3718,N_3762);
and U3884 (N_3884,N_3711,N_3709);
nor U3885 (N_3885,N_3759,N_3754);
or U3886 (N_3886,N_3730,N_3773);
or U3887 (N_3887,N_3764,N_3756);
and U3888 (N_3888,N_3784,N_3750);
nand U3889 (N_3889,N_3710,N_3786);
nor U3890 (N_3890,N_3719,N_3766);
and U3891 (N_3891,N_3719,N_3736);
and U3892 (N_3892,N_3760,N_3725);
and U3893 (N_3893,N_3709,N_3730);
nand U3894 (N_3894,N_3771,N_3723);
nand U3895 (N_3895,N_3701,N_3767);
nor U3896 (N_3896,N_3729,N_3783);
nor U3897 (N_3897,N_3794,N_3798);
and U3898 (N_3898,N_3755,N_3745);
nor U3899 (N_3899,N_3702,N_3730);
or U3900 (N_3900,N_3899,N_3859);
or U3901 (N_3901,N_3841,N_3862);
nor U3902 (N_3902,N_3845,N_3893);
xnor U3903 (N_3903,N_3833,N_3851);
nor U3904 (N_3904,N_3805,N_3882);
nor U3905 (N_3905,N_3883,N_3807);
nand U3906 (N_3906,N_3829,N_3891);
or U3907 (N_3907,N_3898,N_3846);
nand U3908 (N_3908,N_3885,N_3808);
xnor U3909 (N_3909,N_3861,N_3894);
and U3910 (N_3910,N_3800,N_3848);
nor U3911 (N_3911,N_3880,N_3872);
and U3912 (N_3912,N_3876,N_3804);
nor U3913 (N_3913,N_3860,N_3813);
and U3914 (N_3914,N_3884,N_3812);
nor U3915 (N_3915,N_3896,N_3875);
nor U3916 (N_3916,N_3867,N_3881);
nor U3917 (N_3917,N_3887,N_3895);
nor U3918 (N_3918,N_3834,N_3821);
and U3919 (N_3919,N_3826,N_3811);
nor U3920 (N_3920,N_3858,N_3822);
or U3921 (N_3921,N_3863,N_3879);
and U3922 (N_3922,N_3886,N_3832);
or U3923 (N_3923,N_3809,N_3823);
and U3924 (N_3924,N_3870,N_3803);
nor U3925 (N_3925,N_3869,N_3877);
xnor U3926 (N_3926,N_3853,N_3854);
or U3927 (N_3927,N_3888,N_3844);
and U3928 (N_3928,N_3878,N_3892);
nand U3929 (N_3929,N_3868,N_3847);
and U3930 (N_3930,N_3857,N_3818);
nand U3931 (N_3931,N_3897,N_3825);
nand U3932 (N_3932,N_3856,N_3842);
nand U3933 (N_3933,N_3839,N_3850);
and U3934 (N_3934,N_3838,N_3816);
nand U3935 (N_3935,N_3830,N_3843);
and U3936 (N_3936,N_3815,N_3840);
nor U3937 (N_3937,N_3819,N_3866);
xor U3938 (N_3938,N_3873,N_3864);
nand U3939 (N_3939,N_3837,N_3836);
nand U3940 (N_3940,N_3874,N_3814);
xnor U3941 (N_3941,N_3827,N_3831);
nand U3942 (N_3942,N_3865,N_3890);
nand U3943 (N_3943,N_3855,N_3889);
nand U3944 (N_3944,N_3835,N_3817);
and U3945 (N_3945,N_3871,N_3802);
or U3946 (N_3946,N_3806,N_3849);
xor U3947 (N_3947,N_3824,N_3852);
nor U3948 (N_3948,N_3820,N_3810);
xnor U3949 (N_3949,N_3801,N_3828);
or U3950 (N_3950,N_3835,N_3850);
or U3951 (N_3951,N_3817,N_3826);
nand U3952 (N_3952,N_3838,N_3899);
or U3953 (N_3953,N_3808,N_3803);
nand U3954 (N_3954,N_3838,N_3889);
and U3955 (N_3955,N_3846,N_3889);
nand U3956 (N_3956,N_3867,N_3847);
xor U3957 (N_3957,N_3859,N_3882);
nor U3958 (N_3958,N_3826,N_3878);
and U3959 (N_3959,N_3823,N_3859);
and U3960 (N_3960,N_3875,N_3891);
xor U3961 (N_3961,N_3854,N_3807);
nor U3962 (N_3962,N_3899,N_3892);
nand U3963 (N_3963,N_3883,N_3895);
nand U3964 (N_3964,N_3857,N_3864);
nand U3965 (N_3965,N_3857,N_3860);
nor U3966 (N_3966,N_3851,N_3887);
nor U3967 (N_3967,N_3862,N_3874);
or U3968 (N_3968,N_3852,N_3808);
or U3969 (N_3969,N_3804,N_3892);
and U3970 (N_3970,N_3880,N_3831);
and U3971 (N_3971,N_3849,N_3811);
nand U3972 (N_3972,N_3895,N_3808);
xor U3973 (N_3973,N_3827,N_3866);
nand U3974 (N_3974,N_3845,N_3853);
xnor U3975 (N_3975,N_3862,N_3843);
nor U3976 (N_3976,N_3815,N_3871);
nand U3977 (N_3977,N_3869,N_3863);
and U3978 (N_3978,N_3847,N_3842);
or U3979 (N_3979,N_3894,N_3823);
and U3980 (N_3980,N_3882,N_3842);
and U3981 (N_3981,N_3833,N_3829);
or U3982 (N_3982,N_3836,N_3858);
or U3983 (N_3983,N_3877,N_3855);
and U3984 (N_3984,N_3898,N_3840);
xor U3985 (N_3985,N_3807,N_3891);
or U3986 (N_3986,N_3804,N_3808);
nor U3987 (N_3987,N_3898,N_3829);
nand U3988 (N_3988,N_3839,N_3803);
nand U3989 (N_3989,N_3851,N_3824);
nand U3990 (N_3990,N_3825,N_3814);
or U3991 (N_3991,N_3856,N_3827);
or U3992 (N_3992,N_3843,N_3859);
nor U3993 (N_3993,N_3803,N_3898);
nand U3994 (N_3994,N_3848,N_3896);
nor U3995 (N_3995,N_3862,N_3866);
nand U3996 (N_3996,N_3876,N_3800);
nand U3997 (N_3997,N_3885,N_3835);
xor U3998 (N_3998,N_3823,N_3879);
nand U3999 (N_3999,N_3845,N_3877);
and U4000 (N_4000,N_3901,N_3982);
nand U4001 (N_4001,N_3912,N_3972);
and U4002 (N_4002,N_3962,N_3914);
or U4003 (N_4003,N_3963,N_3910);
nor U4004 (N_4004,N_3934,N_3965);
nand U4005 (N_4005,N_3942,N_3992);
nand U4006 (N_4006,N_3954,N_3955);
and U4007 (N_4007,N_3978,N_3967);
nand U4008 (N_4008,N_3921,N_3998);
or U4009 (N_4009,N_3986,N_3930);
nand U4010 (N_4010,N_3993,N_3902);
and U4011 (N_4011,N_3996,N_3915);
or U4012 (N_4012,N_3995,N_3935);
nand U4013 (N_4013,N_3943,N_3984);
and U4014 (N_4014,N_3991,N_3939);
nor U4015 (N_4015,N_3957,N_3906);
nand U4016 (N_4016,N_3948,N_3961);
and U4017 (N_4017,N_3927,N_3917);
and U4018 (N_4018,N_3908,N_3913);
nand U4019 (N_4019,N_3987,N_3969);
nor U4020 (N_4020,N_3966,N_3973);
nand U4021 (N_4021,N_3924,N_3960);
nor U4022 (N_4022,N_3916,N_3947);
nor U4023 (N_4023,N_3980,N_3907);
or U4024 (N_4024,N_3900,N_3951);
nand U4025 (N_4025,N_3926,N_3911);
nand U4026 (N_4026,N_3958,N_3971);
or U4027 (N_4027,N_3952,N_3909);
xnor U4028 (N_4028,N_3929,N_3983);
or U4029 (N_4029,N_3933,N_3985);
xor U4030 (N_4030,N_3932,N_3928);
or U4031 (N_4031,N_3981,N_3977);
or U4032 (N_4032,N_3936,N_3944);
nor U4033 (N_4033,N_3968,N_3923);
and U4034 (N_4034,N_3905,N_3979);
and U4035 (N_4035,N_3903,N_3959);
nor U4036 (N_4036,N_3904,N_3946);
nand U4037 (N_4037,N_3999,N_3920);
and U4038 (N_4038,N_3945,N_3974);
and U4039 (N_4039,N_3997,N_3931);
nand U4040 (N_4040,N_3919,N_3956);
or U4041 (N_4041,N_3976,N_3950);
nor U4042 (N_4042,N_3937,N_3940);
nor U4043 (N_4043,N_3988,N_3964);
nor U4044 (N_4044,N_3925,N_3990);
nand U4045 (N_4045,N_3938,N_3994);
nor U4046 (N_4046,N_3918,N_3953);
or U4047 (N_4047,N_3922,N_3975);
xnor U4048 (N_4048,N_3989,N_3970);
and U4049 (N_4049,N_3949,N_3941);
nor U4050 (N_4050,N_3940,N_3995);
nand U4051 (N_4051,N_3943,N_3925);
or U4052 (N_4052,N_3998,N_3980);
nand U4053 (N_4053,N_3938,N_3992);
and U4054 (N_4054,N_3954,N_3993);
and U4055 (N_4055,N_3949,N_3947);
nor U4056 (N_4056,N_3962,N_3937);
nor U4057 (N_4057,N_3911,N_3952);
and U4058 (N_4058,N_3902,N_3937);
or U4059 (N_4059,N_3902,N_3970);
nor U4060 (N_4060,N_3917,N_3920);
nor U4061 (N_4061,N_3914,N_3948);
xnor U4062 (N_4062,N_3932,N_3938);
nand U4063 (N_4063,N_3928,N_3941);
nand U4064 (N_4064,N_3994,N_3941);
nand U4065 (N_4065,N_3908,N_3904);
nand U4066 (N_4066,N_3932,N_3900);
or U4067 (N_4067,N_3902,N_3947);
nand U4068 (N_4068,N_3976,N_3961);
nor U4069 (N_4069,N_3917,N_3995);
and U4070 (N_4070,N_3932,N_3912);
nand U4071 (N_4071,N_3922,N_3942);
and U4072 (N_4072,N_3970,N_3923);
nor U4073 (N_4073,N_3985,N_3927);
or U4074 (N_4074,N_3931,N_3967);
and U4075 (N_4075,N_3918,N_3911);
nand U4076 (N_4076,N_3954,N_3994);
nand U4077 (N_4077,N_3929,N_3984);
nor U4078 (N_4078,N_3964,N_3921);
nand U4079 (N_4079,N_3900,N_3954);
nand U4080 (N_4080,N_3905,N_3993);
nor U4081 (N_4081,N_3985,N_3981);
and U4082 (N_4082,N_3983,N_3911);
and U4083 (N_4083,N_3944,N_3903);
nand U4084 (N_4084,N_3991,N_3910);
or U4085 (N_4085,N_3968,N_3986);
nor U4086 (N_4086,N_3995,N_3928);
or U4087 (N_4087,N_3965,N_3932);
nand U4088 (N_4088,N_3927,N_3990);
or U4089 (N_4089,N_3903,N_3965);
nor U4090 (N_4090,N_3937,N_3975);
and U4091 (N_4091,N_3980,N_3975);
and U4092 (N_4092,N_3952,N_3944);
or U4093 (N_4093,N_3955,N_3904);
nand U4094 (N_4094,N_3905,N_3942);
nor U4095 (N_4095,N_3994,N_3980);
xor U4096 (N_4096,N_3903,N_3983);
nor U4097 (N_4097,N_3934,N_3954);
or U4098 (N_4098,N_3907,N_3922);
and U4099 (N_4099,N_3957,N_3932);
and U4100 (N_4100,N_4012,N_4028);
nor U4101 (N_4101,N_4070,N_4062);
nor U4102 (N_4102,N_4069,N_4014);
or U4103 (N_4103,N_4046,N_4043);
xor U4104 (N_4104,N_4082,N_4018);
or U4105 (N_4105,N_4057,N_4021);
xor U4106 (N_4106,N_4017,N_4020);
and U4107 (N_4107,N_4010,N_4047);
or U4108 (N_4108,N_4077,N_4097);
and U4109 (N_4109,N_4038,N_4023);
or U4110 (N_4110,N_4074,N_4004);
nand U4111 (N_4111,N_4048,N_4024);
or U4112 (N_4112,N_4054,N_4040);
xnor U4113 (N_4113,N_4005,N_4049);
and U4114 (N_4114,N_4085,N_4008);
nand U4115 (N_4115,N_4051,N_4090);
and U4116 (N_4116,N_4011,N_4019);
nand U4117 (N_4117,N_4061,N_4079);
nor U4118 (N_4118,N_4083,N_4032);
or U4119 (N_4119,N_4072,N_4081);
nand U4120 (N_4120,N_4063,N_4068);
and U4121 (N_4121,N_4089,N_4071);
nand U4122 (N_4122,N_4003,N_4033);
nor U4123 (N_4123,N_4001,N_4073);
nand U4124 (N_4124,N_4042,N_4025);
nand U4125 (N_4125,N_4029,N_4094);
xnor U4126 (N_4126,N_4060,N_4098);
nand U4127 (N_4127,N_4045,N_4092);
and U4128 (N_4128,N_4053,N_4075);
or U4129 (N_4129,N_4056,N_4000);
nand U4130 (N_4130,N_4067,N_4086);
and U4131 (N_4131,N_4091,N_4055);
xnor U4132 (N_4132,N_4022,N_4093);
nand U4133 (N_4133,N_4084,N_4044);
nor U4134 (N_4134,N_4076,N_4095);
or U4135 (N_4135,N_4065,N_4099);
xnor U4136 (N_4136,N_4016,N_4006);
xnor U4137 (N_4137,N_4041,N_4013);
or U4138 (N_4138,N_4080,N_4007);
nor U4139 (N_4139,N_4096,N_4087);
or U4140 (N_4140,N_4009,N_4027);
xor U4141 (N_4141,N_4036,N_4052);
and U4142 (N_4142,N_4088,N_4078);
or U4143 (N_4143,N_4030,N_4039);
nand U4144 (N_4144,N_4050,N_4058);
nor U4145 (N_4145,N_4037,N_4031);
nor U4146 (N_4146,N_4026,N_4059);
nor U4147 (N_4147,N_4034,N_4015);
and U4148 (N_4148,N_4035,N_4002);
or U4149 (N_4149,N_4064,N_4066);
and U4150 (N_4150,N_4008,N_4091);
nor U4151 (N_4151,N_4019,N_4088);
or U4152 (N_4152,N_4066,N_4091);
xor U4153 (N_4153,N_4070,N_4059);
and U4154 (N_4154,N_4072,N_4069);
and U4155 (N_4155,N_4079,N_4059);
or U4156 (N_4156,N_4081,N_4083);
nand U4157 (N_4157,N_4064,N_4080);
nor U4158 (N_4158,N_4077,N_4036);
and U4159 (N_4159,N_4089,N_4005);
nand U4160 (N_4160,N_4053,N_4066);
xor U4161 (N_4161,N_4083,N_4045);
nand U4162 (N_4162,N_4093,N_4024);
nand U4163 (N_4163,N_4085,N_4020);
nand U4164 (N_4164,N_4048,N_4041);
and U4165 (N_4165,N_4075,N_4008);
nor U4166 (N_4166,N_4063,N_4005);
nand U4167 (N_4167,N_4068,N_4099);
nor U4168 (N_4168,N_4098,N_4009);
and U4169 (N_4169,N_4033,N_4034);
nand U4170 (N_4170,N_4055,N_4033);
xor U4171 (N_4171,N_4050,N_4080);
xor U4172 (N_4172,N_4003,N_4023);
or U4173 (N_4173,N_4069,N_4071);
or U4174 (N_4174,N_4029,N_4064);
or U4175 (N_4175,N_4069,N_4068);
nor U4176 (N_4176,N_4065,N_4003);
and U4177 (N_4177,N_4029,N_4077);
nand U4178 (N_4178,N_4033,N_4071);
nand U4179 (N_4179,N_4017,N_4050);
or U4180 (N_4180,N_4072,N_4082);
xor U4181 (N_4181,N_4079,N_4087);
or U4182 (N_4182,N_4000,N_4029);
nor U4183 (N_4183,N_4064,N_4020);
nand U4184 (N_4184,N_4001,N_4057);
nand U4185 (N_4185,N_4014,N_4055);
or U4186 (N_4186,N_4059,N_4061);
nor U4187 (N_4187,N_4070,N_4060);
nor U4188 (N_4188,N_4017,N_4038);
and U4189 (N_4189,N_4081,N_4061);
xnor U4190 (N_4190,N_4018,N_4031);
nand U4191 (N_4191,N_4046,N_4036);
nor U4192 (N_4192,N_4031,N_4069);
xor U4193 (N_4193,N_4073,N_4058);
or U4194 (N_4194,N_4001,N_4090);
nand U4195 (N_4195,N_4044,N_4042);
nor U4196 (N_4196,N_4074,N_4046);
and U4197 (N_4197,N_4002,N_4060);
or U4198 (N_4198,N_4055,N_4093);
xnor U4199 (N_4199,N_4045,N_4004);
and U4200 (N_4200,N_4140,N_4103);
or U4201 (N_4201,N_4178,N_4139);
nor U4202 (N_4202,N_4104,N_4157);
nor U4203 (N_4203,N_4134,N_4102);
nor U4204 (N_4204,N_4137,N_4154);
nand U4205 (N_4205,N_4177,N_4106);
nor U4206 (N_4206,N_4151,N_4182);
nor U4207 (N_4207,N_4181,N_4145);
nor U4208 (N_4208,N_4163,N_4166);
nand U4209 (N_4209,N_4171,N_4195);
xnor U4210 (N_4210,N_4185,N_4127);
nand U4211 (N_4211,N_4101,N_4125);
nand U4212 (N_4212,N_4161,N_4190);
nand U4213 (N_4213,N_4188,N_4148);
nand U4214 (N_4214,N_4122,N_4194);
nand U4215 (N_4215,N_4120,N_4119);
and U4216 (N_4216,N_4128,N_4158);
or U4217 (N_4217,N_4193,N_4117);
nand U4218 (N_4218,N_4116,N_4143);
or U4219 (N_4219,N_4180,N_4115);
nor U4220 (N_4220,N_4108,N_4149);
or U4221 (N_4221,N_4100,N_4113);
nand U4222 (N_4222,N_4136,N_4187);
nand U4223 (N_4223,N_4138,N_4150);
and U4224 (N_4224,N_4162,N_4141);
or U4225 (N_4225,N_4179,N_4105);
nand U4226 (N_4226,N_4114,N_4198);
and U4227 (N_4227,N_4169,N_4152);
nand U4228 (N_4228,N_4155,N_4153);
xnor U4229 (N_4229,N_4191,N_4111);
and U4230 (N_4230,N_4167,N_4110);
or U4231 (N_4231,N_4196,N_4121);
nand U4232 (N_4232,N_4170,N_4147);
xnor U4233 (N_4233,N_4186,N_4164);
and U4234 (N_4234,N_4146,N_4129);
nor U4235 (N_4235,N_4183,N_4197);
xor U4236 (N_4236,N_4130,N_4172);
nand U4237 (N_4237,N_4173,N_4144);
nand U4238 (N_4238,N_4107,N_4156);
xor U4239 (N_4239,N_4123,N_4131);
or U4240 (N_4240,N_4135,N_4174);
nand U4241 (N_4241,N_4168,N_4199);
or U4242 (N_4242,N_4175,N_4142);
nor U4243 (N_4243,N_4126,N_4124);
and U4244 (N_4244,N_4159,N_4184);
or U4245 (N_4245,N_4189,N_4133);
nor U4246 (N_4246,N_4132,N_4109);
nand U4247 (N_4247,N_4160,N_4112);
nand U4248 (N_4248,N_4165,N_4176);
xor U4249 (N_4249,N_4192,N_4118);
xnor U4250 (N_4250,N_4126,N_4112);
and U4251 (N_4251,N_4119,N_4106);
and U4252 (N_4252,N_4121,N_4158);
nor U4253 (N_4253,N_4134,N_4175);
and U4254 (N_4254,N_4198,N_4103);
or U4255 (N_4255,N_4168,N_4116);
and U4256 (N_4256,N_4176,N_4108);
nand U4257 (N_4257,N_4132,N_4196);
nand U4258 (N_4258,N_4111,N_4123);
nand U4259 (N_4259,N_4187,N_4169);
nand U4260 (N_4260,N_4135,N_4104);
or U4261 (N_4261,N_4153,N_4125);
and U4262 (N_4262,N_4185,N_4163);
xor U4263 (N_4263,N_4129,N_4183);
nor U4264 (N_4264,N_4176,N_4173);
nand U4265 (N_4265,N_4173,N_4179);
or U4266 (N_4266,N_4101,N_4155);
or U4267 (N_4267,N_4145,N_4118);
or U4268 (N_4268,N_4103,N_4127);
or U4269 (N_4269,N_4126,N_4160);
nand U4270 (N_4270,N_4195,N_4149);
nor U4271 (N_4271,N_4136,N_4170);
or U4272 (N_4272,N_4103,N_4171);
nand U4273 (N_4273,N_4157,N_4141);
nand U4274 (N_4274,N_4110,N_4185);
nand U4275 (N_4275,N_4144,N_4145);
and U4276 (N_4276,N_4190,N_4102);
and U4277 (N_4277,N_4103,N_4146);
nand U4278 (N_4278,N_4141,N_4136);
nor U4279 (N_4279,N_4193,N_4181);
nor U4280 (N_4280,N_4109,N_4173);
nand U4281 (N_4281,N_4191,N_4101);
nand U4282 (N_4282,N_4166,N_4199);
xnor U4283 (N_4283,N_4179,N_4115);
nor U4284 (N_4284,N_4113,N_4126);
nand U4285 (N_4285,N_4165,N_4156);
or U4286 (N_4286,N_4196,N_4150);
or U4287 (N_4287,N_4131,N_4166);
nor U4288 (N_4288,N_4127,N_4187);
nand U4289 (N_4289,N_4172,N_4163);
or U4290 (N_4290,N_4174,N_4192);
nand U4291 (N_4291,N_4194,N_4179);
nor U4292 (N_4292,N_4120,N_4196);
nor U4293 (N_4293,N_4145,N_4170);
nor U4294 (N_4294,N_4156,N_4184);
or U4295 (N_4295,N_4124,N_4181);
nor U4296 (N_4296,N_4181,N_4195);
xnor U4297 (N_4297,N_4148,N_4163);
nor U4298 (N_4298,N_4182,N_4187);
and U4299 (N_4299,N_4124,N_4152);
or U4300 (N_4300,N_4257,N_4223);
or U4301 (N_4301,N_4261,N_4265);
and U4302 (N_4302,N_4268,N_4273);
or U4303 (N_4303,N_4240,N_4216);
or U4304 (N_4304,N_4299,N_4276);
nor U4305 (N_4305,N_4245,N_4266);
and U4306 (N_4306,N_4281,N_4292);
and U4307 (N_4307,N_4231,N_4278);
nand U4308 (N_4308,N_4235,N_4252);
nor U4309 (N_4309,N_4255,N_4230);
or U4310 (N_4310,N_4237,N_4225);
nand U4311 (N_4311,N_4286,N_4229);
nand U4312 (N_4312,N_4226,N_4213);
or U4313 (N_4313,N_4205,N_4274);
nor U4314 (N_4314,N_4247,N_4239);
xnor U4315 (N_4315,N_4290,N_4233);
nand U4316 (N_4316,N_4207,N_4296);
and U4317 (N_4317,N_4267,N_4293);
nand U4318 (N_4318,N_4297,N_4287);
nor U4319 (N_4319,N_4218,N_4220);
and U4320 (N_4320,N_4241,N_4275);
and U4321 (N_4321,N_4206,N_4242);
nor U4322 (N_4322,N_4211,N_4272);
nand U4323 (N_4323,N_4217,N_4298);
and U4324 (N_4324,N_4219,N_4262);
nor U4325 (N_4325,N_4244,N_4250);
or U4326 (N_4326,N_4212,N_4284);
or U4327 (N_4327,N_4282,N_4283);
and U4328 (N_4328,N_4289,N_4263);
or U4329 (N_4329,N_4285,N_4234);
xnor U4330 (N_4330,N_4248,N_4258);
xnor U4331 (N_4331,N_4204,N_4200);
nor U4332 (N_4332,N_4201,N_4254);
nand U4333 (N_4333,N_4202,N_4221);
nand U4334 (N_4334,N_4222,N_4259);
or U4335 (N_4335,N_4214,N_4277);
or U4336 (N_4336,N_4288,N_4294);
nand U4337 (N_4337,N_4215,N_4228);
nor U4338 (N_4338,N_4227,N_4208);
and U4339 (N_4339,N_4256,N_4246);
nand U4340 (N_4340,N_4236,N_4271);
xor U4341 (N_4341,N_4269,N_4251);
and U4342 (N_4342,N_4249,N_4295);
and U4343 (N_4343,N_4291,N_4260);
nor U4344 (N_4344,N_4232,N_4264);
or U4345 (N_4345,N_4238,N_4280);
nand U4346 (N_4346,N_4270,N_4209);
nand U4347 (N_4347,N_4210,N_4253);
nor U4348 (N_4348,N_4243,N_4203);
or U4349 (N_4349,N_4279,N_4224);
nor U4350 (N_4350,N_4287,N_4241);
and U4351 (N_4351,N_4272,N_4283);
and U4352 (N_4352,N_4208,N_4278);
nand U4353 (N_4353,N_4264,N_4206);
and U4354 (N_4354,N_4299,N_4274);
nand U4355 (N_4355,N_4204,N_4268);
nor U4356 (N_4356,N_4208,N_4265);
nand U4357 (N_4357,N_4287,N_4207);
and U4358 (N_4358,N_4248,N_4200);
and U4359 (N_4359,N_4280,N_4278);
or U4360 (N_4360,N_4247,N_4275);
nand U4361 (N_4361,N_4260,N_4289);
xor U4362 (N_4362,N_4210,N_4268);
nand U4363 (N_4363,N_4292,N_4202);
nor U4364 (N_4364,N_4271,N_4240);
or U4365 (N_4365,N_4293,N_4231);
nor U4366 (N_4366,N_4220,N_4285);
or U4367 (N_4367,N_4291,N_4249);
nor U4368 (N_4368,N_4225,N_4271);
nand U4369 (N_4369,N_4261,N_4226);
nor U4370 (N_4370,N_4272,N_4234);
xor U4371 (N_4371,N_4237,N_4200);
or U4372 (N_4372,N_4212,N_4249);
xor U4373 (N_4373,N_4259,N_4267);
xor U4374 (N_4374,N_4207,N_4242);
xnor U4375 (N_4375,N_4242,N_4246);
or U4376 (N_4376,N_4239,N_4234);
nor U4377 (N_4377,N_4230,N_4278);
or U4378 (N_4378,N_4211,N_4253);
nand U4379 (N_4379,N_4217,N_4200);
nor U4380 (N_4380,N_4285,N_4224);
or U4381 (N_4381,N_4295,N_4204);
or U4382 (N_4382,N_4257,N_4284);
nand U4383 (N_4383,N_4295,N_4262);
nor U4384 (N_4384,N_4239,N_4206);
nor U4385 (N_4385,N_4222,N_4231);
and U4386 (N_4386,N_4277,N_4257);
or U4387 (N_4387,N_4251,N_4295);
xor U4388 (N_4388,N_4244,N_4222);
nor U4389 (N_4389,N_4278,N_4279);
and U4390 (N_4390,N_4271,N_4245);
nand U4391 (N_4391,N_4290,N_4200);
nor U4392 (N_4392,N_4211,N_4208);
nor U4393 (N_4393,N_4278,N_4284);
or U4394 (N_4394,N_4293,N_4265);
nor U4395 (N_4395,N_4296,N_4287);
or U4396 (N_4396,N_4271,N_4272);
or U4397 (N_4397,N_4293,N_4219);
nor U4398 (N_4398,N_4266,N_4240);
and U4399 (N_4399,N_4207,N_4201);
nor U4400 (N_4400,N_4378,N_4344);
xnor U4401 (N_4401,N_4342,N_4396);
xor U4402 (N_4402,N_4386,N_4300);
and U4403 (N_4403,N_4307,N_4366);
and U4404 (N_4404,N_4336,N_4348);
nor U4405 (N_4405,N_4347,N_4355);
and U4406 (N_4406,N_4365,N_4397);
nand U4407 (N_4407,N_4334,N_4343);
xnor U4408 (N_4408,N_4353,N_4338);
or U4409 (N_4409,N_4323,N_4318);
xnor U4410 (N_4410,N_4398,N_4305);
nand U4411 (N_4411,N_4322,N_4390);
or U4412 (N_4412,N_4327,N_4309);
nor U4413 (N_4413,N_4316,N_4384);
nor U4414 (N_4414,N_4364,N_4359);
or U4415 (N_4415,N_4380,N_4360);
and U4416 (N_4416,N_4394,N_4377);
and U4417 (N_4417,N_4385,N_4381);
or U4418 (N_4418,N_4361,N_4310);
or U4419 (N_4419,N_4350,N_4326);
or U4420 (N_4420,N_4363,N_4339);
and U4421 (N_4421,N_4371,N_4328);
nor U4422 (N_4422,N_4372,N_4399);
nor U4423 (N_4423,N_4304,N_4331);
and U4424 (N_4424,N_4302,N_4356);
nand U4425 (N_4425,N_4374,N_4352);
nor U4426 (N_4426,N_4354,N_4325);
nand U4427 (N_4427,N_4392,N_4312);
or U4428 (N_4428,N_4324,N_4341);
nand U4429 (N_4429,N_4345,N_4335);
and U4430 (N_4430,N_4329,N_4391);
xnor U4431 (N_4431,N_4311,N_4373);
or U4432 (N_4432,N_4370,N_4301);
or U4433 (N_4433,N_4349,N_4308);
and U4434 (N_4434,N_4340,N_4314);
nor U4435 (N_4435,N_4382,N_4303);
xor U4436 (N_4436,N_4393,N_4306);
xor U4437 (N_4437,N_4351,N_4337);
or U4438 (N_4438,N_4321,N_4387);
nand U4439 (N_4439,N_4333,N_4379);
xor U4440 (N_4440,N_4315,N_4346);
nand U4441 (N_4441,N_4317,N_4395);
nor U4442 (N_4442,N_4368,N_4362);
and U4443 (N_4443,N_4313,N_4319);
or U4444 (N_4444,N_4376,N_4389);
xnor U4445 (N_4445,N_4375,N_4330);
nand U4446 (N_4446,N_4320,N_4383);
or U4447 (N_4447,N_4388,N_4357);
or U4448 (N_4448,N_4332,N_4367);
and U4449 (N_4449,N_4358,N_4369);
and U4450 (N_4450,N_4334,N_4303);
nor U4451 (N_4451,N_4336,N_4381);
nor U4452 (N_4452,N_4345,N_4369);
and U4453 (N_4453,N_4340,N_4331);
nor U4454 (N_4454,N_4358,N_4356);
and U4455 (N_4455,N_4387,N_4302);
or U4456 (N_4456,N_4383,N_4378);
and U4457 (N_4457,N_4320,N_4398);
nor U4458 (N_4458,N_4360,N_4376);
or U4459 (N_4459,N_4338,N_4371);
or U4460 (N_4460,N_4366,N_4340);
xnor U4461 (N_4461,N_4369,N_4352);
and U4462 (N_4462,N_4363,N_4374);
nand U4463 (N_4463,N_4373,N_4381);
nand U4464 (N_4464,N_4304,N_4357);
and U4465 (N_4465,N_4311,N_4328);
xnor U4466 (N_4466,N_4377,N_4348);
nor U4467 (N_4467,N_4368,N_4317);
nor U4468 (N_4468,N_4314,N_4348);
xnor U4469 (N_4469,N_4329,N_4381);
nand U4470 (N_4470,N_4313,N_4352);
or U4471 (N_4471,N_4374,N_4306);
nand U4472 (N_4472,N_4361,N_4332);
nor U4473 (N_4473,N_4305,N_4372);
nand U4474 (N_4474,N_4300,N_4308);
xnor U4475 (N_4475,N_4329,N_4399);
or U4476 (N_4476,N_4345,N_4381);
and U4477 (N_4477,N_4372,N_4303);
nand U4478 (N_4478,N_4392,N_4379);
xor U4479 (N_4479,N_4390,N_4347);
nor U4480 (N_4480,N_4339,N_4367);
or U4481 (N_4481,N_4346,N_4382);
and U4482 (N_4482,N_4366,N_4371);
xor U4483 (N_4483,N_4347,N_4362);
or U4484 (N_4484,N_4370,N_4356);
nor U4485 (N_4485,N_4329,N_4303);
nor U4486 (N_4486,N_4378,N_4390);
nor U4487 (N_4487,N_4360,N_4352);
nand U4488 (N_4488,N_4308,N_4344);
nand U4489 (N_4489,N_4374,N_4329);
and U4490 (N_4490,N_4349,N_4374);
nand U4491 (N_4491,N_4391,N_4360);
xor U4492 (N_4492,N_4345,N_4365);
xor U4493 (N_4493,N_4331,N_4333);
nor U4494 (N_4494,N_4376,N_4351);
nand U4495 (N_4495,N_4382,N_4356);
xor U4496 (N_4496,N_4325,N_4345);
and U4497 (N_4497,N_4324,N_4300);
and U4498 (N_4498,N_4386,N_4355);
and U4499 (N_4499,N_4302,N_4357);
or U4500 (N_4500,N_4429,N_4434);
or U4501 (N_4501,N_4406,N_4475);
or U4502 (N_4502,N_4454,N_4435);
nand U4503 (N_4503,N_4413,N_4414);
or U4504 (N_4504,N_4415,N_4467);
xor U4505 (N_4505,N_4469,N_4478);
and U4506 (N_4506,N_4452,N_4444);
or U4507 (N_4507,N_4411,N_4439);
and U4508 (N_4508,N_4459,N_4422);
or U4509 (N_4509,N_4492,N_4497);
or U4510 (N_4510,N_4450,N_4499);
and U4511 (N_4511,N_4448,N_4440);
nand U4512 (N_4512,N_4479,N_4419);
or U4513 (N_4513,N_4460,N_4409);
nand U4514 (N_4514,N_4480,N_4437);
nand U4515 (N_4515,N_4423,N_4484);
or U4516 (N_4516,N_4436,N_4490);
and U4517 (N_4517,N_4445,N_4446);
and U4518 (N_4518,N_4416,N_4493);
or U4519 (N_4519,N_4491,N_4458);
and U4520 (N_4520,N_4482,N_4468);
nand U4521 (N_4521,N_4453,N_4473);
nand U4522 (N_4522,N_4485,N_4489);
or U4523 (N_4523,N_4412,N_4476);
and U4524 (N_4524,N_4403,N_4471);
xnor U4525 (N_4525,N_4494,N_4451);
or U4526 (N_4526,N_4456,N_4466);
nand U4527 (N_4527,N_4470,N_4400);
or U4528 (N_4528,N_4421,N_4427);
nor U4529 (N_4529,N_4463,N_4426);
nand U4530 (N_4530,N_4410,N_4474);
or U4531 (N_4531,N_4402,N_4495);
and U4532 (N_4532,N_4449,N_4465);
nor U4533 (N_4533,N_4404,N_4498);
xnor U4534 (N_4534,N_4418,N_4462);
or U4535 (N_4535,N_4447,N_4438);
and U4536 (N_4536,N_4408,N_4483);
or U4537 (N_4537,N_4428,N_4441);
nor U4538 (N_4538,N_4420,N_4481);
nand U4539 (N_4539,N_4425,N_4432);
and U4540 (N_4540,N_4488,N_4496);
xnor U4541 (N_4541,N_4442,N_4443);
nor U4542 (N_4542,N_4401,N_4457);
or U4543 (N_4543,N_4417,N_4433);
and U4544 (N_4544,N_4455,N_4407);
and U4545 (N_4545,N_4430,N_4487);
xor U4546 (N_4546,N_4424,N_4486);
nor U4547 (N_4547,N_4477,N_4431);
nor U4548 (N_4548,N_4472,N_4464);
nor U4549 (N_4549,N_4405,N_4461);
nor U4550 (N_4550,N_4469,N_4460);
nor U4551 (N_4551,N_4456,N_4429);
and U4552 (N_4552,N_4442,N_4411);
nand U4553 (N_4553,N_4413,N_4497);
or U4554 (N_4554,N_4431,N_4451);
or U4555 (N_4555,N_4407,N_4491);
or U4556 (N_4556,N_4459,N_4406);
nand U4557 (N_4557,N_4447,N_4430);
nand U4558 (N_4558,N_4468,N_4475);
or U4559 (N_4559,N_4433,N_4402);
nor U4560 (N_4560,N_4446,N_4462);
or U4561 (N_4561,N_4488,N_4497);
nor U4562 (N_4562,N_4483,N_4423);
nand U4563 (N_4563,N_4413,N_4424);
nand U4564 (N_4564,N_4413,N_4437);
or U4565 (N_4565,N_4407,N_4488);
nor U4566 (N_4566,N_4473,N_4455);
or U4567 (N_4567,N_4447,N_4497);
nor U4568 (N_4568,N_4486,N_4459);
and U4569 (N_4569,N_4460,N_4404);
nand U4570 (N_4570,N_4430,N_4476);
and U4571 (N_4571,N_4442,N_4475);
or U4572 (N_4572,N_4403,N_4402);
nand U4573 (N_4573,N_4442,N_4436);
or U4574 (N_4574,N_4415,N_4409);
or U4575 (N_4575,N_4482,N_4408);
xor U4576 (N_4576,N_4492,N_4432);
xor U4577 (N_4577,N_4477,N_4470);
nand U4578 (N_4578,N_4491,N_4455);
and U4579 (N_4579,N_4484,N_4459);
or U4580 (N_4580,N_4412,N_4456);
or U4581 (N_4581,N_4411,N_4497);
and U4582 (N_4582,N_4406,N_4423);
and U4583 (N_4583,N_4430,N_4435);
nand U4584 (N_4584,N_4432,N_4409);
xnor U4585 (N_4585,N_4487,N_4429);
nand U4586 (N_4586,N_4475,N_4401);
nand U4587 (N_4587,N_4488,N_4435);
nand U4588 (N_4588,N_4421,N_4472);
and U4589 (N_4589,N_4452,N_4473);
xor U4590 (N_4590,N_4424,N_4495);
or U4591 (N_4591,N_4426,N_4440);
nand U4592 (N_4592,N_4432,N_4471);
or U4593 (N_4593,N_4431,N_4437);
or U4594 (N_4594,N_4419,N_4480);
xor U4595 (N_4595,N_4493,N_4400);
nand U4596 (N_4596,N_4477,N_4409);
xor U4597 (N_4597,N_4415,N_4463);
and U4598 (N_4598,N_4490,N_4453);
nor U4599 (N_4599,N_4469,N_4486);
or U4600 (N_4600,N_4501,N_4590);
or U4601 (N_4601,N_4542,N_4579);
nand U4602 (N_4602,N_4541,N_4588);
or U4603 (N_4603,N_4557,N_4528);
and U4604 (N_4604,N_4529,N_4514);
and U4605 (N_4605,N_4537,N_4572);
nor U4606 (N_4606,N_4520,N_4505);
and U4607 (N_4607,N_4521,N_4578);
and U4608 (N_4608,N_4553,N_4536);
or U4609 (N_4609,N_4595,N_4574);
and U4610 (N_4610,N_4547,N_4551);
and U4611 (N_4611,N_4591,N_4575);
or U4612 (N_4612,N_4580,N_4549);
nand U4613 (N_4613,N_4599,N_4518);
and U4614 (N_4614,N_4517,N_4597);
xor U4615 (N_4615,N_4512,N_4568);
nand U4616 (N_4616,N_4534,N_4532);
nand U4617 (N_4617,N_4533,N_4552);
and U4618 (N_4618,N_4524,N_4598);
and U4619 (N_4619,N_4509,N_4594);
and U4620 (N_4620,N_4576,N_4507);
xnor U4621 (N_4621,N_4589,N_4506);
nor U4622 (N_4622,N_4516,N_4531);
or U4623 (N_4623,N_4502,N_4593);
and U4624 (N_4624,N_4592,N_4545);
and U4625 (N_4625,N_4530,N_4561);
and U4626 (N_4626,N_4596,N_4569);
or U4627 (N_4627,N_4559,N_4526);
nor U4628 (N_4628,N_4565,N_4570);
and U4629 (N_4629,N_4513,N_4519);
nor U4630 (N_4630,N_4539,N_4522);
or U4631 (N_4631,N_4581,N_4548);
nand U4632 (N_4632,N_4573,N_4554);
and U4633 (N_4633,N_4571,N_4535);
or U4634 (N_4634,N_4525,N_4586);
or U4635 (N_4635,N_4582,N_4544);
and U4636 (N_4636,N_4511,N_4562);
xnor U4637 (N_4637,N_4503,N_4508);
or U4638 (N_4638,N_4523,N_4550);
nand U4639 (N_4639,N_4563,N_4527);
xnor U4640 (N_4640,N_4583,N_4543);
nand U4641 (N_4641,N_4566,N_4538);
nor U4642 (N_4642,N_4504,N_4560);
nand U4643 (N_4643,N_4540,N_4555);
xnor U4644 (N_4644,N_4567,N_4577);
or U4645 (N_4645,N_4558,N_4584);
nor U4646 (N_4646,N_4510,N_4515);
and U4647 (N_4647,N_4564,N_4587);
nand U4648 (N_4648,N_4500,N_4546);
nor U4649 (N_4649,N_4556,N_4585);
nand U4650 (N_4650,N_4592,N_4535);
and U4651 (N_4651,N_4551,N_4558);
or U4652 (N_4652,N_4526,N_4597);
or U4653 (N_4653,N_4551,N_4507);
and U4654 (N_4654,N_4551,N_4514);
and U4655 (N_4655,N_4537,N_4560);
nor U4656 (N_4656,N_4588,N_4547);
nor U4657 (N_4657,N_4531,N_4555);
nor U4658 (N_4658,N_4534,N_4552);
or U4659 (N_4659,N_4553,N_4580);
or U4660 (N_4660,N_4559,N_4504);
or U4661 (N_4661,N_4586,N_4511);
nand U4662 (N_4662,N_4515,N_4504);
and U4663 (N_4663,N_4571,N_4582);
and U4664 (N_4664,N_4555,N_4511);
nor U4665 (N_4665,N_4552,N_4562);
or U4666 (N_4666,N_4587,N_4508);
nor U4667 (N_4667,N_4535,N_4523);
or U4668 (N_4668,N_4539,N_4591);
or U4669 (N_4669,N_4532,N_4530);
xnor U4670 (N_4670,N_4559,N_4505);
and U4671 (N_4671,N_4506,N_4517);
or U4672 (N_4672,N_4506,N_4551);
and U4673 (N_4673,N_4510,N_4546);
xnor U4674 (N_4674,N_4544,N_4532);
and U4675 (N_4675,N_4524,N_4509);
or U4676 (N_4676,N_4576,N_4567);
nand U4677 (N_4677,N_4539,N_4550);
and U4678 (N_4678,N_4509,N_4547);
or U4679 (N_4679,N_4507,N_4516);
nor U4680 (N_4680,N_4540,N_4504);
nand U4681 (N_4681,N_4598,N_4594);
nand U4682 (N_4682,N_4520,N_4515);
or U4683 (N_4683,N_4567,N_4586);
and U4684 (N_4684,N_4569,N_4592);
nor U4685 (N_4685,N_4567,N_4548);
nand U4686 (N_4686,N_4529,N_4578);
or U4687 (N_4687,N_4563,N_4573);
nor U4688 (N_4688,N_4544,N_4555);
nand U4689 (N_4689,N_4562,N_4570);
nand U4690 (N_4690,N_4521,N_4590);
nor U4691 (N_4691,N_4557,N_4535);
xor U4692 (N_4692,N_4545,N_4507);
nor U4693 (N_4693,N_4582,N_4547);
nor U4694 (N_4694,N_4576,N_4546);
nor U4695 (N_4695,N_4560,N_4539);
or U4696 (N_4696,N_4542,N_4546);
nand U4697 (N_4697,N_4541,N_4511);
or U4698 (N_4698,N_4564,N_4562);
and U4699 (N_4699,N_4531,N_4552);
nor U4700 (N_4700,N_4646,N_4699);
and U4701 (N_4701,N_4685,N_4671);
and U4702 (N_4702,N_4609,N_4628);
and U4703 (N_4703,N_4692,N_4663);
nor U4704 (N_4704,N_4697,N_4686);
or U4705 (N_4705,N_4656,N_4642);
or U4706 (N_4706,N_4620,N_4645);
and U4707 (N_4707,N_4624,N_4636);
nand U4708 (N_4708,N_4629,N_4687);
or U4709 (N_4709,N_4637,N_4660);
and U4710 (N_4710,N_4605,N_4666);
or U4711 (N_4711,N_4675,N_4639);
nand U4712 (N_4712,N_4622,N_4681);
nand U4713 (N_4713,N_4658,N_4649);
xnor U4714 (N_4714,N_4652,N_4662);
or U4715 (N_4715,N_4691,N_4694);
and U4716 (N_4716,N_4618,N_4698);
and U4717 (N_4717,N_4695,N_4643);
nand U4718 (N_4718,N_4661,N_4650);
nand U4719 (N_4719,N_4608,N_4682);
nand U4720 (N_4720,N_4648,N_4654);
xnor U4721 (N_4721,N_4600,N_4630);
and U4722 (N_4722,N_4669,N_4607);
nand U4723 (N_4723,N_4615,N_4623);
and U4724 (N_4724,N_4667,N_4601);
xnor U4725 (N_4725,N_4603,N_4651);
and U4726 (N_4726,N_4673,N_4696);
nand U4727 (N_4727,N_4610,N_4684);
nand U4728 (N_4728,N_4602,N_4640);
nand U4729 (N_4729,N_4647,N_4668);
and U4730 (N_4730,N_4625,N_4659);
or U4731 (N_4731,N_4613,N_4653);
and U4732 (N_4732,N_4690,N_4683);
nor U4733 (N_4733,N_4655,N_4670);
and U4734 (N_4734,N_4635,N_4633);
and U4735 (N_4735,N_4626,N_4606);
nand U4736 (N_4736,N_4611,N_4631);
and U4737 (N_4737,N_4679,N_4680);
or U4738 (N_4738,N_4693,N_4616);
xor U4739 (N_4739,N_4664,N_4619);
or U4740 (N_4740,N_4688,N_4617);
or U4741 (N_4741,N_4634,N_4678);
and U4742 (N_4742,N_4674,N_4604);
or U4743 (N_4743,N_4677,N_4632);
and U4744 (N_4744,N_4644,N_4676);
nand U4745 (N_4745,N_4627,N_4612);
and U4746 (N_4746,N_4657,N_4665);
nor U4747 (N_4747,N_4621,N_4689);
xnor U4748 (N_4748,N_4641,N_4672);
and U4749 (N_4749,N_4638,N_4614);
nor U4750 (N_4750,N_4627,N_4681);
nand U4751 (N_4751,N_4647,N_4665);
and U4752 (N_4752,N_4667,N_4637);
nor U4753 (N_4753,N_4600,N_4615);
nand U4754 (N_4754,N_4647,N_4697);
nand U4755 (N_4755,N_4673,N_4627);
or U4756 (N_4756,N_4622,N_4634);
and U4757 (N_4757,N_4614,N_4646);
or U4758 (N_4758,N_4601,N_4613);
and U4759 (N_4759,N_4607,N_4645);
nor U4760 (N_4760,N_4677,N_4626);
nor U4761 (N_4761,N_4670,N_4657);
nand U4762 (N_4762,N_4616,N_4646);
or U4763 (N_4763,N_4652,N_4624);
nand U4764 (N_4764,N_4635,N_4623);
or U4765 (N_4765,N_4657,N_4605);
nand U4766 (N_4766,N_4654,N_4676);
nand U4767 (N_4767,N_4602,N_4693);
nor U4768 (N_4768,N_4682,N_4652);
nand U4769 (N_4769,N_4668,N_4662);
or U4770 (N_4770,N_4640,N_4686);
nor U4771 (N_4771,N_4666,N_4609);
nand U4772 (N_4772,N_4673,N_4638);
xor U4773 (N_4773,N_4605,N_4663);
nand U4774 (N_4774,N_4602,N_4623);
nand U4775 (N_4775,N_4674,N_4664);
xor U4776 (N_4776,N_4686,N_4683);
nand U4777 (N_4777,N_4623,N_4684);
and U4778 (N_4778,N_4684,N_4671);
or U4779 (N_4779,N_4690,N_4692);
and U4780 (N_4780,N_4659,N_4651);
and U4781 (N_4781,N_4623,N_4607);
nand U4782 (N_4782,N_4656,N_4619);
and U4783 (N_4783,N_4676,N_4655);
or U4784 (N_4784,N_4649,N_4650);
and U4785 (N_4785,N_4641,N_4608);
or U4786 (N_4786,N_4609,N_4646);
and U4787 (N_4787,N_4679,N_4612);
xor U4788 (N_4788,N_4699,N_4621);
and U4789 (N_4789,N_4660,N_4612);
or U4790 (N_4790,N_4642,N_4636);
or U4791 (N_4791,N_4618,N_4603);
nor U4792 (N_4792,N_4687,N_4680);
nand U4793 (N_4793,N_4635,N_4663);
nor U4794 (N_4794,N_4682,N_4609);
nand U4795 (N_4795,N_4668,N_4695);
or U4796 (N_4796,N_4624,N_4634);
or U4797 (N_4797,N_4691,N_4606);
nor U4798 (N_4798,N_4609,N_4664);
nor U4799 (N_4799,N_4635,N_4679);
nor U4800 (N_4800,N_4797,N_4780);
and U4801 (N_4801,N_4751,N_4758);
nor U4802 (N_4802,N_4785,N_4709);
nor U4803 (N_4803,N_4755,N_4774);
xor U4804 (N_4804,N_4783,N_4726);
nor U4805 (N_4805,N_4713,N_4788);
nor U4806 (N_4806,N_4739,N_4706);
and U4807 (N_4807,N_4707,N_4778);
nand U4808 (N_4808,N_4703,N_4757);
nor U4809 (N_4809,N_4743,N_4770);
or U4810 (N_4810,N_4766,N_4710);
nand U4811 (N_4811,N_4712,N_4723);
nand U4812 (N_4812,N_4764,N_4719);
xor U4813 (N_4813,N_4724,N_4704);
or U4814 (N_4814,N_4722,N_4773);
nand U4815 (N_4815,N_4720,N_4776);
and U4816 (N_4816,N_4791,N_4730);
or U4817 (N_4817,N_4716,N_4784);
or U4818 (N_4818,N_4717,N_4789);
nor U4819 (N_4819,N_4782,N_4790);
nand U4820 (N_4820,N_4746,N_4754);
nand U4821 (N_4821,N_4747,N_4744);
nor U4822 (N_4822,N_4761,N_4793);
nand U4823 (N_4823,N_4740,N_4734);
and U4824 (N_4824,N_4763,N_4752);
and U4825 (N_4825,N_4700,N_4737);
nand U4826 (N_4826,N_4714,N_4799);
nor U4827 (N_4827,N_4748,N_4753);
and U4828 (N_4828,N_4798,N_4731);
or U4829 (N_4829,N_4771,N_4777);
and U4830 (N_4830,N_4772,N_4701);
nor U4831 (N_4831,N_4718,N_4745);
and U4832 (N_4832,N_4775,N_4750);
or U4833 (N_4833,N_4749,N_4767);
nand U4834 (N_4834,N_4705,N_4794);
nand U4835 (N_4835,N_4711,N_4728);
xnor U4836 (N_4836,N_4762,N_4742);
nor U4837 (N_4837,N_4738,N_4721);
or U4838 (N_4838,N_4792,N_4795);
or U4839 (N_4839,N_4760,N_4733);
nor U4840 (N_4840,N_4779,N_4725);
nand U4841 (N_4841,N_4715,N_4768);
nand U4842 (N_4842,N_4786,N_4729);
and U4843 (N_4843,N_4769,N_4736);
nor U4844 (N_4844,N_4759,N_4732);
or U4845 (N_4845,N_4735,N_4756);
nor U4846 (N_4846,N_4765,N_4727);
nand U4847 (N_4847,N_4708,N_4781);
and U4848 (N_4848,N_4787,N_4741);
and U4849 (N_4849,N_4702,N_4796);
and U4850 (N_4850,N_4794,N_4723);
nand U4851 (N_4851,N_4710,N_4701);
and U4852 (N_4852,N_4723,N_4725);
and U4853 (N_4853,N_4752,N_4733);
nand U4854 (N_4854,N_4706,N_4761);
or U4855 (N_4855,N_4783,N_4754);
xnor U4856 (N_4856,N_4773,N_4766);
and U4857 (N_4857,N_4715,N_4724);
and U4858 (N_4858,N_4728,N_4754);
nand U4859 (N_4859,N_4723,N_4782);
xnor U4860 (N_4860,N_4722,N_4717);
or U4861 (N_4861,N_4770,N_4739);
and U4862 (N_4862,N_4779,N_4789);
or U4863 (N_4863,N_4737,N_4750);
nor U4864 (N_4864,N_4769,N_4727);
nand U4865 (N_4865,N_4736,N_4770);
nand U4866 (N_4866,N_4745,N_4799);
and U4867 (N_4867,N_4796,N_4776);
and U4868 (N_4868,N_4737,N_4746);
and U4869 (N_4869,N_4780,N_4739);
or U4870 (N_4870,N_4724,N_4743);
or U4871 (N_4871,N_4734,N_4707);
nor U4872 (N_4872,N_4704,N_4708);
and U4873 (N_4873,N_4795,N_4745);
and U4874 (N_4874,N_4733,N_4720);
or U4875 (N_4875,N_4745,N_4797);
nand U4876 (N_4876,N_4748,N_4726);
nand U4877 (N_4877,N_4736,N_4724);
or U4878 (N_4878,N_4745,N_4717);
xnor U4879 (N_4879,N_4709,N_4732);
or U4880 (N_4880,N_4766,N_4799);
or U4881 (N_4881,N_4757,N_4784);
and U4882 (N_4882,N_4781,N_4731);
xor U4883 (N_4883,N_4781,N_4732);
xnor U4884 (N_4884,N_4780,N_4762);
nor U4885 (N_4885,N_4779,N_4756);
nand U4886 (N_4886,N_4719,N_4736);
and U4887 (N_4887,N_4746,N_4738);
or U4888 (N_4888,N_4700,N_4713);
nand U4889 (N_4889,N_4795,N_4711);
and U4890 (N_4890,N_4752,N_4789);
nand U4891 (N_4891,N_4778,N_4751);
nand U4892 (N_4892,N_4722,N_4757);
nand U4893 (N_4893,N_4747,N_4748);
or U4894 (N_4894,N_4799,N_4702);
nand U4895 (N_4895,N_4744,N_4733);
or U4896 (N_4896,N_4707,N_4719);
or U4897 (N_4897,N_4766,N_4793);
or U4898 (N_4898,N_4785,N_4704);
nor U4899 (N_4899,N_4709,N_4798);
nand U4900 (N_4900,N_4890,N_4862);
or U4901 (N_4901,N_4865,N_4821);
or U4902 (N_4902,N_4829,N_4856);
or U4903 (N_4903,N_4843,N_4868);
xnor U4904 (N_4904,N_4886,N_4816);
or U4905 (N_4905,N_4817,N_4827);
xor U4906 (N_4906,N_4830,N_4882);
nand U4907 (N_4907,N_4804,N_4811);
nand U4908 (N_4908,N_4823,N_4833);
and U4909 (N_4909,N_4870,N_4875);
nor U4910 (N_4910,N_4854,N_4845);
and U4911 (N_4911,N_4863,N_4826);
xor U4912 (N_4912,N_4834,N_4807);
or U4913 (N_4913,N_4867,N_4855);
nand U4914 (N_4914,N_4881,N_4879);
nand U4915 (N_4915,N_4898,N_4894);
and U4916 (N_4916,N_4893,N_4841);
nor U4917 (N_4917,N_4869,N_4891);
nand U4918 (N_4918,N_4885,N_4803);
or U4919 (N_4919,N_4859,N_4820);
or U4920 (N_4920,N_4851,N_4848);
and U4921 (N_4921,N_4801,N_4896);
nor U4922 (N_4922,N_4878,N_4805);
nor U4923 (N_4923,N_4889,N_4897);
xor U4924 (N_4924,N_4813,N_4842);
xor U4925 (N_4925,N_4872,N_4800);
and U4926 (N_4926,N_4815,N_4836);
and U4927 (N_4927,N_4835,N_4844);
and U4928 (N_4928,N_4857,N_4887);
nor U4929 (N_4929,N_4831,N_4824);
or U4930 (N_4930,N_4850,N_4884);
or U4931 (N_4931,N_4864,N_4809);
nand U4932 (N_4932,N_4814,N_4822);
or U4933 (N_4933,N_4883,N_4876);
nor U4934 (N_4934,N_4861,N_4874);
and U4935 (N_4935,N_4808,N_4873);
xor U4936 (N_4936,N_4852,N_4860);
nand U4937 (N_4937,N_4810,N_4846);
nand U4938 (N_4938,N_4849,N_4812);
nor U4939 (N_4939,N_4866,N_4828);
nand U4940 (N_4940,N_4892,N_4858);
and U4941 (N_4941,N_4819,N_4806);
nor U4942 (N_4942,N_4818,N_4871);
nor U4943 (N_4943,N_4802,N_4895);
nor U4944 (N_4944,N_4825,N_4847);
nor U4945 (N_4945,N_4837,N_4880);
or U4946 (N_4946,N_4877,N_4838);
nand U4947 (N_4947,N_4840,N_4853);
or U4948 (N_4948,N_4832,N_4888);
nor U4949 (N_4949,N_4839,N_4899);
or U4950 (N_4950,N_4802,N_4887);
or U4951 (N_4951,N_4805,N_4851);
or U4952 (N_4952,N_4862,N_4849);
or U4953 (N_4953,N_4827,N_4858);
xnor U4954 (N_4954,N_4876,N_4808);
and U4955 (N_4955,N_4814,N_4852);
and U4956 (N_4956,N_4883,N_4843);
or U4957 (N_4957,N_4876,N_4821);
or U4958 (N_4958,N_4896,N_4850);
or U4959 (N_4959,N_4834,N_4878);
and U4960 (N_4960,N_4834,N_4853);
nand U4961 (N_4961,N_4817,N_4878);
nor U4962 (N_4962,N_4874,N_4884);
and U4963 (N_4963,N_4802,N_4843);
or U4964 (N_4964,N_4804,N_4832);
and U4965 (N_4965,N_4829,N_4873);
nand U4966 (N_4966,N_4816,N_4808);
or U4967 (N_4967,N_4832,N_4876);
and U4968 (N_4968,N_4873,N_4870);
or U4969 (N_4969,N_4801,N_4869);
nand U4970 (N_4970,N_4880,N_4807);
and U4971 (N_4971,N_4859,N_4829);
nand U4972 (N_4972,N_4856,N_4897);
xor U4973 (N_4973,N_4870,N_4857);
or U4974 (N_4974,N_4808,N_4854);
and U4975 (N_4975,N_4840,N_4821);
xnor U4976 (N_4976,N_4879,N_4866);
and U4977 (N_4977,N_4856,N_4849);
and U4978 (N_4978,N_4849,N_4899);
nand U4979 (N_4979,N_4822,N_4835);
nand U4980 (N_4980,N_4887,N_4854);
or U4981 (N_4981,N_4805,N_4809);
and U4982 (N_4982,N_4814,N_4802);
nor U4983 (N_4983,N_4804,N_4826);
nand U4984 (N_4984,N_4860,N_4845);
and U4985 (N_4985,N_4893,N_4875);
or U4986 (N_4986,N_4809,N_4827);
nand U4987 (N_4987,N_4844,N_4819);
nor U4988 (N_4988,N_4891,N_4818);
nor U4989 (N_4989,N_4834,N_4865);
and U4990 (N_4990,N_4841,N_4847);
and U4991 (N_4991,N_4866,N_4835);
nand U4992 (N_4992,N_4876,N_4860);
or U4993 (N_4993,N_4873,N_4843);
nor U4994 (N_4994,N_4890,N_4821);
and U4995 (N_4995,N_4800,N_4839);
xnor U4996 (N_4996,N_4812,N_4830);
nand U4997 (N_4997,N_4888,N_4882);
nand U4998 (N_4998,N_4865,N_4819);
nand U4999 (N_4999,N_4885,N_4883);
or U5000 (N_5000,N_4921,N_4987);
and U5001 (N_5001,N_4956,N_4979);
or U5002 (N_5002,N_4939,N_4983);
nor U5003 (N_5003,N_4993,N_4914);
or U5004 (N_5004,N_4952,N_4965);
nand U5005 (N_5005,N_4935,N_4949);
nand U5006 (N_5006,N_4948,N_4911);
nand U5007 (N_5007,N_4918,N_4932);
nor U5008 (N_5008,N_4961,N_4907);
nand U5009 (N_5009,N_4902,N_4964);
nor U5010 (N_5010,N_4958,N_4990);
nor U5011 (N_5011,N_4991,N_4904);
or U5012 (N_5012,N_4943,N_4923);
nor U5013 (N_5013,N_4917,N_4915);
or U5014 (N_5014,N_4973,N_4936);
xor U5015 (N_5015,N_4927,N_4909);
and U5016 (N_5016,N_4905,N_4951);
or U5017 (N_5017,N_4963,N_4997);
nor U5018 (N_5018,N_4920,N_4957);
nand U5019 (N_5019,N_4966,N_4994);
nand U5020 (N_5020,N_4933,N_4981);
and U5021 (N_5021,N_4984,N_4998);
nor U5022 (N_5022,N_4922,N_4970);
nor U5023 (N_5023,N_4913,N_4969);
nand U5024 (N_5024,N_4971,N_4985);
nand U5025 (N_5025,N_4988,N_4977);
and U5026 (N_5026,N_4910,N_4975);
xnor U5027 (N_5027,N_4928,N_4938);
xor U5028 (N_5028,N_4912,N_4996);
and U5029 (N_5029,N_4937,N_4900);
or U5030 (N_5030,N_4926,N_4955);
and U5031 (N_5031,N_4929,N_4901);
and U5032 (N_5032,N_4953,N_4992);
nand U5033 (N_5033,N_4989,N_4947);
or U5034 (N_5034,N_4930,N_4903);
and U5035 (N_5035,N_4934,N_4976);
nand U5036 (N_5036,N_4916,N_4974);
or U5037 (N_5037,N_4908,N_4931);
nand U5038 (N_5038,N_4982,N_4906);
or U5039 (N_5039,N_4942,N_4944);
or U5040 (N_5040,N_4959,N_4941);
nor U5041 (N_5041,N_4960,N_4954);
or U5042 (N_5042,N_4986,N_4967);
xor U5043 (N_5043,N_4978,N_4925);
or U5044 (N_5044,N_4950,N_4946);
nand U5045 (N_5045,N_4995,N_4940);
and U5046 (N_5046,N_4962,N_4968);
nand U5047 (N_5047,N_4924,N_4919);
or U5048 (N_5048,N_4999,N_4972);
and U5049 (N_5049,N_4980,N_4945);
nand U5050 (N_5050,N_4969,N_4963);
or U5051 (N_5051,N_4971,N_4987);
nand U5052 (N_5052,N_4943,N_4976);
nand U5053 (N_5053,N_4969,N_4954);
and U5054 (N_5054,N_4959,N_4916);
or U5055 (N_5055,N_4960,N_4921);
nand U5056 (N_5056,N_4922,N_4939);
xnor U5057 (N_5057,N_4902,N_4937);
and U5058 (N_5058,N_4956,N_4997);
xnor U5059 (N_5059,N_4905,N_4949);
nand U5060 (N_5060,N_4998,N_4996);
nand U5061 (N_5061,N_4995,N_4949);
nand U5062 (N_5062,N_4916,N_4927);
nand U5063 (N_5063,N_4999,N_4912);
and U5064 (N_5064,N_4962,N_4931);
nor U5065 (N_5065,N_4974,N_4954);
and U5066 (N_5066,N_4935,N_4974);
nor U5067 (N_5067,N_4987,N_4974);
nand U5068 (N_5068,N_4921,N_4986);
nand U5069 (N_5069,N_4975,N_4982);
nor U5070 (N_5070,N_4945,N_4953);
or U5071 (N_5071,N_4906,N_4913);
or U5072 (N_5072,N_4997,N_4984);
nand U5073 (N_5073,N_4919,N_4938);
and U5074 (N_5074,N_4971,N_4975);
nand U5075 (N_5075,N_4931,N_4960);
or U5076 (N_5076,N_4967,N_4940);
nor U5077 (N_5077,N_4934,N_4919);
or U5078 (N_5078,N_4922,N_4952);
nand U5079 (N_5079,N_4994,N_4991);
and U5080 (N_5080,N_4919,N_4963);
or U5081 (N_5081,N_4940,N_4953);
xnor U5082 (N_5082,N_4914,N_4946);
and U5083 (N_5083,N_4914,N_4943);
nor U5084 (N_5084,N_4963,N_4912);
nand U5085 (N_5085,N_4903,N_4910);
or U5086 (N_5086,N_4991,N_4966);
xnor U5087 (N_5087,N_4956,N_4995);
and U5088 (N_5088,N_4917,N_4923);
nor U5089 (N_5089,N_4921,N_4943);
or U5090 (N_5090,N_4989,N_4913);
nand U5091 (N_5091,N_4961,N_4923);
or U5092 (N_5092,N_4915,N_4986);
nand U5093 (N_5093,N_4972,N_4962);
nor U5094 (N_5094,N_4964,N_4995);
or U5095 (N_5095,N_4913,N_4942);
or U5096 (N_5096,N_4986,N_4929);
and U5097 (N_5097,N_4957,N_4931);
nor U5098 (N_5098,N_4994,N_4951);
nand U5099 (N_5099,N_4975,N_4937);
and U5100 (N_5100,N_5014,N_5059);
xnor U5101 (N_5101,N_5071,N_5001);
or U5102 (N_5102,N_5051,N_5013);
or U5103 (N_5103,N_5037,N_5010);
or U5104 (N_5104,N_5048,N_5046);
or U5105 (N_5105,N_5009,N_5021);
nor U5106 (N_5106,N_5004,N_5073);
nor U5107 (N_5107,N_5050,N_5043);
nor U5108 (N_5108,N_5066,N_5098);
and U5109 (N_5109,N_5076,N_5091);
nor U5110 (N_5110,N_5019,N_5090);
xnor U5111 (N_5111,N_5032,N_5055);
or U5112 (N_5112,N_5062,N_5003);
and U5113 (N_5113,N_5017,N_5082);
nand U5114 (N_5114,N_5027,N_5042);
xor U5115 (N_5115,N_5024,N_5012);
and U5116 (N_5116,N_5023,N_5045);
and U5117 (N_5117,N_5078,N_5083);
or U5118 (N_5118,N_5022,N_5092);
xor U5119 (N_5119,N_5064,N_5065);
xnor U5120 (N_5120,N_5053,N_5028);
nand U5121 (N_5121,N_5077,N_5063);
or U5122 (N_5122,N_5085,N_5084);
or U5123 (N_5123,N_5058,N_5034);
nand U5124 (N_5124,N_5079,N_5087);
nor U5125 (N_5125,N_5038,N_5089);
and U5126 (N_5126,N_5088,N_5093);
or U5127 (N_5127,N_5002,N_5049);
or U5128 (N_5128,N_5018,N_5030);
xor U5129 (N_5129,N_5069,N_5094);
nand U5130 (N_5130,N_5072,N_5075);
or U5131 (N_5131,N_5052,N_5080);
or U5132 (N_5132,N_5097,N_5036);
nand U5133 (N_5133,N_5020,N_5041);
nand U5134 (N_5134,N_5060,N_5086);
nor U5135 (N_5135,N_5015,N_5047);
nor U5136 (N_5136,N_5025,N_5040);
and U5137 (N_5137,N_5029,N_5044);
and U5138 (N_5138,N_5074,N_5031);
nor U5139 (N_5139,N_5005,N_5099);
nor U5140 (N_5140,N_5039,N_5067);
nand U5141 (N_5141,N_5033,N_5070);
nor U5142 (N_5142,N_5016,N_5096);
nor U5143 (N_5143,N_5057,N_5061);
and U5144 (N_5144,N_5054,N_5081);
nor U5145 (N_5145,N_5008,N_5026);
or U5146 (N_5146,N_5056,N_5068);
or U5147 (N_5147,N_5000,N_5095);
xor U5148 (N_5148,N_5035,N_5007);
nand U5149 (N_5149,N_5006,N_5011);
nand U5150 (N_5150,N_5083,N_5066);
and U5151 (N_5151,N_5005,N_5062);
and U5152 (N_5152,N_5069,N_5048);
nand U5153 (N_5153,N_5078,N_5042);
or U5154 (N_5154,N_5008,N_5096);
nor U5155 (N_5155,N_5039,N_5098);
and U5156 (N_5156,N_5071,N_5037);
and U5157 (N_5157,N_5005,N_5070);
nor U5158 (N_5158,N_5059,N_5017);
nand U5159 (N_5159,N_5090,N_5020);
nand U5160 (N_5160,N_5060,N_5035);
nor U5161 (N_5161,N_5081,N_5085);
nand U5162 (N_5162,N_5081,N_5086);
nor U5163 (N_5163,N_5034,N_5069);
nor U5164 (N_5164,N_5021,N_5076);
nand U5165 (N_5165,N_5025,N_5032);
and U5166 (N_5166,N_5015,N_5021);
and U5167 (N_5167,N_5089,N_5085);
nand U5168 (N_5168,N_5038,N_5099);
nand U5169 (N_5169,N_5010,N_5058);
nor U5170 (N_5170,N_5006,N_5046);
nor U5171 (N_5171,N_5067,N_5069);
and U5172 (N_5172,N_5057,N_5072);
nor U5173 (N_5173,N_5097,N_5073);
nand U5174 (N_5174,N_5060,N_5043);
nor U5175 (N_5175,N_5048,N_5053);
nand U5176 (N_5176,N_5053,N_5013);
or U5177 (N_5177,N_5057,N_5099);
nand U5178 (N_5178,N_5080,N_5099);
and U5179 (N_5179,N_5039,N_5089);
or U5180 (N_5180,N_5088,N_5072);
or U5181 (N_5181,N_5094,N_5010);
and U5182 (N_5182,N_5011,N_5058);
nor U5183 (N_5183,N_5015,N_5003);
and U5184 (N_5184,N_5080,N_5058);
nand U5185 (N_5185,N_5009,N_5078);
or U5186 (N_5186,N_5021,N_5032);
nor U5187 (N_5187,N_5049,N_5036);
nand U5188 (N_5188,N_5033,N_5037);
and U5189 (N_5189,N_5062,N_5041);
nor U5190 (N_5190,N_5067,N_5009);
xnor U5191 (N_5191,N_5065,N_5002);
or U5192 (N_5192,N_5091,N_5008);
nand U5193 (N_5193,N_5029,N_5087);
nand U5194 (N_5194,N_5006,N_5042);
nand U5195 (N_5195,N_5046,N_5002);
and U5196 (N_5196,N_5056,N_5070);
nand U5197 (N_5197,N_5092,N_5058);
or U5198 (N_5198,N_5066,N_5096);
nand U5199 (N_5199,N_5016,N_5051);
nor U5200 (N_5200,N_5118,N_5166);
nand U5201 (N_5201,N_5155,N_5105);
nor U5202 (N_5202,N_5115,N_5196);
nor U5203 (N_5203,N_5192,N_5195);
nor U5204 (N_5204,N_5179,N_5127);
and U5205 (N_5205,N_5100,N_5141);
nand U5206 (N_5206,N_5134,N_5157);
or U5207 (N_5207,N_5146,N_5116);
and U5208 (N_5208,N_5128,N_5163);
and U5209 (N_5209,N_5142,N_5193);
xor U5210 (N_5210,N_5185,N_5153);
xor U5211 (N_5211,N_5181,N_5164);
or U5212 (N_5212,N_5188,N_5186);
nand U5213 (N_5213,N_5104,N_5174);
and U5214 (N_5214,N_5159,N_5102);
and U5215 (N_5215,N_5152,N_5150);
nor U5216 (N_5216,N_5167,N_5109);
nand U5217 (N_5217,N_5169,N_5190);
or U5218 (N_5218,N_5162,N_5126);
nand U5219 (N_5219,N_5133,N_5183);
nand U5220 (N_5220,N_5114,N_5199);
xor U5221 (N_5221,N_5101,N_5113);
nand U5222 (N_5222,N_5140,N_5124);
xor U5223 (N_5223,N_5120,N_5117);
or U5224 (N_5224,N_5131,N_5121);
or U5225 (N_5225,N_5106,N_5171);
nor U5226 (N_5226,N_5168,N_5156);
or U5227 (N_5227,N_5191,N_5154);
nor U5228 (N_5228,N_5130,N_5187);
xnor U5229 (N_5229,N_5132,N_5198);
and U5230 (N_5230,N_5138,N_5180);
and U5231 (N_5231,N_5151,N_5158);
and U5232 (N_5232,N_5107,N_5112);
nor U5233 (N_5233,N_5160,N_5123);
nor U5234 (N_5234,N_5176,N_5122);
and U5235 (N_5235,N_5119,N_5194);
or U5236 (N_5236,N_5110,N_5197);
xor U5237 (N_5237,N_5145,N_5125);
nand U5238 (N_5238,N_5170,N_5175);
and U5239 (N_5239,N_5149,N_5182);
or U5240 (N_5240,N_5173,N_5189);
nor U5241 (N_5241,N_5135,N_5111);
or U5242 (N_5242,N_5147,N_5144);
nand U5243 (N_5243,N_5137,N_5139);
and U5244 (N_5244,N_5161,N_5165);
or U5245 (N_5245,N_5177,N_5136);
nor U5246 (N_5246,N_5184,N_5129);
or U5247 (N_5247,N_5143,N_5148);
nor U5248 (N_5248,N_5108,N_5172);
or U5249 (N_5249,N_5103,N_5178);
nand U5250 (N_5250,N_5146,N_5151);
and U5251 (N_5251,N_5164,N_5146);
or U5252 (N_5252,N_5148,N_5139);
or U5253 (N_5253,N_5188,N_5168);
or U5254 (N_5254,N_5189,N_5197);
nand U5255 (N_5255,N_5136,N_5155);
nand U5256 (N_5256,N_5110,N_5141);
and U5257 (N_5257,N_5103,N_5100);
nor U5258 (N_5258,N_5169,N_5179);
nor U5259 (N_5259,N_5158,N_5156);
nand U5260 (N_5260,N_5116,N_5155);
nor U5261 (N_5261,N_5119,N_5110);
nand U5262 (N_5262,N_5160,N_5118);
and U5263 (N_5263,N_5110,N_5158);
or U5264 (N_5264,N_5152,N_5168);
and U5265 (N_5265,N_5143,N_5169);
nor U5266 (N_5266,N_5135,N_5157);
nor U5267 (N_5267,N_5127,N_5133);
and U5268 (N_5268,N_5148,N_5188);
nor U5269 (N_5269,N_5120,N_5190);
and U5270 (N_5270,N_5135,N_5144);
nand U5271 (N_5271,N_5127,N_5163);
and U5272 (N_5272,N_5119,N_5145);
xnor U5273 (N_5273,N_5127,N_5102);
and U5274 (N_5274,N_5182,N_5152);
and U5275 (N_5275,N_5149,N_5193);
and U5276 (N_5276,N_5118,N_5195);
nand U5277 (N_5277,N_5119,N_5175);
or U5278 (N_5278,N_5131,N_5194);
nand U5279 (N_5279,N_5141,N_5118);
xnor U5280 (N_5280,N_5102,N_5101);
or U5281 (N_5281,N_5117,N_5152);
and U5282 (N_5282,N_5131,N_5129);
and U5283 (N_5283,N_5158,N_5102);
and U5284 (N_5284,N_5199,N_5135);
nand U5285 (N_5285,N_5179,N_5165);
or U5286 (N_5286,N_5163,N_5194);
or U5287 (N_5287,N_5180,N_5168);
or U5288 (N_5288,N_5171,N_5128);
and U5289 (N_5289,N_5147,N_5148);
and U5290 (N_5290,N_5142,N_5112);
and U5291 (N_5291,N_5145,N_5185);
xor U5292 (N_5292,N_5156,N_5163);
nand U5293 (N_5293,N_5126,N_5191);
or U5294 (N_5294,N_5141,N_5146);
or U5295 (N_5295,N_5171,N_5140);
or U5296 (N_5296,N_5132,N_5163);
nor U5297 (N_5297,N_5160,N_5124);
nand U5298 (N_5298,N_5125,N_5132);
xnor U5299 (N_5299,N_5148,N_5122);
xnor U5300 (N_5300,N_5282,N_5228);
and U5301 (N_5301,N_5234,N_5236);
nor U5302 (N_5302,N_5298,N_5268);
nor U5303 (N_5303,N_5279,N_5251);
nor U5304 (N_5304,N_5267,N_5212);
nand U5305 (N_5305,N_5208,N_5202);
nand U5306 (N_5306,N_5233,N_5259);
nand U5307 (N_5307,N_5246,N_5248);
or U5308 (N_5308,N_5258,N_5238);
or U5309 (N_5309,N_5222,N_5264);
nand U5310 (N_5310,N_5270,N_5219);
and U5311 (N_5311,N_5213,N_5269);
and U5312 (N_5312,N_5225,N_5257);
nand U5313 (N_5313,N_5244,N_5243);
or U5314 (N_5314,N_5247,N_5278);
or U5315 (N_5315,N_5239,N_5221);
xnor U5316 (N_5316,N_5226,N_5241);
nor U5317 (N_5317,N_5277,N_5266);
nor U5318 (N_5318,N_5200,N_5260);
and U5319 (N_5319,N_5237,N_5276);
nor U5320 (N_5320,N_5292,N_5287);
nand U5321 (N_5321,N_5204,N_5294);
and U5322 (N_5322,N_5209,N_5227);
nor U5323 (N_5323,N_5240,N_5205);
or U5324 (N_5324,N_5274,N_5281);
nand U5325 (N_5325,N_5230,N_5283);
nor U5326 (N_5326,N_5265,N_5290);
or U5327 (N_5327,N_5286,N_5255);
xnor U5328 (N_5328,N_5293,N_5215);
nand U5329 (N_5329,N_5273,N_5245);
nor U5330 (N_5330,N_5210,N_5211);
and U5331 (N_5331,N_5223,N_5297);
nand U5332 (N_5332,N_5235,N_5229);
or U5333 (N_5333,N_5217,N_5284);
or U5334 (N_5334,N_5218,N_5263);
nor U5335 (N_5335,N_5291,N_5206);
or U5336 (N_5336,N_5203,N_5272);
and U5337 (N_5337,N_5242,N_5299);
or U5338 (N_5338,N_5249,N_5250);
and U5339 (N_5339,N_5207,N_5232);
nor U5340 (N_5340,N_5253,N_5261);
nand U5341 (N_5341,N_5252,N_5254);
or U5342 (N_5342,N_5262,N_5271);
and U5343 (N_5343,N_5275,N_5289);
nand U5344 (N_5344,N_5288,N_5231);
and U5345 (N_5345,N_5295,N_5285);
nor U5346 (N_5346,N_5296,N_5216);
nor U5347 (N_5347,N_5220,N_5201);
and U5348 (N_5348,N_5224,N_5214);
nor U5349 (N_5349,N_5256,N_5280);
and U5350 (N_5350,N_5225,N_5280);
nor U5351 (N_5351,N_5289,N_5234);
or U5352 (N_5352,N_5267,N_5292);
nor U5353 (N_5353,N_5223,N_5290);
and U5354 (N_5354,N_5276,N_5265);
nor U5355 (N_5355,N_5278,N_5252);
or U5356 (N_5356,N_5215,N_5259);
xnor U5357 (N_5357,N_5264,N_5210);
nand U5358 (N_5358,N_5295,N_5260);
and U5359 (N_5359,N_5279,N_5203);
and U5360 (N_5360,N_5215,N_5204);
xor U5361 (N_5361,N_5257,N_5243);
and U5362 (N_5362,N_5285,N_5200);
nand U5363 (N_5363,N_5229,N_5277);
nand U5364 (N_5364,N_5237,N_5269);
nor U5365 (N_5365,N_5225,N_5256);
nor U5366 (N_5366,N_5245,N_5220);
xnor U5367 (N_5367,N_5293,N_5246);
and U5368 (N_5368,N_5293,N_5245);
nand U5369 (N_5369,N_5222,N_5238);
nand U5370 (N_5370,N_5296,N_5283);
nor U5371 (N_5371,N_5251,N_5217);
nor U5372 (N_5372,N_5228,N_5236);
or U5373 (N_5373,N_5269,N_5207);
nor U5374 (N_5374,N_5211,N_5249);
nand U5375 (N_5375,N_5225,N_5222);
xnor U5376 (N_5376,N_5261,N_5252);
nand U5377 (N_5377,N_5258,N_5214);
nand U5378 (N_5378,N_5292,N_5285);
or U5379 (N_5379,N_5265,N_5273);
or U5380 (N_5380,N_5260,N_5284);
nor U5381 (N_5381,N_5288,N_5294);
nor U5382 (N_5382,N_5225,N_5235);
nand U5383 (N_5383,N_5212,N_5220);
or U5384 (N_5384,N_5267,N_5247);
or U5385 (N_5385,N_5299,N_5279);
and U5386 (N_5386,N_5201,N_5217);
nor U5387 (N_5387,N_5218,N_5247);
xor U5388 (N_5388,N_5273,N_5220);
nand U5389 (N_5389,N_5278,N_5254);
xnor U5390 (N_5390,N_5266,N_5202);
xor U5391 (N_5391,N_5213,N_5239);
nand U5392 (N_5392,N_5282,N_5200);
or U5393 (N_5393,N_5212,N_5299);
and U5394 (N_5394,N_5280,N_5278);
nand U5395 (N_5395,N_5212,N_5216);
nand U5396 (N_5396,N_5225,N_5263);
or U5397 (N_5397,N_5288,N_5233);
nor U5398 (N_5398,N_5230,N_5251);
nand U5399 (N_5399,N_5234,N_5263);
nand U5400 (N_5400,N_5367,N_5347);
nand U5401 (N_5401,N_5350,N_5356);
and U5402 (N_5402,N_5309,N_5333);
nand U5403 (N_5403,N_5343,N_5324);
or U5404 (N_5404,N_5368,N_5340);
nand U5405 (N_5405,N_5312,N_5355);
nand U5406 (N_5406,N_5311,N_5373);
or U5407 (N_5407,N_5321,N_5375);
nor U5408 (N_5408,N_5337,N_5313);
nand U5409 (N_5409,N_5363,N_5395);
and U5410 (N_5410,N_5354,N_5325);
nor U5411 (N_5411,N_5329,N_5303);
or U5412 (N_5412,N_5314,N_5374);
nand U5413 (N_5413,N_5371,N_5319);
or U5414 (N_5414,N_5351,N_5370);
and U5415 (N_5415,N_5353,N_5360);
and U5416 (N_5416,N_5359,N_5300);
or U5417 (N_5417,N_5331,N_5352);
and U5418 (N_5418,N_5318,N_5381);
and U5419 (N_5419,N_5307,N_5382);
and U5420 (N_5420,N_5339,N_5326);
xor U5421 (N_5421,N_5385,N_5393);
xnor U5422 (N_5422,N_5377,N_5348);
nand U5423 (N_5423,N_5361,N_5323);
nor U5424 (N_5424,N_5304,N_5376);
or U5425 (N_5425,N_5334,N_5383);
nand U5426 (N_5426,N_5328,N_5315);
nand U5427 (N_5427,N_5302,N_5308);
nand U5428 (N_5428,N_5398,N_5338);
and U5429 (N_5429,N_5327,N_5305);
and U5430 (N_5430,N_5380,N_5357);
nor U5431 (N_5431,N_5392,N_5346);
nand U5432 (N_5432,N_5358,N_5399);
or U5433 (N_5433,N_5386,N_5316);
or U5434 (N_5434,N_5394,N_5372);
nor U5435 (N_5435,N_5332,N_5320);
or U5436 (N_5436,N_5389,N_5397);
or U5437 (N_5437,N_5390,N_5366);
or U5438 (N_5438,N_5322,N_5345);
nand U5439 (N_5439,N_5341,N_5317);
and U5440 (N_5440,N_5379,N_5349);
nor U5441 (N_5441,N_5378,N_5388);
nand U5442 (N_5442,N_5330,N_5344);
and U5443 (N_5443,N_5335,N_5306);
and U5444 (N_5444,N_5396,N_5391);
and U5445 (N_5445,N_5362,N_5310);
or U5446 (N_5446,N_5384,N_5301);
or U5447 (N_5447,N_5369,N_5336);
or U5448 (N_5448,N_5342,N_5365);
xor U5449 (N_5449,N_5364,N_5387);
or U5450 (N_5450,N_5376,N_5330);
xnor U5451 (N_5451,N_5318,N_5350);
nand U5452 (N_5452,N_5381,N_5305);
nand U5453 (N_5453,N_5359,N_5379);
nand U5454 (N_5454,N_5306,N_5310);
xnor U5455 (N_5455,N_5372,N_5369);
nand U5456 (N_5456,N_5382,N_5386);
nor U5457 (N_5457,N_5332,N_5373);
or U5458 (N_5458,N_5334,N_5324);
or U5459 (N_5459,N_5330,N_5351);
or U5460 (N_5460,N_5320,N_5377);
xnor U5461 (N_5461,N_5336,N_5307);
xor U5462 (N_5462,N_5367,N_5399);
nand U5463 (N_5463,N_5397,N_5316);
nand U5464 (N_5464,N_5322,N_5365);
nand U5465 (N_5465,N_5351,N_5386);
nor U5466 (N_5466,N_5364,N_5311);
or U5467 (N_5467,N_5350,N_5392);
nor U5468 (N_5468,N_5321,N_5373);
nor U5469 (N_5469,N_5310,N_5315);
nand U5470 (N_5470,N_5308,N_5372);
nor U5471 (N_5471,N_5328,N_5386);
or U5472 (N_5472,N_5386,N_5347);
and U5473 (N_5473,N_5334,N_5326);
and U5474 (N_5474,N_5307,N_5356);
nor U5475 (N_5475,N_5382,N_5394);
nand U5476 (N_5476,N_5390,N_5344);
and U5477 (N_5477,N_5302,N_5393);
nor U5478 (N_5478,N_5346,N_5357);
or U5479 (N_5479,N_5339,N_5322);
and U5480 (N_5480,N_5302,N_5353);
nand U5481 (N_5481,N_5380,N_5354);
and U5482 (N_5482,N_5385,N_5320);
or U5483 (N_5483,N_5326,N_5331);
nand U5484 (N_5484,N_5348,N_5333);
and U5485 (N_5485,N_5377,N_5388);
nand U5486 (N_5486,N_5318,N_5326);
and U5487 (N_5487,N_5310,N_5358);
nor U5488 (N_5488,N_5309,N_5312);
or U5489 (N_5489,N_5348,N_5389);
nor U5490 (N_5490,N_5343,N_5339);
nor U5491 (N_5491,N_5357,N_5359);
nand U5492 (N_5492,N_5353,N_5345);
nand U5493 (N_5493,N_5378,N_5396);
nor U5494 (N_5494,N_5354,N_5333);
and U5495 (N_5495,N_5333,N_5322);
nand U5496 (N_5496,N_5346,N_5300);
nor U5497 (N_5497,N_5355,N_5330);
nor U5498 (N_5498,N_5302,N_5395);
nand U5499 (N_5499,N_5315,N_5399);
and U5500 (N_5500,N_5437,N_5417);
or U5501 (N_5501,N_5425,N_5426);
or U5502 (N_5502,N_5434,N_5440);
and U5503 (N_5503,N_5410,N_5465);
nand U5504 (N_5504,N_5488,N_5414);
or U5505 (N_5505,N_5435,N_5499);
nand U5506 (N_5506,N_5483,N_5462);
and U5507 (N_5507,N_5494,N_5455);
and U5508 (N_5508,N_5421,N_5454);
and U5509 (N_5509,N_5443,N_5447);
or U5510 (N_5510,N_5445,N_5412);
nand U5511 (N_5511,N_5492,N_5469);
nor U5512 (N_5512,N_5419,N_5470);
and U5513 (N_5513,N_5448,N_5403);
and U5514 (N_5514,N_5464,N_5457);
and U5515 (N_5515,N_5407,N_5408);
nand U5516 (N_5516,N_5436,N_5490);
xnor U5517 (N_5517,N_5485,N_5460);
and U5518 (N_5518,N_5486,N_5481);
nand U5519 (N_5519,N_5431,N_5456);
nand U5520 (N_5520,N_5428,N_5480);
xor U5521 (N_5521,N_5438,N_5472);
and U5522 (N_5522,N_5424,N_5415);
and U5523 (N_5523,N_5423,N_5430);
nor U5524 (N_5524,N_5405,N_5487);
or U5525 (N_5525,N_5420,N_5433);
nor U5526 (N_5526,N_5422,N_5432);
nor U5527 (N_5527,N_5476,N_5402);
or U5528 (N_5528,N_5461,N_5495);
nand U5529 (N_5529,N_5466,N_5450);
or U5530 (N_5530,N_5400,N_5498);
xor U5531 (N_5531,N_5413,N_5484);
and U5532 (N_5532,N_5429,N_5439);
nor U5533 (N_5533,N_5444,N_5467);
nor U5534 (N_5534,N_5453,N_5489);
and U5535 (N_5535,N_5404,N_5416);
or U5536 (N_5536,N_5475,N_5478);
nand U5537 (N_5537,N_5474,N_5446);
nor U5538 (N_5538,N_5427,N_5497);
or U5539 (N_5539,N_5442,N_5452);
nand U5540 (N_5540,N_5418,N_5451);
or U5541 (N_5541,N_5449,N_5401);
nor U5542 (N_5542,N_5441,N_5473);
xor U5543 (N_5543,N_5463,N_5458);
and U5544 (N_5544,N_5406,N_5477);
or U5545 (N_5545,N_5493,N_5482);
nor U5546 (N_5546,N_5409,N_5468);
nor U5547 (N_5547,N_5496,N_5459);
nor U5548 (N_5548,N_5411,N_5471);
and U5549 (N_5549,N_5491,N_5479);
or U5550 (N_5550,N_5437,N_5445);
nor U5551 (N_5551,N_5450,N_5441);
or U5552 (N_5552,N_5455,N_5463);
nor U5553 (N_5553,N_5480,N_5416);
or U5554 (N_5554,N_5423,N_5479);
or U5555 (N_5555,N_5442,N_5477);
or U5556 (N_5556,N_5446,N_5445);
nor U5557 (N_5557,N_5457,N_5467);
or U5558 (N_5558,N_5474,N_5440);
and U5559 (N_5559,N_5458,N_5422);
xnor U5560 (N_5560,N_5497,N_5453);
xor U5561 (N_5561,N_5429,N_5478);
and U5562 (N_5562,N_5442,N_5449);
nand U5563 (N_5563,N_5433,N_5475);
and U5564 (N_5564,N_5464,N_5460);
and U5565 (N_5565,N_5436,N_5419);
and U5566 (N_5566,N_5480,N_5474);
and U5567 (N_5567,N_5410,N_5409);
nor U5568 (N_5568,N_5415,N_5468);
or U5569 (N_5569,N_5471,N_5489);
and U5570 (N_5570,N_5403,N_5437);
or U5571 (N_5571,N_5478,N_5497);
nand U5572 (N_5572,N_5432,N_5463);
nor U5573 (N_5573,N_5496,N_5437);
and U5574 (N_5574,N_5461,N_5408);
and U5575 (N_5575,N_5478,N_5441);
or U5576 (N_5576,N_5452,N_5482);
or U5577 (N_5577,N_5490,N_5455);
and U5578 (N_5578,N_5419,N_5401);
nor U5579 (N_5579,N_5403,N_5463);
nor U5580 (N_5580,N_5428,N_5451);
and U5581 (N_5581,N_5432,N_5466);
and U5582 (N_5582,N_5489,N_5434);
and U5583 (N_5583,N_5465,N_5412);
xnor U5584 (N_5584,N_5487,N_5484);
nor U5585 (N_5585,N_5465,N_5469);
nand U5586 (N_5586,N_5419,N_5409);
xor U5587 (N_5587,N_5454,N_5418);
xor U5588 (N_5588,N_5448,N_5401);
nor U5589 (N_5589,N_5421,N_5476);
and U5590 (N_5590,N_5484,N_5499);
nor U5591 (N_5591,N_5439,N_5445);
or U5592 (N_5592,N_5447,N_5462);
xor U5593 (N_5593,N_5406,N_5405);
nand U5594 (N_5594,N_5406,N_5449);
and U5595 (N_5595,N_5476,N_5407);
nor U5596 (N_5596,N_5441,N_5403);
and U5597 (N_5597,N_5445,N_5409);
nor U5598 (N_5598,N_5465,N_5478);
nor U5599 (N_5599,N_5446,N_5461);
nor U5600 (N_5600,N_5580,N_5508);
xor U5601 (N_5601,N_5559,N_5573);
and U5602 (N_5602,N_5545,N_5560);
and U5603 (N_5603,N_5529,N_5564);
nand U5604 (N_5604,N_5527,N_5504);
nand U5605 (N_5605,N_5522,N_5579);
and U5606 (N_5606,N_5551,N_5543);
nor U5607 (N_5607,N_5541,N_5590);
or U5608 (N_5608,N_5571,N_5501);
xnor U5609 (N_5609,N_5505,N_5544);
and U5610 (N_5610,N_5586,N_5570);
nor U5611 (N_5611,N_5567,N_5502);
nor U5612 (N_5612,N_5547,N_5526);
nor U5613 (N_5613,N_5563,N_5548);
or U5614 (N_5614,N_5528,N_5511);
nor U5615 (N_5615,N_5574,N_5537);
or U5616 (N_5616,N_5503,N_5514);
nor U5617 (N_5617,N_5558,N_5517);
and U5618 (N_5618,N_5577,N_5583);
and U5619 (N_5619,N_5532,N_5513);
or U5620 (N_5620,N_5582,N_5523);
or U5621 (N_5621,N_5596,N_5510);
nor U5622 (N_5622,N_5569,N_5540);
xor U5623 (N_5623,N_5515,N_5598);
nand U5624 (N_5624,N_5500,N_5561);
nor U5625 (N_5625,N_5506,N_5562);
nor U5626 (N_5626,N_5599,N_5524);
and U5627 (N_5627,N_5566,N_5549);
or U5628 (N_5628,N_5509,N_5578);
nor U5629 (N_5629,N_5591,N_5581);
nor U5630 (N_5630,N_5539,N_5585);
nand U5631 (N_5631,N_5530,N_5531);
or U5632 (N_5632,N_5518,N_5546);
nand U5633 (N_5633,N_5588,N_5584);
and U5634 (N_5634,N_5525,N_5587);
nor U5635 (N_5635,N_5557,N_5593);
xor U5636 (N_5636,N_5572,N_5507);
xnor U5637 (N_5637,N_5553,N_5589);
or U5638 (N_5638,N_5550,N_5536);
nand U5639 (N_5639,N_5552,N_5594);
xnor U5640 (N_5640,N_5568,N_5512);
or U5641 (N_5641,N_5592,N_5595);
or U5642 (N_5642,N_5576,N_5597);
and U5643 (N_5643,N_5575,N_5519);
and U5644 (N_5644,N_5534,N_5555);
and U5645 (N_5645,N_5565,N_5556);
nand U5646 (N_5646,N_5533,N_5538);
xor U5647 (N_5647,N_5520,N_5521);
nand U5648 (N_5648,N_5535,N_5516);
nand U5649 (N_5649,N_5542,N_5554);
nand U5650 (N_5650,N_5583,N_5508);
nor U5651 (N_5651,N_5580,N_5531);
or U5652 (N_5652,N_5507,N_5573);
nand U5653 (N_5653,N_5567,N_5507);
and U5654 (N_5654,N_5575,N_5577);
nor U5655 (N_5655,N_5540,N_5516);
xnor U5656 (N_5656,N_5588,N_5565);
or U5657 (N_5657,N_5520,N_5577);
xnor U5658 (N_5658,N_5586,N_5580);
and U5659 (N_5659,N_5575,N_5535);
and U5660 (N_5660,N_5577,N_5598);
or U5661 (N_5661,N_5548,N_5571);
and U5662 (N_5662,N_5541,N_5588);
or U5663 (N_5663,N_5547,N_5515);
or U5664 (N_5664,N_5545,N_5522);
xnor U5665 (N_5665,N_5541,N_5524);
or U5666 (N_5666,N_5554,N_5507);
or U5667 (N_5667,N_5592,N_5500);
or U5668 (N_5668,N_5503,N_5567);
and U5669 (N_5669,N_5544,N_5566);
nor U5670 (N_5670,N_5520,N_5546);
or U5671 (N_5671,N_5532,N_5506);
or U5672 (N_5672,N_5591,N_5536);
xor U5673 (N_5673,N_5573,N_5524);
or U5674 (N_5674,N_5557,N_5599);
nand U5675 (N_5675,N_5571,N_5517);
or U5676 (N_5676,N_5596,N_5501);
nand U5677 (N_5677,N_5514,N_5527);
and U5678 (N_5678,N_5573,N_5543);
or U5679 (N_5679,N_5574,N_5527);
xor U5680 (N_5680,N_5585,N_5511);
or U5681 (N_5681,N_5584,N_5518);
nor U5682 (N_5682,N_5568,N_5584);
and U5683 (N_5683,N_5566,N_5508);
nand U5684 (N_5684,N_5577,N_5570);
nor U5685 (N_5685,N_5541,N_5523);
or U5686 (N_5686,N_5578,N_5554);
or U5687 (N_5687,N_5505,N_5540);
or U5688 (N_5688,N_5518,N_5553);
nor U5689 (N_5689,N_5568,N_5580);
and U5690 (N_5690,N_5558,N_5569);
nor U5691 (N_5691,N_5515,N_5570);
nand U5692 (N_5692,N_5512,N_5522);
and U5693 (N_5693,N_5535,N_5541);
xnor U5694 (N_5694,N_5575,N_5573);
xor U5695 (N_5695,N_5568,N_5517);
and U5696 (N_5696,N_5526,N_5557);
xor U5697 (N_5697,N_5558,N_5577);
nand U5698 (N_5698,N_5550,N_5582);
xnor U5699 (N_5699,N_5584,N_5556);
and U5700 (N_5700,N_5611,N_5606);
nand U5701 (N_5701,N_5616,N_5675);
and U5702 (N_5702,N_5655,N_5660);
or U5703 (N_5703,N_5625,N_5632);
nor U5704 (N_5704,N_5637,N_5644);
and U5705 (N_5705,N_5649,N_5638);
or U5706 (N_5706,N_5678,N_5605);
or U5707 (N_5707,N_5630,N_5610);
and U5708 (N_5708,N_5691,N_5657);
and U5709 (N_5709,N_5602,N_5696);
xor U5710 (N_5710,N_5658,N_5670);
nor U5711 (N_5711,N_5651,N_5667);
or U5712 (N_5712,N_5687,N_5623);
nand U5713 (N_5713,N_5618,N_5617);
and U5714 (N_5714,N_5626,N_5677);
and U5715 (N_5715,N_5604,N_5645);
nor U5716 (N_5716,N_5689,N_5662);
nand U5717 (N_5717,N_5674,N_5659);
xor U5718 (N_5718,N_5679,N_5698);
or U5719 (N_5719,N_5631,N_5682);
nand U5720 (N_5720,N_5614,N_5695);
xor U5721 (N_5721,N_5684,N_5664);
nand U5722 (N_5722,N_5633,N_5673);
and U5723 (N_5723,N_5676,N_5681);
nor U5724 (N_5724,N_5622,N_5671);
and U5725 (N_5725,N_5634,N_5619);
or U5726 (N_5726,N_5690,N_5652);
and U5727 (N_5727,N_5600,N_5686);
nand U5728 (N_5728,N_5680,N_5612);
or U5729 (N_5729,N_5646,N_5665);
nor U5730 (N_5730,N_5661,N_5685);
nand U5731 (N_5731,N_5615,N_5621);
nor U5732 (N_5732,N_5636,N_5663);
nand U5733 (N_5733,N_5643,N_5603);
or U5734 (N_5734,N_5628,N_5692);
and U5735 (N_5735,N_5647,N_5648);
nand U5736 (N_5736,N_5697,N_5607);
nor U5737 (N_5737,N_5627,N_5641);
and U5738 (N_5738,N_5653,N_5699);
or U5739 (N_5739,N_5683,N_5666);
xor U5740 (N_5740,N_5669,N_5629);
and U5741 (N_5741,N_5688,N_5693);
and U5742 (N_5742,N_5609,N_5601);
and U5743 (N_5743,N_5650,N_5608);
nand U5744 (N_5744,N_5640,N_5635);
or U5745 (N_5745,N_5620,N_5642);
nor U5746 (N_5746,N_5624,N_5654);
nor U5747 (N_5747,N_5613,N_5672);
nor U5748 (N_5748,N_5639,N_5694);
or U5749 (N_5749,N_5668,N_5656);
and U5750 (N_5750,N_5697,N_5663);
and U5751 (N_5751,N_5666,N_5641);
nor U5752 (N_5752,N_5648,N_5630);
or U5753 (N_5753,N_5678,N_5632);
nand U5754 (N_5754,N_5661,N_5669);
nor U5755 (N_5755,N_5605,N_5634);
and U5756 (N_5756,N_5635,N_5626);
or U5757 (N_5757,N_5671,N_5673);
and U5758 (N_5758,N_5676,N_5671);
and U5759 (N_5759,N_5619,N_5616);
and U5760 (N_5760,N_5672,N_5620);
or U5761 (N_5761,N_5630,N_5645);
nand U5762 (N_5762,N_5640,N_5672);
and U5763 (N_5763,N_5605,N_5614);
nand U5764 (N_5764,N_5639,N_5681);
nand U5765 (N_5765,N_5680,N_5653);
and U5766 (N_5766,N_5603,N_5611);
nor U5767 (N_5767,N_5635,N_5680);
or U5768 (N_5768,N_5642,N_5659);
nand U5769 (N_5769,N_5644,N_5679);
nor U5770 (N_5770,N_5637,N_5639);
or U5771 (N_5771,N_5665,N_5603);
nand U5772 (N_5772,N_5684,N_5668);
nand U5773 (N_5773,N_5622,N_5667);
nand U5774 (N_5774,N_5660,N_5600);
and U5775 (N_5775,N_5687,N_5625);
and U5776 (N_5776,N_5640,N_5665);
xnor U5777 (N_5777,N_5694,N_5647);
or U5778 (N_5778,N_5676,N_5608);
xor U5779 (N_5779,N_5652,N_5671);
nand U5780 (N_5780,N_5697,N_5647);
nand U5781 (N_5781,N_5675,N_5619);
or U5782 (N_5782,N_5693,N_5660);
nor U5783 (N_5783,N_5669,N_5647);
or U5784 (N_5784,N_5621,N_5671);
nor U5785 (N_5785,N_5614,N_5650);
or U5786 (N_5786,N_5652,N_5646);
nor U5787 (N_5787,N_5643,N_5628);
and U5788 (N_5788,N_5606,N_5676);
nor U5789 (N_5789,N_5635,N_5641);
nor U5790 (N_5790,N_5645,N_5624);
and U5791 (N_5791,N_5616,N_5615);
or U5792 (N_5792,N_5664,N_5652);
or U5793 (N_5793,N_5683,N_5638);
nor U5794 (N_5794,N_5676,N_5620);
or U5795 (N_5795,N_5630,N_5662);
nor U5796 (N_5796,N_5656,N_5601);
and U5797 (N_5797,N_5688,N_5697);
nand U5798 (N_5798,N_5695,N_5658);
and U5799 (N_5799,N_5689,N_5601);
nor U5800 (N_5800,N_5797,N_5744);
nor U5801 (N_5801,N_5747,N_5774);
and U5802 (N_5802,N_5746,N_5700);
or U5803 (N_5803,N_5734,N_5729);
or U5804 (N_5804,N_5712,N_5783);
nand U5805 (N_5805,N_5759,N_5788);
nand U5806 (N_5806,N_5726,N_5762);
nor U5807 (N_5807,N_5778,N_5754);
or U5808 (N_5808,N_5767,N_5764);
or U5809 (N_5809,N_5745,N_5785);
nor U5810 (N_5810,N_5756,N_5735);
and U5811 (N_5811,N_5707,N_5704);
nor U5812 (N_5812,N_5740,N_5776);
and U5813 (N_5813,N_5741,N_5793);
nand U5814 (N_5814,N_5718,N_5792);
and U5815 (N_5815,N_5781,N_5730);
or U5816 (N_5816,N_5722,N_5736);
and U5817 (N_5817,N_5703,N_5752);
and U5818 (N_5818,N_5705,N_5763);
or U5819 (N_5819,N_5782,N_5775);
nor U5820 (N_5820,N_5711,N_5766);
nor U5821 (N_5821,N_5780,N_5714);
and U5822 (N_5822,N_5749,N_5750);
nand U5823 (N_5823,N_5765,N_5768);
nand U5824 (N_5824,N_5738,N_5733);
and U5825 (N_5825,N_5739,N_5760);
xnor U5826 (N_5826,N_5732,N_5757);
nor U5827 (N_5827,N_5743,N_5779);
or U5828 (N_5828,N_5773,N_5710);
or U5829 (N_5829,N_5709,N_5701);
nand U5830 (N_5830,N_5784,N_5716);
xor U5831 (N_5831,N_5724,N_5795);
nor U5832 (N_5832,N_5708,N_5751);
nand U5833 (N_5833,N_5731,N_5723);
nand U5834 (N_5834,N_5758,N_5720);
and U5835 (N_5835,N_5748,N_5727);
and U5836 (N_5836,N_5799,N_5769);
nor U5837 (N_5837,N_5717,N_5786);
and U5838 (N_5838,N_5787,N_5753);
nor U5839 (N_5839,N_5702,N_5770);
nor U5840 (N_5840,N_5772,N_5728);
and U5841 (N_5841,N_5755,N_5777);
nor U5842 (N_5842,N_5790,N_5798);
and U5843 (N_5843,N_5713,N_5721);
nor U5844 (N_5844,N_5737,N_5706);
and U5845 (N_5845,N_5719,N_5789);
nand U5846 (N_5846,N_5761,N_5742);
nand U5847 (N_5847,N_5796,N_5771);
nand U5848 (N_5848,N_5791,N_5725);
xnor U5849 (N_5849,N_5715,N_5794);
nand U5850 (N_5850,N_5776,N_5736);
and U5851 (N_5851,N_5716,N_5760);
nand U5852 (N_5852,N_5722,N_5755);
nor U5853 (N_5853,N_5731,N_5790);
and U5854 (N_5854,N_5771,N_5749);
nand U5855 (N_5855,N_5705,N_5769);
and U5856 (N_5856,N_5733,N_5732);
and U5857 (N_5857,N_5759,N_5725);
or U5858 (N_5858,N_5715,N_5713);
nand U5859 (N_5859,N_5747,N_5716);
and U5860 (N_5860,N_5726,N_5775);
or U5861 (N_5861,N_5798,N_5704);
or U5862 (N_5862,N_5750,N_5738);
and U5863 (N_5863,N_5724,N_5727);
nor U5864 (N_5864,N_5770,N_5708);
xnor U5865 (N_5865,N_5742,N_5717);
and U5866 (N_5866,N_5794,N_5752);
and U5867 (N_5867,N_5730,N_5745);
nand U5868 (N_5868,N_5739,N_5772);
or U5869 (N_5869,N_5705,N_5751);
nor U5870 (N_5870,N_5704,N_5749);
or U5871 (N_5871,N_5733,N_5722);
and U5872 (N_5872,N_5776,N_5748);
and U5873 (N_5873,N_5764,N_5703);
nand U5874 (N_5874,N_5772,N_5753);
nor U5875 (N_5875,N_5731,N_5791);
or U5876 (N_5876,N_5736,N_5724);
and U5877 (N_5877,N_5776,N_5730);
or U5878 (N_5878,N_5758,N_5741);
nand U5879 (N_5879,N_5725,N_5777);
xor U5880 (N_5880,N_5757,N_5746);
and U5881 (N_5881,N_5736,N_5737);
and U5882 (N_5882,N_5730,N_5737);
nand U5883 (N_5883,N_5736,N_5767);
or U5884 (N_5884,N_5760,N_5735);
nor U5885 (N_5885,N_5730,N_5772);
nor U5886 (N_5886,N_5771,N_5756);
and U5887 (N_5887,N_5742,N_5702);
xor U5888 (N_5888,N_5742,N_5797);
or U5889 (N_5889,N_5748,N_5756);
nor U5890 (N_5890,N_5713,N_5743);
nand U5891 (N_5891,N_5702,N_5774);
and U5892 (N_5892,N_5757,N_5770);
nor U5893 (N_5893,N_5791,N_5771);
nand U5894 (N_5894,N_5729,N_5736);
nand U5895 (N_5895,N_5789,N_5721);
nand U5896 (N_5896,N_5738,N_5723);
nor U5897 (N_5897,N_5782,N_5798);
nand U5898 (N_5898,N_5795,N_5769);
nand U5899 (N_5899,N_5747,N_5794);
nand U5900 (N_5900,N_5841,N_5856);
nor U5901 (N_5901,N_5879,N_5885);
or U5902 (N_5902,N_5817,N_5823);
nand U5903 (N_5903,N_5897,N_5862);
xor U5904 (N_5904,N_5848,N_5826);
nor U5905 (N_5905,N_5873,N_5857);
or U5906 (N_5906,N_5800,N_5837);
nand U5907 (N_5907,N_5812,N_5859);
and U5908 (N_5908,N_5863,N_5819);
nand U5909 (N_5909,N_5836,N_5886);
nor U5910 (N_5910,N_5874,N_5840);
nand U5911 (N_5911,N_5811,N_5883);
nand U5912 (N_5912,N_5864,N_5843);
nor U5913 (N_5913,N_5896,N_5875);
nor U5914 (N_5914,N_5832,N_5894);
nand U5915 (N_5915,N_5866,N_5824);
and U5916 (N_5916,N_5818,N_5820);
and U5917 (N_5917,N_5816,N_5876);
nor U5918 (N_5918,N_5870,N_5880);
xor U5919 (N_5919,N_5833,N_5899);
or U5920 (N_5920,N_5829,N_5850);
nor U5921 (N_5921,N_5898,N_5821);
nor U5922 (N_5922,N_5893,N_5887);
nand U5923 (N_5923,N_5834,N_5828);
nor U5924 (N_5924,N_5854,N_5849);
and U5925 (N_5925,N_5889,N_5867);
and U5926 (N_5926,N_5804,N_5831);
xor U5927 (N_5927,N_5814,N_5861);
and U5928 (N_5928,N_5847,N_5835);
xor U5929 (N_5929,N_5860,N_5853);
nor U5930 (N_5930,N_5807,N_5822);
nor U5931 (N_5931,N_5810,N_5825);
or U5932 (N_5932,N_5808,N_5872);
nor U5933 (N_5933,N_5868,N_5844);
nand U5934 (N_5934,N_5881,N_5869);
or U5935 (N_5935,N_5882,N_5827);
nand U5936 (N_5936,N_5878,N_5851);
nand U5937 (N_5937,N_5813,N_5865);
nand U5938 (N_5938,N_5805,N_5888);
nor U5939 (N_5939,N_5855,N_5803);
and U5940 (N_5940,N_5801,N_5895);
and U5941 (N_5941,N_5892,N_5842);
and U5942 (N_5942,N_5838,N_5815);
and U5943 (N_5943,N_5839,N_5877);
and U5944 (N_5944,N_5802,N_5830);
and U5945 (N_5945,N_5890,N_5806);
and U5946 (N_5946,N_5845,N_5891);
nor U5947 (N_5947,N_5852,N_5884);
or U5948 (N_5948,N_5858,N_5871);
and U5949 (N_5949,N_5809,N_5846);
nand U5950 (N_5950,N_5801,N_5865);
and U5951 (N_5951,N_5835,N_5848);
or U5952 (N_5952,N_5869,N_5823);
or U5953 (N_5953,N_5879,N_5882);
nor U5954 (N_5954,N_5841,N_5850);
nand U5955 (N_5955,N_5849,N_5800);
xor U5956 (N_5956,N_5837,N_5852);
nor U5957 (N_5957,N_5880,N_5891);
nor U5958 (N_5958,N_5865,N_5860);
nand U5959 (N_5959,N_5828,N_5820);
xnor U5960 (N_5960,N_5844,N_5872);
nor U5961 (N_5961,N_5892,N_5879);
nand U5962 (N_5962,N_5821,N_5883);
or U5963 (N_5963,N_5864,N_5880);
nor U5964 (N_5964,N_5854,N_5868);
and U5965 (N_5965,N_5839,N_5893);
and U5966 (N_5966,N_5864,N_5845);
nor U5967 (N_5967,N_5899,N_5894);
xor U5968 (N_5968,N_5845,N_5859);
or U5969 (N_5969,N_5846,N_5865);
and U5970 (N_5970,N_5877,N_5824);
nor U5971 (N_5971,N_5802,N_5885);
xnor U5972 (N_5972,N_5804,N_5814);
or U5973 (N_5973,N_5871,N_5850);
nand U5974 (N_5974,N_5804,N_5875);
and U5975 (N_5975,N_5815,N_5839);
or U5976 (N_5976,N_5879,N_5807);
nand U5977 (N_5977,N_5855,N_5887);
xnor U5978 (N_5978,N_5819,N_5852);
nand U5979 (N_5979,N_5803,N_5825);
nand U5980 (N_5980,N_5837,N_5858);
or U5981 (N_5981,N_5834,N_5847);
nand U5982 (N_5982,N_5846,N_5845);
nand U5983 (N_5983,N_5825,N_5855);
or U5984 (N_5984,N_5878,N_5870);
xnor U5985 (N_5985,N_5824,N_5834);
or U5986 (N_5986,N_5850,N_5849);
nor U5987 (N_5987,N_5820,N_5870);
nor U5988 (N_5988,N_5811,N_5815);
xor U5989 (N_5989,N_5848,N_5881);
nor U5990 (N_5990,N_5830,N_5825);
or U5991 (N_5991,N_5808,N_5825);
or U5992 (N_5992,N_5837,N_5878);
or U5993 (N_5993,N_5886,N_5842);
or U5994 (N_5994,N_5833,N_5818);
nand U5995 (N_5995,N_5861,N_5842);
or U5996 (N_5996,N_5894,N_5843);
or U5997 (N_5997,N_5806,N_5874);
or U5998 (N_5998,N_5868,N_5846);
nor U5999 (N_5999,N_5881,N_5835);
and U6000 (N_6000,N_5960,N_5962);
or U6001 (N_6001,N_5991,N_5986);
xnor U6002 (N_6002,N_5992,N_5993);
and U6003 (N_6003,N_5952,N_5908);
nor U6004 (N_6004,N_5968,N_5983);
or U6005 (N_6005,N_5918,N_5917);
and U6006 (N_6006,N_5916,N_5940);
nand U6007 (N_6007,N_5963,N_5927);
nand U6008 (N_6008,N_5928,N_5939);
xor U6009 (N_6009,N_5921,N_5988);
xnor U6010 (N_6010,N_5914,N_5995);
and U6011 (N_6011,N_5965,N_5910);
or U6012 (N_6012,N_5959,N_5938);
nand U6013 (N_6013,N_5957,N_5905);
and U6014 (N_6014,N_5976,N_5947);
or U6015 (N_6015,N_5904,N_5943);
nor U6016 (N_6016,N_5982,N_5901);
and U6017 (N_6017,N_5969,N_5989);
and U6018 (N_6018,N_5998,N_5966);
nand U6019 (N_6019,N_5984,N_5937);
nand U6020 (N_6020,N_5994,N_5941);
nand U6021 (N_6021,N_5932,N_5931);
xnor U6022 (N_6022,N_5985,N_5956);
and U6023 (N_6023,N_5949,N_5946);
nand U6024 (N_6024,N_5999,N_5955);
or U6025 (N_6025,N_5922,N_5974);
or U6026 (N_6026,N_5951,N_5944);
and U6027 (N_6027,N_5933,N_5923);
or U6028 (N_6028,N_5906,N_5913);
nor U6029 (N_6029,N_5911,N_5924);
xor U6030 (N_6030,N_5996,N_5990);
or U6031 (N_6031,N_5971,N_5981);
and U6032 (N_6032,N_5978,N_5970);
or U6033 (N_6033,N_5934,N_5958);
or U6034 (N_6034,N_5907,N_5987);
nand U6035 (N_6035,N_5936,N_5920);
nand U6036 (N_6036,N_5961,N_5953);
xor U6037 (N_6037,N_5919,N_5972);
nor U6038 (N_6038,N_5997,N_5950);
or U6039 (N_6039,N_5980,N_5929);
nor U6040 (N_6040,N_5973,N_5954);
nand U6041 (N_6041,N_5926,N_5900);
or U6042 (N_6042,N_5964,N_5903);
nor U6043 (N_6043,N_5915,N_5977);
nand U6044 (N_6044,N_5912,N_5967);
and U6045 (N_6045,N_5925,N_5909);
and U6046 (N_6046,N_5942,N_5902);
nand U6047 (N_6047,N_5935,N_5979);
nor U6048 (N_6048,N_5945,N_5948);
nor U6049 (N_6049,N_5975,N_5930);
xor U6050 (N_6050,N_5926,N_5949);
or U6051 (N_6051,N_5989,N_5922);
nor U6052 (N_6052,N_5977,N_5964);
or U6053 (N_6053,N_5919,N_5974);
nor U6054 (N_6054,N_5970,N_5905);
nand U6055 (N_6055,N_5983,N_5989);
nor U6056 (N_6056,N_5913,N_5975);
nand U6057 (N_6057,N_5974,N_5902);
nand U6058 (N_6058,N_5903,N_5975);
or U6059 (N_6059,N_5985,N_5981);
nand U6060 (N_6060,N_5945,N_5940);
nor U6061 (N_6061,N_5994,N_5911);
or U6062 (N_6062,N_5975,N_5989);
and U6063 (N_6063,N_5945,N_5967);
xnor U6064 (N_6064,N_5960,N_5900);
and U6065 (N_6065,N_5958,N_5976);
or U6066 (N_6066,N_5992,N_5994);
nor U6067 (N_6067,N_5967,N_5924);
nor U6068 (N_6068,N_5929,N_5983);
nor U6069 (N_6069,N_5932,N_5905);
and U6070 (N_6070,N_5947,N_5988);
and U6071 (N_6071,N_5976,N_5908);
and U6072 (N_6072,N_5942,N_5925);
or U6073 (N_6073,N_5998,N_5980);
nor U6074 (N_6074,N_5997,N_5906);
nand U6075 (N_6075,N_5997,N_5908);
and U6076 (N_6076,N_5912,N_5986);
or U6077 (N_6077,N_5992,N_5938);
or U6078 (N_6078,N_5926,N_5907);
xnor U6079 (N_6079,N_5990,N_5925);
nand U6080 (N_6080,N_5921,N_5964);
or U6081 (N_6081,N_5961,N_5989);
xnor U6082 (N_6082,N_5992,N_5959);
xor U6083 (N_6083,N_5911,N_5955);
and U6084 (N_6084,N_5951,N_5964);
xor U6085 (N_6085,N_5922,N_5929);
and U6086 (N_6086,N_5986,N_5932);
and U6087 (N_6087,N_5986,N_5985);
nand U6088 (N_6088,N_5989,N_5982);
or U6089 (N_6089,N_5943,N_5972);
xnor U6090 (N_6090,N_5905,N_5943);
xor U6091 (N_6091,N_5984,N_5906);
nand U6092 (N_6092,N_5937,N_5947);
nand U6093 (N_6093,N_5946,N_5972);
nand U6094 (N_6094,N_5925,N_5991);
nor U6095 (N_6095,N_5976,N_5985);
xnor U6096 (N_6096,N_5919,N_5979);
nand U6097 (N_6097,N_5914,N_5942);
nor U6098 (N_6098,N_5968,N_5921);
nand U6099 (N_6099,N_5929,N_5958);
and U6100 (N_6100,N_6001,N_6055);
and U6101 (N_6101,N_6056,N_6087);
xor U6102 (N_6102,N_6060,N_6019);
or U6103 (N_6103,N_6012,N_6070);
nand U6104 (N_6104,N_6036,N_6043);
and U6105 (N_6105,N_6091,N_6015);
nand U6106 (N_6106,N_6008,N_6089);
nor U6107 (N_6107,N_6074,N_6052);
xor U6108 (N_6108,N_6062,N_6026);
nor U6109 (N_6109,N_6025,N_6009);
nor U6110 (N_6110,N_6076,N_6078);
nor U6111 (N_6111,N_6046,N_6048);
nand U6112 (N_6112,N_6040,N_6013);
xor U6113 (N_6113,N_6083,N_6094);
nor U6114 (N_6114,N_6017,N_6051);
and U6115 (N_6115,N_6058,N_6042);
xor U6116 (N_6116,N_6098,N_6059);
and U6117 (N_6117,N_6080,N_6086);
nand U6118 (N_6118,N_6095,N_6049);
or U6119 (N_6119,N_6021,N_6081);
and U6120 (N_6120,N_6041,N_6023);
and U6121 (N_6121,N_6084,N_6085);
or U6122 (N_6122,N_6016,N_6075);
and U6123 (N_6123,N_6011,N_6033);
and U6124 (N_6124,N_6037,N_6050);
and U6125 (N_6125,N_6020,N_6027);
nand U6126 (N_6126,N_6096,N_6018);
or U6127 (N_6127,N_6079,N_6038);
nor U6128 (N_6128,N_6061,N_6082);
nor U6129 (N_6129,N_6093,N_6031);
or U6130 (N_6130,N_6006,N_6063);
or U6131 (N_6131,N_6088,N_6034);
nand U6132 (N_6132,N_6092,N_6028);
xnor U6133 (N_6133,N_6029,N_6090);
nor U6134 (N_6134,N_6053,N_6054);
nand U6135 (N_6135,N_6064,N_6071);
or U6136 (N_6136,N_6068,N_6072);
nor U6137 (N_6137,N_6000,N_6099);
nand U6138 (N_6138,N_6057,N_6069);
nor U6139 (N_6139,N_6066,N_6045);
nand U6140 (N_6140,N_6097,N_6044);
nor U6141 (N_6141,N_6003,N_6039);
nand U6142 (N_6142,N_6005,N_6065);
xnor U6143 (N_6143,N_6024,N_6067);
nand U6144 (N_6144,N_6007,N_6030);
nand U6145 (N_6145,N_6077,N_6022);
nor U6146 (N_6146,N_6073,N_6010);
nand U6147 (N_6147,N_6035,N_6004);
nand U6148 (N_6148,N_6002,N_6014);
or U6149 (N_6149,N_6032,N_6047);
nor U6150 (N_6150,N_6092,N_6029);
nand U6151 (N_6151,N_6028,N_6090);
nor U6152 (N_6152,N_6023,N_6091);
nor U6153 (N_6153,N_6023,N_6075);
nor U6154 (N_6154,N_6029,N_6088);
nand U6155 (N_6155,N_6036,N_6019);
nand U6156 (N_6156,N_6056,N_6010);
nand U6157 (N_6157,N_6008,N_6043);
and U6158 (N_6158,N_6017,N_6047);
xnor U6159 (N_6159,N_6096,N_6036);
nand U6160 (N_6160,N_6000,N_6049);
nand U6161 (N_6161,N_6070,N_6004);
nor U6162 (N_6162,N_6071,N_6053);
nand U6163 (N_6163,N_6002,N_6029);
nand U6164 (N_6164,N_6084,N_6094);
or U6165 (N_6165,N_6062,N_6018);
nor U6166 (N_6166,N_6031,N_6084);
nand U6167 (N_6167,N_6072,N_6073);
or U6168 (N_6168,N_6026,N_6008);
or U6169 (N_6169,N_6044,N_6059);
nand U6170 (N_6170,N_6071,N_6006);
xor U6171 (N_6171,N_6097,N_6000);
nor U6172 (N_6172,N_6059,N_6065);
and U6173 (N_6173,N_6013,N_6069);
and U6174 (N_6174,N_6018,N_6006);
or U6175 (N_6175,N_6011,N_6084);
or U6176 (N_6176,N_6033,N_6006);
nor U6177 (N_6177,N_6062,N_6076);
nand U6178 (N_6178,N_6082,N_6039);
or U6179 (N_6179,N_6004,N_6087);
and U6180 (N_6180,N_6062,N_6028);
nand U6181 (N_6181,N_6021,N_6072);
xnor U6182 (N_6182,N_6006,N_6009);
or U6183 (N_6183,N_6088,N_6044);
xnor U6184 (N_6184,N_6013,N_6070);
or U6185 (N_6185,N_6017,N_6009);
nor U6186 (N_6186,N_6007,N_6065);
nor U6187 (N_6187,N_6033,N_6016);
and U6188 (N_6188,N_6044,N_6015);
nor U6189 (N_6189,N_6066,N_6074);
or U6190 (N_6190,N_6087,N_6034);
and U6191 (N_6191,N_6092,N_6051);
or U6192 (N_6192,N_6099,N_6067);
and U6193 (N_6193,N_6091,N_6088);
nor U6194 (N_6194,N_6086,N_6059);
and U6195 (N_6195,N_6083,N_6086);
and U6196 (N_6196,N_6066,N_6008);
nand U6197 (N_6197,N_6020,N_6057);
and U6198 (N_6198,N_6076,N_6051);
or U6199 (N_6199,N_6070,N_6066);
and U6200 (N_6200,N_6174,N_6181);
nand U6201 (N_6201,N_6185,N_6175);
and U6202 (N_6202,N_6121,N_6131);
nand U6203 (N_6203,N_6178,N_6106);
nor U6204 (N_6204,N_6173,N_6136);
xnor U6205 (N_6205,N_6144,N_6129);
and U6206 (N_6206,N_6114,N_6192);
or U6207 (N_6207,N_6111,N_6142);
nor U6208 (N_6208,N_6120,N_6145);
and U6209 (N_6209,N_6118,N_6198);
nand U6210 (N_6210,N_6119,N_6189);
and U6211 (N_6211,N_6128,N_6122);
and U6212 (N_6212,N_6127,N_6191);
or U6213 (N_6213,N_6133,N_6168);
or U6214 (N_6214,N_6182,N_6167);
nor U6215 (N_6215,N_6154,N_6170);
nor U6216 (N_6216,N_6140,N_6103);
and U6217 (N_6217,N_6172,N_6196);
or U6218 (N_6218,N_6148,N_6125);
or U6219 (N_6219,N_6104,N_6108);
nor U6220 (N_6220,N_6153,N_6187);
nand U6221 (N_6221,N_6179,N_6156);
or U6222 (N_6222,N_6116,N_6124);
nand U6223 (N_6223,N_6162,N_6183);
and U6224 (N_6224,N_6161,N_6113);
nand U6225 (N_6225,N_6107,N_6177);
nand U6226 (N_6226,N_6115,N_6110);
nor U6227 (N_6227,N_6195,N_6188);
or U6228 (N_6228,N_6130,N_6147);
nand U6229 (N_6229,N_6180,N_6126);
or U6230 (N_6230,N_6109,N_6151);
or U6231 (N_6231,N_6143,N_6135);
nand U6232 (N_6232,N_6163,N_6141);
nor U6233 (N_6233,N_6197,N_6102);
or U6234 (N_6234,N_6164,N_6123);
or U6235 (N_6235,N_6112,N_6134);
nand U6236 (N_6236,N_6165,N_6194);
nor U6237 (N_6237,N_6160,N_6159);
nand U6238 (N_6238,N_6166,N_6138);
nor U6239 (N_6239,N_6139,N_6199);
or U6240 (N_6240,N_6186,N_6150);
nor U6241 (N_6241,N_6152,N_6193);
xnor U6242 (N_6242,N_6101,N_6169);
or U6243 (N_6243,N_6157,N_6190);
nand U6244 (N_6244,N_6100,N_6137);
nor U6245 (N_6245,N_6158,N_6105);
nor U6246 (N_6246,N_6176,N_6184);
or U6247 (N_6247,N_6171,N_6132);
nand U6248 (N_6248,N_6146,N_6149);
xnor U6249 (N_6249,N_6155,N_6117);
nand U6250 (N_6250,N_6171,N_6121);
or U6251 (N_6251,N_6110,N_6152);
nand U6252 (N_6252,N_6111,N_6140);
and U6253 (N_6253,N_6152,N_6183);
or U6254 (N_6254,N_6164,N_6196);
nor U6255 (N_6255,N_6146,N_6113);
nand U6256 (N_6256,N_6147,N_6166);
and U6257 (N_6257,N_6146,N_6179);
and U6258 (N_6258,N_6160,N_6193);
or U6259 (N_6259,N_6181,N_6175);
xor U6260 (N_6260,N_6198,N_6147);
and U6261 (N_6261,N_6126,N_6157);
or U6262 (N_6262,N_6158,N_6173);
nor U6263 (N_6263,N_6134,N_6184);
nand U6264 (N_6264,N_6177,N_6111);
nand U6265 (N_6265,N_6138,N_6195);
nand U6266 (N_6266,N_6198,N_6129);
nand U6267 (N_6267,N_6184,N_6143);
nand U6268 (N_6268,N_6116,N_6189);
or U6269 (N_6269,N_6118,N_6148);
and U6270 (N_6270,N_6190,N_6108);
and U6271 (N_6271,N_6199,N_6172);
or U6272 (N_6272,N_6101,N_6191);
or U6273 (N_6273,N_6173,N_6182);
xor U6274 (N_6274,N_6107,N_6172);
and U6275 (N_6275,N_6155,N_6125);
or U6276 (N_6276,N_6121,N_6130);
nand U6277 (N_6277,N_6160,N_6142);
nand U6278 (N_6278,N_6136,N_6109);
or U6279 (N_6279,N_6118,N_6106);
nand U6280 (N_6280,N_6133,N_6130);
nor U6281 (N_6281,N_6159,N_6168);
nor U6282 (N_6282,N_6195,N_6100);
and U6283 (N_6283,N_6113,N_6157);
and U6284 (N_6284,N_6189,N_6177);
and U6285 (N_6285,N_6198,N_6179);
or U6286 (N_6286,N_6140,N_6112);
or U6287 (N_6287,N_6147,N_6101);
nor U6288 (N_6288,N_6150,N_6107);
nand U6289 (N_6289,N_6157,N_6103);
nand U6290 (N_6290,N_6161,N_6120);
nand U6291 (N_6291,N_6126,N_6134);
xnor U6292 (N_6292,N_6185,N_6197);
nor U6293 (N_6293,N_6125,N_6192);
nor U6294 (N_6294,N_6163,N_6192);
nand U6295 (N_6295,N_6145,N_6196);
and U6296 (N_6296,N_6187,N_6182);
nand U6297 (N_6297,N_6120,N_6134);
or U6298 (N_6298,N_6165,N_6110);
nor U6299 (N_6299,N_6108,N_6142);
and U6300 (N_6300,N_6252,N_6200);
and U6301 (N_6301,N_6211,N_6244);
or U6302 (N_6302,N_6268,N_6229);
or U6303 (N_6303,N_6223,N_6214);
nand U6304 (N_6304,N_6277,N_6243);
and U6305 (N_6305,N_6248,N_6296);
xnor U6306 (N_6306,N_6208,N_6276);
nor U6307 (N_6307,N_6215,N_6281);
or U6308 (N_6308,N_6267,N_6206);
nand U6309 (N_6309,N_6201,N_6263);
nor U6310 (N_6310,N_6259,N_6235);
and U6311 (N_6311,N_6234,N_6290);
nand U6312 (N_6312,N_6239,N_6210);
nor U6313 (N_6313,N_6291,N_6212);
or U6314 (N_6314,N_6240,N_6288);
nor U6315 (N_6315,N_6238,N_6219);
nand U6316 (N_6316,N_6286,N_6285);
and U6317 (N_6317,N_6230,N_6204);
and U6318 (N_6318,N_6292,N_6287);
nor U6319 (N_6319,N_6218,N_6258);
nand U6320 (N_6320,N_6222,N_6203);
or U6321 (N_6321,N_6241,N_6233);
and U6322 (N_6322,N_6272,N_6246);
and U6323 (N_6323,N_6298,N_6250);
and U6324 (N_6324,N_6217,N_6232);
or U6325 (N_6325,N_6245,N_6236);
and U6326 (N_6326,N_6265,N_6266);
or U6327 (N_6327,N_6224,N_6255);
and U6328 (N_6328,N_6269,N_6271);
nor U6329 (N_6329,N_6247,N_6216);
or U6330 (N_6330,N_6284,N_6279);
nor U6331 (N_6331,N_6270,N_6221);
and U6332 (N_6332,N_6228,N_6282);
nor U6333 (N_6333,N_6262,N_6294);
nand U6334 (N_6334,N_6205,N_6249);
nand U6335 (N_6335,N_6227,N_6209);
or U6336 (N_6336,N_6251,N_6220);
nor U6337 (N_6337,N_6280,N_6256);
or U6338 (N_6338,N_6295,N_6231);
nor U6339 (N_6339,N_6260,N_6299);
or U6340 (N_6340,N_6297,N_6264);
or U6341 (N_6341,N_6278,N_6213);
xnor U6342 (N_6342,N_6237,N_6261);
and U6343 (N_6343,N_6275,N_6253);
nor U6344 (N_6344,N_6273,N_6202);
or U6345 (N_6345,N_6242,N_6226);
nor U6346 (N_6346,N_6225,N_6254);
nor U6347 (N_6347,N_6274,N_6207);
nor U6348 (N_6348,N_6283,N_6289);
or U6349 (N_6349,N_6257,N_6293);
and U6350 (N_6350,N_6232,N_6261);
nand U6351 (N_6351,N_6285,N_6252);
nor U6352 (N_6352,N_6214,N_6244);
and U6353 (N_6353,N_6260,N_6215);
nor U6354 (N_6354,N_6275,N_6278);
xor U6355 (N_6355,N_6207,N_6215);
and U6356 (N_6356,N_6204,N_6227);
xnor U6357 (N_6357,N_6218,N_6207);
nor U6358 (N_6358,N_6254,N_6224);
nand U6359 (N_6359,N_6230,N_6290);
or U6360 (N_6360,N_6275,N_6202);
nor U6361 (N_6361,N_6262,N_6256);
nor U6362 (N_6362,N_6271,N_6299);
or U6363 (N_6363,N_6296,N_6278);
nor U6364 (N_6364,N_6283,N_6278);
nand U6365 (N_6365,N_6273,N_6231);
nor U6366 (N_6366,N_6217,N_6241);
and U6367 (N_6367,N_6254,N_6281);
nor U6368 (N_6368,N_6256,N_6206);
nand U6369 (N_6369,N_6238,N_6216);
and U6370 (N_6370,N_6293,N_6200);
nor U6371 (N_6371,N_6264,N_6224);
nand U6372 (N_6372,N_6224,N_6231);
nand U6373 (N_6373,N_6269,N_6275);
nor U6374 (N_6374,N_6245,N_6239);
xnor U6375 (N_6375,N_6231,N_6293);
nand U6376 (N_6376,N_6209,N_6270);
nor U6377 (N_6377,N_6273,N_6209);
or U6378 (N_6378,N_6286,N_6209);
or U6379 (N_6379,N_6233,N_6276);
and U6380 (N_6380,N_6230,N_6243);
or U6381 (N_6381,N_6210,N_6201);
and U6382 (N_6382,N_6268,N_6226);
nand U6383 (N_6383,N_6234,N_6229);
or U6384 (N_6384,N_6274,N_6247);
or U6385 (N_6385,N_6266,N_6228);
or U6386 (N_6386,N_6244,N_6297);
nor U6387 (N_6387,N_6275,N_6246);
nand U6388 (N_6388,N_6226,N_6286);
nand U6389 (N_6389,N_6211,N_6282);
nor U6390 (N_6390,N_6201,N_6279);
or U6391 (N_6391,N_6212,N_6202);
or U6392 (N_6392,N_6242,N_6209);
and U6393 (N_6393,N_6252,N_6240);
nand U6394 (N_6394,N_6200,N_6204);
xnor U6395 (N_6395,N_6297,N_6256);
nand U6396 (N_6396,N_6228,N_6275);
nor U6397 (N_6397,N_6289,N_6247);
nand U6398 (N_6398,N_6243,N_6257);
or U6399 (N_6399,N_6212,N_6235);
xor U6400 (N_6400,N_6353,N_6380);
and U6401 (N_6401,N_6361,N_6317);
nor U6402 (N_6402,N_6392,N_6347);
nand U6403 (N_6403,N_6391,N_6388);
nor U6404 (N_6404,N_6372,N_6377);
nand U6405 (N_6405,N_6384,N_6370);
nand U6406 (N_6406,N_6333,N_6307);
or U6407 (N_6407,N_6332,N_6302);
xnor U6408 (N_6408,N_6312,N_6327);
xnor U6409 (N_6409,N_6330,N_6357);
nor U6410 (N_6410,N_6321,N_6319);
or U6411 (N_6411,N_6364,N_6356);
xnor U6412 (N_6412,N_6352,N_6366);
nand U6413 (N_6413,N_6395,N_6315);
nor U6414 (N_6414,N_6320,N_6339);
nand U6415 (N_6415,N_6371,N_6351);
or U6416 (N_6416,N_6349,N_6382);
nor U6417 (N_6417,N_6341,N_6399);
and U6418 (N_6418,N_6304,N_6363);
and U6419 (N_6419,N_6335,N_6389);
and U6420 (N_6420,N_6331,N_6368);
or U6421 (N_6421,N_6326,N_6369);
or U6422 (N_6422,N_6311,N_6316);
nor U6423 (N_6423,N_6359,N_6346);
nor U6424 (N_6424,N_6367,N_6398);
xnor U6425 (N_6425,N_6314,N_6378);
xor U6426 (N_6426,N_6343,N_6325);
xnor U6427 (N_6427,N_6387,N_6396);
nor U6428 (N_6428,N_6334,N_6358);
xnor U6429 (N_6429,N_6328,N_6375);
and U6430 (N_6430,N_6301,N_6303);
or U6431 (N_6431,N_6348,N_6338);
and U6432 (N_6432,N_6362,N_6322);
nor U6433 (N_6433,N_6374,N_6365);
nor U6434 (N_6434,N_6324,N_6323);
or U6435 (N_6435,N_6397,N_6390);
nor U6436 (N_6436,N_6393,N_6305);
and U6437 (N_6437,N_6342,N_6376);
and U6438 (N_6438,N_6373,N_6360);
or U6439 (N_6439,N_6394,N_6329);
nor U6440 (N_6440,N_6385,N_6354);
xnor U6441 (N_6441,N_6306,N_6386);
nor U6442 (N_6442,N_6381,N_6355);
and U6443 (N_6443,N_6340,N_6336);
xor U6444 (N_6444,N_6300,N_6379);
and U6445 (N_6445,N_6318,N_6309);
and U6446 (N_6446,N_6337,N_6344);
and U6447 (N_6447,N_6350,N_6313);
and U6448 (N_6448,N_6345,N_6308);
nor U6449 (N_6449,N_6310,N_6383);
xor U6450 (N_6450,N_6373,N_6320);
nor U6451 (N_6451,N_6333,N_6341);
and U6452 (N_6452,N_6324,N_6361);
nor U6453 (N_6453,N_6362,N_6316);
nor U6454 (N_6454,N_6303,N_6357);
nand U6455 (N_6455,N_6360,N_6348);
nor U6456 (N_6456,N_6398,N_6358);
nor U6457 (N_6457,N_6377,N_6362);
nand U6458 (N_6458,N_6363,N_6300);
xnor U6459 (N_6459,N_6371,N_6301);
nor U6460 (N_6460,N_6353,N_6318);
or U6461 (N_6461,N_6315,N_6351);
and U6462 (N_6462,N_6330,N_6399);
nor U6463 (N_6463,N_6391,N_6315);
or U6464 (N_6464,N_6347,N_6321);
and U6465 (N_6465,N_6343,N_6356);
nand U6466 (N_6466,N_6363,N_6373);
nand U6467 (N_6467,N_6310,N_6384);
nor U6468 (N_6468,N_6309,N_6358);
nand U6469 (N_6469,N_6332,N_6320);
nor U6470 (N_6470,N_6305,N_6374);
nor U6471 (N_6471,N_6327,N_6369);
nand U6472 (N_6472,N_6323,N_6314);
nor U6473 (N_6473,N_6398,N_6355);
or U6474 (N_6474,N_6396,N_6353);
nand U6475 (N_6475,N_6329,N_6361);
xor U6476 (N_6476,N_6369,N_6334);
nor U6477 (N_6477,N_6300,N_6359);
and U6478 (N_6478,N_6352,N_6334);
nor U6479 (N_6479,N_6356,N_6374);
nor U6480 (N_6480,N_6349,N_6343);
xor U6481 (N_6481,N_6376,N_6372);
and U6482 (N_6482,N_6381,N_6360);
nand U6483 (N_6483,N_6362,N_6351);
nor U6484 (N_6484,N_6359,N_6382);
or U6485 (N_6485,N_6313,N_6330);
and U6486 (N_6486,N_6355,N_6346);
nor U6487 (N_6487,N_6335,N_6340);
nor U6488 (N_6488,N_6396,N_6364);
and U6489 (N_6489,N_6300,N_6323);
xnor U6490 (N_6490,N_6380,N_6379);
and U6491 (N_6491,N_6387,N_6336);
and U6492 (N_6492,N_6301,N_6347);
nand U6493 (N_6493,N_6323,N_6308);
nand U6494 (N_6494,N_6391,N_6381);
or U6495 (N_6495,N_6362,N_6386);
nor U6496 (N_6496,N_6342,N_6337);
nor U6497 (N_6497,N_6345,N_6356);
or U6498 (N_6498,N_6316,N_6378);
or U6499 (N_6499,N_6326,N_6360);
nand U6500 (N_6500,N_6483,N_6406);
nand U6501 (N_6501,N_6442,N_6436);
or U6502 (N_6502,N_6461,N_6487);
xnor U6503 (N_6503,N_6451,N_6429);
and U6504 (N_6504,N_6493,N_6432);
and U6505 (N_6505,N_6481,N_6486);
and U6506 (N_6506,N_6435,N_6467);
nor U6507 (N_6507,N_6434,N_6413);
or U6508 (N_6508,N_6439,N_6446);
nor U6509 (N_6509,N_6407,N_6460);
xnor U6510 (N_6510,N_6492,N_6458);
nand U6511 (N_6511,N_6482,N_6445);
or U6512 (N_6512,N_6449,N_6447);
and U6513 (N_6513,N_6485,N_6465);
nand U6514 (N_6514,N_6433,N_6471);
nand U6515 (N_6515,N_6414,N_6453);
nor U6516 (N_6516,N_6480,N_6416);
nor U6517 (N_6517,N_6495,N_6464);
nand U6518 (N_6518,N_6424,N_6450);
nor U6519 (N_6519,N_6409,N_6468);
xnor U6520 (N_6520,N_6403,N_6420);
nand U6521 (N_6521,N_6473,N_6422);
xor U6522 (N_6522,N_6443,N_6497);
and U6523 (N_6523,N_6428,N_6425);
and U6524 (N_6524,N_6401,N_6457);
nand U6525 (N_6525,N_6417,N_6455);
or U6526 (N_6526,N_6421,N_6454);
or U6527 (N_6527,N_6459,N_6405);
nor U6528 (N_6528,N_6489,N_6476);
nand U6529 (N_6529,N_6404,N_6470);
nand U6530 (N_6530,N_6430,N_6415);
and U6531 (N_6531,N_6426,N_6466);
or U6532 (N_6532,N_6488,N_6494);
or U6533 (N_6533,N_6469,N_6478);
and U6534 (N_6534,N_6498,N_6472);
and U6535 (N_6535,N_6477,N_6423);
and U6536 (N_6536,N_6400,N_6463);
nand U6537 (N_6537,N_6475,N_6419);
nor U6538 (N_6538,N_6499,N_6490);
and U6539 (N_6539,N_6411,N_6456);
and U6540 (N_6540,N_6448,N_6479);
and U6541 (N_6541,N_6484,N_6431);
and U6542 (N_6542,N_6412,N_6441);
nand U6543 (N_6543,N_6491,N_6418);
nand U6544 (N_6544,N_6402,N_6410);
and U6545 (N_6545,N_6462,N_6408);
or U6546 (N_6546,N_6474,N_6444);
nand U6547 (N_6547,N_6452,N_6440);
nand U6548 (N_6548,N_6427,N_6438);
or U6549 (N_6549,N_6437,N_6496);
nand U6550 (N_6550,N_6410,N_6491);
and U6551 (N_6551,N_6415,N_6412);
or U6552 (N_6552,N_6480,N_6447);
or U6553 (N_6553,N_6495,N_6424);
nor U6554 (N_6554,N_6403,N_6466);
and U6555 (N_6555,N_6415,N_6433);
nand U6556 (N_6556,N_6479,N_6486);
or U6557 (N_6557,N_6453,N_6441);
nand U6558 (N_6558,N_6445,N_6475);
and U6559 (N_6559,N_6464,N_6480);
xnor U6560 (N_6560,N_6406,N_6455);
and U6561 (N_6561,N_6450,N_6481);
and U6562 (N_6562,N_6420,N_6452);
nor U6563 (N_6563,N_6439,N_6426);
nor U6564 (N_6564,N_6499,N_6482);
and U6565 (N_6565,N_6483,N_6484);
xor U6566 (N_6566,N_6472,N_6414);
and U6567 (N_6567,N_6425,N_6467);
and U6568 (N_6568,N_6486,N_6428);
or U6569 (N_6569,N_6457,N_6460);
and U6570 (N_6570,N_6488,N_6417);
nor U6571 (N_6571,N_6402,N_6419);
nor U6572 (N_6572,N_6495,N_6406);
or U6573 (N_6573,N_6478,N_6425);
or U6574 (N_6574,N_6491,N_6499);
and U6575 (N_6575,N_6409,N_6486);
nand U6576 (N_6576,N_6471,N_6406);
and U6577 (N_6577,N_6485,N_6403);
nor U6578 (N_6578,N_6437,N_6482);
nand U6579 (N_6579,N_6421,N_6480);
nand U6580 (N_6580,N_6481,N_6457);
nor U6581 (N_6581,N_6492,N_6431);
and U6582 (N_6582,N_6497,N_6421);
xnor U6583 (N_6583,N_6492,N_6475);
nand U6584 (N_6584,N_6431,N_6481);
nand U6585 (N_6585,N_6435,N_6446);
nand U6586 (N_6586,N_6427,N_6472);
nor U6587 (N_6587,N_6472,N_6433);
nor U6588 (N_6588,N_6422,N_6423);
or U6589 (N_6589,N_6465,N_6408);
or U6590 (N_6590,N_6458,N_6437);
nand U6591 (N_6591,N_6414,N_6468);
and U6592 (N_6592,N_6494,N_6476);
or U6593 (N_6593,N_6433,N_6430);
nand U6594 (N_6594,N_6419,N_6454);
nor U6595 (N_6595,N_6434,N_6402);
or U6596 (N_6596,N_6410,N_6470);
and U6597 (N_6597,N_6448,N_6498);
nand U6598 (N_6598,N_6450,N_6418);
or U6599 (N_6599,N_6466,N_6418);
nand U6600 (N_6600,N_6562,N_6561);
nand U6601 (N_6601,N_6524,N_6515);
and U6602 (N_6602,N_6567,N_6598);
and U6603 (N_6603,N_6597,N_6507);
nor U6604 (N_6604,N_6539,N_6521);
or U6605 (N_6605,N_6506,N_6547);
nor U6606 (N_6606,N_6595,N_6588);
or U6607 (N_6607,N_6555,N_6579);
and U6608 (N_6608,N_6581,N_6585);
nand U6609 (N_6609,N_6552,N_6560);
or U6610 (N_6610,N_6578,N_6540);
nand U6611 (N_6611,N_6593,N_6544);
nor U6612 (N_6612,N_6501,N_6538);
or U6613 (N_6613,N_6528,N_6545);
nand U6614 (N_6614,N_6565,N_6594);
or U6615 (N_6615,N_6549,N_6550);
and U6616 (N_6616,N_6577,N_6527);
xor U6617 (N_6617,N_6502,N_6546);
or U6618 (N_6618,N_6576,N_6542);
or U6619 (N_6619,N_6520,N_6529);
nor U6620 (N_6620,N_6551,N_6556);
nor U6621 (N_6621,N_6514,N_6510);
and U6622 (N_6622,N_6512,N_6503);
and U6623 (N_6623,N_6500,N_6523);
nand U6624 (N_6624,N_6508,N_6573);
and U6625 (N_6625,N_6548,N_6589);
and U6626 (N_6626,N_6533,N_6554);
nor U6627 (N_6627,N_6509,N_6591);
or U6628 (N_6628,N_6504,N_6558);
and U6629 (N_6629,N_6519,N_6557);
nand U6630 (N_6630,N_6570,N_6522);
nand U6631 (N_6631,N_6564,N_6568);
or U6632 (N_6632,N_6559,N_6536);
nand U6633 (N_6633,N_6580,N_6513);
nor U6634 (N_6634,N_6571,N_6583);
and U6635 (N_6635,N_6525,N_6505);
nor U6636 (N_6636,N_6596,N_6517);
and U6637 (N_6637,N_6518,N_6569);
nand U6638 (N_6638,N_6590,N_6541);
and U6639 (N_6639,N_6535,N_6531);
and U6640 (N_6640,N_6566,N_6574);
or U6641 (N_6641,N_6563,N_6575);
and U6642 (N_6642,N_6532,N_6526);
nor U6643 (N_6643,N_6582,N_6553);
nor U6644 (N_6644,N_6511,N_6534);
or U6645 (N_6645,N_6516,N_6584);
nand U6646 (N_6646,N_6530,N_6586);
nor U6647 (N_6647,N_6587,N_6592);
nor U6648 (N_6648,N_6572,N_6599);
and U6649 (N_6649,N_6543,N_6537);
and U6650 (N_6650,N_6556,N_6579);
and U6651 (N_6651,N_6500,N_6581);
xnor U6652 (N_6652,N_6566,N_6598);
nand U6653 (N_6653,N_6557,N_6572);
nor U6654 (N_6654,N_6522,N_6507);
nor U6655 (N_6655,N_6541,N_6501);
nand U6656 (N_6656,N_6574,N_6597);
nor U6657 (N_6657,N_6546,N_6593);
and U6658 (N_6658,N_6507,N_6523);
or U6659 (N_6659,N_6510,N_6526);
and U6660 (N_6660,N_6512,N_6546);
or U6661 (N_6661,N_6568,N_6593);
xor U6662 (N_6662,N_6599,N_6543);
nand U6663 (N_6663,N_6572,N_6583);
and U6664 (N_6664,N_6516,N_6543);
nand U6665 (N_6665,N_6581,N_6571);
and U6666 (N_6666,N_6580,N_6574);
xnor U6667 (N_6667,N_6536,N_6532);
nor U6668 (N_6668,N_6527,N_6528);
nand U6669 (N_6669,N_6580,N_6526);
or U6670 (N_6670,N_6547,N_6571);
and U6671 (N_6671,N_6593,N_6586);
xor U6672 (N_6672,N_6549,N_6502);
or U6673 (N_6673,N_6551,N_6500);
or U6674 (N_6674,N_6545,N_6518);
nor U6675 (N_6675,N_6503,N_6535);
or U6676 (N_6676,N_6560,N_6556);
or U6677 (N_6677,N_6563,N_6564);
or U6678 (N_6678,N_6545,N_6591);
xor U6679 (N_6679,N_6528,N_6504);
nand U6680 (N_6680,N_6545,N_6589);
or U6681 (N_6681,N_6500,N_6590);
nand U6682 (N_6682,N_6503,N_6570);
nor U6683 (N_6683,N_6574,N_6564);
or U6684 (N_6684,N_6576,N_6590);
nand U6685 (N_6685,N_6544,N_6547);
and U6686 (N_6686,N_6536,N_6520);
xnor U6687 (N_6687,N_6528,N_6593);
or U6688 (N_6688,N_6529,N_6562);
and U6689 (N_6689,N_6536,N_6524);
nor U6690 (N_6690,N_6571,N_6596);
nor U6691 (N_6691,N_6584,N_6583);
xnor U6692 (N_6692,N_6576,N_6589);
and U6693 (N_6693,N_6507,N_6548);
or U6694 (N_6694,N_6595,N_6535);
nor U6695 (N_6695,N_6578,N_6526);
xnor U6696 (N_6696,N_6542,N_6592);
and U6697 (N_6697,N_6549,N_6531);
or U6698 (N_6698,N_6560,N_6500);
nor U6699 (N_6699,N_6571,N_6572);
or U6700 (N_6700,N_6604,N_6639);
and U6701 (N_6701,N_6684,N_6618);
nor U6702 (N_6702,N_6681,N_6624);
and U6703 (N_6703,N_6678,N_6653);
nor U6704 (N_6704,N_6637,N_6670);
nor U6705 (N_6705,N_6654,N_6652);
nor U6706 (N_6706,N_6697,N_6640);
xor U6707 (N_6707,N_6683,N_6685);
or U6708 (N_6708,N_6661,N_6628);
or U6709 (N_6709,N_6603,N_6658);
and U6710 (N_6710,N_6611,N_6675);
or U6711 (N_6711,N_6691,N_6606);
or U6712 (N_6712,N_6600,N_6664);
and U6713 (N_6713,N_6620,N_6690);
xnor U6714 (N_6714,N_6659,N_6662);
and U6715 (N_6715,N_6650,N_6614);
nand U6716 (N_6716,N_6644,N_6605);
nand U6717 (N_6717,N_6655,N_6607);
or U6718 (N_6718,N_6680,N_6689);
and U6719 (N_6719,N_6673,N_6613);
nand U6720 (N_6720,N_6622,N_6609);
or U6721 (N_6721,N_6674,N_6641);
nand U6722 (N_6722,N_6698,N_6676);
nand U6723 (N_6723,N_6660,N_6647);
and U6724 (N_6724,N_6645,N_6646);
or U6725 (N_6725,N_6672,N_6631);
and U6726 (N_6726,N_6634,N_6610);
or U6727 (N_6727,N_6696,N_6617);
nor U6728 (N_6728,N_6651,N_6668);
nand U6729 (N_6729,N_6623,N_6671);
and U6730 (N_6730,N_6635,N_6643);
nand U6731 (N_6731,N_6693,N_6669);
and U6732 (N_6732,N_6677,N_6612);
and U6733 (N_6733,N_6648,N_6615);
or U6734 (N_6734,N_6666,N_6688);
or U6735 (N_6735,N_6679,N_6619);
and U6736 (N_6736,N_6694,N_6616);
or U6737 (N_6737,N_6687,N_6699);
xnor U6738 (N_6738,N_6663,N_6667);
and U6739 (N_6739,N_6627,N_6692);
or U6740 (N_6740,N_6630,N_6649);
nand U6741 (N_6741,N_6629,N_6638);
nor U6742 (N_6742,N_6642,N_6695);
or U6743 (N_6743,N_6657,N_6682);
and U6744 (N_6744,N_6665,N_6625);
nand U6745 (N_6745,N_6601,N_6608);
and U6746 (N_6746,N_6621,N_6686);
nor U6747 (N_6747,N_6602,N_6632);
nand U6748 (N_6748,N_6633,N_6626);
nand U6749 (N_6749,N_6636,N_6656);
or U6750 (N_6750,N_6641,N_6604);
xor U6751 (N_6751,N_6601,N_6672);
nor U6752 (N_6752,N_6616,N_6685);
nand U6753 (N_6753,N_6649,N_6621);
nand U6754 (N_6754,N_6697,N_6677);
nor U6755 (N_6755,N_6642,N_6604);
nand U6756 (N_6756,N_6645,N_6680);
nand U6757 (N_6757,N_6682,N_6639);
and U6758 (N_6758,N_6603,N_6681);
and U6759 (N_6759,N_6684,N_6662);
nor U6760 (N_6760,N_6650,N_6668);
or U6761 (N_6761,N_6606,N_6673);
nor U6762 (N_6762,N_6608,N_6645);
xor U6763 (N_6763,N_6634,N_6622);
nand U6764 (N_6764,N_6614,N_6632);
or U6765 (N_6765,N_6659,N_6669);
xnor U6766 (N_6766,N_6617,N_6654);
nor U6767 (N_6767,N_6663,N_6609);
and U6768 (N_6768,N_6604,N_6673);
or U6769 (N_6769,N_6657,N_6664);
nand U6770 (N_6770,N_6615,N_6604);
nand U6771 (N_6771,N_6641,N_6644);
nor U6772 (N_6772,N_6634,N_6692);
and U6773 (N_6773,N_6654,N_6683);
nor U6774 (N_6774,N_6601,N_6600);
nand U6775 (N_6775,N_6695,N_6638);
nand U6776 (N_6776,N_6668,N_6638);
nor U6777 (N_6777,N_6667,N_6695);
nor U6778 (N_6778,N_6674,N_6655);
and U6779 (N_6779,N_6699,N_6607);
xnor U6780 (N_6780,N_6665,N_6650);
xnor U6781 (N_6781,N_6642,N_6658);
and U6782 (N_6782,N_6619,N_6645);
nand U6783 (N_6783,N_6607,N_6660);
xnor U6784 (N_6784,N_6641,N_6618);
xnor U6785 (N_6785,N_6672,N_6690);
and U6786 (N_6786,N_6668,N_6643);
xnor U6787 (N_6787,N_6671,N_6613);
nor U6788 (N_6788,N_6620,N_6676);
nor U6789 (N_6789,N_6654,N_6646);
nand U6790 (N_6790,N_6676,N_6691);
xnor U6791 (N_6791,N_6699,N_6671);
nor U6792 (N_6792,N_6604,N_6699);
xnor U6793 (N_6793,N_6660,N_6629);
and U6794 (N_6794,N_6626,N_6691);
nor U6795 (N_6795,N_6661,N_6657);
or U6796 (N_6796,N_6637,N_6698);
nand U6797 (N_6797,N_6665,N_6638);
or U6798 (N_6798,N_6657,N_6630);
nand U6799 (N_6799,N_6681,N_6684);
and U6800 (N_6800,N_6774,N_6765);
xor U6801 (N_6801,N_6786,N_6712);
and U6802 (N_6802,N_6776,N_6771);
and U6803 (N_6803,N_6716,N_6795);
and U6804 (N_6804,N_6740,N_6794);
nand U6805 (N_6805,N_6785,N_6767);
nand U6806 (N_6806,N_6721,N_6792);
nand U6807 (N_6807,N_6722,N_6715);
or U6808 (N_6808,N_6798,N_6702);
and U6809 (N_6809,N_6743,N_6700);
xor U6810 (N_6810,N_6723,N_6766);
and U6811 (N_6811,N_6783,N_6752);
or U6812 (N_6812,N_6762,N_6727);
or U6813 (N_6813,N_6737,N_6761);
and U6814 (N_6814,N_6724,N_6741);
or U6815 (N_6815,N_6789,N_6755);
nand U6816 (N_6816,N_6784,N_6747);
xor U6817 (N_6817,N_6754,N_6729);
or U6818 (N_6818,N_6750,N_6760);
xor U6819 (N_6819,N_6701,N_6710);
and U6820 (N_6820,N_6772,N_6757);
xor U6821 (N_6821,N_6705,N_6709);
nor U6822 (N_6822,N_6781,N_6732);
nor U6823 (N_6823,N_6748,N_6773);
and U6824 (N_6824,N_6726,N_6720);
and U6825 (N_6825,N_6742,N_6735);
nand U6826 (N_6826,N_6770,N_6731);
nor U6827 (N_6827,N_6769,N_6706);
nor U6828 (N_6828,N_6707,N_6734);
xnor U6829 (N_6829,N_6746,N_6793);
or U6830 (N_6830,N_6780,N_6744);
or U6831 (N_6831,N_6796,N_6758);
or U6832 (N_6832,N_6708,N_6749);
nand U6833 (N_6833,N_6791,N_6704);
nand U6834 (N_6834,N_6790,N_6779);
nand U6835 (N_6835,N_6736,N_6745);
nand U6836 (N_6836,N_6717,N_6703);
or U6837 (N_6837,N_6718,N_6787);
and U6838 (N_6838,N_6764,N_6788);
nand U6839 (N_6839,N_6753,N_6763);
nand U6840 (N_6840,N_6728,N_6725);
nor U6841 (N_6841,N_6756,N_6778);
or U6842 (N_6842,N_6719,N_6782);
or U6843 (N_6843,N_6768,N_6739);
and U6844 (N_6844,N_6797,N_6751);
and U6845 (N_6845,N_6799,N_6711);
or U6846 (N_6846,N_6730,N_6714);
nand U6847 (N_6847,N_6775,N_6738);
nor U6848 (N_6848,N_6713,N_6733);
or U6849 (N_6849,N_6777,N_6759);
or U6850 (N_6850,N_6734,N_6737);
or U6851 (N_6851,N_6764,N_6781);
or U6852 (N_6852,N_6753,N_6777);
and U6853 (N_6853,N_6702,N_6711);
or U6854 (N_6854,N_6703,N_6775);
nand U6855 (N_6855,N_6793,N_6742);
and U6856 (N_6856,N_6729,N_6747);
nor U6857 (N_6857,N_6777,N_6794);
and U6858 (N_6858,N_6754,N_6721);
xor U6859 (N_6859,N_6724,N_6734);
nor U6860 (N_6860,N_6706,N_6742);
and U6861 (N_6861,N_6768,N_6762);
nand U6862 (N_6862,N_6710,N_6796);
or U6863 (N_6863,N_6712,N_6702);
or U6864 (N_6864,N_6706,N_6757);
or U6865 (N_6865,N_6776,N_6792);
or U6866 (N_6866,N_6735,N_6769);
or U6867 (N_6867,N_6784,N_6743);
nor U6868 (N_6868,N_6789,N_6760);
or U6869 (N_6869,N_6773,N_6785);
nor U6870 (N_6870,N_6725,N_6771);
and U6871 (N_6871,N_6749,N_6735);
nor U6872 (N_6872,N_6771,N_6780);
nor U6873 (N_6873,N_6730,N_6704);
or U6874 (N_6874,N_6760,N_6778);
nor U6875 (N_6875,N_6745,N_6702);
or U6876 (N_6876,N_6748,N_6792);
nor U6877 (N_6877,N_6707,N_6771);
or U6878 (N_6878,N_6744,N_6749);
xnor U6879 (N_6879,N_6743,N_6761);
nand U6880 (N_6880,N_6772,N_6704);
or U6881 (N_6881,N_6717,N_6707);
and U6882 (N_6882,N_6776,N_6760);
nand U6883 (N_6883,N_6782,N_6786);
nor U6884 (N_6884,N_6768,N_6731);
nand U6885 (N_6885,N_6743,N_6788);
xnor U6886 (N_6886,N_6772,N_6780);
xor U6887 (N_6887,N_6716,N_6748);
and U6888 (N_6888,N_6797,N_6798);
nand U6889 (N_6889,N_6767,N_6766);
or U6890 (N_6890,N_6757,N_6782);
and U6891 (N_6891,N_6770,N_6715);
nand U6892 (N_6892,N_6749,N_6777);
or U6893 (N_6893,N_6718,N_6767);
nor U6894 (N_6894,N_6777,N_6768);
nor U6895 (N_6895,N_6718,N_6799);
nand U6896 (N_6896,N_6760,N_6744);
and U6897 (N_6897,N_6725,N_6766);
and U6898 (N_6898,N_6742,N_6783);
or U6899 (N_6899,N_6708,N_6703);
or U6900 (N_6900,N_6891,N_6865);
or U6901 (N_6901,N_6825,N_6864);
and U6902 (N_6902,N_6871,N_6873);
nand U6903 (N_6903,N_6875,N_6821);
xor U6904 (N_6904,N_6877,N_6886);
xor U6905 (N_6905,N_6890,N_6850);
and U6906 (N_6906,N_6817,N_6870);
nor U6907 (N_6907,N_6862,N_6881);
or U6908 (N_6908,N_6805,N_6880);
and U6909 (N_6909,N_6897,N_6895);
and U6910 (N_6910,N_6868,N_6872);
or U6911 (N_6911,N_6853,N_6848);
or U6912 (N_6912,N_6854,N_6827);
nand U6913 (N_6913,N_6815,N_6836);
or U6914 (N_6914,N_6894,N_6849);
and U6915 (N_6915,N_6896,N_6866);
and U6916 (N_6916,N_6861,N_6832);
xnor U6917 (N_6917,N_6822,N_6892);
or U6918 (N_6918,N_6835,N_6879);
nor U6919 (N_6919,N_6814,N_6811);
and U6920 (N_6920,N_6878,N_6869);
nor U6921 (N_6921,N_6874,N_6813);
nor U6922 (N_6922,N_6838,N_6842);
and U6923 (N_6923,N_6820,N_6834);
and U6924 (N_6924,N_6804,N_6843);
nor U6925 (N_6925,N_6831,N_6851);
xor U6926 (N_6926,N_6801,N_6856);
xnor U6927 (N_6927,N_6826,N_6837);
nand U6928 (N_6928,N_6887,N_6845);
nand U6929 (N_6929,N_6858,N_6806);
and U6930 (N_6930,N_6860,N_6882);
and U6931 (N_6931,N_6828,N_6807);
xnor U6932 (N_6932,N_6884,N_6840);
or U6933 (N_6933,N_6839,N_6898);
nor U6934 (N_6934,N_6819,N_6803);
and U6935 (N_6935,N_6802,N_6818);
xor U6936 (N_6936,N_6885,N_6867);
xnor U6937 (N_6937,N_6859,N_6808);
and U6938 (N_6938,N_6833,N_6824);
xnor U6939 (N_6939,N_6889,N_6899);
nor U6940 (N_6940,N_6812,N_6893);
and U6941 (N_6941,N_6876,N_6810);
or U6942 (N_6942,N_6829,N_6888);
nand U6943 (N_6943,N_6809,N_6846);
and U6944 (N_6944,N_6830,N_6823);
or U6945 (N_6945,N_6800,N_6841);
nor U6946 (N_6946,N_6847,N_6883);
nor U6947 (N_6947,N_6816,N_6852);
nand U6948 (N_6948,N_6857,N_6844);
nand U6949 (N_6949,N_6863,N_6855);
nand U6950 (N_6950,N_6883,N_6866);
and U6951 (N_6951,N_6884,N_6824);
nor U6952 (N_6952,N_6896,N_6892);
xor U6953 (N_6953,N_6807,N_6858);
or U6954 (N_6954,N_6869,N_6802);
nand U6955 (N_6955,N_6844,N_6805);
or U6956 (N_6956,N_6866,N_6885);
and U6957 (N_6957,N_6895,N_6887);
nor U6958 (N_6958,N_6863,N_6848);
and U6959 (N_6959,N_6844,N_6899);
nand U6960 (N_6960,N_6859,N_6819);
nand U6961 (N_6961,N_6875,N_6811);
nand U6962 (N_6962,N_6813,N_6855);
or U6963 (N_6963,N_6867,N_6846);
xor U6964 (N_6964,N_6862,N_6879);
nor U6965 (N_6965,N_6860,N_6870);
xnor U6966 (N_6966,N_6898,N_6818);
nor U6967 (N_6967,N_6884,N_6896);
nand U6968 (N_6968,N_6871,N_6846);
nor U6969 (N_6969,N_6805,N_6814);
nand U6970 (N_6970,N_6833,N_6851);
and U6971 (N_6971,N_6822,N_6852);
nand U6972 (N_6972,N_6818,N_6875);
or U6973 (N_6973,N_6818,N_6883);
or U6974 (N_6974,N_6804,N_6800);
and U6975 (N_6975,N_6897,N_6894);
nor U6976 (N_6976,N_6889,N_6823);
xnor U6977 (N_6977,N_6870,N_6853);
nand U6978 (N_6978,N_6856,N_6809);
or U6979 (N_6979,N_6888,N_6862);
and U6980 (N_6980,N_6895,N_6803);
and U6981 (N_6981,N_6847,N_6870);
or U6982 (N_6982,N_6845,N_6815);
and U6983 (N_6983,N_6852,N_6818);
or U6984 (N_6984,N_6841,N_6847);
nor U6985 (N_6985,N_6876,N_6862);
or U6986 (N_6986,N_6899,N_6851);
nor U6987 (N_6987,N_6838,N_6855);
nand U6988 (N_6988,N_6818,N_6891);
and U6989 (N_6989,N_6863,N_6838);
nor U6990 (N_6990,N_6814,N_6809);
nor U6991 (N_6991,N_6825,N_6813);
and U6992 (N_6992,N_6813,N_6863);
nor U6993 (N_6993,N_6867,N_6803);
or U6994 (N_6994,N_6862,N_6825);
and U6995 (N_6995,N_6855,N_6893);
and U6996 (N_6996,N_6870,N_6844);
or U6997 (N_6997,N_6888,N_6841);
nand U6998 (N_6998,N_6857,N_6800);
or U6999 (N_6999,N_6845,N_6869);
nor U7000 (N_7000,N_6976,N_6915);
nor U7001 (N_7001,N_6919,N_6939);
or U7002 (N_7002,N_6946,N_6958);
nor U7003 (N_7003,N_6955,N_6905);
nand U7004 (N_7004,N_6925,N_6933);
nand U7005 (N_7005,N_6952,N_6970);
and U7006 (N_7006,N_6916,N_6960);
xnor U7007 (N_7007,N_6931,N_6956);
nor U7008 (N_7008,N_6950,N_6977);
and U7009 (N_7009,N_6954,N_6938);
nand U7010 (N_7010,N_6963,N_6949);
and U7011 (N_7011,N_6914,N_6959);
or U7012 (N_7012,N_6923,N_6997);
xnor U7013 (N_7013,N_6918,N_6943);
nand U7014 (N_7014,N_6992,N_6922);
or U7015 (N_7015,N_6927,N_6989);
and U7016 (N_7016,N_6967,N_6951);
nor U7017 (N_7017,N_6944,N_6953);
and U7018 (N_7018,N_6978,N_6924);
nor U7019 (N_7019,N_6962,N_6913);
and U7020 (N_7020,N_6966,N_6921);
xnor U7021 (N_7021,N_6971,N_6920);
or U7022 (N_7022,N_6961,N_6906);
nand U7023 (N_7023,N_6993,N_6983);
nor U7024 (N_7024,N_6935,N_6900);
nand U7025 (N_7025,N_6903,N_6928);
xor U7026 (N_7026,N_6907,N_6937);
and U7027 (N_7027,N_6979,N_6910);
nor U7028 (N_7028,N_6912,N_6988);
or U7029 (N_7029,N_6996,N_6941);
nand U7030 (N_7030,N_6990,N_6929);
nand U7031 (N_7031,N_6999,N_6981);
and U7032 (N_7032,N_6908,N_6995);
or U7033 (N_7033,N_6984,N_6926);
and U7034 (N_7034,N_6957,N_6980);
nor U7035 (N_7035,N_6942,N_6975);
and U7036 (N_7036,N_6968,N_6986);
nand U7037 (N_7037,N_6982,N_6904);
nand U7038 (N_7038,N_6936,N_6917);
and U7039 (N_7039,N_6901,N_6930);
xor U7040 (N_7040,N_6964,N_6945);
nor U7041 (N_7041,N_6991,N_6973);
and U7042 (N_7042,N_6974,N_6985);
or U7043 (N_7043,N_6947,N_6909);
nor U7044 (N_7044,N_6932,N_6987);
nand U7045 (N_7045,N_6998,N_6934);
nand U7046 (N_7046,N_6911,N_6965);
and U7047 (N_7047,N_6972,N_6994);
or U7048 (N_7048,N_6940,N_6948);
xnor U7049 (N_7049,N_6902,N_6969);
or U7050 (N_7050,N_6952,N_6976);
xor U7051 (N_7051,N_6945,N_6925);
nand U7052 (N_7052,N_6934,N_6949);
nor U7053 (N_7053,N_6917,N_6997);
xnor U7054 (N_7054,N_6946,N_6903);
and U7055 (N_7055,N_6931,N_6949);
nor U7056 (N_7056,N_6991,N_6985);
or U7057 (N_7057,N_6926,N_6907);
nor U7058 (N_7058,N_6931,N_6932);
or U7059 (N_7059,N_6916,N_6985);
xor U7060 (N_7060,N_6934,N_6923);
xor U7061 (N_7061,N_6950,N_6933);
xnor U7062 (N_7062,N_6977,N_6963);
or U7063 (N_7063,N_6961,N_6985);
or U7064 (N_7064,N_6962,N_6911);
or U7065 (N_7065,N_6989,N_6921);
or U7066 (N_7066,N_6977,N_6952);
nor U7067 (N_7067,N_6989,N_6976);
nand U7068 (N_7068,N_6900,N_6927);
and U7069 (N_7069,N_6905,N_6959);
and U7070 (N_7070,N_6936,N_6929);
nand U7071 (N_7071,N_6963,N_6987);
nand U7072 (N_7072,N_6998,N_6925);
and U7073 (N_7073,N_6925,N_6965);
xor U7074 (N_7074,N_6907,N_6909);
and U7075 (N_7075,N_6909,N_6912);
nand U7076 (N_7076,N_6977,N_6913);
nor U7077 (N_7077,N_6946,N_6959);
and U7078 (N_7078,N_6966,N_6918);
xnor U7079 (N_7079,N_6971,N_6930);
nand U7080 (N_7080,N_6934,N_6916);
nor U7081 (N_7081,N_6903,N_6986);
or U7082 (N_7082,N_6906,N_6921);
or U7083 (N_7083,N_6907,N_6978);
or U7084 (N_7084,N_6986,N_6941);
nor U7085 (N_7085,N_6900,N_6924);
or U7086 (N_7086,N_6928,N_6953);
and U7087 (N_7087,N_6934,N_6991);
or U7088 (N_7088,N_6900,N_6962);
and U7089 (N_7089,N_6951,N_6931);
nor U7090 (N_7090,N_6977,N_6951);
nor U7091 (N_7091,N_6946,N_6909);
xnor U7092 (N_7092,N_6997,N_6951);
xnor U7093 (N_7093,N_6985,N_6995);
and U7094 (N_7094,N_6911,N_6950);
nand U7095 (N_7095,N_6970,N_6909);
nor U7096 (N_7096,N_6955,N_6967);
nor U7097 (N_7097,N_6927,N_6901);
or U7098 (N_7098,N_6961,N_6902);
nand U7099 (N_7099,N_6925,N_6990);
nor U7100 (N_7100,N_7045,N_7003);
nor U7101 (N_7101,N_7046,N_7006);
nand U7102 (N_7102,N_7082,N_7015);
nor U7103 (N_7103,N_7073,N_7020);
nor U7104 (N_7104,N_7000,N_7063);
and U7105 (N_7105,N_7005,N_7089);
nor U7106 (N_7106,N_7001,N_7077);
or U7107 (N_7107,N_7023,N_7024);
nand U7108 (N_7108,N_7016,N_7075);
or U7109 (N_7109,N_7038,N_7097);
nand U7110 (N_7110,N_7028,N_7088);
xnor U7111 (N_7111,N_7030,N_7065);
and U7112 (N_7112,N_7004,N_7011);
and U7113 (N_7113,N_7056,N_7050);
or U7114 (N_7114,N_7047,N_7029);
nand U7115 (N_7115,N_7092,N_7080);
nor U7116 (N_7116,N_7019,N_7086);
nand U7117 (N_7117,N_7009,N_7002);
nor U7118 (N_7118,N_7062,N_7012);
nand U7119 (N_7119,N_7051,N_7074);
or U7120 (N_7120,N_7078,N_7070);
nor U7121 (N_7121,N_7098,N_7007);
nor U7122 (N_7122,N_7053,N_7044);
xnor U7123 (N_7123,N_7049,N_7060);
or U7124 (N_7124,N_7034,N_7081);
nand U7125 (N_7125,N_7036,N_7043);
nand U7126 (N_7126,N_7042,N_7087);
and U7127 (N_7127,N_7061,N_7066);
nor U7128 (N_7128,N_7025,N_7010);
nand U7129 (N_7129,N_7058,N_7059);
and U7130 (N_7130,N_7027,N_7055);
or U7131 (N_7131,N_7041,N_7048);
nor U7132 (N_7132,N_7071,N_7018);
nor U7133 (N_7133,N_7052,N_7054);
nor U7134 (N_7134,N_7068,N_7013);
xor U7135 (N_7135,N_7090,N_7033);
and U7136 (N_7136,N_7099,N_7031);
nor U7137 (N_7137,N_7094,N_7039);
or U7138 (N_7138,N_7021,N_7069);
nand U7139 (N_7139,N_7084,N_7008);
and U7140 (N_7140,N_7091,N_7064);
and U7141 (N_7141,N_7096,N_7093);
nand U7142 (N_7142,N_7040,N_7095);
or U7143 (N_7143,N_7014,N_7076);
xor U7144 (N_7144,N_7017,N_7035);
nand U7145 (N_7145,N_7067,N_7032);
nor U7146 (N_7146,N_7022,N_7026);
nand U7147 (N_7147,N_7079,N_7085);
and U7148 (N_7148,N_7072,N_7083);
or U7149 (N_7149,N_7057,N_7037);
or U7150 (N_7150,N_7048,N_7004);
nand U7151 (N_7151,N_7059,N_7095);
nor U7152 (N_7152,N_7024,N_7084);
nor U7153 (N_7153,N_7059,N_7057);
xnor U7154 (N_7154,N_7044,N_7038);
nor U7155 (N_7155,N_7096,N_7091);
or U7156 (N_7156,N_7046,N_7090);
or U7157 (N_7157,N_7020,N_7032);
or U7158 (N_7158,N_7095,N_7039);
xor U7159 (N_7159,N_7077,N_7076);
or U7160 (N_7160,N_7022,N_7065);
or U7161 (N_7161,N_7055,N_7079);
nor U7162 (N_7162,N_7002,N_7060);
or U7163 (N_7163,N_7047,N_7012);
nor U7164 (N_7164,N_7006,N_7022);
nor U7165 (N_7165,N_7021,N_7051);
and U7166 (N_7166,N_7055,N_7059);
nor U7167 (N_7167,N_7080,N_7043);
nor U7168 (N_7168,N_7042,N_7074);
and U7169 (N_7169,N_7030,N_7001);
nor U7170 (N_7170,N_7038,N_7053);
or U7171 (N_7171,N_7098,N_7012);
or U7172 (N_7172,N_7036,N_7006);
and U7173 (N_7173,N_7085,N_7086);
and U7174 (N_7174,N_7023,N_7050);
or U7175 (N_7175,N_7087,N_7049);
nand U7176 (N_7176,N_7039,N_7093);
and U7177 (N_7177,N_7026,N_7030);
and U7178 (N_7178,N_7088,N_7011);
or U7179 (N_7179,N_7018,N_7020);
or U7180 (N_7180,N_7013,N_7006);
nor U7181 (N_7181,N_7043,N_7024);
nor U7182 (N_7182,N_7012,N_7099);
xor U7183 (N_7183,N_7063,N_7051);
and U7184 (N_7184,N_7053,N_7094);
and U7185 (N_7185,N_7084,N_7061);
and U7186 (N_7186,N_7063,N_7084);
xnor U7187 (N_7187,N_7065,N_7043);
nor U7188 (N_7188,N_7084,N_7064);
or U7189 (N_7189,N_7087,N_7008);
xnor U7190 (N_7190,N_7006,N_7054);
nand U7191 (N_7191,N_7020,N_7061);
nand U7192 (N_7192,N_7073,N_7099);
and U7193 (N_7193,N_7071,N_7050);
nor U7194 (N_7194,N_7073,N_7008);
or U7195 (N_7195,N_7036,N_7041);
and U7196 (N_7196,N_7065,N_7067);
or U7197 (N_7197,N_7004,N_7026);
and U7198 (N_7198,N_7054,N_7004);
nand U7199 (N_7199,N_7085,N_7098);
nor U7200 (N_7200,N_7168,N_7175);
nand U7201 (N_7201,N_7193,N_7108);
or U7202 (N_7202,N_7166,N_7137);
nor U7203 (N_7203,N_7163,N_7125);
or U7204 (N_7204,N_7116,N_7107);
and U7205 (N_7205,N_7105,N_7135);
or U7206 (N_7206,N_7190,N_7120);
nand U7207 (N_7207,N_7159,N_7113);
nand U7208 (N_7208,N_7161,N_7188);
and U7209 (N_7209,N_7134,N_7132);
and U7210 (N_7210,N_7141,N_7173);
and U7211 (N_7211,N_7152,N_7148);
nand U7212 (N_7212,N_7154,N_7104);
or U7213 (N_7213,N_7197,N_7124);
or U7214 (N_7214,N_7167,N_7151);
and U7215 (N_7215,N_7187,N_7102);
nand U7216 (N_7216,N_7160,N_7100);
nor U7217 (N_7217,N_7142,N_7191);
nand U7218 (N_7218,N_7118,N_7199);
or U7219 (N_7219,N_7195,N_7112);
xnor U7220 (N_7220,N_7181,N_7189);
xor U7221 (N_7221,N_7128,N_7180);
nand U7222 (N_7222,N_7101,N_7194);
nor U7223 (N_7223,N_7174,N_7184);
or U7224 (N_7224,N_7103,N_7133);
nand U7225 (N_7225,N_7121,N_7153);
or U7226 (N_7226,N_7170,N_7143);
or U7227 (N_7227,N_7129,N_7158);
xnor U7228 (N_7228,N_7126,N_7140);
nand U7229 (N_7229,N_7119,N_7186);
or U7230 (N_7230,N_7178,N_7145);
xor U7231 (N_7231,N_7117,N_7165);
and U7232 (N_7232,N_7149,N_7110);
or U7233 (N_7233,N_7138,N_7162);
nor U7234 (N_7234,N_7183,N_7144);
or U7235 (N_7235,N_7156,N_7182);
and U7236 (N_7236,N_7171,N_7127);
xor U7237 (N_7237,N_7109,N_7155);
nand U7238 (N_7238,N_7192,N_7177);
nand U7239 (N_7239,N_7146,N_7106);
nor U7240 (N_7240,N_7179,N_7164);
nand U7241 (N_7241,N_7123,N_7150);
or U7242 (N_7242,N_7196,N_7122);
xor U7243 (N_7243,N_7198,N_7136);
nor U7244 (N_7244,N_7130,N_7115);
or U7245 (N_7245,N_7111,N_7169);
nand U7246 (N_7246,N_7147,N_7185);
xnor U7247 (N_7247,N_7114,N_7172);
or U7248 (N_7248,N_7131,N_7139);
and U7249 (N_7249,N_7157,N_7176);
or U7250 (N_7250,N_7136,N_7122);
nand U7251 (N_7251,N_7112,N_7181);
nor U7252 (N_7252,N_7154,N_7137);
xnor U7253 (N_7253,N_7132,N_7122);
and U7254 (N_7254,N_7154,N_7183);
or U7255 (N_7255,N_7172,N_7147);
xor U7256 (N_7256,N_7102,N_7146);
nand U7257 (N_7257,N_7136,N_7180);
nand U7258 (N_7258,N_7103,N_7154);
or U7259 (N_7259,N_7153,N_7161);
or U7260 (N_7260,N_7184,N_7108);
nor U7261 (N_7261,N_7126,N_7106);
and U7262 (N_7262,N_7181,N_7109);
or U7263 (N_7263,N_7188,N_7179);
and U7264 (N_7264,N_7168,N_7143);
nand U7265 (N_7265,N_7182,N_7195);
nand U7266 (N_7266,N_7199,N_7198);
or U7267 (N_7267,N_7199,N_7178);
nand U7268 (N_7268,N_7132,N_7176);
nor U7269 (N_7269,N_7138,N_7125);
and U7270 (N_7270,N_7113,N_7120);
and U7271 (N_7271,N_7143,N_7162);
nand U7272 (N_7272,N_7185,N_7139);
nand U7273 (N_7273,N_7120,N_7143);
or U7274 (N_7274,N_7140,N_7165);
or U7275 (N_7275,N_7188,N_7178);
nand U7276 (N_7276,N_7155,N_7137);
and U7277 (N_7277,N_7193,N_7130);
nand U7278 (N_7278,N_7130,N_7197);
and U7279 (N_7279,N_7108,N_7135);
or U7280 (N_7280,N_7145,N_7181);
or U7281 (N_7281,N_7151,N_7197);
nand U7282 (N_7282,N_7150,N_7162);
or U7283 (N_7283,N_7119,N_7168);
or U7284 (N_7284,N_7116,N_7169);
and U7285 (N_7285,N_7194,N_7100);
and U7286 (N_7286,N_7189,N_7114);
nor U7287 (N_7287,N_7141,N_7194);
xnor U7288 (N_7288,N_7190,N_7109);
nor U7289 (N_7289,N_7104,N_7109);
or U7290 (N_7290,N_7139,N_7177);
and U7291 (N_7291,N_7182,N_7157);
and U7292 (N_7292,N_7113,N_7112);
and U7293 (N_7293,N_7145,N_7148);
and U7294 (N_7294,N_7184,N_7164);
nand U7295 (N_7295,N_7122,N_7155);
nor U7296 (N_7296,N_7175,N_7154);
or U7297 (N_7297,N_7166,N_7120);
or U7298 (N_7298,N_7120,N_7134);
or U7299 (N_7299,N_7145,N_7149);
or U7300 (N_7300,N_7249,N_7212);
nor U7301 (N_7301,N_7285,N_7288);
xor U7302 (N_7302,N_7201,N_7280);
or U7303 (N_7303,N_7269,N_7275);
nor U7304 (N_7304,N_7264,N_7298);
nand U7305 (N_7305,N_7241,N_7223);
and U7306 (N_7306,N_7245,N_7239);
or U7307 (N_7307,N_7290,N_7224);
and U7308 (N_7308,N_7268,N_7218);
nor U7309 (N_7309,N_7236,N_7279);
nand U7310 (N_7310,N_7206,N_7217);
xnor U7311 (N_7311,N_7247,N_7276);
nand U7312 (N_7312,N_7274,N_7211);
and U7313 (N_7313,N_7281,N_7273);
nand U7314 (N_7314,N_7238,N_7230);
or U7315 (N_7315,N_7265,N_7233);
and U7316 (N_7316,N_7294,N_7295);
nand U7317 (N_7317,N_7237,N_7222);
or U7318 (N_7318,N_7244,N_7254);
or U7319 (N_7319,N_7248,N_7221);
xor U7320 (N_7320,N_7257,N_7256);
nand U7321 (N_7321,N_7200,N_7287);
nor U7322 (N_7322,N_7210,N_7251);
nor U7323 (N_7323,N_7231,N_7293);
and U7324 (N_7324,N_7243,N_7260);
or U7325 (N_7325,N_7271,N_7216);
or U7326 (N_7326,N_7208,N_7297);
nor U7327 (N_7327,N_7246,N_7215);
or U7328 (N_7328,N_7299,N_7240);
and U7329 (N_7329,N_7284,N_7255);
and U7330 (N_7330,N_7266,N_7213);
or U7331 (N_7331,N_7250,N_7272);
and U7332 (N_7332,N_7270,N_7226);
nor U7333 (N_7333,N_7291,N_7282);
nand U7334 (N_7334,N_7289,N_7209);
and U7335 (N_7335,N_7202,N_7235);
nor U7336 (N_7336,N_7259,N_7227);
nand U7337 (N_7337,N_7253,N_7204);
or U7338 (N_7338,N_7234,N_7263);
nand U7339 (N_7339,N_7267,N_7232);
nor U7340 (N_7340,N_7228,N_7214);
nor U7341 (N_7341,N_7252,N_7277);
or U7342 (N_7342,N_7242,N_7225);
or U7343 (N_7343,N_7229,N_7296);
or U7344 (N_7344,N_7286,N_7220);
and U7345 (N_7345,N_7292,N_7205);
nand U7346 (N_7346,N_7262,N_7283);
and U7347 (N_7347,N_7219,N_7258);
nor U7348 (N_7348,N_7207,N_7203);
nor U7349 (N_7349,N_7278,N_7261);
nor U7350 (N_7350,N_7297,N_7291);
and U7351 (N_7351,N_7244,N_7246);
and U7352 (N_7352,N_7221,N_7211);
and U7353 (N_7353,N_7218,N_7253);
nor U7354 (N_7354,N_7288,N_7205);
xnor U7355 (N_7355,N_7253,N_7283);
nand U7356 (N_7356,N_7232,N_7202);
nand U7357 (N_7357,N_7288,N_7213);
nand U7358 (N_7358,N_7283,N_7285);
or U7359 (N_7359,N_7206,N_7210);
or U7360 (N_7360,N_7280,N_7269);
xnor U7361 (N_7361,N_7276,N_7260);
xor U7362 (N_7362,N_7211,N_7257);
nor U7363 (N_7363,N_7213,N_7208);
nor U7364 (N_7364,N_7274,N_7226);
or U7365 (N_7365,N_7278,N_7247);
nor U7366 (N_7366,N_7273,N_7253);
or U7367 (N_7367,N_7209,N_7208);
or U7368 (N_7368,N_7246,N_7270);
nor U7369 (N_7369,N_7217,N_7270);
or U7370 (N_7370,N_7274,N_7212);
or U7371 (N_7371,N_7282,N_7292);
nand U7372 (N_7372,N_7280,N_7232);
nor U7373 (N_7373,N_7222,N_7223);
nor U7374 (N_7374,N_7205,N_7203);
nand U7375 (N_7375,N_7245,N_7263);
and U7376 (N_7376,N_7222,N_7266);
and U7377 (N_7377,N_7222,N_7254);
and U7378 (N_7378,N_7204,N_7252);
or U7379 (N_7379,N_7278,N_7275);
or U7380 (N_7380,N_7200,N_7205);
nor U7381 (N_7381,N_7211,N_7260);
nand U7382 (N_7382,N_7229,N_7223);
nor U7383 (N_7383,N_7242,N_7210);
nand U7384 (N_7384,N_7246,N_7260);
xor U7385 (N_7385,N_7233,N_7252);
nand U7386 (N_7386,N_7265,N_7299);
xnor U7387 (N_7387,N_7269,N_7245);
or U7388 (N_7388,N_7281,N_7255);
nand U7389 (N_7389,N_7263,N_7253);
or U7390 (N_7390,N_7286,N_7293);
and U7391 (N_7391,N_7265,N_7280);
or U7392 (N_7392,N_7296,N_7214);
nand U7393 (N_7393,N_7224,N_7271);
nor U7394 (N_7394,N_7296,N_7227);
or U7395 (N_7395,N_7209,N_7282);
nor U7396 (N_7396,N_7288,N_7251);
nand U7397 (N_7397,N_7204,N_7276);
nand U7398 (N_7398,N_7257,N_7284);
or U7399 (N_7399,N_7290,N_7203);
or U7400 (N_7400,N_7362,N_7396);
nor U7401 (N_7401,N_7391,N_7310);
or U7402 (N_7402,N_7304,N_7343);
nand U7403 (N_7403,N_7351,N_7346);
nor U7404 (N_7404,N_7341,N_7366);
nand U7405 (N_7405,N_7360,N_7393);
and U7406 (N_7406,N_7395,N_7317);
xnor U7407 (N_7407,N_7368,N_7348);
nor U7408 (N_7408,N_7370,N_7301);
nor U7409 (N_7409,N_7325,N_7354);
nand U7410 (N_7410,N_7327,N_7384);
nand U7411 (N_7411,N_7381,N_7388);
xor U7412 (N_7412,N_7329,N_7355);
nand U7413 (N_7413,N_7353,N_7392);
and U7414 (N_7414,N_7363,N_7385);
xor U7415 (N_7415,N_7323,N_7345);
or U7416 (N_7416,N_7383,N_7364);
nor U7417 (N_7417,N_7365,N_7379);
or U7418 (N_7418,N_7372,N_7303);
nor U7419 (N_7419,N_7386,N_7330);
xnor U7420 (N_7420,N_7359,N_7335);
nand U7421 (N_7421,N_7397,N_7340);
nor U7422 (N_7422,N_7306,N_7350);
nand U7423 (N_7423,N_7349,N_7336);
nor U7424 (N_7424,N_7314,N_7389);
nor U7425 (N_7425,N_7376,N_7394);
and U7426 (N_7426,N_7390,N_7382);
nand U7427 (N_7427,N_7369,N_7357);
and U7428 (N_7428,N_7321,N_7358);
and U7429 (N_7429,N_7352,N_7375);
and U7430 (N_7430,N_7328,N_7344);
nor U7431 (N_7431,N_7378,N_7322);
or U7432 (N_7432,N_7367,N_7361);
or U7433 (N_7433,N_7347,N_7356);
or U7434 (N_7434,N_7320,N_7316);
and U7435 (N_7435,N_7318,N_7334);
nor U7436 (N_7436,N_7339,N_7331);
and U7437 (N_7437,N_7326,N_7319);
or U7438 (N_7438,N_7373,N_7371);
nor U7439 (N_7439,N_7338,N_7300);
nand U7440 (N_7440,N_7309,N_7342);
nand U7441 (N_7441,N_7377,N_7387);
and U7442 (N_7442,N_7337,N_7374);
nor U7443 (N_7443,N_7307,N_7302);
or U7444 (N_7444,N_7399,N_7305);
xnor U7445 (N_7445,N_7311,N_7332);
and U7446 (N_7446,N_7313,N_7333);
or U7447 (N_7447,N_7312,N_7308);
and U7448 (N_7448,N_7398,N_7315);
xor U7449 (N_7449,N_7380,N_7324);
nand U7450 (N_7450,N_7387,N_7355);
and U7451 (N_7451,N_7337,N_7314);
nand U7452 (N_7452,N_7371,N_7351);
nor U7453 (N_7453,N_7336,N_7327);
or U7454 (N_7454,N_7352,N_7343);
and U7455 (N_7455,N_7351,N_7358);
nand U7456 (N_7456,N_7373,N_7324);
nand U7457 (N_7457,N_7314,N_7344);
xnor U7458 (N_7458,N_7308,N_7367);
nand U7459 (N_7459,N_7398,N_7349);
nor U7460 (N_7460,N_7318,N_7375);
or U7461 (N_7461,N_7308,N_7355);
xor U7462 (N_7462,N_7336,N_7386);
or U7463 (N_7463,N_7394,N_7359);
nand U7464 (N_7464,N_7374,N_7339);
and U7465 (N_7465,N_7340,N_7333);
and U7466 (N_7466,N_7362,N_7353);
or U7467 (N_7467,N_7366,N_7356);
nor U7468 (N_7468,N_7328,N_7374);
or U7469 (N_7469,N_7377,N_7351);
and U7470 (N_7470,N_7308,N_7347);
xnor U7471 (N_7471,N_7330,N_7314);
and U7472 (N_7472,N_7383,N_7321);
and U7473 (N_7473,N_7331,N_7307);
or U7474 (N_7474,N_7317,N_7342);
nor U7475 (N_7475,N_7367,N_7309);
and U7476 (N_7476,N_7348,N_7330);
and U7477 (N_7477,N_7377,N_7390);
xor U7478 (N_7478,N_7339,N_7328);
nand U7479 (N_7479,N_7331,N_7376);
and U7480 (N_7480,N_7340,N_7392);
nand U7481 (N_7481,N_7389,N_7359);
and U7482 (N_7482,N_7374,N_7359);
nor U7483 (N_7483,N_7398,N_7343);
nor U7484 (N_7484,N_7384,N_7349);
nand U7485 (N_7485,N_7378,N_7311);
nor U7486 (N_7486,N_7313,N_7346);
nand U7487 (N_7487,N_7334,N_7382);
nor U7488 (N_7488,N_7328,N_7391);
or U7489 (N_7489,N_7399,N_7383);
nand U7490 (N_7490,N_7387,N_7304);
and U7491 (N_7491,N_7316,N_7373);
nand U7492 (N_7492,N_7308,N_7360);
and U7493 (N_7493,N_7325,N_7312);
and U7494 (N_7494,N_7373,N_7356);
nand U7495 (N_7495,N_7336,N_7352);
or U7496 (N_7496,N_7322,N_7383);
nor U7497 (N_7497,N_7315,N_7327);
and U7498 (N_7498,N_7333,N_7324);
nand U7499 (N_7499,N_7356,N_7339);
nand U7500 (N_7500,N_7427,N_7473);
nand U7501 (N_7501,N_7464,N_7492);
nand U7502 (N_7502,N_7414,N_7404);
and U7503 (N_7503,N_7424,N_7444);
nand U7504 (N_7504,N_7488,N_7409);
and U7505 (N_7505,N_7449,N_7425);
and U7506 (N_7506,N_7432,N_7418);
or U7507 (N_7507,N_7417,N_7495);
or U7508 (N_7508,N_7437,N_7471);
xor U7509 (N_7509,N_7420,N_7481);
nor U7510 (N_7510,N_7462,N_7469);
nand U7511 (N_7511,N_7459,N_7408);
and U7512 (N_7512,N_7443,N_7419);
or U7513 (N_7513,N_7407,N_7478);
xor U7514 (N_7514,N_7465,N_7458);
and U7515 (N_7515,N_7453,N_7402);
nand U7516 (N_7516,N_7493,N_7450);
nor U7517 (N_7517,N_7479,N_7440);
nor U7518 (N_7518,N_7476,N_7496);
nand U7519 (N_7519,N_7470,N_7415);
and U7520 (N_7520,N_7498,N_7456);
nor U7521 (N_7521,N_7494,N_7423);
or U7522 (N_7522,N_7436,N_7400);
nor U7523 (N_7523,N_7477,N_7486);
or U7524 (N_7524,N_7438,N_7412);
and U7525 (N_7525,N_7410,N_7451);
or U7526 (N_7526,N_7446,N_7475);
or U7527 (N_7527,N_7499,N_7483);
or U7528 (N_7528,N_7445,N_7441);
xnor U7529 (N_7529,N_7463,N_7466);
nand U7530 (N_7530,N_7411,N_7480);
nor U7531 (N_7531,N_7439,N_7487);
and U7532 (N_7532,N_7497,N_7430);
or U7533 (N_7533,N_7442,N_7467);
nor U7534 (N_7534,N_7472,N_7448);
xor U7535 (N_7535,N_7447,N_7434);
xor U7536 (N_7536,N_7482,N_7429);
xnor U7537 (N_7537,N_7421,N_7413);
xnor U7538 (N_7538,N_7457,N_7433);
nor U7539 (N_7539,N_7485,N_7490);
xor U7540 (N_7540,N_7403,N_7401);
nand U7541 (N_7541,N_7422,N_7416);
and U7542 (N_7542,N_7431,N_7428);
and U7543 (N_7543,N_7474,N_7406);
xnor U7544 (N_7544,N_7405,N_7468);
or U7545 (N_7545,N_7455,N_7452);
xor U7546 (N_7546,N_7489,N_7454);
and U7547 (N_7547,N_7426,N_7461);
nor U7548 (N_7548,N_7491,N_7460);
or U7549 (N_7549,N_7435,N_7484);
and U7550 (N_7550,N_7487,N_7458);
nor U7551 (N_7551,N_7402,N_7406);
or U7552 (N_7552,N_7499,N_7417);
nor U7553 (N_7553,N_7432,N_7423);
and U7554 (N_7554,N_7491,N_7455);
nand U7555 (N_7555,N_7447,N_7439);
xor U7556 (N_7556,N_7480,N_7451);
xnor U7557 (N_7557,N_7408,N_7422);
nor U7558 (N_7558,N_7474,N_7417);
nor U7559 (N_7559,N_7408,N_7467);
and U7560 (N_7560,N_7487,N_7440);
or U7561 (N_7561,N_7440,N_7422);
nand U7562 (N_7562,N_7441,N_7408);
xor U7563 (N_7563,N_7409,N_7413);
or U7564 (N_7564,N_7469,N_7443);
nand U7565 (N_7565,N_7439,N_7474);
nor U7566 (N_7566,N_7412,N_7452);
xor U7567 (N_7567,N_7497,N_7459);
nor U7568 (N_7568,N_7405,N_7462);
xnor U7569 (N_7569,N_7400,N_7416);
nand U7570 (N_7570,N_7452,N_7437);
xnor U7571 (N_7571,N_7462,N_7473);
xnor U7572 (N_7572,N_7453,N_7436);
or U7573 (N_7573,N_7472,N_7432);
nor U7574 (N_7574,N_7463,N_7404);
or U7575 (N_7575,N_7450,N_7440);
nor U7576 (N_7576,N_7452,N_7451);
or U7577 (N_7577,N_7419,N_7420);
xnor U7578 (N_7578,N_7402,N_7463);
and U7579 (N_7579,N_7410,N_7425);
nand U7580 (N_7580,N_7430,N_7498);
or U7581 (N_7581,N_7428,N_7433);
and U7582 (N_7582,N_7419,N_7466);
xnor U7583 (N_7583,N_7409,N_7433);
and U7584 (N_7584,N_7433,N_7479);
nor U7585 (N_7585,N_7423,N_7421);
or U7586 (N_7586,N_7472,N_7412);
nand U7587 (N_7587,N_7413,N_7456);
and U7588 (N_7588,N_7480,N_7437);
nand U7589 (N_7589,N_7416,N_7483);
or U7590 (N_7590,N_7447,N_7484);
and U7591 (N_7591,N_7429,N_7402);
or U7592 (N_7592,N_7476,N_7432);
nand U7593 (N_7593,N_7452,N_7440);
nand U7594 (N_7594,N_7452,N_7465);
nor U7595 (N_7595,N_7405,N_7414);
or U7596 (N_7596,N_7463,N_7449);
nand U7597 (N_7597,N_7456,N_7417);
or U7598 (N_7598,N_7402,N_7498);
nor U7599 (N_7599,N_7494,N_7470);
and U7600 (N_7600,N_7593,N_7562);
or U7601 (N_7601,N_7541,N_7516);
or U7602 (N_7602,N_7544,N_7522);
or U7603 (N_7603,N_7503,N_7557);
or U7604 (N_7604,N_7547,N_7533);
nand U7605 (N_7605,N_7502,N_7517);
nand U7606 (N_7606,N_7577,N_7550);
nor U7607 (N_7607,N_7596,N_7564);
nand U7608 (N_7608,N_7597,N_7589);
and U7609 (N_7609,N_7584,N_7583);
nor U7610 (N_7610,N_7580,N_7598);
nor U7611 (N_7611,N_7594,N_7542);
nor U7612 (N_7612,N_7520,N_7552);
nor U7613 (N_7613,N_7530,N_7571);
nor U7614 (N_7614,N_7560,N_7534);
nor U7615 (N_7615,N_7590,N_7506);
or U7616 (N_7616,N_7510,N_7511);
xor U7617 (N_7617,N_7586,N_7585);
nand U7618 (N_7618,N_7543,N_7500);
or U7619 (N_7619,N_7574,N_7521);
and U7620 (N_7620,N_7519,N_7587);
nor U7621 (N_7621,N_7592,N_7568);
nand U7622 (N_7622,N_7537,N_7561);
nor U7623 (N_7623,N_7555,N_7532);
nand U7624 (N_7624,N_7549,N_7575);
xor U7625 (N_7625,N_7536,N_7515);
nor U7626 (N_7626,N_7553,N_7525);
and U7627 (N_7627,N_7591,N_7539);
or U7628 (N_7628,N_7527,N_7529);
nor U7629 (N_7629,N_7588,N_7578);
or U7630 (N_7630,N_7559,N_7566);
and U7631 (N_7631,N_7512,N_7582);
or U7632 (N_7632,N_7545,N_7509);
or U7633 (N_7633,N_7565,N_7556);
or U7634 (N_7634,N_7548,N_7507);
or U7635 (N_7635,N_7567,N_7523);
xor U7636 (N_7636,N_7595,N_7526);
nand U7637 (N_7637,N_7524,N_7570);
nor U7638 (N_7638,N_7599,N_7579);
or U7639 (N_7639,N_7531,N_7528);
nor U7640 (N_7640,N_7538,N_7572);
nor U7641 (N_7641,N_7501,N_7508);
or U7642 (N_7642,N_7504,N_7540);
and U7643 (N_7643,N_7514,N_7518);
or U7644 (N_7644,N_7551,N_7513);
nor U7645 (N_7645,N_7558,N_7563);
or U7646 (N_7646,N_7554,N_7569);
or U7647 (N_7647,N_7535,N_7546);
and U7648 (N_7648,N_7573,N_7576);
or U7649 (N_7649,N_7505,N_7581);
nand U7650 (N_7650,N_7559,N_7524);
and U7651 (N_7651,N_7551,N_7567);
nand U7652 (N_7652,N_7529,N_7525);
or U7653 (N_7653,N_7561,N_7593);
nand U7654 (N_7654,N_7506,N_7571);
or U7655 (N_7655,N_7555,N_7556);
and U7656 (N_7656,N_7593,N_7597);
nor U7657 (N_7657,N_7502,N_7589);
nor U7658 (N_7658,N_7535,N_7522);
or U7659 (N_7659,N_7553,N_7570);
nor U7660 (N_7660,N_7565,N_7551);
nor U7661 (N_7661,N_7507,N_7579);
and U7662 (N_7662,N_7517,N_7576);
nand U7663 (N_7663,N_7550,N_7513);
xor U7664 (N_7664,N_7505,N_7593);
nor U7665 (N_7665,N_7544,N_7576);
or U7666 (N_7666,N_7568,N_7538);
and U7667 (N_7667,N_7561,N_7573);
nand U7668 (N_7668,N_7514,N_7574);
and U7669 (N_7669,N_7581,N_7592);
xor U7670 (N_7670,N_7519,N_7511);
nor U7671 (N_7671,N_7522,N_7505);
and U7672 (N_7672,N_7519,N_7523);
nand U7673 (N_7673,N_7538,N_7524);
nand U7674 (N_7674,N_7561,N_7591);
nor U7675 (N_7675,N_7507,N_7557);
nor U7676 (N_7676,N_7554,N_7577);
and U7677 (N_7677,N_7508,N_7585);
nand U7678 (N_7678,N_7565,N_7503);
or U7679 (N_7679,N_7501,N_7533);
nor U7680 (N_7680,N_7585,N_7539);
nand U7681 (N_7681,N_7571,N_7511);
nand U7682 (N_7682,N_7593,N_7534);
and U7683 (N_7683,N_7573,N_7522);
nand U7684 (N_7684,N_7561,N_7596);
and U7685 (N_7685,N_7517,N_7554);
and U7686 (N_7686,N_7579,N_7511);
and U7687 (N_7687,N_7516,N_7501);
or U7688 (N_7688,N_7537,N_7596);
and U7689 (N_7689,N_7584,N_7579);
and U7690 (N_7690,N_7516,N_7535);
or U7691 (N_7691,N_7542,N_7506);
nor U7692 (N_7692,N_7512,N_7571);
nand U7693 (N_7693,N_7580,N_7548);
or U7694 (N_7694,N_7539,N_7555);
or U7695 (N_7695,N_7513,N_7547);
or U7696 (N_7696,N_7552,N_7529);
and U7697 (N_7697,N_7546,N_7582);
xnor U7698 (N_7698,N_7526,N_7597);
or U7699 (N_7699,N_7575,N_7561);
nand U7700 (N_7700,N_7663,N_7636);
and U7701 (N_7701,N_7667,N_7695);
nand U7702 (N_7702,N_7614,N_7600);
and U7703 (N_7703,N_7603,N_7666);
and U7704 (N_7704,N_7664,N_7659);
and U7705 (N_7705,N_7647,N_7672);
and U7706 (N_7706,N_7698,N_7625);
nor U7707 (N_7707,N_7681,N_7601);
nor U7708 (N_7708,N_7612,N_7627);
and U7709 (N_7709,N_7609,N_7649);
and U7710 (N_7710,N_7617,N_7602);
nand U7711 (N_7711,N_7629,N_7646);
nor U7712 (N_7712,N_7678,N_7679);
nand U7713 (N_7713,N_7615,N_7616);
and U7714 (N_7714,N_7651,N_7669);
and U7715 (N_7715,N_7608,N_7691);
and U7716 (N_7716,N_7622,N_7611);
and U7717 (N_7717,N_7640,N_7641);
nor U7718 (N_7718,N_7673,N_7638);
and U7719 (N_7719,N_7630,N_7668);
or U7720 (N_7720,N_7653,N_7631);
xnor U7721 (N_7721,N_7676,N_7632);
nand U7722 (N_7722,N_7605,N_7686);
or U7723 (N_7723,N_7635,N_7670);
and U7724 (N_7724,N_7692,N_7656);
nand U7725 (N_7725,N_7637,N_7690);
and U7726 (N_7726,N_7604,N_7623);
nor U7727 (N_7727,N_7675,N_7677);
nand U7728 (N_7728,N_7657,N_7644);
nand U7729 (N_7729,N_7658,N_7682);
nand U7730 (N_7730,N_7610,N_7694);
nor U7731 (N_7731,N_7639,N_7606);
and U7732 (N_7732,N_7642,N_7693);
or U7733 (N_7733,N_7643,N_7619);
nor U7734 (N_7734,N_7624,N_7645);
and U7735 (N_7735,N_7628,N_7618);
nand U7736 (N_7736,N_7684,N_7633);
nor U7737 (N_7737,N_7662,N_7687);
nor U7738 (N_7738,N_7683,N_7648);
or U7739 (N_7739,N_7661,N_7660);
nor U7740 (N_7740,N_7685,N_7650);
nand U7741 (N_7741,N_7620,N_7652);
or U7742 (N_7742,N_7680,N_7621);
nand U7743 (N_7743,N_7689,N_7634);
or U7744 (N_7744,N_7696,N_7665);
nand U7745 (N_7745,N_7626,N_7699);
or U7746 (N_7746,N_7655,N_7671);
and U7747 (N_7747,N_7613,N_7654);
and U7748 (N_7748,N_7697,N_7674);
xor U7749 (N_7749,N_7607,N_7688);
or U7750 (N_7750,N_7657,N_7634);
and U7751 (N_7751,N_7632,N_7652);
nor U7752 (N_7752,N_7670,N_7634);
xnor U7753 (N_7753,N_7669,N_7609);
nand U7754 (N_7754,N_7640,N_7654);
nand U7755 (N_7755,N_7683,N_7665);
and U7756 (N_7756,N_7683,N_7681);
and U7757 (N_7757,N_7696,N_7648);
nand U7758 (N_7758,N_7696,N_7687);
or U7759 (N_7759,N_7630,N_7643);
and U7760 (N_7760,N_7653,N_7676);
or U7761 (N_7761,N_7630,N_7695);
or U7762 (N_7762,N_7611,N_7608);
and U7763 (N_7763,N_7611,N_7613);
xor U7764 (N_7764,N_7691,N_7634);
nor U7765 (N_7765,N_7679,N_7636);
nand U7766 (N_7766,N_7678,N_7655);
nor U7767 (N_7767,N_7632,N_7644);
nand U7768 (N_7768,N_7628,N_7619);
or U7769 (N_7769,N_7605,N_7612);
and U7770 (N_7770,N_7658,N_7617);
nor U7771 (N_7771,N_7641,N_7608);
nand U7772 (N_7772,N_7672,N_7659);
or U7773 (N_7773,N_7605,N_7601);
nand U7774 (N_7774,N_7680,N_7657);
or U7775 (N_7775,N_7639,N_7656);
nand U7776 (N_7776,N_7686,N_7693);
or U7777 (N_7777,N_7680,N_7688);
nand U7778 (N_7778,N_7693,N_7608);
xnor U7779 (N_7779,N_7664,N_7666);
and U7780 (N_7780,N_7649,N_7668);
or U7781 (N_7781,N_7677,N_7622);
or U7782 (N_7782,N_7606,N_7632);
nor U7783 (N_7783,N_7620,N_7670);
nor U7784 (N_7784,N_7633,N_7692);
xor U7785 (N_7785,N_7610,N_7615);
and U7786 (N_7786,N_7694,N_7622);
nor U7787 (N_7787,N_7601,N_7644);
or U7788 (N_7788,N_7649,N_7653);
nand U7789 (N_7789,N_7665,N_7667);
nor U7790 (N_7790,N_7639,N_7629);
or U7791 (N_7791,N_7673,N_7654);
and U7792 (N_7792,N_7658,N_7636);
nand U7793 (N_7793,N_7690,N_7697);
or U7794 (N_7794,N_7654,N_7696);
and U7795 (N_7795,N_7661,N_7611);
nor U7796 (N_7796,N_7648,N_7657);
and U7797 (N_7797,N_7690,N_7650);
or U7798 (N_7798,N_7694,N_7666);
nand U7799 (N_7799,N_7636,N_7624);
nand U7800 (N_7800,N_7757,N_7725);
nor U7801 (N_7801,N_7766,N_7702);
nand U7802 (N_7802,N_7719,N_7754);
and U7803 (N_7803,N_7734,N_7764);
nor U7804 (N_7804,N_7755,N_7771);
nor U7805 (N_7805,N_7762,N_7718);
nor U7806 (N_7806,N_7770,N_7739);
nor U7807 (N_7807,N_7714,N_7751);
and U7808 (N_7808,N_7788,N_7794);
nor U7809 (N_7809,N_7767,N_7727);
xnor U7810 (N_7810,N_7744,N_7756);
nand U7811 (N_7811,N_7785,N_7704);
and U7812 (N_7812,N_7779,N_7736);
nand U7813 (N_7813,N_7763,N_7772);
or U7814 (N_7814,N_7765,N_7781);
or U7815 (N_7815,N_7724,N_7769);
and U7816 (N_7816,N_7748,N_7708);
nand U7817 (N_7817,N_7715,N_7791);
and U7818 (N_7818,N_7717,N_7795);
xor U7819 (N_7819,N_7720,N_7790);
nor U7820 (N_7820,N_7740,N_7732);
nand U7821 (N_7821,N_7777,N_7760);
nand U7822 (N_7822,N_7759,N_7733);
xor U7823 (N_7823,N_7706,N_7793);
nand U7824 (N_7824,N_7792,N_7709);
nor U7825 (N_7825,N_7703,N_7742);
or U7826 (N_7826,N_7743,N_7773);
nand U7827 (N_7827,N_7726,N_7721);
and U7828 (N_7828,N_7745,N_7747);
or U7829 (N_7829,N_7737,N_7716);
nor U7830 (N_7830,N_7746,N_7768);
and U7831 (N_7831,N_7784,N_7701);
or U7832 (N_7832,N_7700,N_7713);
xnor U7833 (N_7833,N_7728,N_7796);
nor U7834 (N_7834,N_7707,N_7723);
nor U7835 (N_7835,N_7731,N_7753);
and U7836 (N_7836,N_7758,N_7735);
nand U7837 (N_7837,N_7749,N_7730);
nand U7838 (N_7838,N_7750,N_7776);
nand U7839 (N_7839,N_7778,N_7761);
xor U7840 (N_7840,N_7705,N_7710);
and U7841 (N_7841,N_7774,N_7775);
or U7842 (N_7842,N_7729,N_7786);
nand U7843 (N_7843,N_7711,N_7787);
nor U7844 (N_7844,N_7722,N_7798);
nor U7845 (N_7845,N_7752,N_7712);
nand U7846 (N_7846,N_7789,N_7799);
and U7847 (N_7847,N_7783,N_7782);
xnor U7848 (N_7848,N_7738,N_7780);
or U7849 (N_7849,N_7797,N_7741);
nand U7850 (N_7850,N_7755,N_7708);
nand U7851 (N_7851,N_7796,N_7731);
xor U7852 (N_7852,N_7777,N_7772);
or U7853 (N_7853,N_7721,N_7705);
or U7854 (N_7854,N_7792,N_7793);
and U7855 (N_7855,N_7796,N_7780);
nand U7856 (N_7856,N_7733,N_7731);
and U7857 (N_7857,N_7706,N_7770);
nor U7858 (N_7858,N_7788,N_7719);
and U7859 (N_7859,N_7749,N_7783);
or U7860 (N_7860,N_7794,N_7787);
nor U7861 (N_7861,N_7799,N_7729);
and U7862 (N_7862,N_7763,N_7706);
or U7863 (N_7863,N_7799,N_7758);
nor U7864 (N_7864,N_7737,N_7760);
nor U7865 (N_7865,N_7723,N_7714);
or U7866 (N_7866,N_7709,N_7716);
nor U7867 (N_7867,N_7720,N_7762);
xor U7868 (N_7868,N_7743,N_7784);
and U7869 (N_7869,N_7741,N_7756);
nand U7870 (N_7870,N_7706,N_7745);
nand U7871 (N_7871,N_7718,N_7735);
nand U7872 (N_7872,N_7781,N_7727);
or U7873 (N_7873,N_7794,N_7779);
nand U7874 (N_7874,N_7751,N_7771);
nor U7875 (N_7875,N_7754,N_7737);
nor U7876 (N_7876,N_7706,N_7708);
or U7877 (N_7877,N_7709,N_7764);
nand U7878 (N_7878,N_7795,N_7785);
or U7879 (N_7879,N_7780,N_7708);
nand U7880 (N_7880,N_7752,N_7745);
and U7881 (N_7881,N_7785,N_7727);
nand U7882 (N_7882,N_7707,N_7753);
nand U7883 (N_7883,N_7738,N_7782);
nor U7884 (N_7884,N_7799,N_7767);
or U7885 (N_7885,N_7785,N_7791);
nor U7886 (N_7886,N_7706,N_7750);
and U7887 (N_7887,N_7737,N_7790);
nand U7888 (N_7888,N_7774,N_7748);
or U7889 (N_7889,N_7727,N_7782);
nor U7890 (N_7890,N_7786,N_7739);
nor U7891 (N_7891,N_7721,N_7715);
and U7892 (N_7892,N_7718,N_7785);
nand U7893 (N_7893,N_7753,N_7741);
or U7894 (N_7894,N_7776,N_7785);
nor U7895 (N_7895,N_7791,N_7752);
and U7896 (N_7896,N_7776,N_7775);
nand U7897 (N_7897,N_7713,N_7738);
nand U7898 (N_7898,N_7747,N_7769);
nor U7899 (N_7899,N_7791,N_7761);
or U7900 (N_7900,N_7860,N_7802);
nor U7901 (N_7901,N_7815,N_7830);
nand U7902 (N_7902,N_7866,N_7881);
nand U7903 (N_7903,N_7890,N_7885);
nor U7904 (N_7904,N_7827,N_7809);
nand U7905 (N_7905,N_7803,N_7872);
and U7906 (N_7906,N_7850,N_7818);
nor U7907 (N_7907,N_7873,N_7897);
or U7908 (N_7908,N_7804,N_7858);
or U7909 (N_7909,N_7822,N_7807);
nand U7910 (N_7910,N_7842,N_7859);
and U7911 (N_7911,N_7870,N_7849);
nor U7912 (N_7912,N_7886,N_7864);
nor U7913 (N_7913,N_7848,N_7820);
xor U7914 (N_7914,N_7835,N_7874);
nand U7915 (N_7915,N_7898,N_7896);
nor U7916 (N_7916,N_7862,N_7857);
or U7917 (N_7917,N_7892,N_7816);
or U7918 (N_7918,N_7891,N_7868);
xnor U7919 (N_7919,N_7819,N_7888);
and U7920 (N_7920,N_7847,N_7829);
nor U7921 (N_7921,N_7841,N_7801);
nor U7922 (N_7922,N_7882,N_7811);
nand U7923 (N_7923,N_7840,N_7812);
nor U7924 (N_7924,N_7861,N_7853);
and U7925 (N_7925,N_7877,N_7814);
xor U7926 (N_7926,N_7837,N_7887);
or U7927 (N_7927,N_7883,N_7832);
nand U7928 (N_7928,N_7894,N_7863);
nand U7929 (N_7929,N_7813,N_7893);
nand U7930 (N_7930,N_7834,N_7889);
or U7931 (N_7931,N_7838,N_7851);
and U7932 (N_7932,N_7867,N_7854);
and U7933 (N_7933,N_7839,N_7856);
and U7934 (N_7934,N_7831,N_7810);
nand U7935 (N_7935,N_7895,N_7869);
and U7936 (N_7936,N_7800,N_7836);
nor U7937 (N_7937,N_7844,N_7855);
xor U7938 (N_7938,N_7821,N_7843);
xor U7939 (N_7939,N_7852,N_7865);
xnor U7940 (N_7940,N_7880,N_7876);
and U7941 (N_7941,N_7806,N_7871);
nand U7942 (N_7942,N_7899,N_7824);
and U7943 (N_7943,N_7823,N_7878);
or U7944 (N_7944,N_7825,N_7875);
or U7945 (N_7945,N_7884,N_7879);
and U7946 (N_7946,N_7845,N_7833);
and U7947 (N_7947,N_7808,N_7828);
and U7948 (N_7948,N_7817,N_7846);
xor U7949 (N_7949,N_7826,N_7805);
nand U7950 (N_7950,N_7875,N_7821);
or U7951 (N_7951,N_7801,N_7845);
or U7952 (N_7952,N_7834,N_7892);
xor U7953 (N_7953,N_7833,N_7806);
nor U7954 (N_7954,N_7881,N_7841);
xnor U7955 (N_7955,N_7875,N_7884);
and U7956 (N_7956,N_7801,N_7837);
nand U7957 (N_7957,N_7826,N_7807);
xnor U7958 (N_7958,N_7896,N_7883);
nand U7959 (N_7959,N_7844,N_7859);
nor U7960 (N_7960,N_7826,N_7882);
xor U7961 (N_7961,N_7837,N_7892);
and U7962 (N_7962,N_7857,N_7889);
and U7963 (N_7963,N_7817,N_7840);
and U7964 (N_7964,N_7893,N_7896);
or U7965 (N_7965,N_7877,N_7819);
and U7966 (N_7966,N_7825,N_7866);
and U7967 (N_7967,N_7827,N_7818);
and U7968 (N_7968,N_7844,N_7815);
xor U7969 (N_7969,N_7800,N_7897);
xnor U7970 (N_7970,N_7806,N_7841);
nor U7971 (N_7971,N_7884,N_7849);
nor U7972 (N_7972,N_7857,N_7870);
nand U7973 (N_7973,N_7800,N_7879);
or U7974 (N_7974,N_7822,N_7886);
nand U7975 (N_7975,N_7884,N_7827);
and U7976 (N_7976,N_7895,N_7848);
nor U7977 (N_7977,N_7844,N_7890);
nand U7978 (N_7978,N_7859,N_7823);
nand U7979 (N_7979,N_7867,N_7853);
or U7980 (N_7980,N_7854,N_7805);
xor U7981 (N_7981,N_7853,N_7817);
or U7982 (N_7982,N_7813,N_7879);
nand U7983 (N_7983,N_7870,N_7830);
and U7984 (N_7984,N_7811,N_7804);
nand U7985 (N_7985,N_7887,N_7824);
nor U7986 (N_7986,N_7848,N_7812);
nor U7987 (N_7987,N_7850,N_7836);
or U7988 (N_7988,N_7861,N_7820);
and U7989 (N_7989,N_7810,N_7814);
or U7990 (N_7990,N_7862,N_7899);
or U7991 (N_7991,N_7839,N_7808);
or U7992 (N_7992,N_7843,N_7803);
nand U7993 (N_7993,N_7808,N_7835);
xnor U7994 (N_7994,N_7805,N_7815);
or U7995 (N_7995,N_7893,N_7837);
and U7996 (N_7996,N_7859,N_7890);
xnor U7997 (N_7997,N_7816,N_7844);
and U7998 (N_7998,N_7868,N_7827);
and U7999 (N_7999,N_7819,N_7878);
nand U8000 (N_8000,N_7922,N_7901);
and U8001 (N_8001,N_7941,N_7976);
nor U8002 (N_8002,N_7962,N_7977);
nand U8003 (N_8003,N_7903,N_7955);
nand U8004 (N_8004,N_7988,N_7948);
or U8005 (N_8005,N_7943,N_7917);
nand U8006 (N_8006,N_7942,N_7950);
nor U8007 (N_8007,N_7927,N_7907);
and U8008 (N_8008,N_7952,N_7945);
xnor U8009 (N_8009,N_7986,N_7937);
and U8010 (N_8010,N_7929,N_7919);
nand U8011 (N_8011,N_7908,N_7914);
nand U8012 (N_8012,N_7956,N_7969);
xnor U8013 (N_8013,N_7909,N_7981);
and U8014 (N_8014,N_7925,N_7918);
nor U8015 (N_8015,N_7989,N_7999);
nand U8016 (N_8016,N_7970,N_7972);
or U8017 (N_8017,N_7900,N_7973);
and U8018 (N_8018,N_7939,N_7985);
nand U8019 (N_8019,N_7931,N_7930);
nand U8020 (N_8020,N_7996,N_7957);
or U8021 (N_8021,N_7951,N_7947);
or U8022 (N_8022,N_7997,N_7983);
nor U8023 (N_8023,N_7993,N_7953);
or U8024 (N_8024,N_7932,N_7949);
nand U8025 (N_8025,N_7906,N_7958);
and U8026 (N_8026,N_7936,N_7912);
xnor U8027 (N_8027,N_7974,N_7926);
and U8028 (N_8028,N_7959,N_7995);
nand U8029 (N_8029,N_7928,N_7913);
and U8030 (N_8030,N_7984,N_7966);
or U8031 (N_8031,N_7946,N_7975);
nand U8032 (N_8032,N_7987,N_7965);
nor U8033 (N_8033,N_7979,N_7991);
nand U8034 (N_8034,N_7938,N_7924);
and U8035 (N_8035,N_7992,N_7916);
nor U8036 (N_8036,N_7982,N_7944);
or U8037 (N_8037,N_7921,N_7933);
or U8038 (N_8038,N_7994,N_7967);
and U8039 (N_8039,N_7954,N_7964);
nand U8040 (N_8040,N_7904,N_7980);
or U8041 (N_8041,N_7978,N_7910);
and U8042 (N_8042,N_7911,N_7963);
nor U8043 (N_8043,N_7990,N_7902);
nor U8044 (N_8044,N_7920,N_7905);
or U8045 (N_8045,N_7923,N_7934);
nor U8046 (N_8046,N_7935,N_7968);
and U8047 (N_8047,N_7961,N_7940);
or U8048 (N_8048,N_7971,N_7960);
nor U8049 (N_8049,N_7915,N_7998);
and U8050 (N_8050,N_7992,N_7954);
xor U8051 (N_8051,N_7971,N_7958);
nand U8052 (N_8052,N_7911,N_7932);
and U8053 (N_8053,N_7910,N_7991);
or U8054 (N_8054,N_7919,N_7935);
nand U8055 (N_8055,N_7964,N_7956);
nand U8056 (N_8056,N_7982,N_7994);
nand U8057 (N_8057,N_7926,N_7984);
nor U8058 (N_8058,N_7904,N_7957);
and U8059 (N_8059,N_7912,N_7913);
nor U8060 (N_8060,N_7968,N_7944);
or U8061 (N_8061,N_7938,N_7993);
or U8062 (N_8062,N_7990,N_7992);
nor U8063 (N_8063,N_7956,N_7959);
nor U8064 (N_8064,N_7939,N_7962);
nand U8065 (N_8065,N_7949,N_7945);
or U8066 (N_8066,N_7993,N_7957);
and U8067 (N_8067,N_7988,N_7919);
xor U8068 (N_8068,N_7900,N_7976);
nor U8069 (N_8069,N_7991,N_7983);
xnor U8070 (N_8070,N_7956,N_7971);
or U8071 (N_8071,N_7979,N_7954);
xor U8072 (N_8072,N_7912,N_7996);
nor U8073 (N_8073,N_7902,N_7955);
nand U8074 (N_8074,N_7981,N_7960);
and U8075 (N_8075,N_7946,N_7974);
or U8076 (N_8076,N_7997,N_7920);
xnor U8077 (N_8077,N_7977,N_7980);
and U8078 (N_8078,N_7904,N_7948);
nand U8079 (N_8079,N_7962,N_7980);
and U8080 (N_8080,N_7986,N_7918);
and U8081 (N_8081,N_7922,N_7996);
nor U8082 (N_8082,N_7927,N_7934);
nand U8083 (N_8083,N_7945,N_7911);
and U8084 (N_8084,N_7916,N_7961);
or U8085 (N_8085,N_7972,N_7959);
nand U8086 (N_8086,N_7914,N_7988);
and U8087 (N_8087,N_7985,N_7923);
and U8088 (N_8088,N_7976,N_7975);
and U8089 (N_8089,N_7910,N_7921);
nand U8090 (N_8090,N_7920,N_7982);
or U8091 (N_8091,N_7943,N_7959);
or U8092 (N_8092,N_7968,N_7927);
and U8093 (N_8093,N_7908,N_7938);
nor U8094 (N_8094,N_7963,N_7906);
xnor U8095 (N_8095,N_7979,N_7957);
xor U8096 (N_8096,N_7932,N_7939);
nor U8097 (N_8097,N_7906,N_7937);
nor U8098 (N_8098,N_7947,N_7900);
nand U8099 (N_8099,N_7991,N_7992);
and U8100 (N_8100,N_8005,N_8052);
nand U8101 (N_8101,N_8048,N_8046);
and U8102 (N_8102,N_8086,N_8028);
xnor U8103 (N_8103,N_8054,N_8049);
nor U8104 (N_8104,N_8080,N_8050);
and U8105 (N_8105,N_8061,N_8074);
or U8106 (N_8106,N_8081,N_8036);
nor U8107 (N_8107,N_8065,N_8075);
and U8108 (N_8108,N_8014,N_8082);
nor U8109 (N_8109,N_8042,N_8066);
nor U8110 (N_8110,N_8084,N_8015);
nor U8111 (N_8111,N_8009,N_8033);
and U8112 (N_8112,N_8023,N_8022);
and U8113 (N_8113,N_8092,N_8039);
nand U8114 (N_8114,N_8000,N_8097);
nand U8115 (N_8115,N_8063,N_8071);
xor U8116 (N_8116,N_8011,N_8002);
nand U8117 (N_8117,N_8057,N_8090);
nor U8118 (N_8118,N_8016,N_8067);
nand U8119 (N_8119,N_8085,N_8013);
nand U8120 (N_8120,N_8055,N_8034);
nor U8121 (N_8121,N_8051,N_8026);
or U8122 (N_8122,N_8091,N_8038);
and U8123 (N_8123,N_8087,N_8025);
or U8124 (N_8124,N_8072,N_8064);
and U8125 (N_8125,N_8068,N_8032);
nor U8126 (N_8126,N_8044,N_8098);
nor U8127 (N_8127,N_8010,N_8088);
xnor U8128 (N_8128,N_8073,N_8012);
nor U8129 (N_8129,N_8037,N_8008);
nor U8130 (N_8130,N_8030,N_8062);
or U8131 (N_8131,N_8093,N_8070);
nor U8132 (N_8132,N_8056,N_8004);
and U8133 (N_8133,N_8017,N_8076);
nand U8134 (N_8134,N_8060,N_8096);
nor U8135 (N_8135,N_8024,N_8007);
xnor U8136 (N_8136,N_8058,N_8099);
nor U8137 (N_8137,N_8003,N_8095);
nor U8138 (N_8138,N_8040,N_8006);
nor U8139 (N_8139,N_8089,N_8069);
xor U8140 (N_8140,N_8035,N_8027);
nor U8141 (N_8141,N_8020,N_8018);
nand U8142 (N_8142,N_8094,N_8001);
nor U8143 (N_8143,N_8053,N_8059);
xnor U8144 (N_8144,N_8029,N_8043);
or U8145 (N_8145,N_8083,N_8021);
or U8146 (N_8146,N_8047,N_8041);
or U8147 (N_8147,N_8031,N_8078);
or U8148 (N_8148,N_8077,N_8045);
nor U8149 (N_8149,N_8019,N_8079);
nor U8150 (N_8150,N_8044,N_8077);
and U8151 (N_8151,N_8025,N_8019);
nand U8152 (N_8152,N_8062,N_8058);
xor U8153 (N_8153,N_8034,N_8006);
nor U8154 (N_8154,N_8078,N_8022);
nor U8155 (N_8155,N_8091,N_8014);
nor U8156 (N_8156,N_8092,N_8074);
nor U8157 (N_8157,N_8090,N_8004);
nand U8158 (N_8158,N_8046,N_8067);
or U8159 (N_8159,N_8009,N_8090);
xnor U8160 (N_8160,N_8006,N_8092);
nor U8161 (N_8161,N_8095,N_8037);
nor U8162 (N_8162,N_8007,N_8025);
nand U8163 (N_8163,N_8075,N_8068);
and U8164 (N_8164,N_8042,N_8088);
nand U8165 (N_8165,N_8008,N_8097);
nor U8166 (N_8166,N_8031,N_8062);
or U8167 (N_8167,N_8010,N_8031);
xor U8168 (N_8168,N_8053,N_8073);
xor U8169 (N_8169,N_8029,N_8030);
nor U8170 (N_8170,N_8041,N_8076);
xnor U8171 (N_8171,N_8046,N_8034);
nor U8172 (N_8172,N_8093,N_8057);
nor U8173 (N_8173,N_8023,N_8092);
or U8174 (N_8174,N_8039,N_8023);
and U8175 (N_8175,N_8012,N_8009);
or U8176 (N_8176,N_8037,N_8018);
or U8177 (N_8177,N_8066,N_8085);
nand U8178 (N_8178,N_8004,N_8083);
or U8179 (N_8179,N_8089,N_8035);
or U8180 (N_8180,N_8075,N_8066);
nor U8181 (N_8181,N_8021,N_8011);
nor U8182 (N_8182,N_8041,N_8039);
or U8183 (N_8183,N_8001,N_8027);
xnor U8184 (N_8184,N_8079,N_8083);
and U8185 (N_8185,N_8028,N_8043);
nand U8186 (N_8186,N_8038,N_8037);
nand U8187 (N_8187,N_8042,N_8033);
and U8188 (N_8188,N_8035,N_8080);
nor U8189 (N_8189,N_8047,N_8053);
or U8190 (N_8190,N_8001,N_8075);
or U8191 (N_8191,N_8086,N_8099);
nand U8192 (N_8192,N_8074,N_8032);
and U8193 (N_8193,N_8013,N_8007);
and U8194 (N_8194,N_8081,N_8082);
nand U8195 (N_8195,N_8041,N_8098);
and U8196 (N_8196,N_8012,N_8030);
nor U8197 (N_8197,N_8045,N_8024);
nor U8198 (N_8198,N_8051,N_8009);
and U8199 (N_8199,N_8055,N_8049);
nor U8200 (N_8200,N_8157,N_8105);
or U8201 (N_8201,N_8166,N_8140);
and U8202 (N_8202,N_8113,N_8141);
nand U8203 (N_8203,N_8182,N_8180);
nand U8204 (N_8204,N_8162,N_8153);
xnor U8205 (N_8205,N_8174,N_8123);
or U8206 (N_8206,N_8164,N_8172);
or U8207 (N_8207,N_8171,N_8159);
nand U8208 (N_8208,N_8181,N_8104);
nor U8209 (N_8209,N_8184,N_8132);
and U8210 (N_8210,N_8160,N_8173);
and U8211 (N_8211,N_8103,N_8117);
nor U8212 (N_8212,N_8185,N_8142);
and U8213 (N_8213,N_8102,N_8150);
and U8214 (N_8214,N_8110,N_8115);
nor U8215 (N_8215,N_8175,N_8138);
or U8216 (N_8216,N_8177,N_8167);
and U8217 (N_8217,N_8116,N_8129);
nand U8218 (N_8218,N_8196,N_8198);
nor U8219 (N_8219,N_8120,N_8109);
nand U8220 (N_8220,N_8146,N_8191);
nand U8221 (N_8221,N_8128,N_8137);
nor U8222 (N_8222,N_8118,N_8139);
nor U8223 (N_8223,N_8189,N_8168);
nor U8224 (N_8224,N_8188,N_8163);
nand U8225 (N_8225,N_8156,N_8122);
and U8226 (N_8226,N_8183,N_8127);
or U8227 (N_8227,N_8158,N_8161);
nor U8228 (N_8228,N_8195,N_8179);
nand U8229 (N_8229,N_8147,N_8145);
nand U8230 (N_8230,N_8165,N_8199);
and U8231 (N_8231,N_8190,N_8112);
nor U8232 (N_8232,N_8111,N_8192);
or U8233 (N_8233,N_8149,N_8126);
nor U8234 (N_8234,N_8197,N_8152);
and U8235 (N_8235,N_8101,N_8134);
nor U8236 (N_8236,N_8154,N_8100);
or U8237 (N_8237,N_8124,N_8121);
or U8238 (N_8238,N_8133,N_8136);
and U8239 (N_8239,N_8114,N_8186);
nor U8240 (N_8240,N_8178,N_8130);
and U8241 (N_8241,N_8194,N_8143);
and U8242 (N_8242,N_8170,N_8144);
nor U8243 (N_8243,N_8106,N_8151);
nand U8244 (N_8244,N_8107,N_8125);
or U8245 (N_8245,N_8148,N_8176);
nor U8246 (N_8246,N_8193,N_8155);
nor U8247 (N_8247,N_8187,N_8169);
and U8248 (N_8248,N_8119,N_8131);
nand U8249 (N_8249,N_8135,N_8108);
or U8250 (N_8250,N_8108,N_8124);
nor U8251 (N_8251,N_8190,N_8192);
nor U8252 (N_8252,N_8128,N_8182);
xnor U8253 (N_8253,N_8143,N_8191);
or U8254 (N_8254,N_8147,N_8188);
or U8255 (N_8255,N_8120,N_8136);
or U8256 (N_8256,N_8159,N_8149);
nand U8257 (N_8257,N_8174,N_8155);
and U8258 (N_8258,N_8130,N_8111);
and U8259 (N_8259,N_8140,N_8125);
or U8260 (N_8260,N_8183,N_8147);
xor U8261 (N_8261,N_8198,N_8146);
nor U8262 (N_8262,N_8130,N_8190);
and U8263 (N_8263,N_8118,N_8194);
nand U8264 (N_8264,N_8128,N_8105);
xor U8265 (N_8265,N_8149,N_8102);
nor U8266 (N_8266,N_8132,N_8188);
nor U8267 (N_8267,N_8197,N_8108);
nor U8268 (N_8268,N_8152,N_8114);
or U8269 (N_8269,N_8116,N_8130);
and U8270 (N_8270,N_8127,N_8194);
nor U8271 (N_8271,N_8153,N_8110);
or U8272 (N_8272,N_8176,N_8144);
nand U8273 (N_8273,N_8126,N_8150);
nand U8274 (N_8274,N_8132,N_8173);
and U8275 (N_8275,N_8173,N_8135);
and U8276 (N_8276,N_8163,N_8111);
nor U8277 (N_8277,N_8104,N_8117);
nand U8278 (N_8278,N_8104,N_8174);
or U8279 (N_8279,N_8171,N_8113);
or U8280 (N_8280,N_8170,N_8112);
nor U8281 (N_8281,N_8153,N_8167);
nand U8282 (N_8282,N_8113,N_8129);
or U8283 (N_8283,N_8110,N_8176);
and U8284 (N_8284,N_8118,N_8187);
nand U8285 (N_8285,N_8105,N_8162);
nor U8286 (N_8286,N_8144,N_8100);
xor U8287 (N_8287,N_8146,N_8101);
nand U8288 (N_8288,N_8117,N_8168);
nand U8289 (N_8289,N_8191,N_8137);
or U8290 (N_8290,N_8145,N_8137);
and U8291 (N_8291,N_8155,N_8180);
nor U8292 (N_8292,N_8174,N_8152);
nor U8293 (N_8293,N_8158,N_8156);
nand U8294 (N_8294,N_8196,N_8132);
xnor U8295 (N_8295,N_8118,N_8137);
nor U8296 (N_8296,N_8145,N_8111);
xor U8297 (N_8297,N_8153,N_8121);
and U8298 (N_8298,N_8181,N_8120);
nand U8299 (N_8299,N_8179,N_8128);
nand U8300 (N_8300,N_8260,N_8265);
nor U8301 (N_8301,N_8292,N_8220);
and U8302 (N_8302,N_8296,N_8270);
nor U8303 (N_8303,N_8299,N_8225);
nor U8304 (N_8304,N_8238,N_8208);
or U8305 (N_8305,N_8274,N_8261);
or U8306 (N_8306,N_8281,N_8224);
or U8307 (N_8307,N_8259,N_8207);
and U8308 (N_8308,N_8269,N_8257);
or U8309 (N_8309,N_8293,N_8201);
and U8310 (N_8310,N_8249,N_8278);
nand U8311 (N_8311,N_8233,N_8230);
nand U8312 (N_8312,N_8277,N_8285);
nand U8313 (N_8313,N_8222,N_8240);
nand U8314 (N_8314,N_8203,N_8241);
nand U8315 (N_8315,N_8227,N_8243);
nor U8316 (N_8316,N_8275,N_8219);
nor U8317 (N_8317,N_8213,N_8264);
nand U8318 (N_8318,N_8256,N_8286);
or U8319 (N_8319,N_8202,N_8221);
or U8320 (N_8320,N_8237,N_8223);
and U8321 (N_8321,N_8295,N_8284);
and U8322 (N_8322,N_8282,N_8287);
nand U8323 (N_8323,N_8267,N_8239);
or U8324 (N_8324,N_8288,N_8247);
nand U8325 (N_8325,N_8210,N_8217);
nand U8326 (N_8326,N_8266,N_8268);
or U8327 (N_8327,N_8228,N_8234);
or U8328 (N_8328,N_8200,N_8253);
or U8329 (N_8329,N_8216,N_8211);
nand U8330 (N_8330,N_8258,N_8279);
xor U8331 (N_8331,N_8205,N_8272);
and U8332 (N_8332,N_8242,N_8215);
nor U8333 (N_8333,N_8289,N_8214);
nor U8334 (N_8334,N_8229,N_8232);
nand U8335 (N_8335,N_8248,N_8276);
nand U8336 (N_8336,N_8218,N_8235);
nand U8337 (N_8337,N_8290,N_8244);
and U8338 (N_8338,N_8236,N_8273);
or U8339 (N_8339,N_8204,N_8226);
and U8340 (N_8340,N_8298,N_8212);
xor U8341 (N_8341,N_8262,N_8231);
xnor U8342 (N_8342,N_8209,N_8246);
nor U8343 (N_8343,N_8297,N_8255);
nand U8344 (N_8344,N_8283,N_8263);
nor U8345 (N_8345,N_8251,N_8254);
xor U8346 (N_8346,N_8252,N_8271);
nand U8347 (N_8347,N_8294,N_8206);
nor U8348 (N_8348,N_8245,N_8280);
or U8349 (N_8349,N_8250,N_8291);
or U8350 (N_8350,N_8237,N_8226);
and U8351 (N_8351,N_8261,N_8209);
xor U8352 (N_8352,N_8256,N_8215);
nand U8353 (N_8353,N_8295,N_8218);
nor U8354 (N_8354,N_8292,N_8219);
nand U8355 (N_8355,N_8273,N_8244);
nor U8356 (N_8356,N_8263,N_8287);
nand U8357 (N_8357,N_8244,N_8275);
nand U8358 (N_8358,N_8203,N_8205);
nand U8359 (N_8359,N_8251,N_8265);
and U8360 (N_8360,N_8212,N_8225);
and U8361 (N_8361,N_8298,N_8254);
xnor U8362 (N_8362,N_8283,N_8284);
and U8363 (N_8363,N_8270,N_8222);
or U8364 (N_8364,N_8203,N_8211);
and U8365 (N_8365,N_8294,N_8256);
and U8366 (N_8366,N_8249,N_8241);
nand U8367 (N_8367,N_8223,N_8257);
and U8368 (N_8368,N_8271,N_8266);
or U8369 (N_8369,N_8234,N_8250);
nor U8370 (N_8370,N_8204,N_8225);
nand U8371 (N_8371,N_8243,N_8238);
and U8372 (N_8372,N_8233,N_8249);
nand U8373 (N_8373,N_8200,N_8294);
or U8374 (N_8374,N_8263,N_8239);
or U8375 (N_8375,N_8273,N_8234);
and U8376 (N_8376,N_8294,N_8211);
xnor U8377 (N_8377,N_8200,N_8281);
nand U8378 (N_8378,N_8299,N_8292);
and U8379 (N_8379,N_8258,N_8263);
and U8380 (N_8380,N_8233,N_8269);
nor U8381 (N_8381,N_8234,N_8275);
nor U8382 (N_8382,N_8212,N_8270);
nand U8383 (N_8383,N_8214,N_8215);
nor U8384 (N_8384,N_8224,N_8213);
and U8385 (N_8385,N_8255,N_8230);
nand U8386 (N_8386,N_8252,N_8246);
and U8387 (N_8387,N_8260,N_8250);
and U8388 (N_8388,N_8274,N_8258);
or U8389 (N_8389,N_8258,N_8229);
nand U8390 (N_8390,N_8256,N_8291);
or U8391 (N_8391,N_8294,N_8220);
or U8392 (N_8392,N_8215,N_8255);
and U8393 (N_8393,N_8283,N_8298);
or U8394 (N_8394,N_8227,N_8245);
or U8395 (N_8395,N_8272,N_8254);
and U8396 (N_8396,N_8251,N_8286);
nor U8397 (N_8397,N_8277,N_8271);
nand U8398 (N_8398,N_8228,N_8204);
and U8399 (N_8399,N_8220,N_8244);
nor U8400 (N_8400,N_8303,N_8330);
and U8401 (N_8401,N_8386,N_8313);
and U8402 (N_8402,N_8380,N_8385);
and U8403 (N_8403,N_8323,N_8331);
nor U8404 (N_8404,N_8325,N_8389);
nor U8405 (N_8405,N_8314,N_8304);
nand U8406 (N_8406,N_8375,N_8382);
and U8407 (N_8407,N_8376,N_8337);
and U8408 (N_8408,N_8377,N_8362);
and U8409 (N_8409,N_8366,N_8394);
xnor U8410 (N_8410,N_8347,N_8332);
and U8411 (N_8411,N_8356,N_8398);
or U8412 (N_8412,N_8348,N_8317);
and U8413 (N_8413,N_8343,N_8378);
or U8414 (N_8414,N_8360,N_8396);
nor U8415 (N_8415,N_8300,N_8354);
nand U8416 (N_8416,N_8383,N_8310);
nor U8417 (N_8417,N_8312,N_8335);
nor U8418 (N_8418,N_8399,N_8324);
nor U8419 (N_8419,N_8365,N_8326);
and U8420 (N_8420,N_8372,N_8315);
xnor U8421 (N_8421,N_8363,N_8357);
nor U8422 (N_8422,N_8334,N_8327);
or U8423 (N_8423,N_8319,N_8374);
or U8424 (N_8424,N_8373,N_8328);
nand U8425 (N_8425,N_8390,N_8336);
xor U8426 (N_8426,N_8395,N_8381);
nor U8427 (N_8427,N_8345,N_8338);
or U8428 (N_8428,N_8309,N_8369);
and U8429 (N_8429,N_8387,N_8393);
nand U8430 (N_8430,N_8397,N_8371);
nand U8431 (N_8431,N_8350,N_8322);
or U8432 (N_8432,N_8392,N_8388);
nand U8433 (N_8433,N_8341,N_8329);
and U8434 (N_8434,N_8361,N_8391);
nand U8435 (N_8435,N_8301,N_8379);
and U8436 (N_8436,N_8307,N_8384);
nand U8437 (N_8437,N_8305,N_8306);
or U8438 (N_8438,N_8318,N_8358);
or U8439 (N_8439,N_8339,N_8342);
nand U8440 (N_8440,N_8344,N_8368);
nand U8441 (N_8441,N_8364,N_8340);
and U8442 (N_8442,N_8359,N_8352);
and U8443 (N_8443,N_8367,N_8355);
and U8444 (N_8444,N_8308,N_8316);
nand U8445 (N_8445,N_8346,N_8321);
nor U8446 (N_8446,N_8311,N_8349);
nand U8447 (N_8447,N_8370,N_8320);
nand U8448 (N_8448,N_8333,N_8351);
or U8449 (N_8449,N_8302,N_8353);
nand U8450 (N_8450,N_8351,N_8349);
and U8451 (N_8451,N_8392,N_8344);
and U8452 (N_8452,N_8321,N_8388);
nand U8453 (N_8453,N_8399,N_8375);
xor U8454 (N_8454,N_8382,N_8316);
or U8455 (N_8455,N_8396,N_8328);
or U8456 (N_8456,N_8324,N_8304);
xnor U8457 (N_8457,N_8376,N_8347);
or U8458 (N_8458,N_8394,N_8375);
and U8459 (N_8459,N_8368,N_8309);
nand U8460 (N_8460,N_8345,N_8337);
nor U8461 (N_8461,N_8317,N_8338);
or U8462 (N_8462,N_8385,N_8364);
nor U8463 (N_8463,N_8330,N_8341);
nand U8464 (N_8464,N_8373,N_8375);
or U8465 (N_8465,N_8317,N_8311);
nand U8466 (N_8466,N_8358,N_8385);
xor U8467 (N_8467,N_8389,N_8340);
nand U8468 (N_8468,N_8376,N_8303);
nand U8469 (N_8469,N_8325,N_8387);
nand U8470 (N_8470,N_8387,N_8376);
nor U8471 (N_8471,N_8326,N_8378);
xnor U8472 (N_8472,N_8397,N_8366);
or U8473 (N_8473,N_8310,N_8355);
and U8474 (N_8474,N_8383,N_8326);
and U8475 (N_8475,N_8350,N_8307);
nand U8476 (N_8476,N_8321,N_8328);
nor U8477 (N_8477,N_8330,N_8394);
nand U8478 (N_8478,N_8393,N_8302);
nand U8479 (N_8479,N_8307,N_8329);
nand U8480 (N_8480,N_8381,N_8355);
nand U8481 (N_8481,N_8372,N_8314);
nor U8482 (N_8482,N_8341,N_8332);
and U8483 (N_8483,N_8308,N_8367);
and U8484 (N_8484,N_8383,N_8389);
and U8485 (N_8485,N_8350,N_8327);
and U8486 (N_8486,N_8341,N_8339);
nor U8487 (N_8487,N_8378,N_8353);
or U8488 (N_8488,N_8353,N_8308);
xor U8489 (N_8489,N_8382,N_8351);
nor U8490 (N_8490,N_8312,N_8316);
nor U8491 (N_8491,N_8347,N_8326);
nor U8492 (N_8492,N_8346,N_8364);
nor U8493 (N_8493,N_8316,N_8349);
or U8494 (N_8494,N_8327,N_8393);
nor U8495 (N_8495,N_8328,N_8313);
and U8496 (N_8496,N_8374,N_8358);
nor U8497 (N_8497,N_8379,N_8335);
nor U8498 (N_8498,N_8396,N_8373);
or U8499 (N_8499,N_8314,N_8366);
and U8500 (N_8500,N_8424,N_8470);
and U8501 (N_8501,N_8433,N_8477);
xor U8502 (N_8502,N_8482,N_8496);
xnor U8503 (N_8503,N_8420,N_8407);
nand U8504 (N_8504,N_8411,N_8471);
and U8505 (N_8505,N_8475,N_8488);
or U8506 (N_8506,N_8435,N_8403);
and U8507 (N_8507,N_8416,N_8493);
nor U8508 (N_8508,N_8401,N_8423);
xnor U8509 (N_8509,N_8485,N_8434);
nor U8510 (N_8510,N_8427,N_8418);
nand U8511 (N_8511,N_8480,N_8442);
nand U8512 (N_8512,N_8458,N_8445);
nor U8513 (N_8513,N_8492,N_8473);
nor U8514 (N_8514,N_8455,N_8464);
and U8515 (N_8515,N_8422,N_8443);
nor U8516 (N_8516,N_8454,N_8481);
nand U8517 (N_8517,N_8487,N_8486);
nand U8518 (N_8518,N_8456,N_8429);
nand U8519 (N_8519,N_8465,N_8446);
or U8520 (N_8520,N_8400,N_8436);
or U8521 (N_8521,N_8404,N_8415);
xor U8522 (N_8522,N_8406,N_8438);
and U8523 (N_8523,N_8457,N_8426);
or U8524 (N_8524,N_8450,N_8484);
or U8525 (N_8525,N_8462,N_8444);
xor U8526 (N_8526,N_8490,N_8421);
or U8527 (N_8527,N_8408,N_8483);
or U8528 (N_8528,N_8494,N_8437);
nor U8529 (N_8529,N_8453,N_8409);
or U8530 (N_8530,N_8402,N_8447);
nor U8531 (N_8531,N_8468,N_8466);
or U8532 (N_8532,N_8451,N_8441);
nor U8533 (N_8533,N_8491,N_8495);
and U8534 (N_8534,N_8417,N_8413);
or U8535 (N_8535,N_8474,N_8472);
xor U8536 (N_8536,N_8431,N_8432);
nor U8537 (N_8537,N_8461,N_8405);
and U8538 (N_8538,N_8476,N_8410);
xnor U8539 (N_8539,N_8430,N_8440);
or U8540 (N_8540,N_8412,N_8479);
and U8541 (N_8541,N_8428,N_8469);
or U8542 (N_8542,N_8452,N_8439);
nor U8543 (N_8543,N_8489,N_8425);
and U8544 (N_8544,N_8448,N_8478);
and U8545 (N_8545,N_8467,N_8498);
and U8546 (N_8546,N_8460,N_8463);
nor U8547 (N_8547,N_8499,N_8459);
or U8548 (N_8548,N_8419,N_8497);
nor U8549 (N_8549,N_8449,N_8414);
or U8550 (N_8550,N_8401,N_8436);
nor U8551 (N_8551,N_8459,N_8468);
nand U8552 (N_8552,N_8411,N_8464);
xnor U8553 (N_8553,N_8412,N_8474);
and U8554 (N_8554,N_8430,N_8486);
or U8555 (N_8555,N_8448,N_8420);
or U8556 (N_8556,N_8424,N_8455);
xnor U8557 (N_8557,N_8461,N_8443);
or U8558 (N_8558,N_8409,N_8440);
or U8559 (N_8559,N_8464,N_8462);
and U8560 (N_8560,N_8495,N_8410);
nor U8561 (N_8561,N_8475,N_8474);
and U8562 (N_8562,N_8493,N_8414);
nor U8563 (N_8563,N_8470,N_8419);
or U8564 (N_8564,N_8473,N_8412);
xnor U8565 (N_8565,N_8444,N_8460);
or U8566 (N_8566,N_8493,N_8433);
and U8567 (N_8567,N_8408,N_8472);
nand U8568 (N_8568,N_8431,N_8455);
nor U8569 (N_8569,N_8417,N_8493);
and U8570 (N_8570,N_8497,N_8479);
nand U8571 (N_8571,N_8455,N_8410);
nor U8572 (N_8572,N_8431,N_8438);
nand U8573 (N_8573,N_8472,N_8403);
and U8574 (N_8574,N_8417,N_8465);
or U8575 (N_8575,N_8451,N_8476);
xnor U8576 (N_8576,N_8454,N_8459);
and U8577 (N_8577,N_8403,N_8450);
xor U8578 (N_8578,N_8442,N_8482);
xnor U8579 (N_8579,N_8409,N_8444);
nor U8580 (N_8580,N_8449,N_8486);
nand U8581 (N_8581,N_8421,N_8418);
nand U8582 (N_8582,N_8458,N_8495);
or U8583 (N_8583,N_8443,N_8473);
nor U8584 (N_8584,N_8444,N_8496);
nor U8585 (N_8585,N_8444,N_8400);
xnor U8586 (N_8586,N_8437,N_8439);
xor U8587 (N_8587,N_8497,N_8476);
xor U8588 (N_8588,N_8402,N_8429);
or U8589 (N_8589,N_8425,N_8412);
nand U8590 (N_8590,N_8424,N_8406);
or U8591 (N_8591,N_8433,N_8463);
or U8592 (N_8592,N_8488,N_8445);
and U8593 (N_8593,N_8489,N_8456);
or U8594 (N_8594,N_8471,N_8480);
nand U8595 (N_8595,N_8434,N_8427);
nand U8596 (N_8596,N_8453,N_8415);
nand U8597 (N_8597,N_8472,N_8455);
nand U8598 (N_8598,N_8424,N_8483);
nand U8599 (N_8599,N_8413,N_8427);
nand U8600 (N_8600,N_8536,N_8505);
xnor U8601 (N_8601,N_8502,N_8573);
nor U8602 (N_8602,N_8576,N_8586);
or U8603 (N_8603,N_8588,N_8533);
nor U8604 (N_8604,N_8561,N_8577);
nand U8605 (N_8605,N_8593,N_8500);
and U8606 (N_8606,N_8567,N_8504);
or U8607 (N_8607,N_8558,N_8524);
or U8608 (N_8608,N_8572,N_8544);
and U8609 (N_8609,N_8590,N_8569);
nor U8610 (N_8610,N_8597,N_8591);
and U8611 (N_8611,N_8522,N_8506);
nor U8612 (N_8612,N_8552,N_8582);
nand U8613 (N_8613,N_8555,N_8589);
nand U8614 (N_8614,N_8532,N_8512);
nand U8615 (N_8615,N_8540,N_8546);
nor U8616 (N_8616,N_8548,N_8580);
nand U8617 (N_8617,N_8517,N_8518);
nand U8618 (N_8618,N_8543,N_8519);
nand U8619 (N_8619,N_8515,N_8538);
or U8620 (N_8620,N_8514,N_8581);
and U8621 (N_8621,N_8553,N_8551);
nand U8622 (N_8622,N_8531,N_8564);
or U8623 (N_8623,N_8501,N_8545);
nand U8624 (N_8624,N_8584,N_8583);
nor U8625 (N_8625,N_8575,N_8598);
nand U8626 (N_8626,N_8513,N_8563);
nor U8627 (N_8627,N_8559,N_8556);
and U8628 (N_8628,N_8579,N_8535);
nand U8629 (N_8629,N_8596,N_8539);
nand U8630 (N_8630,N_8510,N_8578);
nand U8631 (N_8631,N_8521,N_8520);
and U8632 (N_8632,N_8527,N_8587);
or U8633 (N_8633,N_8537,N_8550);
nor U8634 (N_8634,N_8523,N_8560);
xnor U8635 (N_8635,N_8547,N_8507);
nor U8636 (N_8636,N_8528,N_8599);
nor U8637 (N_8637,N_8534,N_8595);
and U8638 (N_8638,N_8554,N_8594);
nor U8639 (N_8639,N_8562,N_8565);
or U8640 (N_8640,N_8530,N_8585);
or U8641 (N_8641,N_8557,N_8571);
nor U8642 (N_8642,N_8503,N_8525);
or U8643 (N_8643,N_8509,N_8529);
nand U8644 (N_8644,N_8542,N_8541);
nor U8645 (N_8645,N_8511,N_8549);
or U8646 (N_8646,N_8592,N_8574);
nor U8647 (N_8647,N_8568,N_8516);
nor U8648 (N_8648,N_8526,N_8566);
nor U8649 (N_8649,N_8508,N_8570);
and U8650 (N_8650,N_8507,N_8568);
nand U8651 (N_8651,N_8519,N_8536);
xor U8652 (N_8652,N_8579,N_8529);
and U8653 (N_8653,N_8501,N_8540);
xor U8654 (N_8654,N_8577,N_8597);
and U8655 (N_8655,N_8506,N_8523);
or U8656 (N_8656,N_8598,N_8531);
nor U8657 (N_8657,N_8577,N_8540);
or U8658 (N_8658,N_8544,N_8523);
nor U8659 (N_8659,N_8536,N_8533);
or U8660 (N_8660,N_8515,N_8504);
and U8661 (N_8661,N_8539,N_8501);
or U8662 (N_8662,N_8518,N_8502);
nand U8663 (N_8663,N_8540,N_8596);
or U8664 (N_8664,N_8582,N_8587);
and U8665 (N_8665,N_8566,N_8569);
nor U8666 (N_8666,N_8500,N_8521);
or U8667 (N_8667,N_8517,N_8504);
nand U8668 (N_8668,N_8508,N_8571);
nand U8669 (N_8669,N_8555,N_8543);
nand U8670 (N_8670,N_8565,N_8525);
and U8671 (N_8671,N_8579,N_8550);
nor U8672 (N_8672,N_8580,N_8574);
nand U8673 (N_8673,N_8578,N_8550);
nand U8674 (N_8674,N_8523,N_8522);
nor U8675 (N_8675,N_8589,N_8581);
or U8676 (N_8676,N_8551,N_8519);
nand U8677 (N_8677,N_8541,N_8527);
and U8678 (N_8678,N_8553,N_8517);
xnor U8679 (N_8679,N_8570,N_8512);
nor U8680 (N_8680,N_8563,N_8596);
nor U8681 (N_8681,N_8532,N_8523);
nor U8682 (N_8682,N_8505,N_8588);
or U8683 (N_8683,N_8575,N_8554);
or U8684 (N_8684,N_8569,N_8551);
nand U8685 (N_8685,N_8522,N_8598);
nor U8686 (N_8686,N_8500,N_8599);
xor U8687 (N_8687,N_8551,N_8584);
nor U8688 (N_8688,N_8537,N_8544);
nor U8689 (N_8689,N_8508,N_8562);
nor U8690 (N_8690,N_8513,N_8516);
nand U8691 (N_8691,N_8563,N_8503);
and U8692 (N_8692,N_8535,N_8537);
and U8693 (N_8693,N_8512,N_8559);
nor U8694 (N_8694,N_8534,N_8502);
nor U8695 (N_8695,N_8517,N_8527);
and U8696 (N_8696,N_8590,N_8592);
xnor U8697 (N_8697,N_8575,N_8510);
nor U8698 (N_8698,N_8524,N_8561);
nand U8699 (N_8699,N_8538,N_8510);
nand U8700 (N_8700,N_8681,N_8605);
nand U8701 (N_8701,N_8634,N_8601);
nor U8702 (N_8702,N_8614,N_8649);
or U8703 (N_8703,N_8629,N_8622);
nand U8704 (N_8704,N_8621,N_8635);
nand U8705 (N_8705,N_8647,N_8626);
nor U8706 (N_8706,N_8664,N_8662);
nor U8707 (N_8707,N_8625,N_8666);
and U8708 (N_8708,N_8610,N_8640);
or U8709 (N_8709,N_8620,N_8643);
nand U8710 (N_8710,N_8637,N_8656);
xor U8711 (N_8711,N_8683,N_8676);
or U8712 (N_8712,N_8693,N_8657);
or U8713 (N_8713,N_8630,N_8663);
or U8714 (N_8714,N_8609,N_8668);
and U8715 (N_8715,N_8651,N_8680);
nor U8716 (N_8716,N_8636,N_8603);
nor U8717 (N_8717,N_8642,N_8624);
and U8718 (N_8718,N_8646,N_8616);
or U8719 (N_8719,N_8691,N_8644);
nor U8720 (N_8720,N_8687,N_8698);
or U8721 (N_8721,N_8632,N_8623);
nor U8722 (N_8722,N_8655,N_8678);
and U8723 (N_8723,N_8611,N_8694);
xor U8724 (N_8724,N_8653,N_8665);
nor U8725 (N_8725,N_8602,N_8679);
nor U8726 (N_8726,N_8695,N_8689);
and U8727 (N_8727,N_8650,N_8669);
or U8728 (N_8728,N_8652,N_8600);
and U8729 (N_8729,N_8670,N_8682);
and U8730 (N_8730,N_8692,N_8627);
and U8731 (N_8731,N_8671,N_8638);
and U8732 (N_8732,N_8639,N_8615);
or U8733 (N_8733,N_8612,N_8606);
nor U8734 (N_8734,N_8667,N_8631);
nor U8735 (N_8735,N_8613,N_8633);
and U8736 (N_8736,N_8673,N_8608);
nand U8737 (N_8737,N_8628,N_8618);
and U8738 (N_8738,N_8685,N_8675);
or U8739 (N_8739,N_8696,N_8674);
and U8740 (N_8740,N_8661,N_8648);
nor U8741 (N_8741,N_8617,N_8641);
and U8742 (N_8742,N_8604,N_8686);
nor U8743 (N_8743,N_8688,N_8697);
nand U8744 (N_8744,N_8660,N_8619);
or U8745 (N_8745,N_8659,N_8690);
nor U8746 (N_8746,N_8607,N_8677);
and U8747 (N_8747,N_8654,N_8645);
nand U8748 (N_8748,N_8684,N_8672);
and U8749 (N_8749,N_8658,N_8699);
or U8750 (N_8750,N_8621,N_8681);
xnor U8751 (N_8751,N_8635,N_8667);
nand U8752 (N_8752,N_8676,N_8642);
or U8753 (N_8753,N_8662,N_8612);
xor U8754 (N_8754,N_8666,N_8651);
nand U8755 (N_8755,N_8615,N_8638);
nand U8756 (N_8756,N_8646,N_8663);
or U8757 (N_8757,N_8698,N_8652);
and U8758 (N_8758,N_8600,N_8691);
nor U8759 (N_8759,N_8635,N_8613);
nor U8760 (N_8760,N_8663,N_8679);
nand U8761 (N_8761,N_8659,N_8695);
or U8762 (N_8762,N_8673,N_8669);
or U8763 (N_8763,N_8664,N_8685);
nor U8764 (N_8764,N_8627,N_8606);
nor U8765 (N_8765,N_8686,N_8687);
and U8766 (N_8766,N_8674,N_8656);
and U8767 (N_8767,N_8637,N_8600);
nor U8768 (N_8768,N_8606,N_8682);
or U8769 (N_8769,N_8639,N_8643);
nand U8770 (N_8770,N_8631,N_8616);
nor U8771 (N_8771,N_8624,N_8638);
and U8772 (N_8772,N_8604,N_8667);
nand U8773 (N_8773,N_8686,N_8600);
nand U8774 (N_8774,N_8624,N_8660);
or U8775 (N_8775,N_8680,N_8615);
or U8776 (N_8776,N_8663,N_8616);
and U8777 (N_8777,N_8655,N_8697);
and U8778 (N_8778,N_8600,N_8661);
xor U8779 (N_8779,N_8699,N_8666);
nor U8780 (N_8780,N_8671,N_8647);
nor U8781 (N_8781,N_8625,N_8633);
nor U8782 (N_8782,N_8651,N_8636);
or U8783 (N_8783,N_8669,N_8640);
and U8784 (N_8784,N_8672,N_8600);
or U8785 (N_8785,N_8672,N_8682);
nand U8786 (N_8786,N_8650,N_8677);
xnor U8787 (N_8787,N_8696,N_8627);
nand U8788 (N_8788,N_8693,N_8624);
nand U8789 (N_8789,N_8655,N_8649);
nand U8790 (N_8790,N_8618,N_8657);
or U8791 (N_8791,N_8614,N_8629);
nor U8792 (N_8792,N_8648,N_8621);
and U8793 (N_8793,N_8648,N_8606);
nand U8794 (N_8794,N_8625,N_8675);
nor U8795 (N_8795,N_8676,N_8684);
xnor U8796 (N_8796,N_8640,N_8614);
nor U8797 (N_8797,N_8641,N_8624);
nand U8798 (N_8798,N_8675,N_8630);
nor U8799 (N_8799,N_8660,N_8623);
or U8800 (N_8800,N_8704,N_8705);
nand U8801 (N_8801,N_8724,N_8756);
or U8802 (N_8802,N_8733,N_8731);
and U8803 (N_8803,N_8711,N_8735);
and U8804 (N_8804,N_8761,N_8774);
nand U8805 (N_8805,N_8775,N_8776);
nor U8806 (N_8806,N_8741,N_8760);
or U8807 (N_8807,N_8751,N_8771);
and U8808 (N_8808,N_8764,N_8719);
nor U8809 (N_8809,N_8739,N_8700);
xnor U8810 (N_8810,N_8795,N_8754);
nand U8811 (N_8811,N_8755,N_8791);
nor U8812 (N_8812,N_8786,N_8792);
nor U8813 (N_8813,N_8777,N_8785);
nor U8814 (N_8814,N_8799,N_8757);
nor U8815 (N_8815,N_8714,N_8706);
nand U8816 (N_8816,N_8726,N_8709);
nand U8817 (N_8817,N_8727,N_8703);
nor U8818 (N_8818,N_8770,N_8758);
xnor U8819 (N_8819,N_8766,N_8748);
nor U8820 (N_8820,N_8710,N_8794);
or U8821 (N_8821,N_8718,N_8720);
or U8822 (N_8822,N_8716,N_8702);
nand U8823 (N_8823,N_8749,N_8715);
xnor U8824 (N_8824,N_8717,N_8784);
or U8825 (N_8825,N_8750,N_8778);
and U8826 (N_8826,N_8763,N_8781);
xor U8827 (N_8827,N_8740,N_8729);
or U8828 (N_8828,N_8722,N_8787);
or U8829 (N_8829,N_8789,N_8707);
xnor U8830 (N_8830,N_8747,N_8745);
nand U8831 (N_8831,N_8732,N_8768);
and U8832 (N_8832,N_8780,N_8738);
nor U8833 (N_8833,N_8742,N_8752);
nand U8834 (N_8834,N_8772,N_8753);
nor U8835 (N_8835,N_8798,N_8782);
nand U8836 (N_8836,N_8762,N_8765);
or U8837 (N_8837,N_8779,N_8797);
nor U8838 (N_8838,N_8723,N_8783);
nor U8839 (N_8839,N_8708,N_8728);
xor U8840 (N_8840,N_8713,N_8769);
nand U8841 (N_8841,N_8790,N_8793);
nand U8842 (N_8842,N_8744,N_8736);
xor U8843 (N_8843,N_8773,N_8746);
nand U8844 (N_8844,N_8796,N_8734);
nand U8845 (N_8845,N_8725,N_8767);
and U8846 (N_8846,N_8730,N_8701);
or U8847 (N_8847,N_8737,N_8788);
or U8848 (N_8848,N_8712,N_8721);
and U8849 (N_8849,N_8759,N_8743);
nor U8850 (N_8850,N_8789,N_8744);
xnor U8851 (N_8851,N_8737,N_8756);
nor U8852 (N_8852,N_8700,N_8702);
and U8853 (N_8853,N_8716,N_8755);
nor U8854 (N_8854,N_8724,N_8765);
or U8855 (N_8855,N_8751,N_8777);
nand U8856 (N_8856,N_8709,N_8797);
nand U8857 (N_8857,N_8789,N_8716);
nand U8858 (N_8858,N_8719,N_8706);
and U8859 (N_8859,N_8767,N_8789);
nand U8860 (N_8860,N_8775,N_8788);
or U8861 (N_8861,N_8740,N_8755);
and U8862 (N_8862,N_8791,N_8701);
nor U8863 (N_8863,N_8785,N_8743);
or U8864 (N_8864,N_8790,N_8750);
xor U8865 (N_8865,N_8763,N_8720);
nand U8866 (N_8866,N_8727,N_8766);
nor U8867 (N_8867,N_8748,N_8712);
and U8868 (N_8868,N_8753,N_8707);
or U8869 (N_8869,N_8755,N_8748);
xnor U8870 (N_8870,N_8715,N_8781);
or U8871 (N_8871,N_8723,N_8754);
or U8872 (N_8872,N_8764,N_8758);
nor U8873 (N_8873,N_8782,N_8724);
nor U8874 (N_8874,N_8753,N_8754);
nor U8875 (N_8875,N_8713,N_8755);
and U8876 (N_8876,N_8709,N_8737);
nand U8877 (N_8877,N_8721,N_8702);
or U8878 (N_8878,N_8755,N_8753);
and U8879 (N_8879,N_8797,N_8756);
nand U8880 (N_8880,N_8733,N_8718);
and U8881 (N_8881,N_8705,N_8700);
nor U8882 (N_8882,N_8726,N_8798);
nand U8883 (N_8883,N_8703,N_8766);
or U8884 (N_8884,N_8743,N_8788);
nand U8885 (N_8885,N_8742,N_8780);
nand U8886 (N_8886,N_8775,N_8760);
xor U8887 (N_8887,N_8756,N_8766);
and U8888 (N_8888,N_8751,N_8708);
nand U8889 (N_8889,N_8730,N_8752);
nand U8890 (N_8890,N_8717,N_8747);
nor U8891 (N_8891,N_8743,N_8711);
nand U8892 (N_8892,N_8793,N_8732);
xnor U8893 (N_8893,N_8749,N_8779);
or U8894 (N_8894,N_8721,N_8730);
and U8895 (N_8895,N_8785,N_8706);
or U8896 (N_8896,N_8724,N_8774);
and U8897 (N_8897,N_8752,N_8775);
nand U8898 (N_8898,N_8782,N_8774);
or U8899 (N_8899,N_8729,N_8753);
and U8900 (N_8900,N_8871,N_8885);
nor U8901 (N_8901,N_8806,N_8842);
nor U8902 (N_8902,N_8831,N_8835);
nand U8903 (N_8903,N_8839,N_8808);
or U8904 (N_8904,N_8815,N_8888);
nor U8905 (N_8905,N_8850,N_8862);
nor U8906 (N_8906,N_8893,N_8848);
or U8907 (N_8907,N_8890,N_8813);
xnor U8908 (N_8908,N_8856,N_8870);
and U8909 (N_8909,N_8823,N_8843);
and U8910 (N_8910,N_8891,N_8887);
and U8911 (N_8911,N_8899,N_8880);
nand U8912 (N_8912,N_8837,N_8804);
xor U8913 (N_8913,N_8827,N_8829);
nor U8914 (N_8914,N_8853,N_8859);
nand U8915 (N_8915,N_8828,N_8894);
nor U8916 (N_8916,N_8864,N_8852);
or U8917 (N_8917,N_8802,N_8879);
or U8918 (N_8918,N_8834,N_8874);
xor U8919 (N_8919,N_8872,N_8858);
or U8920 (N_8920,N_8857,N_8810);
nor U8921 (N_8921,N_8861,N_8803);
or U8922 (N_8922,N_8836,N_8824);
or U8923 (N_8923,N_8840,N_8849);
nor U8924 (N_8924,N_8881,N_8897);
nor U8925 (N_8925,N_8801,N_8882);
or U8926 (N_8926,N_8886,N_8876);
or U8927 (N_8927,N_8868,N_8832);
nand U8928 (N_8928,N_8817,N_8812);
nand U8929 (N_8929,N_8809,N_8807);
nor U8930 (N_8930,N_8811,N_8826);
nor U8931 (N_8931,N_8825,N_8866);
nand U8932 (N_8932,N_8883,N_8821);
nand U8933 (N_8933,N_8898,N_8896);
and U8934 (N_8934,N_8865,N_8884);
nand U8935 (N_8935,N_8863,N_8854);
or U8936 (N_8936,N_8873,N_8895);
nor U8937 (N_8937,N_8818,N_8867);
nor U8938 (N_8938,N_8855,N_8819);
and U8939 (N_8939,N_8800,N_8841);
and U8940 (N_8940,N_8845,N_8830);
or U8941 (N_8941,N_8851,N_8878);
nor U8942 (N_8942,N_8822,N_8889);
and U8943 (N_8943,N_8860,N_8869);
nor U8944 (N_8944,N_8838,N_8892);
and U8945 (N_8945,N_8816,N_8846);
nand U8946 (N_8946,N_8847,N_8814);
or U8947 (N_8947,N_8820,N_8875);
nand U8948 (N_8948,N_8844,N_8877);
nand U8949 (N_8949,N_8833,N_8805);
nand U8950 (N_8950,N_8809,N_8834);
xor U8951 (N_8951,N_8810,N_8849);
nand U8952 (N_8952,N_8879,N_8860);
nand U8953 (N_8953,N_8840,N_8830);
nor U8954 (N_8954,N_8820,N_8805);
or U8955 (N_8955,N_8821,N_8834);
nand U8956 (N_8956,N_8856,N_8868);
and U8957 (N_8957,N_8848,N_8842);
nand U8958 (N_8958,N_8878,N_8837);
and U8959 (N_8959,N_8832,N_8835);
nor U8960 (N_8960,N_8852,N_8832);
nand U8961 (N_8961,N_8836,N_8896);
nand U8962 (N_8962,N_8866,N_8839);
or U8963 (N_8963,N_8840,N_8815);
or U8964 (N_8964,N_8853,N_8833);
or U8965 (N_8965,N_8873,N_8876);
nand U8966 (N_8966,N_8861,N_8872);
nor U8967 (N_8967,N_8802,N_8885);
and U8968 (N_8968,N_8883,N_8826);
nor U8969 (N_8969,N_8809,N_8805);
nor U8970 (N_8970,N_8806,N_8824);
nand U8971 (N_8971,N_8838,N_8846);
nor U8972 (N_8972,N_8898,N_8845);
nor U8973 (N_8973,N_8858,N_8856);
and U8974 (N_8974,N_8849,N_8808);
or U8975 (N_8975,N_8868,N_8848);
nor U8976 (N_8976,N_8883,N_8879);
and U8977 (N_8977,N_8878,N_8811);
nand U8978 (N_8978,N_8856,N_8807);
or U8979 (N_8979,N_8822,N_8806);
or U8980 (N_8980,N_8851,N_8887);
and U8981 (N_8981,N_8801,N_8800);
or U8982 (N_8982,N_8898,N_8804);
nand U8983 (N_8983,N_8852,N_8834);
or U8984 (N_8984,N_8898,N_8853);
nand U8985 (N_8985,N_8810,N_8862);
nor U8986 (N_8986,N_8818,N_8804);
nand U8987 (N_8987,N_8866,N_8831);
xor U8988 (N_8988,N_8865,N_8818);
and U8989 (N_8989,N_8874,N_8809);
or U8990 (N_8990,N_8833,N_8804);
nand U8991 (N_8991,N_8808,N_8840);
or U8992 (N_8992,N_8856,N_8837);
nand U8993 (N_8993,N_8804,N_8897);
nor U8994 (N_8994,N_8885,N_8814);
nand U8995 (N_8995,N_8808,N_8812);
nor U8996 (N_8996,N_8899,N_8810);
xnor U8997 (N_8997,N_8870,N_8889);
xnor U8998 (N_8998,N_8858,N_8881);
nand U8999 (N_8999,N_8813,N_8836);
or U9000 (N_9000,N_8995,N_8937);
and U9001 (N_9001,N_8967,N_8948);
and U9002 (N_9002,N_8946,N_8984);
nor U9003 (N_9003,N_8936,N_8963);
nor U9004 (N_9004,N_8979,N_8959);
nor U9005 (N_9005,N_8933,N_8998);
xnor U9006 (N_9006,N_8908,N_8918);
nor U9007 (N_9007,N_8966,N_8921);
xnor U9008 (N_9008,N_8954,N_8925);
xor U9009 (N_9009,N_8935,N_8983);
and U9010 (N_9010,N_8997,N_8960);
xnor U9011 (N_9011,N_8944,N_8957);
nand U9012 (N_9012,N_8977,N_8938);
nand U9013 (N_9013,N_8927,N_8996);
and U9014 (N_9014,N_8905,N_8934);
and U9015 (N_9015,N_8914,N_8973);
and U9016 (N_9016,N_8987,N_8949);
and U9017 (N_9017,N_8974,N_8950);
nand U9018 (N_9018,N_8971,N_8906);
or U9019 (N_9019,N_8951,N_8992);
nor U9020 (N_9020,N_8917,N_8912);
nand U9021 (N_9021,N_8962,N_8991);
or U9022 (N_9022,N_8956,N_8961);
nor U9023 (N_9023,N_8982,N_8980);
and U9024 (N_9024,N_8952,N_8939);
nand U9025 (N_9025,N_8907,N_8940);
nor U9026 (N_9026,N_8994,N_8981);
nor U9027 (N_9027,N_8989,N_8976);
xnor U9028 (N_9028,N_8986,N_8926);
and U9029 (N_9029,N_8932,N_8985);
nand U9030 (N_9030,N_8910,N_8958);
and U9031 (N_9031,N_8928,N_8941);
xor U9032 (N_9032,N_8902,N_8901);
or U9033 (N_9033,N_8943,N_8913);
nor U9034 (N_9034,N_8955,N_8978);
and U9035 (N_9035,N_8975,N_8923);
xnor U9036 (N_9036,N_8964,N_8942);
nand U9037 (N_9037,N_8900,N_8969);
and U9038 (N_9038,N_8965,N_8911);
nor U9039 (N_9039,N_8990,N_8903);
nor U9040 (N_9040,N_8945,N_8947);
nand U9041 (N_9041,N_8920,N_8924);
or U9042 (N_9042,N_8909,N_8919);
xor U9043 (N_9043,N_8929,N_8968);
and U9044 (N_9044,N_8930,N_8922);
nand U9045 (N_9045,N_8988,N_8993);
or U9046 (N_9046,N_8915,N_8916);
nand U9047 (N_9047,N_8972,N_8970);
and U9048 (N_9048,N_8953,N_8904);
nand U9049 (N_9049,N_8931,N_8999);
or U9050 (N_9050,N_8968,N_8983);
nor U9051 (N_9051,N_8903,N_8979);
nor U9052 (N_9052,N_8930,N_8929);
nor U9053 (N_9053,N_8983,N_8921);
xor U9054 (N_9054,N_8984,N_8956);
nand U9055 (N_9055,N_8968,N_8962);
nand U9056 (N_9056,N_8998,N_8926);
nand U9057 (N_9057,N_8953,N_8960);
nand U9058 (N_9058,N_8943,N_8940);
nand U9059 (N_9059,N_8972,N_8953);
and U9060 (N_9060,N_8904,N_8965);
xnor U9061 (N_9061,N_8955,N_8993);
nor U9062 (N_9062,N_8918,N_8936);
nand U9063 (N_9063,N_8971,N_8946);
and U9064 (N_9064,N_8902,N_8967);
nor U9065 (N_9065,N_8980,N_8998);
and U9066 (N_9066,N_8905,N_8958);
nand U9067 (N_9067,N_8993,N_8963);
or U9068 (N_9068,N_8992,N_8910);
xnor U9069 (N_9069,N_8941,N_8934);
nor U9070 (N_9070,N_8909,N_8956);
nor U9071 (N_9071,N_8936,N_8969);
nand U9072 (N_9072,N_8997,N_8921);
xnor U9073 (N_9073,N_8964,N_8928);
and U9074 (N_9074,N_8900,N_8918);
or U9075 (N_9075,N_8979,N_8920);
nand U9076 (N_9076,N_8944,N_8928);
nand U9077 (N_9077,N_8981,N_8917);
or U9078 (N_9078,N_8981,N_8991);
nand U9079 (N_9079,N_8979,N_8992);
or U9080 (N_9080,N_8979,N_8942);
or U9081 (N_9081,N_8983,N_8906);
and U9082 (N_9082,N_8986,N_8923);
nand U9083 (N_9083,N_8950,N_8933);
nor U9084 (N_9084,N_8902,N_8949);
and U9085 (N_9085,N_8935,N_8926);
or U9086 (N_9086,N_8972,N_8967);
nor U9087 (N_9087,N_8916,N_8928);
nand U9088 (N_9088,N_8975,N_8945);
nor U9089 (N_9089,N_8989,N_8908);
and U9090 (N_9090,N_8980,N_8984);
nor U9091 (N_9091,N_8981,N_8951);
or U9092 (N_9092,N_8989,N_8913);
or U9093 (N_9093,N_8981,N_8919);
nand U9094 (N_9094,N_8916,N_8981);
and U9095 (N_9095,N_8928,N_8930);
and U9096 (N_9096,N_8922,N_8942);
or U9097 (N_9097,N_8903,N_8959);
and U9098 (N_9098,N_8955,N_8943);
nor U9099 (N_9099,N_8947,N_8941);
nor U9100 (N_9100,N_9019,N_9001);
nor U9101 (N_9101,N_9004,N_9005);
nor U9102 (N_9102,N_9016,N_9050);
nor U9103 (N_9103,N_9012,N_9045);
nor U9104 (N_9104,N_9011,N_9015);
nor U9105 (N_9105,N_9067,N_9039);
nand U9106 (N_9106,N_9053,N_9082);
and U9107 (N_9107,N_9020,N_9021);
or U9108 (N_9108,N_9090,N_9041);
and U9109 (N_9109,N_9033,N_9089);
nand U9110 (N_9110,N_9065,N_9032);
and U9111 (N_9111,N_9042,N_9069);
xnor U9112 (N_9112,N_9068,N_9071);
and U9113 (N_9113,N_9025,N_9029);
or U9114 (N_9114,N_9098,N_9034);
nor U9115 (N_9115,N_9056,N_9066);
or U9116 (N_9116,N_9072,N_9076);
and U9117 (N_9117,N_9008,N_9002);
nand U9118 (N_9118,N_9023,N_9092);
nor U9119 (N_9119,N_9070,N_9075);
nand U9120 (N_9120,N_9073,N_9055);
xor U9121 (N_9121,N_9049,N_9086);
nand U9122 (N_9122,N_9094,N_9063);
nor U9123 (N_9123,N_9026,N_9051);
nand U9124 (N_9124,N_9085,N_9038);
and U9125 (N_9125,N_9091,N_9077);
nand U9126 (N_9126,N_9013,N_9095);
or U9127 (N_9127,N_9080,N_9027);
and U9128 (N_9128,N_9030,N_9059);
and U9129 (N_9129,N_9018,N_9031);
or U9130 (N_9130,N_9014,N_9093);
and U9131 (N_9131,N_9064,N_9052);
and U9132 (N_9132,N_9079,N_9007);
nand U9133 (N_9133,N_9010,N_9044);
nor U9134 (N_9134,N_9060,N_9047);
nand U9135 (N_9135,N_9083,N_9048);
and U9136 (N_9136,N_9061,N_9078);
xor U9137 (N_9137,N_9054,N_9024);
and U9138 (N_9138,N_9000,N_9040);
or U9139 (N_9139,N_9099,N_9036);
nor U9140 (N_9140,N_9022,N_9097);
nor U9141 (N_9141,N_9046,N_9003);
xnor U9142 (N_9142,N_9057,N_9074);
and U9143 (N_9143,N_9009,N_9084);
and U9144 (N_9144,N_9096,N_9017);
and U9145 (N_9145,N_9006,N_9062);
xor U9146 (N_9146,N_9087,N_9081);
nor U9147 (N_9147,N_9028,N_9088);
and U9148 (N_9148,N_9043,N_9058);
nand U9149 (N_9149,N_9037,N_9035);
or U9150 (N_9150,N_9078,N_9003);
xor U9151 (N_9151,N_9043,N_9067);
nor U9152 (N_9152,N_9023,N_9052);
and U9153 (N_9153,N_9025,N_9081);
nand U9154 (N_9154,N_9062,N_9057);
nor U9155 (N_9155,N_9051,N_9071);
nand U9156 (N_9156,N_9031,N_9006);
or U9157 (N_9157,N_9017,N_9039);
xor U9158 (N_9158,N_9091,N_9002);
and U9159 (N_9159,N_9048,N_9098);
xor U9160 (N_9160,N_9029,N_9088);
nor U9161 (N_9161,N_9031,N_9016);
nand U9162 (N_9162,N_9098,N_9076);
nand U9163 (N_9163,N_9069,N_9044);
and U9164 (N_9164,N_9001,N_9081);
or U9165 (N_9165,N_9020,N_9056);
nand U9166 (N_9166,N_9006,N_9073);
or U9167 (N_9167,N_9083,N_9024);
nand U9168 (N_9168,N_9032,N_9011);
and U9169 (N_9169,N_9046,N_9092);
nand U9170 (N_9170,N_9001,N_9045);
and U9171 (N_9171,N_9087,N_9049);
and U9172 (N_9172,N_9063,N_9046);
or U9173 (N_9173,N_9007,N_9049);
or U9174 (N_9174,N_9063,N_9080);
nor U9175 (N_9175,N_9096,N_9058);
nor U9176 (N_9176,N_9002,N_9079);
xnor U9177 (N_9177,N_9034,N_9006);
nand U9178 (N_9178,N_9051,N_9079);
nor U9179 (N_9179,N_9063,N_9022);
nor U9180 (N_9180,N_9020,N_9035);
nor U9181 (N_9181,N_9009,N_9049);
nand U9182 (N_9182,N_9048,N_9023);
and U9183 (N_9183,N_9036,N_9006);
nand U9184 (N_9184,N_9083,N_9093);
or U9185 (N_9185,N_9039,N_9097);
nand U9186 (N_9186,N_9062,N_9075);
nor U9187 (N_9187,N_9048,N_9032);
xor U9188 (N_9188,N_9008,N_9080);
nand U9189 (N_9189,N_9026,N_9065);
nor U9190 (N_9190,N_9077,N_9084);
nor U9191 (N_9191,N_9000,N_9072);
nand U9192 (N_9192,N_9059,N_9070);
nand U9193 (N_9193,N_9032,N_9004);
or U9194 (N_9194,N_9056,N_9082);
and U9195 (N_9195,N_9062,N_9083);
or U9196 (N_9196,N_9082,N_9062);
and U9197 (N_9197,N_9099,N_9021);
or U9198 (N_9198,N_9039,N_9035);
nor U9199 (N_9199,N_9079,N_9052);
nand U9200 (N_9200,N_9186,N_9182);
and U9201 (N_9201,N_9129,N_9165);
and U9202 (N_9202,N_9114,N_9116);
nor U9203 (N_9203,N_9195,N_9101);
nor U9204 (N_9204,N_9173,N_9183);
and U9205 (N_9205,N_9139,N_9127);
or U9206 (N_9206,N_9174,N_9196);
nor U9207 (N_9207,N_9110,N_9179);
and U9208 (N_9208,N_9131,N_9170);
nand U9209 (N_9209,N_9176,N_9118);
xnor U9210 (N_9210,N_9146,N_9148);
and U9211 (N_9211,N_9159,N_9137);
or U9212 (N_9212,N_9119,N_9162);
or U9213 (N_9213,N_9198,N_9171);
or U9214 (N_9214,N_9193,N_9152);
and U9215 (N_9215,N_9142,N_9163);
nor U9216 (N_9216,N_9167,N_9168);
nand U9217 (N_9217,N_9124,N_9197);
nor U9218 (N_9218,N_9185,N_9134);
and U9219 (N_9219,N_9180,N_9192);
nand U9220 (N_9220,N_9156,N_9194);
nor U9221 (N_9221,N_9128,N_9100);
nor U9222 (N_9222,N_9135,N_9199);
nor U9223 (N_9223,N_9138,N_9191);
xor U9224 (N_9224,N_9147,N_9141);
xnor U9225 (N_9225,N_9158,N_9155);
nor U9226 (N_9226,N_9166,N_9175);
or U9227 (N_9227,N_9161,N_9190);
nand U9228 (N_9228,N_9123,N_9130);
nor U9229 (N_9229,N_9177,N_9187);
and U9230 (N_9230,N_9122,N_9136);
nand U9231 (N_9231,N_9104,N_9149);
nor U9232 (N_9232,N_9111,N_9132);
or U9233 (N_9233,N_9188,N_9184);
xnor U9234 (N_9234,N_9153,N_9150);
nor U9235 (N_9235,N_9108,N_9144);
nand U9236 (N_9236,N_9154,N_9151);
nor U9237 (N_9237,N_9113,N_9157);
and U9238 (N_9238,N_9125,N_9160);
or U9239 (N_9239,N_9105,N_9103);
nand U9240 (N_9240,N_9189,N_9164);
nand U9241 (N_9241,N_9145,N_9133);
or U9242 (N_9242,N_9126,N_9169);
nand U9243 (N_9243,N_9109,N_9115);
and U9244 (N_9244,N_9107,N_9143);
and U9245 (N_9245,N_9178,N_9172);
or U9246 (N_9246,N_9117,N_9120);
nand U9247 (N_9247,N_9112,N_9181);
or U9248 (N_9248,N_9106,N_9121);
or U9249 (N_9249,N_9140,N_9102);
and U9250 (N_9250,N_9138,N_9156);
nand U9251 (N_9251,N_9101,N_9170);
xnor U9252 (N_9252,N_9118,N_9143);
or U9253 (N_9253,N_9153,N_9110);
and U9254 (N_9254,N_9118,N_9174);
nand U9255 (N_9255,N_9173,N_9116);
or U9256 (N_9256,N_9158,N_9107);
xnor U9257 (N_9257,N_9149,N_9166);
nand U9258 (N_9258,N_9133,N_9157);
nor U9259 (N_9259,N_9161,N_9137);
nand U9260 (N_9260,N_9104,N_9159);
xor U9261 (N_9261,N_9144,N_9110);
or U9262 (N_9262,N_9148,N_9177);
nand U9263 (N_9263,N_9113,N_9170);
nor U9264 (N_9264,N_9141,N_9112);
xnor U9265 (N_9265,N_9126,N_9124);
nand U9266 (N_9266,N_9158,N_9150);
nand U9267 (N_9267,N_9150,N_9115);
or U9268 (N_9268,N_9148,N_9124);
nand U9269 (N_9269,N_9156,N_9199);
and U9270 (N_9270,N_9129,N_9166);
and U9271 (N_9271,N_9161,N_9186);
and U9272 (N_9272,N_9174,N_9168);
nor U9273 (N_9273,N_9151,N_9184);
or U9274 (N_9274,N_9109,N_9117);
and U9275 (N_9275,N_9198,N_9168);
nand U9276 (N_9276,N_9183,N_9102);
nor U9277 (N_9277,N_9137,N_9186);
nand U9278 (N_9278,N_9141,N_9152);
nand U9279 (N_9279,N_9106,N_9136);
nand U9280 (N_9280,N_9127,N_9133);
xor U9281 (N_9281,N_9199,N_9195);
and U9282 (N_9282,N_9114,N_9141);
or U9283 (N_9283,N_9195,N_9128);
xnor U9284 (N_9284,N_9196,N_9187);
xor U9285 (N_9285,N_9133,N_9198);
or U9286 (N_9286,N_9161,N_9127);
or U9287 (N_9287,N_9197,N_9132);
and U9288 (N_9288,N_9133,N_9121);
nor U9289 (N_9289,N_9149,N_9183);
nor U9290 (N_9290,N_9195,N_9187);
nand U9291 (N_9291,N_9184,N_9172);
or U9292 (N_9292,N_9126,N_9188);
nand U9293 (N_9293,N_9163,N_9106);
nand U9294 (N_9294,N_9159,N_9128);
or U9295 (N_9295,N_9178,N_9179);
nor U9296 (N_9296,N_9175,N_9155);
and U9297 (N_9297,N_9125,N_9197);
or U9298 (N_9298,N_9184,N_9135);
and U9299 (N_9299,N_9160,N_9106);
or U9300 (N_9300,N_9270,N_9205);
and U9301 (N_9301,N_9289,N_9213);
or U9302 (N_9302,N_9257,N_9259);
nand U9303 (N_9303,N_9214,N_9255);
or U9304 (N_9304,N_9287,N_9238);
or U9305 (N_9305,N_9277,N_9272);
xor U9306 (N_9306,N_9285,N_9219);
nand U9307 (N_9307,N_9252,N_9281);
nand U9308 (N_9308,N_9210,N_9286);
nor U9309 (N_9309,N_9245,N_9282);
or U9310 (N_9310,N_9273,N_9283);
and U9311 (N_9311,N_9296,N_9254);
nand U9312 (N_9312,N_9200,N_9222);
nor U9313 (N_9313,N_9269,N_9231);
nand U9314 (N_9314,N_9223,N_9256);
and U9315 (N_9315,N_9244,N_9203);
xnor U9316 (N_9316,N_9229,N_9266);
and U9317 (N_9317,N_9261,N_9260);
nand U9318 (N_9318,N_9209,N_9239);
nand U9319 (N_9319,N_9251,N_9233);
nand U9320 (N_9320,N_9204,N_9284);
nand U9321 (N_9321,N_9232,N_9237);
nor U9322 (N_9322,N_9242,N_9211);
nor U9323 (N_9323,N_9274,N_9243);
or U9324 (N_9324,N_9208,N_9299);
and U9325 (N_9325,N_9276,N_9297);
nor U9326 (N_9326,N_9224,N_9298);
and U9327 (N_9327,N_9241,N_9258);
xor U9328 (N_9328,N_9250,N_9268);
nand U9329 (N_9329,N_9288,N_9236);
and U9330 (N_9330,N_9212,N_9294);
or U9331 (N_9331,N_9240,N_9265);
nand U9332 (N_9332,N_9206,N_9218);
nand U9333 (N_9333,N_9225,N_9278);
nand U9334 (N_9334,N_9291,N_9247);
or U9335 (N_9335,N_9249,N_9263);
xnor U9336 (N_9336,N_9275,N_9267);
and U9337 (N_9337,N_9216,N_9279);
or U9338 (N_9338,N_9226,N_9264);
nand U9339 (N_9339,N_9271,N_9248);
nor U9340 (N_9340,N_9290,N_9207);
or U9341 (N_9341,N_9201,N_9221);
nor U9342 (N_9342,N_9293,N_9262);
nand U9343 (N_9343,N_9215,N_9228);
nor U9344 (N_9344,N_9295,N_9227);
nor U9345 (N_9345,N_9253,N_9292);
xnor U9346 (N_9346,N_9217,N_9202);
nor U9347 (N_9347,N_9234,N_9235);
nand U9348 (N_9348,N_9280,N_9246);
and U9349 (N_9349,N_9220,N_9230);
nor U9350 (N_9350,N_9250,N_9291);
nor U9351 (N_9351,N_9264,N_9282);
nor U9352 (N_9352,N_9230,N_9225);
and U9353 (N_9353,N_9266,N_9264);
nor U9354 (N_9354,N_9292,N_9210);
xor U9355 (N_9355,N_9226,N_9258);
and U9356 (N_9356,N_9295,N_9266);
nor U9357 (N_9357,N_9280,N_9255);
nand U9358 (N_9358,N_9275,N_9271);
nand U9359 (N_9359,N_9222,N_9234);
and U9360 (N_9360,N_9266,N_9227);
nand U9361 (N_9361,N_9238,N_9246);
nand U9362 (N_9362,N_9275,N_9245);
nor U9363 (N_9363,N_9238,N_9237);
and U9364 (N_9364,N_9280,N_9271);
nor U9365 (N_9365,N_9245,N_9208);
or U9366 (N_9366,N_9248,N_9279);
and U9367 (N_9367,N_9234,N_9284);
or U9368 (N_9368,N_9267,N_9278);
nor U9369 (N_9369,N_9262,N_9288);
nand U9370 (N_9370,N_9272,N_9290);
or U9371 (N_9371,N_9263,N_9271);
and U9372 (N_9372,N_9254,N_9219);
nand U9373 (N_9373,N_9228,N_9268);
or U9374 (N_9374,N_9256,N_9277);
and U9375 (N_9375,N_9256,N_9215);
or U9376 (N_9376,N_9213,N_9211);
or U9377 (N_9377,N_9232,N_9279);
xnor U9378 (N_9378,N_9231,N_9236);
xor U9379 (N_9379,N_9208,N_9225);
or U9380 (N_9380,N_9232,N_9274);
and U9381 (N_9381,N_9287,N_9262);
nor U9382 (N_9382,N_9238,N_9274);
nand U9383 (N_9383,N_9260,N_9238);
nor U9384 (N_9384,N_9210,N_9271);
nor U9385 (N_9385,N_9236,N_9208);
and U9386 (N_9386,N_9263,N_9238);
xor U9387 (N_9387,N_9224,N_9267);
and U9388 (N_9388,N_9260,N_9257);
and U9389 (N_9389,N_9232,N_9293);
nor U9390 (N_9390,N_9247,N_9211);
nand U9391 (N_9391,N_9212,N_9269);
or U9392 (N_9392,N_9275,N_9295);
and U9393 (N_9393,N_9257,N_9234);
nand U9394 (N_9394,N_9262,N_9211);
or U9395 (N_9395,N_9290,N_9291);
or U9396 (N_9396,N_9247,N_9217);
xor U9397 (N_9397,N_9251,N_9264);
nand U9398 (N_9398,N_9225,N_9200);
nor U9399 (N_9399,N_9205,N_9235);
and U9400 (N_9400,N_9331,N_9333);
nor U9401 (N_9401,N_9316,N_9320);
xor U9402 (N_9402,N_9392,N_9358);
nand U9403 (N_9403,N_9344,N_9343);
nand U9404 (N_9404,N_9351,N_9317);
nand U9405 (N_9405,N_9349,N_9309);
nand U9406 (N_9406,N_9345,N_9366);
nor U9407 (N_9407,N_9312,N_9368);
nand U9408 (N_9408,N_9360,N_9336);
and U9409 (N_9409,N_9319,N_9308);
nand U9410 (N_9410,N_9363,N_9340);
nor U9411 (N_9411,N_9322,N_9387);
nor U9412 (N_9412,N_9323,N_9304);
and U9413 (N_9413,N_9381,N_9357);
xor U9414 (N_9414,N_9395,N_9325);
and U9415 (N_9415,N_9394,N_9382);
nand U9416 (N_9416,N_9384,N_9307);
xor U9417 (N_9417,N_9399,N_9342);
nor U9418 (N_9418,N_9378,N_9377);
xnor U9419 (N_9419,N_9372,N_9332);
nor U9420 (N_9420,N_9356,N_9367);
nor U9421 (N_9421,N_9396,N_9301);
xnor U9422 (N_9422,N_9305,N_9389);
nor U9423 (N_9423,N_9339,N_9365);
or U9424 (N_9424,N_9306,N_9390);
and U9425 (N_9425,N_9329,N_9373);
nand U9426 (N_9426,N_9354,N_9353);
nor U9427 (N_9427,N_9327,N_9310);
and U9428 (N_9428,N_9311,N_9386);
nor U9429 (N_9429,N_9313,N_9303);
xnor U9430 (N_9430,N_9338,N_9350);
nand U9431 (N_9431,N_9324,N_9346);
or U9432 (N_9432,N_9374,N_9328);
or U9433 (N_9433,N_9337,N_9383);
and U9434 (N_9434,N_9398,N_9326);
nor U9435 (N_9435,N_9361,N_9380);
or U9436 (N_9436,N_9391,N_9359);
nand U9437 (N_9437,N_9379,N_9388);
and U9438 (N_9438,N_9334,N_9371);
and U9439 (N_9439,N_9369,N_9321);
or U9440 (N_9440,N_9330,N_9352);
and U9441 (N_9441,N_9315,N_9300);
nand U9442 (N_9442,N_9355,N_9376);
nor U9443 (N_9443,N_9341,N_9347);
nand U9444 (N_9444,N_9348,N_9364);
nor U9445 (N_9445,N_9393,N_9318);
nand U9446 (N_9446,N_9385,N_9375);
xnor U9447 (N_9447,N_9397,N_9314);
or U9448 (N_9448,N_9335,N_9302);
nand U9449 (N_9449,N_9370,N_9362);
and U9450 (N_9450,N_9388,N_9323);
and U9451 (N_9451,N_9377,N_9383);
or U9452 (N_9452,N_9303,N_9363);
or U9453 (N_9453,N_9377,N_9321);
or U9454 (N_9454,N_9310,N_9336);
and U9455 (N_9455,N_9385,N_9344);
and U9456 (N_9456,N_9338,N_9347);
nor U9457 (N_9457,N_9322,N_9365);
nand U9458 (N_9458,N_9398,N_9323);
nand U9459 (N_9459,N_9378,N_9367);
xnor U9460 (N_9460,N_9310,N_9315);
nor U9461 (N_9461,N_9317,N_9326);
and U9462 (N_9462,N_9322,N_9393);
and U9463 (N_9463,N_9309,N_9346);
or U9464 (N_9464,N_9352,N_9300);
or U9465 (N_9465,N_9338,N_9323);
nand U9466 (N_9466,N_9317,N_9361);
and U9467 (N_9467,N_9388,N_9304);
xor U9468 (N_9468,N_9308,N_9348);
xor U9469 (N_9469,N_9316,N_9345);
or U9470 (N_9470,N_9353,N_9356);
and U9471 (N_9471,N_9385,N_9347);
and U9472 (N_9472,N_9353,N_9302);
nand U9473 (N_9473,N_9310,N_9306);
and U9474 (N_9474,N_9390,N_9326);
or U9475 (N_9475,N_9310,N_9329);
and U9476 (N_9476,N_9315,N_9305);
nand U9477 (N_9477,N_9366,N_9349);
and U9478 (N_9478,N_9344,N_9395);
and U9479 (N_9479,N_9328,N_9373);
or U9480 (N_9480,N_9389,N_9386);
or U9481 (N_9481,N_9388,N_9301);
and U9482 (N_9482,N_9301,N_9311);
or U9483 (N_9483,N_9352,N_9336);
or U9484 (N_9484,N_9325,N_9381);
nand U9485 (N_9485,N_9367,N_9336);
or U9486 (N_9486,N_9320,N_9334);
nor U9487 (N_9487,N_9391,N_9373);
nand U9488 (N_9488,N_9378,N_9334);
and U9489 (N_9489,N_9331,N_9356);
nand U9490 (N_9490,N_9344,N_9366);
or U9491 (N_9491,N_9356,N_9377);
xnor U9492 (N_9492,N_9370,N_9318);
nor U9493 (N_9493,N_9340,N_9317);
nand U9494 (N_9494,N_9346,N_9322);
nor U9495 (N_9495,N_9346,N_9380);
nor U9496 (N_9496,N_9381,N_9327);
nor U9497 (N_9497,N_9357,N_9354);
and U9498 (N_9498,N_9344,N_9373);
nand U9499 (N_9499,N_9322,N_9308);
or U9500 (N_9500,N_9491,N_9430);
and U9501 (N_9501,N_9400,N_9499);
nor U9502 (N_9502,N_9484,N_9427);
or U9503 (N_9503,N_9417,N_9439);
and U9504 (N_9504,N_9404,N_9468);
nor U9505 (N_9505,N_9460,N_9421);
nor U9506 (N_9506,N_9432,N_9428);
nor U9507 (N_9507,N_9426,N_9408);
nand U9508 (N_9508,N_9459,N_9476);
nand U9509 (N_9509,N_9475,N_9447);
and U9510 (N_9510,N_9470,N_9441);
nand U9511 (N_9511,N_9465,N_9446);
nor U9512 (N_9512,N_9495,N_9486);
nor U9513 (N_9513,N_9483,N_9497);
nand U9514 (N_9514,N_9452,N_9418);
nand U9515 (N_9515,N_9451,N_9487);
and U9516 (N_9516,N_9401,N_9478);
or U9517 (N_9517,N_9431,N_9489);
nor U9518 (N_9518,N_9458,N_9409);
or U9519 (N_9519,N_9469,N_9467);
and U9520 (N_9520,N_9498,N_9482);
nand U9521 (N_9521,N_9454,N_9410);
nand U9522 (N_9522,N_9425,N_9402);
nand U9523 (N_9523,N_9413,N_9436);
or U9524 (N_9524,N_9435,N_9445);
or U9525 (N_9525,N_9456,N_9429);
or U9526 (N_9526,N_9477,N_9472);
nor U9527 (N_9527,N_9416,N_9464);
nand U9528 (N_9528,N_9405,N_9423);
or U9529 (N_9529,N_9480,N_9412);
nor U9530 (N_9530,N_9474,N_9466);
nor U9531 (N_9531,N_9449,N_9453);
and U9532 (N_9532,N_9450,N_9485);
or U9533 (N_9533,N_9481,N_9492);
or U9534 (N_9534,N_9411,N_9406);
nor U9535 (N_9535,N_9494,N_9471);
and U9536 (N_9536,N_9479,N_9414);
nand U9537 (N_9537,N_9440,N_9493);
and U9538 (N_9538,N_9461,N_9437);
nand U9539 (N_9539,N_9443,N_9420);
nor U9540 (N_9540,N_9434,N_9422);
or U9541 (N_9541,N_9415,N_9463);
and U9542 (N_9542,N_9424,N_9448);
nand U9543 (N_9543,N_9442,N_9407);
nand U9544 (N_9544,N_9496,N_9403);
xnor U9545 (N_9545,N_9419,N_9433);
xnor U9546 (N_9546,N_9457,N_9490);
nor U9547 (N_9547,N_9488,N_9462);
and U9548 (N_9548,N_9473,N_9438);
nor U9549 (N_9549,N_9455,N_9444);
nor U9550 (N_9550,N_9471,N_9496);
or U9551 (N_9551,N_9412,N_9440);
nand U9552 (N_9552,N_9464,N_9462);
and U9553 (N_9553,N_9424,N_9495);
and U9554 (N_9554,N_9483,N_9447);
nor U9555 (N_9555,N_9478,N_9409);
nor U9556 (N_9556,N_9437,N_9426);
nor U9557 (N_9557,N_9408,N_9454);
nor U9558 (N_9558,N_9408,N_9407);
nor U9559 (N_9559,N_9490,N_9446);
nand U9560 (N_9560,N_9444,N_9461);
nand U9561 (N_9561,N_9499,N_9482);
or U9562 (N_9562,N_9481,N_9442);
or U9563 (N_9563,N_9432,N_9442);
and U9564 (N_9564,N_9481,N_9409);
nor U9565 (N_9565,N_9418,N_9466);
nor U9566 (N_9566,N_9449,N_9425);
nand U9567 (N_9567,N_9442,N_9402);
nand U9568 (N_9568,N_9414,N_9419);
xor U9569 (N_9569,N_9479,N_9454);
or U9570 (N_9570,N_9455,N_9434);
or U9571 (N_9571,N_9428,N_9435);
or U9572 (N_9572,N_9463,N_9453);
and U9573 (N_9573,N_9419,N_9492);
nor U9574 (N_9574,N_9499,N_9413);
or U9575 (N_9575,N_9421,N_9439);
and U9576 (N_9576,N_9436,N_9434);
and U9577 (N_9577,N_9475,N_9487);
nand U9578 (N_9578,N_9402,N_9450);
or U9579 (N_9579,N_9408,N_9422);
or U9580 (N_9580,N_9412,N_9448);
or U9581 (N_9581,N_9473,N_9462);
nor U9582 (N_9582,N_9425,N_9462);
nor U9583 (N_9583,N_9405,N_9411);
nand U9584 (N_9584,N_9472,N_9421);
nor U9585 (N_9585,N_9475,N_9405);
or U9586 (N_9586,N_9407,N_9466);
nor U9587 (N_9587,N_9438,N_9413);
or U9588 (N_9588,N_9409,N_9462);
nor U9589 (N_9589,N_9474,N_9448);
nor U9590 (N_9590,N_9400,N_9434);
nand U9591 (N_9591,N_9452,N_9428);
nand U9592 (N_9592,N_9471,N_9432);
nor U9593 (N_9593,N_9466,N_9435);
or U9594 (N_9594,N_9469,N_9474);
or U9595 (N_9595,N_9499,N_9468);
nand U9596 (N_9596,N_9474,N_9478);
or U9597 (N_9597,N_9484,N_9422);
nor U9598 (N_9598,N_9446,N_9431);
nand U9599 (N_9599,N_9404,N_9456);
nor U9600 (N_9600,N_9597,N_9524);
nand U9601 (N_9601,N_9564,N_9539);
xnor U9602 (N_9602,N_9589,N_9575);
nor U9603 (N_9603,N_9565,N_9540);
and U9604 (N_9604,N_9504,N_9557);
and U9605 (N_9605,N_9576,N_9598);
and U9606 (N_9606,N_9570,N_9535);
xor U9607 (N_9607,N_9568,N_9596);
or U9608 (N_9608,N_9595,N_9543);
and U9609 (N_9609,N_9549,N_9534);
and U9610 (N_9610,N_9551,N_9523);
and U9611 (N_9611,N_9542,N_9517);
or U9612 (N_9612,N_9558,N_9591);
xor U9613 (N_9613,N_9544,N_9548);
or U9614 (N_9614,N_9514,N_9559);
and U9615 (N_9615,N_9560,N_9506);
nand U9616 (N_9616,N_9521,N_9580);
nand U9617 (N_9617,N_9553,N_9546);
and U9618 (N_9618,N_9563,N_9511);
xor U9619 (N_9619,N_9577,N_9538);
or U9620 (N_9620,N_9578,N_9522);
xor U9621 (N_9621,N_9574,N_9516);
nand U9622 (N_9622,N_9592,N_9550);
xor U9623 (N_9623,N_9507,N_9527);
and U9624 (N_9624,N_9573,N_9541);
and U9625 (N_9625,N_9533,N_9505);
nand U9626 (N_9626,N_9552,N_9536);
nand U9627 (N_9627,N_9566,N_9518);
xor U9628 (N_9628,N_9512,N_9581);
and U9629 (N_9629,N_9502,N_9556);
or U9630 (N_9630,N_9579,N_9567);
nor U9631 (N_9631,N_9586,N_9525);
nor U9632 (N_9632,N_9500,N_9554);
xnor U9633 (N_9633,N_9594,N_9513);
nor U9634 (N_9634,N_9508,N_9571);
xor U9635 (N_9635,N_9545,N_9562);
and U9636 (N_9636,N_9530,N_9584);
nand U9637 (N_9637,N_9590,N_9555);
nor U9638 (N_9638,N_9531,N_9526);
and U9639 (N_9639,N_9582,N_9529);
nand U9640 (N_9640,N_9515,N_9561);
nand U9641 (N_9641,N_9583,N_9587);
and U9642 (N_9642,N_9572,N_9547);
or U9643 (N_9643,N_9519,N_9510);
or U9644 (N_9644,N_9593,N_9503);
nand U9645 (N_9645,N_9588,N_9532);
xor U9646 (N_9646,N_9509,N_9528);
nand U9647 (N_9647,N_9599,N_9501);
and U9648 (N_9648,N_9569,N_9520);
nor U9649 (N_9649,N_9585,N_9537);
or U9650 (N_9650,N_9527,N_9536);
nand U9651 (N_9651,N_9507,N_9557);
or U9652 (N_9652,N_9564,N_9538);
xnor U9653 (N_9653,N_9525,N_9532);
nand U9654 (N_9654,N_9527,N_9571);
nand U9655 (N_9655,N_9577,N_9570);
nand U9656 (N_9656,N_9523,N_9517);
nor U9657 (N_9657,N_9557,N_9538);
and U9658 (N_9658,N_9525,N_9555);
nor U9659 (N_9659,N_9576,N_9552);
nor U9660 (N_9660,N_9523,N_9590);
xnor U9661 (N_9661,N_9504,N_9570);
or U9662 (N_9662,N_9543,N_9541);
nor U9663 (N_9663,N_9519,N_9554);
or U9664 (N_9664,N_9558,N_9586);
nand U9665 (N_9665,N_9510,N_9552);
nand U9666 (N_9666,N_9538,N_9526);
or U9667 (N_9667,N_9583,N_9507);
nor U9668 (N_9668,N_9582,N_9512);
xnor U9669 (N_9669,N_9553,N_9540);
nor U9670 (N_9670,N_9505,N_9581);
nand U9671 (N_9671,N_9534,N_9535);
nand U9672 (N_9672,N_9565,N_9570);
nor U9673 (N_9673,N_9544,N_9515);
and U9674 (N_9674,N_9564,N_9503);
nor U9675 (N_9675,N_9594,N_9524);
xor U9676 (N_9676,N_9568,N_9543);
or U9677 (N_9677,N_9520,N_9596);
xor U9678 (N_9678,N_9594,N_9595);
and U9679 (N_9679,N_9568,N_9500);
or U9680 (N_9680,N_9557,N_9595);
nor U9681 (N_9681,N_9580,N_9549);
and U9682 (N_9682,N_9553,N_9505);
and U9683 (N_9683,N_9501,N_9544);
xor U9684 (N_9684,N_9516,N_9528);
or U9685 (N_9685,N_9521,N_9537);
nor U9686 (N_9686,N_9551,N_9581);
and U9687 (N_9687,N_9505,N_9510);
and U9688 (N_9688,N_9510,N_9548);
or U9689 (N_9689,N_9595,N_9570);
nand U9690 (N_9690,N_9587,N_9506);
nand U9691 (N_9691,N_9586,N_9530);
or U9692 (N_9692,N_9512,N_9538);
nor U9693 (N_9693,N_9573,N_9592);
or U9694 (N_9694,N_9568,N_9572);
nand U9695 (N_9695,N_9545,N_9572);
xor U9696 (N_9696,N_9590,N_9534);
and U9697 (N_9697,N_9582,N_9551);
nand U9698 (N_9698,N_9513,N_9570);
nand U9699 (N_9699,N_9580,N_9553);
or U9700 (N_9700,N_9639,N_9662);
nor U9701 (N_9701,N_9637,N_9686);
nor U9702 (N_9702,N_9698,N_9624);
xor U9703 (N_9703,N_9646,N_9631);
nor U9704 (N_9704,N_9622,N_9685);
nor U9705 (N_9705,N_9649,N_9640);
and U9706 (N_9706,N_9605,N_9677);
nand U9707 (N_9707,N_9652,N_9656);
and U9708 (N_9708,N_9654,N_9651);
and U9709 (N_9709,N_9611,N_9665);
nor U9710 (N_9710,N_9653,N_9642);
and U9711 (N_9711,N_9666,N_9647);
nand U9712 (N_9712,N_9683,N_9658);
xnor U9713 (N_9713,N_9607,N_9641);
nand U9714 (N_9714,N_9634,N_9603);
nor U9715 (N_9715,N_9601,N_9648);
or U9716 (N_9716,N_9676,N_9674);
nor U9717 (N_9717,N_9678,N_9673);
nand U9718 (N_9718,N_9661,N_9664);
nand U9719 (N_9719,N_9663,N_9696);
nand U9720 (N_9720,N_9645,N_9687);
nor U9721 (N_9721,N_9660,N_9657);
or U9722 (N_9722,N_9621,N_9667);
nor U9723 (N_9723,N_9638,N_9623);
nand U9724 (N_9724,N_9606,N_9632);
nand U9725 (N_9725,N_9689,N_9612);
or U9726 (N_9726,N_9688,N_9681);
nor U9727 (N_9727,N_9616,N_9694);
or U9728 (N_9728,N_9615,N_9644);
nand U9729 (N_9729,N_9618,N_9655);
and U9730 (N_9730,N_9680,N_9609);
and U9731 (N_9731,N_9608,N_9697);
or U9732 (N_9732,N_9633,N_9675);
and U9733 (N_9733,N_9636,N_9668);
nor U9734 (N_9734,N_9692,N_9614);
nand U9735 (N_9735,N_9691,N_9684);
xor U9736 (N_9736,N_9650,N_9604);
and U9737 (N_9737,N_9629,N_9643);
or U9738 (N_9738,N_9672,N_9635);
nand U9739 (N_9739,N_9619,N_9625);
nor U9740 (N_9740,N_9679,N_9600);
or U9741 (N_9741,N_9693,N_9659);
or U9742 (N_9742,N_9613,N_9670);
nor U9743 (N_9743,N_9626,N_9669);
nand U9744 (N_9744,N_9627,N_9671);
nand U9745 (N_9745,N_9630,N_9628);
nand U9746 (N_9746,N_9682,N_9690);
nand U9747 (N_9747,N_9602,N_9620);
nand U9748 (N_9748,N_9617,N_9610);
nand U9749 (N_9749,N_9699,N_9695);
xor U9750 (N_9750,N_9667,N_9609);
or U9751 (N_9751,N_9686,N_9602);
xnor U9752 (N_9752,N_9634,N_9602);
nand U9753 (N_9753,N_9679,N_9665);
or U9754 (N_9754,N_9694,N_9615);
nand U9755 (N_9755,N_9645,N_9648);
nand U9756 (N_9756,N_9648,N_9653);
nand U9757 (N_9757,N_9653,N_9623);
xnor U9758 (N_9758,N_9630,N_9611);
nand U9759 (N_9759,N_9650,N_9654);
and U9760 (N_9760,N_9617,N_9655);
nor U9761 (N_9761,N_9634,N_9661);
nor U9762 (N_9762,N_9697,N_9659);
nand U9763 (N_9763,N_9651,N_9689);
or U9764 (N_9764,N_9696,N_9662);
nor U9765 (N_9765,N_9623,N_9671);
nand U9766 (N_9766,N_9614,N_9638);
nand U9767 (N_9767,N_9608,N_9629);
nand U9768 (N_9768,N_9609,N_9686);
and U9769 (N_9769,N_9685,N_9667);
and U9770 (N_9770,N_9635,N_9639);
nor U9771 (N_9771,N_9654,N_9653);
and U9772 (N_9772,N_9650,N_9616);
nor U9773 (N_9773,N_9673,N_9681);
nor U9774 (N_9774,N_9688,N_9661);
nor U9775 (N_9775,N_9687,N_9688);
nand U9776 (N_9776,N_9676,N_9657);
or U9777 (N_9777,N_9693,N_9633);
nand U9778 (N_9778,N_9693,N_9653);
nor U9779 (N_9779,N_9651,N_9605);
nand U9780 (N_9780,N_9682,N_9679);
nor U9781 (N_9781,N_9665,N_9608);
and U9782 (N_9782,N_9637,N_9667);
nand U9783 (N_9783,N_9648,N_9654);
nor U9784 (N_9784,N_9647,N_9682);
xnor U9785 (N_9785,N_9620,N_9615);
nand U9786 (N_9786,N_9620,N_9600);
xor U9787 (N_9787,N_9643,N_9695);
nand U9788 (N_9788,N_9634,N_9635);
or U9789 (N_9789,N_9652,N_9604);
xor U9790 (N_9790,N_9619,N_9605);
nand U9791 (N_9791,N_9635,N_9613);
nor U9792 (N_9792,N_9638,N_9642);
nor U9793 (N_9793,N_9630,N_9619);
nand U9794 (N_9794,N_9675,N_9648);
or U9795 (N_9795,N_9609,N_9691);
or U9796 (N_9796,N_9643,N_9685);
or U9797 (N_9797,N_9688,N_9666);
nor U9798 (N_9798,N_9615,N_9643);
nor U9799 (N_9799,N_9621,N_9674);
nand U9800 (N_9800,N_9720,N_9770);
or U9801 (N_9801,N_9705,N_9724);
and U9802 (N_9802,N_9757,N_9725);
nor U9803 (N_9803,N_9774,N_9728);
xnor U9804 (N_9804,N_9733,N_9749);
and U9805 (N_9805,N_9798,N_9708);
nand U9806 (N_9806,N_9716,N_9755);
nand U9807 (N_9807,N_9775,N_9727);
or U9808 (N_9808,N_9793,N_9717);
and U9809 (N_9809,N_9769,N_9737);
xor U9810 (N_9810,N_9796,N_9799);
and U9811 (N_9811,N_9702,N_9759);
nand U9812 (N_9812,N_9712,N_9711);
xor U9813 (N_9813,N_9714,N_9732);
nor U9814 (N_9814,N_9776,N_9772);
nand U9815 (N_9815,N_9742,N_9768);
nor U9816 (N_9816,N_9771,N_9762);
or U9817 (N_9817,N_9751,N_9789);
xor U9818 (N_9818,N_9758,N_9753);
and U9819 (N_9819,N_9773,N_9763);
nor U9820 (N_9820,N_9704,N_9765);
and U9821 (N_9821,N_9752,N_9736);
and U9822 (N_9822,N_9795,N_9760);
nor U9823 (N_9823,N_9788,N_9747);
nor U9824 (N_9824,N_9744,N_9734);
or U9825 (N_9825,N_9791,N_9780);
nor U9826 (N_9826,N_9722,N_9746);
and U9827 (N_9827,N_9787,N_9782);
xor U9828 (N_9828,N_9745,N_9735);
nor U9829 (N_9829,N_9738,N_9777);
nand U9830 (N_9830,N_9743,N_9764);
or U9831 (N_9831,N_9721,N_9726);
and U9832 (N_9832,N_9785,N_9794);
and U9833 (N_9833,N_9754,N_9739);
and U9834 (N_9834,N_9713,N_9792);
or U9835 (N_9835,N_9797,N_9701);
xnor U9836 (N_9836,N_9748,N_9784);
or U9837 (N_9837,N_9786,N_9700);
nor U9838 (N_9838,N_9766,N_9731);
or U9839 (N_9839,N_9715,N_9709);
nand U9840 (N_9840,N_9779,N_9761);
or U9841 (N_9841,N_9756,N_9719);
nor U9842 (N_9842,N_9718,N_9778);
nand U9843 (N_9843,N_9790,N_9750);
and U9844 (N_9844,N_9703,N_9740);
or U9845 (N_9845,N_9729,N_9781);
nand U9846 (N_9846,N_9710,N_9706);
or U9847 (N_9847,N_9730,N_9707);
xnor U9848 (N_9848,N_9783,N_9767);
nand U9849 (N_9849,N_9741,N_9723);
nor U9850 (N_9850,N_9732,N_9705);
nor U9851 (N_9851,N_9744,N_9711);
nand U9852 (N_9852,N_9774,N_9786);
xor U9853 (N_9853,N_9724,N_9728);
nor U9854 (N_9854,N_9791,N_9703);
nand U9855 (N_9855,N_9735,N_9720);
and U9856 (N_9856,N_9778,N_9775);
and U9857 (N_9857,N_9768,N_9723);
nor U9858 (N_9858,N_9798,N_9710);
nor U9859 (N_9859,N_9737,N_9741);
or U9860 (N_9860,N_9725,N_9793);
nor U9861 (N_9861,N_9744,N_9729);
and U9862 (N_9862,N_9720,N_9739);
nand U9863 (N_9863,N_9752,N_9759);
nand U9864 (N_9864,N_9721,N_9780);
nand U9865 (N_9865,N_9703,N_9781);
nor U9866 (N_9866,N_9741,N_9763);
xor U9867 (N_9867,N_9791,N_9702);
nand U9868 (N_9868,N_9784,N_9704);
or U9869 (N_9869,N_9777,N_9769);
nand U9870 (N_9870,N_9774,N_9782);
and U9871 (N_9871,N_9723,N_9707);
nand U9872 (N_9872,N_9781,N_9704);
nand U9873 (N_9873,N_9757,N_9763);
nor U9874 (N_9874,N_9787,N_9711);
nand U9875 (N_9875,N_9772,N_9787);
nand U9876 (N_9876,N_9736,N_9745);
and U9877 (N_9877,N_9726,N_9713);
and U9878 (N_9878,N_9776,N_9788);
xnor U9879 (N_9879,N_9709,N_9757);
nand U9880 (N_9880,N_9743,N_9750);
or U9881 (N_9881,N_9709,N_9797);
and U9882 (N_9882,N_9717,N_9745);
and U9883 (N_9883,N_9756,N_9794);
and U9884 (N_9884,N_9762,N_9768);
or U9885 (N_9885,N_9780,N_9738);
or U9886 (N_9886,N_9751,N_9757);
xnor U9887 (N_9887,N_9724,N_9709);
nor U9888 (N_9888,N_9747,N_9740);
or U9889 (N_9889,N_9793,N_9761);
and U9890 (N_9890,N_9703,N_9735);
and U9891 (N_9891,N_9720,N_9799);
or U9892 (N_9892,N_9754,N_9765);
nor U9893 (N_9893,N_9712,N_9730);
or U9894 (N_9894,N_9725,N_9777);
or U9895 (N_9895,N_9753,N_9708);
and U9896 (N_9896,N_9720,N_9709);
or U9897 (N_9897,N_9701,N_9789);
and U9898 (N_9898,N_9710,N_9784);
nor U9899 (N_9899,N_9777,N_9760);
nor U9900 (N_9900,N_9841,N_9872);
nor U9901 (N_9901,N_9851,N_9822);
nor U9902 (N_9902,N_9850,N_9857);
nor U9903 (N_9903,N_9848,N_9801);
nand U9904 (N_9904,N_9837,N_9889);
and U9905 (N_9905,N_9821,N_9805);
xor U9906 (N_9906,N_9880,N_9860);
nor U9907 (N_9907,N_9864,N_9881);
or U9908 (N_9908,N_9847,N_9849);
or U9909 (N_9909,N_9818,N_9843);
xnor U9910 (N_9910,N_9867,N_9884);
xor U9911 (N_9911,N_9898,N_9809);
or U9912 (N_9912,N_9856,N_9861);
or U9913 (N_9913,N_9874,N_9883);
nor U9914 (N_9914,N_9854,N_9887);
nor U9915 (N_9915,N_9892,N_9834);
nor U9916 (N_9916,N_9811,N_9815);
or U9917 (N_9917,N_9835,N_9804);
nand U9918 (N_9918,N_9807,N_9895);
or U9919 (N_9919,N_9899,N_9840);
and U9920 (N_9920,N_9871,N_9877);
or U9921 (N_9921,N_9838,N_9875);
or U9922 (N_9922,N_9820,N_9812);
nor U9923 (N_9923,N_9819,N_9814);
nor U9924 (N_9924,N_9845,N_9882);
nand U9925 (N_9925,N_9865,N_9816);
nand U9926 (N_9926,N_9808,N_9886);
or U9927 (N_9927,N_9855,N_9817);
nand U9928 (N_9928,N_9852,N_9894);
nand U9929 (N_9929,N_9866,N_9828);
nand U9930 (N_9930,N_9893,N_9813);
and U9931 (N_9931,N_9885,N_9833);
xor U9932 (N_9932,N_9862,N_9890);
or U9933 (N_9933,N_9810,N_9836);
nor U9934 (N_9934,N_9824,N_9823);
nand U9935 (N_9935,N_9839,N_9827);
xnor U9936 (N_9936,N_9846,N_9829);
xor U9937 (N_9937,N_9897,N_9858);
and U9938 (N_9938,N_9879,N_9870);
nor U9939 (N_9939,N_9878,N_9868);
and U9940 (N_9940,N_9888,N_9853);
nand U9941 (N_9941,N_9876,N_9844);
nor U9942 (N_9942,N_9830,N_9825);
nor U9943 (N_9943,N_9896,N_9863);
nor U9944 (N_9944,N_9800,N_9802);
or U9945 (N_9945,N_9859,N_9826);
or U9946 (N_9946,N_9832,N_9891);
or U9947 (N_9947,N_9806,N_9842);
and U9948 (N_9948,N_9869,N_9831);
and U9949 (N_9949,N_9873,N_9803);
nand U9950 (N_9950,N_9881,N_9890);
and U9951 (N_9951,N_9859,N_9860);
nor U9952 (N_9952,N_9888,N_9802);
or U9953 (N_9953,N_9826,N_9878);
nor U9954 (N_9954,N_9801,N_9845);
and U9955 (N_9955,N_9841,N_9888);
and U9956 (N_9956,N_9808,N_9893);
or U9957 (N_9957,N_9876,N_9868);
or U9958 (N_9958,N_9867,N_9830);
nand U9959 (N_9959,N_9825,N_9814);
and U9960 (N_9960,N_9810,N_9896);
nand U9961 (N_9961,N_9863,N_9861);
or U9962 (N_9962,N_9887,N_9839);
xor U9963 (N_9963,N_9818,N_9898);
and U9964 (N_9964,N_9877,N_9858);
nand U9965 (N_9965,N_9851,N_9897);
nor U9966 (N_9966,N_9805,N_9845);
or U9967 (N_9967,N_9864,N_9839);
or U9968 (N_9968,N_9835,N_9873);
nor U9969 (N_9969,N_9833,N_9804);
nor U9970 (N_9970,N_9854,N_9878);
nand U9971 (N_9971,N_9883,N_9895);
nand U9972 (N_9972,N_9842,N_9803);
xnor U9973 (N_9973,N_9834,N_9819);
or U9974 (N_9974,N_9881,N_9842);
nand U9975 (N_9975,N_9853,N_9885);
nor U9976 (N_9976,N_9807,N_9884);
nand U9977 (N_9977,N_9889,N_9838);
nor U9978 (N_9978,N_9888,N_9842);
or U9979 (N_9979,N_9872,N_9837);
and U9980 (N_9980,N_9856,N_9838);
nand U9981 (N_9981,N_9805,N_9880);
and U9982 (N_9982,N_9876,N_9845);
nand U9983 (N_9983,N_9800,N_9878);
nand U9984 (N_9984,N_9844,N_9803);
or U9985 (N_9985,N_9881,N_9897);
or U9986 (N_9986,N_9806,N_9854);
nor U9987 (N_9987,N_9886,N_9859);
or U9988 (N_9988,N_9852,N_9890);
nor U9989 (N_9989,N_9885,N_9808);
and U9990 (N_9990,N_9896,N_9856);
nor U9991 (N_9991,N_9833,N_9834);
and U9992 (N_9992,N_9892,N_9816);
xor U9993 (N_9993,N_9863,N_9823);
and U9994 (N_9994,N_9805,N_9812);
and U9995 (N_9995,N_9873,N_9898);
and U9996 (N_9996,N_9875,N_9842);
or U9997 (N_9997,N_9823,N_9862);
or U9998 (N_9998,N_9825,N_9865);
nor U9999 (N_9999,N_9822,N_9871);
nand UO_0 (O_0,N_9943,N_9931);
or UO_1 (O_1,N_9906,N_9941);
or UO_2 (O_2,N_9917,N_9970);
xor UO_3 (O_3,N_9932,N_9912);
nor UO_4 (O_4,N_9983,N_9947);
and UO_5 (O_5,N_9937,N_9997);
and UO_6 (O_6,N_9989,N_9910);
xnor UO_7 (O_7,N_9938,N_9998);
nand UO_8 (O_8,N_9969,N_9979);
and UO_9 (O_9,N_9935,N_9950);
nor UO_10 (O_10,N_9918,N_9958);
and UO_11 (O_11,N_9934,N_9920);
nor UO_12 (O_12,N_9963,N_9996);
and UO_13 (O_13,N_9921,N_9953);
nand UO_14 (O_14,N_9913,N_9976);
nand UO_15 (O_15,N_9954,N_9914);
and UO_16 (O_16,N_9901,N_9999);
nor UO_17 (O_17,N_9929,N_9940);
nand UO_18 (O_18,N_9975,N_9967);
or UO_19 (O_19,N_9986,N_9987);
or UO_20 (O_20,N_9984,N_9994);
xor UO_21 (O_21,N_9946,N_9911);
nor UO_22 (O_22,N_9991,N_9919);
or UO_23 (O_23,N_9985,N_9971);
xor UO_24 (O_24,N_9908,N_9952);
nand UO_25 (O_25,N_9949,N_9992);
xor UO_26 (O_26,N_9942,N_9903);
nand UO_27 (O_27,N_9928,N_9962);
and UO_28 (O_28,N_9981,N_9982);
xor UO_29 (O_29,N_9965,N_9955);
xor UO_30 (O_30,N_9904,N_9995);
and UO_31 (O_31,N_9916,N_9907);
nor UO_32 (O_32,N_9966,N_9915);
and UO_33 (O_33,N_9972,N_9980);
nor UO_34 (O_34,N_9964,N_9905);
nand UO_35 (O_35,N_9993,N_9944);
nand UO_36 (O_36,N_9930,N_9974);
nor UO_37 (O_37,N_9925,N_9936);
nand UO_38 (O_38,N_9939,N_9961);
or UO_39 (O_39,N_9923,N_9960);
or UO_40 (O_40,N_9924,N_9927);
or UO_41 (O_41,N_9951,N_9990);
xor UO_42 (O_42,N_9988,N_9978);
nor UO_43 (O_43,N_9977,N_9968);
nand UO_44 (O_44,N_9900,N_9945);
xor UO_45 (O_45,N_9926,N_9922);
or UO_46 (O_46,N_9956,N_9948);
and UO_47 (O_47,N_9973,N_9909);
or UO_48 (O_48,N_9933,N_9902);
or UO_49 (O_49,N_9959,N_9957);
nand UO_50 (O_50,N_9952,N_9993);
and UO_51 (O_51,N_9955,N_9956);
nor UO_52 (O_52,N_9919,N_9975);
nor UO_53 (O_53,N_9915,N_9986);
and UO_54 (O_54,N_9929,N_9971);
nand UO_55 (O_55,N_9998,N_9978);
or UO_56 (O_56,N_9913,N_9938);
nor UO_57 (O_57,N_9977,N_9949);
and UO_58 (O_58,N_9914,N_9990);
and UO_59 (O_59,N_9999,N_9972);
or UO_60 (O_60,N_9945,N_9956);
and UO_61 (O_61,N_9985,N_9935);
nand UO_62 (O_62,N_9900,N_9964);
or UO_63 (O_63,N_9902,N_9966);
or UO_64 (O_64,N_9970,N_9910);
nand UO_65 (O_65,N_9983,N_9998);
and UO_66 (O_66,N_9926,N_9939);
nor UO_67 (O_67,N_9901,N_9972);
or UO_68 (O_68,N_9938,N_9920);
and UO_69 (O_69,N_9931,N_9997);
and UO_70 (O_70,N_9962,N_9936);
nor UO_71 (O_71,N_9944,N_9920);
xor UO_72 (O_72,N_9941,N_9931);
nand UO_73 (O_73,N_9969,N_9956);
nand UO_74 (O_74,N_9928,N_9919);
nor UO_75 (O_75,N_9903,N_9927);
nor UO_76 (O_76,N_9918,N_9900);
or UO_77 (O_77,N_9911,N_9941);
nor UO_78 (O_78,N_9964,N_9971);
and UO_79 (O_79,N_9963,N_9991);
and UO_80 (O_80,N_9939,N_9929);
or UO_81 (O_81,N_9949,N_9940);
or UO_82 (O_82,N_9990,N_9964);
or UO_83 (O_83,N_9905,N_9970);
and UO_84 (O_84,N_9923,N_9908);
nor UO_85 (O_85,N_9932,N_9991);
nor UO_86 (O_86,N_9968,N_9994);
nor UO_87 (O_87,N_9956,N_9993);
nor UO_88 (O_88,N_9962,N_9925);
or UO_89 (O_89,N_9994,N_9919);
or UO_90 (O_90,N_9945,N_9905);
nor UO_91 (O_91,N_9969,N_9937);
nand UO_92 (O_92,N_9910,N_9927);
or UO_93 (O_93,N_9970,N_9946);
or UO_94 (O_94,N_9996,N_9922);
nand UO_95 (O_95,N_9930,N_9969);
xor UO_96 (O_96,N_9967,N_9966);
and UO_97 (O_97,N_9917,N_9988);
nor UO_98 (O_98,N_9982,N_9916);
and UO_99 (O_99,N_9933,N_9976);
nor UO_100 (O_100,N_9946,N_9902);
nor UO_101 (O_101,N_9942,N_9943);
nand UO_102 (O_102,N_9944,N_9918);
and UO_103 (O_103,N_9919,N_9940);
nand UO_104 (O_104,N_9915,N_9960);
and UO_105 (O_105,N_9907,N_9977);
xnor UO_106 (O_106,N_9908,N_9983);
nor UO_107 (O_107,N_9921,N_9952);
nand UO_108 (O_108,N_9945,N_9997);
xor UO_109 (O_109,N_9959,N_9955);
and UO_110 (O_110,N_9919,N_9999);
nor UO_111 (O_111,N_9936,N_9983);
nand UO_112 (O_112,N_9963,N_9990);
or UO_113 (O_113,N_9984,N_9926);
or UO_114 (O_114,N_9906,N_9911);
nand UO_115 (O_115,N_9957,N_9981);
xor UO_116 (O_116,N_9967,N_9935);
nand UO_117 (O_117,N_9993,N_9950);
and UO_118 (O_118,N_9903,N_9961);
and UO_119 (O_119,N_9972,N_9918);
and UO_120 (O_120,N_9938,N_9911);
and UO_121 (O_121,N_9906,N_9992);
and UO_122 (O_122,N_9939,N_9946);
nand UO_123 (O_123,N_9916,N_9974);
xor UO_124 (O_124,N_9907,N_9908);
nor UO_125 (O_125,N_9927,N_9981);
and UO_126 (O_126,N_9903,N_9997);
nand UO_127 (O_127,N_9956,N_9954);
nor UO_128 (O_128,N_9918,N_9964);
or UO_129 (O_129,N_9936,N_9987);
nor UO_130 (O_130,N_9922,N_9972);
nor UO_131 (O_131,N_9993,N_9930);
xnor UO_132 (O_132,N_9979,N_9913);
and UO_133 (O_133,N_9952,N_9919);
or UO_134 (O_134,N_9938,N_9994);
or UO_135 (O_135,N_9956,N_9970);
nor UO_136 (O_136,N_9922,N_9969);
nor UO_137 (O_137,N_9986,N_9962);
and UO_138 (O_138,N_9990,N_9910);
nand UO_139 (O_139,N_9904,N_9928);
nand UO_140 (O_140,N_9933,N_9934);
nor UO_141 (O_141,N_9952,N_9990);
and UO_142 (O_142,N_9978,N_9961);
nor UO_143 (O_143,N_9974,N_9951);
or UO_144 (O_144,N_9939,N_9913);
nor UO_145 (O_145,N_9972,N_9995);
nand UO_146 (O_146,N_9917,N_9967);
nor UO_147 (O_147,N_9991,N_9903);
nor UO_148 (O_148,N_9925,N_9932);
nand UO_149 (O_149,N_9906,N_9998);
or UO_150 (O_150,N_9932,N_9918);
nor UO_151 (O_151,N_9983,N_9945);
nor UO_152 (O_152,N_9904,N_9961);
nor UO_153 (O_153,N_9926,N_9986);
nor UO_154 (O_154,N_9996,N_9965);
nor UO_155 (O_155,N_9979,N_9957);
xnor UO_156 (O_156,N_9911,N_9926);
or UO_157 (O_157,N_9936,N_9953);
nor UO_158 (O_158,N_9918,N_9978);
and UO_159 (O_159,N_9947,N_9961);
nor UO_160 (O_160,N_9924,N_9941);
and UO_161 (O_161,N_9972,N_9988);
and UO_162 (O_162,N_9925,N_9922);
nor UO_163 (O_163,N_9933,N_9916);
nor UO_164 (O_164,N_9908,N_9970);
nand UO_165 (O_165,N_9966,N_9920);
or UO_166 (O_166,N_9980,N_9962);
xor UO_167 (O_167,N_9909,N_9993);
xnor UO_168 (O_168,N_9939,N_9907);
xnor UO_169 (O_169,N_9941,N_9988);
nand UO_170 (O_170,N_9934,N_9935);
or UO_171 (O_171,N_9931,N_9985);
xnor UO_172 (O_172,N_9924,N_9969);
or UO_173 (O_173,N_9913,N_9928);
and UO_174 (O_174,N_9909,N_9982);
nand UO_175 (O_175,N_9909,N_9990);
nand UO_176 (O_176,N_9949,N_9948);
and UO_177 (O_177,N_9986,N_9983);
xor UO_178 (O_178,N_9970,N_9966);
nand UO_179 (O_179,N_9913,N_9948);
nand UO_180 (O_180,N_9924,N_9913);
xnor UO_181 (O_181,N_9958,N_9997);
and UO_182 (O_182,N_9922,N_9958);
nor UO_183 (O_183,N_9943,N_9996);
nor UO_184 (O_184,N_9925,N_9990);
or UO_185 (O_185,N_9911,N_9962);
nand UO_186 (O_186,N_9921,N_9963);
nor UO_187 (O_187,N_9947,N_9982);
and UO_188 (O_188,N_9926,N_9929);
nor UO_189 (O_189,N_9912,N_9968);
or UO_190 (O_190,N_9921,N_9915);
nor UO_191 (O_191,N_9923,N_9957);
nand UO_192 (O_192,N_9997,N_9979);
and UO_193 (O_193,N_9925,N_9927);
nor UO_194 (O_194,N_9935,N_9918);
nor UO_195 (O_195,N_9977,N_9917);
nand UO_196 (O_196,N_9993,N_9988);
or UO_197 (O_197,N_9999,N_9974);
nand UO_198 (O_198,N_9994,N_9929);
and UO_199 (O_199,N_9925,N_9959);
or UO_200 (O_200,N_9956,N_9989);
and UO_201 (O_201,N_9933,N_9977);
nor UO_202 (O_202,N_9998,N_9988);
nor UO_203 (O_203,N_9945,N_9976);
xnor UO_204 (O_204,N_9929,N_9923);
xor UO_205 (O_205,N_9963,N_9999);
nor UO_206 (O_206,N_9981,N_9939);
nand UO_207 (O_207,N_9995,N_9959);
and UO_208 (O_208,N_9972,N_9974);
xor UO_209 (O_209,N_9952,N_9962);
nor UO_210 (O_210,N_9975,N_9946);
or UO_211 (O_211,N_9993,N_9919);
and UO_212 (O_212,N_9982,N_9965);
nor UO_213 (O_213,N_9952,N_9941);
xor UO_214 (O_214,N_9973,N_9946);
nor UO_215 (O_215,N_9934,N_9989);
nor UO_216 (O_216,N_9974,N_9960);
xnor UO_217 (O_217,N_9973,N_9979);
or UO_218 (O_218,N_9941,N_9912);
nor UO_219 (O_219,N_9968,N_9931);
or UO_220 (O_220,N_9979,N_9962);
nand UO_221 (O_221,N_9964,N_9917);
or UO_222 (O_222,N_9960,N_9995);
nand UO_223 (O_223,N_9933,N_9914);
nand UO_224 (O_224,N_9972,N_9916);
and UO_225 (O_225,N_9998,N_9957);
and UO_226 (O_226,N_9910,N_9957);
and UO_227 (O_227,N_9942,N_9958);
and UO_228 (O_228,N_9920,N_9913);
or UO_229 (O_229,N_9963,N_9952);
nor UO_230 (O_230,N_9977,N_9973);
nor UO_231 (O_231,N_9900,N_9901);
or UO_232 (O_232,N_9935,N_9958);
or UO_233 (O_233,N_9923,N_9928);
nand UO_234 (O_234,N_9934,N_9957);
nor UO_235 (O_235,N_9960,N_9977);
nand UO_236 (O_236,N_9993,N_9904);
nand UO_237 (O_237,N_9948,N_9987);
nor UO_238 (O_238,N_9996,N_9951);
and UO_239 (O_239,N_9953,N_9965);
nand UO_240 (O_240,N_9992,N_9952);
nor UO_241 (O_241,N_9937,N_9964);
xor UO_242 (O_242,N_9974,N_9928);
or UO_243 (O_243,N_9913,N_9930);
and UO_244 (O_244,N_9975,N_9985);
or UO_245 (O_245,N_9959,N_9974);
and UO_246 (O_246,N_9935,N_9951);
nand UO_247 (O_247,N_9975,N_9970);
or UO_248 (O_248,N_9963,N_9972);
or UO_249 (O_249,N_9983,N_9928);
or UO_250 (O_250,N_9992,N_9946);
xor UO_251 (O_251,N_9954,N_9983);
xor UO_252 (O_252,N_9959,N_9914);
nor UO_253 (O_253,N_9983,N_9904);
and UO_254 (O_254,N_9931,N_9945);
nand UO_255 (O_255,N_9970,N_9909);
or UO_256 (O_256,N_9901,N_9913);
xnor UO_257 (O_257,N_9907,N_9923);
nand UO_258 (O_258,N_9912,N_9939);
nor UO_259 (O_259,N_9929,N_9953);
or UO_260 (O_260,N_9902,N_9909);
or UO_261 (O_261,N_9937,N_9933);
nand UO_262 (O_262,N_9908,N_9905);
and UO_263 (O_263,N_9909,N_9985);
nand UO_264 (O_264,N_9987,N_9961);
nor UO_265 (O_265,N_9975,N_9982);
nand UO_266 (O_266,N_9953,N_9912);
or UO_267 (O_267,N_9903,N_9901);
nor UO_268 (O_268,N_9927,N_9957);
and UO_269 (O_269,N_9955,N_9930);
nand UO_270 (O_270,N_9937,N_9957);
nand UO_271 (O_271,N_9906,N_9904);
and UO_272 (O_272,N_9935,N_9987);
and UO_273 (O_273,N_9966,N_9901);
xnor UO_274 (O_274,N_9907,N_9928);
nand UO_275 (O_275,N_9931,N_9930);
xor UO_276 (O_276,N_9908,N_9964);
and UO_277 (O_277,N_9977,N_9981);
and UO_278 (O_278,N_9965,N_9957);
nor UO_279 (O_279,N_9915,N_9995);
nor UO_280 (O_280,N_9947,N_9907);
or UO_281 (O_281,N_9949,N_9985);
or UO_282 (O_282,N_9924,N_9978);
and UO_283 (O_283,N_9940,N_9983);
nand UO_284 (O_284,N_9964,N_9931);
and UO_285 (O_285,N_9957,N_9958);
nor UO_286 (O_286,N_9980,N_9947);
nor UO_287 (O_287,N_9922,N_9966);
nor UO_288 (O_288,N_9932,N_9945);
nor UO_289 (O_289,N_9902,N_9989);
or UO_290 (O_290,N_9955,N_9907);
nor UO_291 (O_291,N_9954,N_9904);
or UO_292 (O_292,N_9922,N_9990);
nor UO_293 (O_293,N_9927,N_9949);
or UO_294 (O_294,N_9983,N_9952);
or UO_295 (O_295,N_9940,N_9939);
nor UO_296 (O_296,N_9976,N_9957);
xnor UO_297 (O_297,N_9963,N_9930);
nor UO_298 (O_298,N_9930,N_9914);
or UO_299 (O_299,N_9972,N_9943);
nand UO_300 (O_300,N_9925,N_9961);
xnor UO_301 (O_301,N_9998,N_9939);
nor UO_302 (O_302,N_9997,N_9946);
or UO_303 (O_303,N_9985,N_9979);
nand UO_304 (O_304,N_9975,N_9988);
or UO_305 (O_305,N_9977,N_9963);
and UO_306 (O_306,N_9986,N_9904);
nor UO_307 (O_307,N_9906,N_9994);
nand UO_308 (O_308,N_9927,N_9914);
or UO_309 (O_309,N_9970,N_9985);
and UO_310 (O_310,N_9996,N_9950);
nand UO_311 (O_311,N_9970,N_9984);
nand UO_312 (O_312,N_9996,N_9959);
and UO_313 (O_313,N_9997,N_9940);
nor UO_314 (O_314,N_9903,N_9909);
or UO_315 (O_315,N_9991,N_9958);
xor UO_316 (O_316,N_9976,N_9964);
nand UO_317 (O_317,N_9986,N_9908);
and UO_318 (O_318,N_9912,N_9973);
and UO_319 (O_319,N_9922,N_9979);
nand UO_320 (O_320,N_9917,N_9924);
nand UO_321 (O_321,N_9947,N_9968);
nand UO_322 (O_322,N_9976,N_9983);
and UO_323 (O_323,N_9986,N_9959);
nor UO_324 (O_324,N_9936,N_9902);
xor UO_325 (O_325,N_9958,N_9912);
and UO_326 (O_326,N_9914,N_9936);
nand UO_327 (O_327,N_9993,N_9925);
nand UO_328 (O_328,N_9959,N_9964);
or UO_329 (O_329,N_9981,N_9984);
xor UO_330 (O_330,N_9952,N_9988);
nor UO_331 (O_331,N_9911,N_9992);
or UO_332 (O_332,N_9926,N_9976);
xor UO_333 (O_333,N_9963,N_9986);
and UO_334 (O_334,N_9938,N_9907);
xor UO_335 (O_335,N_9975,N_9901);
nor UO_336 (O_336,N_9929,N_9998);
or UO_337 (O_337,N_9918,N_9906);
nand UO_338 (O_338,N_9960,N_9914);
and UO_339 (O_339,N_9965,N_9910);
or UO_340 (O_340,N_9935,N_9925);
or UO_341 (O_341,N_9921,N_9945);
or UO_342 (O_342,N_9973,N_9925);
and UO_343 (O_343,N_9960,N_9924);
nor UO_344 (O_344,N_9995,N_9966);
nand UO_345 (O_345,N_9995,N_9990);
and UO_346 (O_346,N_9978,N_9968);
nor UO_347 (O_347,N_9981,N_9974);
nor UO_348 (O_348,N_9926,N_9989);
and UO_349 (O_349,N_9901,N_9959);
and UO_350 (O_350,N_9909,N_9943);
and UO_351 (O_351,N_9922,N_9962);
or UO_352 (O_352,N_9923,N_9950);
nand UO_353 (O_353,N_9955,N_9969);
nand UO_354 (O_354,N_9905,N_9978);
and UO_355 (O_355,N_9933,N_9998);
nor UO_356 (O_356,N_9948,N_9912);
and UO_357 (O_357,N_9956,N_9944);
nand UO_358 (O_358,N_9993,N_9996);
or UO_359 (O_359,N_9958,N_9939);
or UO_360 (O_360,N_9953,N_9920);
nand UO_361 (O_361,N_9934,N_9906);
and UO_362 (O_362,N_9928,N_9921);
or UO_363 (O_363,N_9974,N_9903);
and UO_364 (O_364,N_9974,N_9971);
nor UO_365 (O_365,N_9915,N_9913);
xnor UO_366 (O_366,N_9953,N_9959);
and UO_367 (O_367,N_9953,N_9902);
and UO_368 (O_368,N_9976,N_9910);
xor UO_369 (O_369,N_9998,N_9923);
xnor UO_370 (O_370,N_9993,N_9912);
and UO_371 (O_371,N_9977,N_9934);
xnor UO_372 (O_372,N_9997,N_9950);
or UO_373 (O_373,N_9934,N_9922);
and UO_374 (O_374,N_9959,N_9927);
or UO_375 (O_375,N_9942,N_9960);
and UO_376 (O_376,N_9992,N_9921);
xnor UO_377 (O_377,N_9955,N_9921);
xnor UO_378 (O_378,N_9910,N_9950);
and UO_379 (O_379,N_9965,N_9945);
nand UO_380 (O_380,N_9952,N_9928);
or UO_381 (O_381,N_9940,N_9917);
and UO_382 (O_382,N_9977,N_9987);
or UO_383 (O_383,N_9971,N_9970);
xnor UO_384 (O_384,N_9987,N_9991);
and UO_385 (O_385,N_9976,N_9966);
nand UO_386 (O_386,N_9917,N_9931);
nor UO_387 (O_387,N_9981,N_9951);
and UO_388 (O_388,N_9932,N_9958);
or UO_389 (O_389,N_9926,N_9933);
and UO_390 (O_390,N_9933,N_9944);
or UO_391 (O_391,N_9991,N_9900);
and UO_392 (O_392,N_9935,N_9944);
and UO_393 (O_393,N_9920,N_9981);
or UO_394 (O_394,N_9935,N_9917);
nand UO_395 (O_395,N_9973,N_9932);
or UO_396 (O_396,N_9981,N_9914);
nor UO_397 (O_397,N_9998,N_9919);
or UO_398 (O_398,N_9950,N_9928);
and UO_399 (O_399,N_9963,N_9965);
or UO_400 (O_400,N_9953,N_9906);
nor UO_401 (O_401,N_9937,N_9992);
xor UO_402 (O_402,N_9940,N_9942);
nand UO_403 (O_403,N_9917,N_9993);
or UO_404 (O_404,N_9976,N_9917);
or UO_405 (O_405,N_9908,N_9971);
xnor UO_406 (O_406,N_9949,N_9995);
and UO_407 (O_407,N_9938,N_9921);
or UO_408 (O_408,N_9951,N_9932);
or UO_409 (O_409,N_9979,N_9983);
nor UO_410 (O_410,N_9906,N_9901);
or UO_411 (O_411,N_9949,N_9939);
and UO_412 (O_412,N_9958,N_9931);
nor UO_413 (O_413,N_9958,N_9990);
and UO_414 (O_414,N_9955,N_9966);
nand UO_415 (O_415,N_9952,N_9989);
and UO_416 (O_416,N_9935,N_9922);
nor UO_417 (O_417,N_9939,N_9994);
nor UO_418 (O_418,N_9913,N_9943);
nor UO_419 (O_419,N_9943,N_9952);
or UO_420 (O_420,N_9962,N_9944);
xor UO_421 (O_421,N_9947,N_9937);
and UO_422 (O_422,N_9940,N_9950);
xor UO_423 (O_423,N_9972,N_9907);
nand UO_424 (O_424,N_9954,N_9910);
xor UO_425 (O_425,N_9935,N_9983);
xor UO_426 (O_426,N_9913,N_9992);
or UO_427 (O_427,N_9953,N_9926);
nor UO_428 (O_428,N_9975,N_9918);
and UO_429 (O_429,N_9948,N_9917);
or UO_430 (O_430,N_9929,N_9937);
or UO_431 (O_431,N_9916,N_9992);
nor UO_432 (O_432,N_9907,N_9949);
nor UO_433 (O_433,N_9930,N_9952);
nor UO_434 (O_434,N_9970,N_9943);
xnor UO_435 (O_435,N_9954,N_9934);
nand UO_436 (O_436,N_9996,N_9936);
and UO_437 (O_437,N_9942,N_9938);
nor UO_438 (O_438,N_9933,N_9987);
or UO_439 (O_439,N_9916,N_9999);
or UO_440 (O_440,N_9960,N_9941);
or UO_441 (O_441,N_9949,N_9903);
nand UO_442 (O_442,N_9942,N_9928);
or UO_443 (O_443,N_9931,N_9940);
nand UO_444 (O_444,N_9973,N_9997);
nand UO_445 (O_445,N_9952,N_9971);
or UO_446 (O_446,N_9943,N_9948);
nor UO_447 (O_447,N_9900,N_9933);
or UO_448 (O_448,N_9927,N_9980);
or UO_449 (O_449,N_9912,N_9916);
nor UO_450 (O_450,N_9978,N_9944);
and UO_451 (O_451,N_9948,N_9945);
nand UO_452 (O_452,N_9953,N_9976);
and UO_453 (O_453,N_9954,N_9965);
nor UO_454 (O_454,N_9949,N_9993);
or UO_455 (O_455,N_9992,N_9930);
nor UO_456 (O_456,N_9978,N_9991);
nand UO_457 (O_457,N_9963,N_9970);
and UO_458 (O_458,N_9958,N_9924);
or UO_459 (O_459,N_9981,N_9916);
xnor UO_460 (O_460,N_9999,N_9997);
and UO_461 (O_461,N_9976,N_9932);
nor UO_462 (O_462,N_9995,N_9982);
nor UO_463 (O_463,N_9957,N_9945);
xnor UO_464 (O_464,N_9940,N_9971);
or UO_465 (O_465,N_9994,N_9964);
nor UO_466 (O_466,N_9992,N_9923);
nand UO_467 (O_467,N_9950,N_9995);
nand UO_468 (O_468,N_9904,N_9939);
nand UO_469 (O_469,N_9936,N_9926);
nor UO_470 (O_470,N_9948,N_9915);
nor UO_471 (O_471,N_9957,N_9919);
or UO_472 (O_472,N_9937,N_9914);
nand UO_473 (O_473,N_9976,N_9998);
or UO_474 (O_474,N_9972,N_9940);
or UO_475 (O_475,N_9900,N_9911);
or UO_476 (O_476,N_9996,N_9980);
nand UO_477 (O_477,N_9955,N_9939);
nand UO_478 (O_478,N_9922,N_9994);
nor UO_479 (O_479,N_9942,N_9989);
or UO_480 (O_480,N_9920,N_9975);
nor UO_481 (O_481,N_9987,N_9937);
nand UO_482 (O_482,N_9938,N_9904);
nor UO_483 (O_483,N_9922,N_9975);
nand UO_484 (O_484,N_9903,N_9940);
xnor UO_485 (O_485,N_9994,N_9972);
nand UO_486 (O_486,N_9974,N_9914);
or UO_487 (O_487,N_9931,N_9956);
nand UO_488 (O_488,N_9994,N_9997);
or UO_489 (O_489,N_9963,N_9903);
xnor UO_490 (O_490,N_9980,N_9939);
nand UO_491 (O_491,N_9956,N_9979);
xor UO_492 (O_492,N_9925,N_9960);
or UO_493 (O_493,N_9910,N_9962);
nor UO_494 (O_494,N_9979,N_9914);
and UO_495 (O_495,N_9937,N_9968);
and UO_496 (O_496,N_9927,N_9922);
nand UO_497 (O_497,N_9919,N_9929);
nand UO_498 (O_498,N_9965,N_9929);
nor UO_499 (O_499,N_9949,N_9964);
nand UO_500 (O_500,N_9929,N_9909);
nand UO_501 (O_501,N_9938,N_9977);
nand UO_502 (O_502,N_9969,N_9981);
and UO_503 (O_503,N_9942,N_9996);
or UO_504 (O_504,N_9980,N_9917);
and UO_505 (O_505,N_9929,N_9991);
nor UO_506 (O_506,N_9944,N_9958);
nand UO_507 (O_507,N_9976,N_9999);
and UO_508 (O_508,N_9963,N_9962);
or UO_509 (O_509,N_9904,N_9916);
nor UO_510 (O_510,N_9915,N_9925);
nor UO_511 (O_511,N_9914,N_9918);
nand UO_512 (O_512,N_9931,N_9911);
and UO_513 (O_513,N_9933,N_9959);
or UO_514 (O_514,N_9911,N_9940);
nand UO_515 (O_515,N_9902,N_9973);
and UO_516 (O_516,N_9963,N_9920);
nor UO_517 (O_517,N_9968,N_9922);
xnor UO_518 (O_518,N_9988,N_9946);
nand UO_519 (O_519,N_9996,N_9966);
nor UO_520 (O_520,N_9929,N_9966);
or UO_521 (O_521,N_9970,N_9902);
and UO_522 (O_522,N_9924,N_9995);
and UO_523 (O_523,N_9957,N_9940);
nor UO_524 (O_524,N_9976,N_9925);
and UO_525 (O_525,N_9992,N_9920);
or UO_526 (O_526,N_9980,N_9905);
and UO_527 (O_527,N_9983,N_9920);
and UO_528 (O_528,N_9950,N_9998);
or UO_529 (O_529,N_9910,N_9959);
and UO_530 (O_530,N_9974,N_9940);
or UO_531 (O_531,N_9958,N_9926);
xor UO_532 (O_532,N_9937,N_9945);
or UO_533 (O_533,N_9914,N_9901);
and UO_534 (O_534,N_9949,N_9996);
and UO_535 (O_535,N_9997,N_9919);
or UO_536 (O_536,N_9925,N_9955);
xor UO_537 (O_537,N_9933,N_9903);
xor UO_538 (O_538,N_9975,N_9977);
nor UO_539 (O_539,N_9974,N_9965);
or UO_540 (O_540,N_9950,N_9992);
or UO_541 (O_541,N_9992,N_9956);
nand UO_542 (O_542,N_9963,N_9904);
and UO_543 (O_543,N_9948,N_9933);
or UO_544 (O_544,N_9960,N_9943);
xnor UO_545 (O_545,N_9999,N_9928);
or UO_546 (O_546,N_9906,N_9944);
or UO_547 (O_547,N_9966,N_9977);
nor UO_548 (O_548,N_9923,N_9981);
nor UO_549 (O_549,N_9972,N_9966);
nand UO_550 (O_550,N_9908,N_9925);
nand UO_551 (O_551,N_9908,N_9928);
nand UO_552 (O_552,N_9978,N_9909);
nand UO_553 (O_553,N_9957,N_9912);
or UO_554 (O_554,N_9950,N_9981);
or UO_555 (O_555,N_9913,N_9921);
or UO_556 (O_556,N_9953,N_9901);
nand UO_557 (O_557,N_9934,N_9910);
or UO_558 (O_558,N_9965,N_9991);
and UO_559 (O_559,N_9902,N_9948);
nor UO_560 (O_560,N_9932,N_9944);
nand UO_561 (O_561,N_9981,N_9947);
nand UO_562 (O_562,N_9990,N_9967);
nand UO_563 (O_563,N_9990,N_9998);
xor UO_564 (O_564,N_9944,N_9903);
nand UO_565 (O_565,N_9933,N_9963);
or UO_566 (O_566,N_9975,N_9991);
or UO_567 (O_567,N_9956,N_9991);
nor UO_568 (O_568,N_9999,N_9937);
nor UO_569 (O_569,N_9939,N_9925);
nand UO_570 (O_570,N_9979,N_9938);
nand UO_571 (O_571,N_9967,N_9908);
and UO_572 (O_572,N_9967,N_9929);
xor UO_573 (O_573,N_9968,N_9982);
nor UO_574 (O_574,N_9917,N_9991);
and UO_575 (O_575,N_9914,N_9973);
or UO_576 (O_576,N_9904,N_9991);
nand UO_577 (O_577,N_9962,N_9989);
or UO_578 (O_578,N_9968,N_9980);
nor UO_579 (O_579,N_9905,N_9930);
or UO_580 (O_580,N_9923,N_9938);
nand UO_581 (O_581,N_9942,N_9926);
nand UO_582 (O_582,N_9910,N_9923);
and UO_583 (O_583,N_9928,N_9977);
nand UO_584 (O_584,N_9940,N_9924);
nor UO_585 (O_585,N_9903,N_9938);
and UO_586 (O_586,N_9935,N_9926);
and UO_587 (O_587,N_9997,N_9908);
nand UO_588 (O_588,N_9996,N_9962);
nand UO_589 (O_589,N_9975,N_9905);
nor UO_590 (O_590,N_9927,N_9985);
nand UO_591 (O_591,N_9940,N_9937);
nor UO_592 (O_592,N_9976,N_9901);
xnor UO_593 (O_593,N_9923,N_9921);
or UO_594 (O_594,N_9916,N_9908);
nor UO_595 (O_595,N_9903,N_9906);
xor UO_596 (O_596,N_9991,N_9960);
or UO_597 (O_597,N_9996,N_9901);
nor UO_598 (O_598,N_9936,N_9904);
nor UO_599 (O_599,N_9928,N_9930);
nor UO_600 (O_600,N_9988,N_9989);
nor UO_601 (O_601,N_9977,N_9992);
or UO_602 (O_602,N_9976,N_9974);
or UO_603 (O_603,N_9927,N_9934);
and UO_604 (O_604,N_9900,N_9920);
or UO_605 (O_605,N_9905,N_9984);
nor UO_606 (O_606,N_9905,N_9913);
or UO_607 (O_607,N_9942,N_9964);
nor UO_608 (O_608,N_9910,N_9900);
or UO_609 (O_609,N_9940,N_9909);
and UO_610 (O_610,N_9909,N_9959);
and UO_611 (O_611,N_9969,N_9950);
or UO_612 (O_612,N_9998,N_9908);
xor UO_613 (O_613,N_9951,N_9940);
or UO_614 (O_614,N_9926,N_9947);
nor UO_615 (O_615,N_9986,N_9913);
and UO_616 (O_616,N_9940,N_9916);
and UO_617 (O_617,N_9973,N_9956);
xnor UO_618 (O_618,N_9988,N_9932);
and UO_619 (O_619,N_9998,N_9941);
or UO_620 (O_620,N_9997,N_9965);
or UO_621 (O_621,N_9913,N_9909);
nand UO_622 (O_622,N_9996,N_9939);
nor UO_623 (O_623,N_9962,N_9931);
or UO_624 (O_624,N_9927,N_9976);
and UO_625 (O_625,N_9911,N_9939);
and UO_626 (O_626,N_9975,N_9914);
or UO_627 (O_627,N_9964,N_9960);
nand UO_628 (O_628,N_9953,N_9908);
or UO_629 (O_629,N_9935,N_9977);
xor UO_630 (O_630,N_9943,N_9904);
nand UO_631 (O_631,N_9961,N_9910);
nor UO_632 (O_632,N_9906,N_9962);
xnor UO_633 (O_633,N_9912,N_9987);
nand UO_634 (O_634,N_9905,N_9956);
or UO_635 (O_635,N_9946,N_9977);
or UO_636 (O_636,N_9989,N_9959);
and UO_637 (O_637,N_9967,N_9937);
and UO_638 (O_638,N_9967,N_9999);
nor UO_639 (O_639,N_9920,N_9922);
xor UO_640 (O_640,N_9944,N_9938);
xnor UO_641 (O_641,N_9908,N_9972);
or UO_642 (O_642,N_9974,N_9991);
or UO_643 (O_643,N_9966,N_9986);
and UO_644 (O_644,N_9939,N_9984);
and UO_645 (O_645,N_9967,N_9921);
xnor UO_646 (O_646,N_9900,N_9908);
nor UO_647 (O_647,N_9950,N_9902);
nand UO_648 (O_648,N_9998,N_9945);
or UO_649 (O_649,N_9994,N_9951);
or UO_650 (O_650,N_9963,N_9981);
or UO_651 (O_651,N_9923,N_9954);
or UO_652 (O_652,N_9948,N_9989);
nand UO_653 (O_653,N_9953,N_9980);
and UO_654 (O_654,N_9967,N_9900);
nor UO_655 (O_655,N_9975,N_9936);
or UO_656 (O_656,N_9914,N_9939);
xnor UO_657 (O_657,N_9917,N_9927);
nand UO_658 (O_658,N_9982,N_9908);
xor UO_659 (O_659,N_9902,N_9994);
and UO_660 (O_660,N_9945,N_9930);
xor UO_661 (O_661,N_9938,N_9936);
or UO_662 (O_662,N_9983,N_9968);
nand UO_663 (O_663,N_9979,N_9945);
nor UO_664 (O_664,N_9931,N_9986);
xnor UO_665 (O_665,N_9913,N_9972);
nand UO_666 (O_666,N_9915,N_9943);
and UO_667 (O_667,N_9920,N_9970);
and UO_668 (O_668,N_9955,N_9963);
and UO_669 (O_669,N_9913,N_9978);
nor UO_670 (O_670,N_9979,N_9993);
xor UO_671 (O_671,N_9951,N_9933);
nor UO_672 (O_672,N_9969,N_9954);
xnor UO_673 (O_673,N_9957,N_9933);
nand UO_674 (O_674,N_9951,N_9942);
or UO_675 (O_675,N_9968,N_9962);
or UO_676 (O_676,N_9956,N_9901);
xnor UO_677 (O_677,N_9958,N_9920);
and UO_678 (O_678,N_9922,N_9908);
nor UO_679 (O_679,N_9995,N_9925);
and UO_680 (O_680,N_9995,N_9937);
nor UO_681 (O_681,N_9926,N_9950);
or UO_682 (O_682,N_9926,N_9966);
and UO_683 (O_683,N_9910,N_9928);
nor UO_684 (O_684,N_9959,N_9956);
and UO_685 (O_685,N_9915,N_9936);
nand UO_686 (O_686,N_9958,N_9927);
or UO_687 (O_687,N_9920,N_9973);
and UO_688 (O_688,N_9949,N_9978);
nand UO_689 (O_689,N_9928,N_9955);
nor UO_690 (O_690,N_9936,N_9985);
xnor UO_691 (O_691,N_9904,N_9979);
nor UO_692 (O_692,N_9985,N_9917);
xnor UO_693 (O_693,N_9927,N_9939);
and UO_694 (O_694,N_9906,N_9942);
and UO_695 (O_695,N_9925,N_9987);
and UO_696 (O_696,N_9945,N_9973);
nand UO_697 (O_697,N_9944,N_9925);
nor UO_698 (O_698,N_9999,N_9952);
or UO_699 (O_699,N_9901,N_9990);
or UO_700 (O_700,N_9923,N_9941);
nor UO_701 (O_701,N_9919,N_9923);
or UO_702 (O_702,N_9988,N_9928);
and UO_703 (O_703,N_9988,N_9904);
or UO_704 (O_704,N_9999,N_9932);
or UO_705 (O_705,N_9917,N_9969);
nor UO_706 (O_706,N_9927,N_9931);
and UO_707 (O_707,N_9961,N_9946);
and UO_708 (O_708,N_9902,N_9934);
nand UO_709 (O_709,N_9985,N_9922);
and UO_710 (O_710,N_9933,N_9931);
or UO_711 (O_711,N_9992,N_9957);
and UO_712 (O_712,N_9995,N_9991);
nand UO_713 (O_713,N_9945,N_9982);
nand UO_714 (O_714,N_9917,N_9926);
xnor UO_715 (O_715,N_9993,N_9968);
or UO_716 (O_716,N_9935,N_9909);
and UO_717 (O_717,N_9918,N_9999);
nand UO_718 (O_718,N_9942,N_9986);
xor UO_719 (O_719,N_9965,N_9985);
or UO_720 (O_720,N_9986,N_9923);
xor UO_721 (O_721,N_9932,N_9961);
or UO_722 (O_722,N_9921,N_9993);
nand UO_723 (O_723,N_9928,N_9967);
or UO_724 (O_724,N_9956,N_9940);
and UO_725 (O_725,N_9934,N_9900);
and UO_726 (O_726,N_9989,N_9993);
nor UO_727 (O_727,N_9904,N_9978);
or UO_728 (O_728,N_9950,N_9978);
or UO_729 (O_729,N_9981,N_9958);
and UO_730 (O_730,N_9951,N_9961);
and UO_731 (O_731,N_9955,N_9977);
nor UO_732 (O_732,N_9932,N_9980);
or UO_733 (O_733,N_9978,N_9947);
or UO_734 (O_734,N_9909,N_9941);
xor UO_735 (O_735,N_9939,N_9909);
or UO_736 (O_736,N_9937,N_9902);
xnor UO_737 (O_737,N_9978,N_9925);
xnor UO_738 (O_738,N_9953,N_9966);
and UO_739 (O_739,N_9903,N_9988);
nor UO_740 (O_740,N_9963,N_9913);
and UO_741 (O_741,N_9951,N_9914);
xor UO_742 (O_742,N_9999,N_9958);
nand UO_743 (O_743,N_9945,N_9995);
xor UO_744 (O_744,N_9994,N_9974);
nor UO_745 (O_745,N_9964,N_9977);
nor UO_746 (O_746,N_9990,N_9971);
nand UO_747 (O_747,N_9903,N_9919);
xnor UO_748 (O_748,N_9951,N_9985);
and UO_749 (O_749,N_9928,N_9927);
xor UO_750 (O_750,N_9951,N_9972);
or UO_751 (O_751,N_9949,N_9958);
and UO_752 (O_752,N_9977,N_9990);
and UO_753 (O_753,N_9941,N_9948);
nand UO_754 (O_754,N_9961,N_9999);
nand UO_755 (O_755,N_9942,N_9962);
nor UO_756 (O_756,N_9979,N_9988);
or UO_757 (O_757,N_9902,N_9992);
nand UO_758 (O_758,N_9908,N_9935);
and UO_759 (O_759,N_9989,N_9947);
xor UO_760 (O_760,N_9964,N_9932);
or UO_761 (O_761,N_9905,N_9944);
nand UO_762 (O_762,N_9906,N_9919);
or UO_763 (O_763,N_9939,N_9990);
nand UO_764 (O_764,N_9933,N_9979);
nor UO_765 (O_765,N_9912,N_9991);
or UO_766 (O_766,N_9926,N_9973);
nand UO_767 (O_767,N_9943,N_9951);
or UO_768 (O_768,N_9909,N_9919);
and UO_769 (O_769,N_9993,N_9935);
xor UO_770 (O_770,N_9988,N_9959);
xnor UO_771 (O_771,N_9983,N_9917);
nand UO_772 (O_772,N_9998,N_9943);
and UO_773 (O_773,N_9915,N_9999);
xnor UO_774 (O_774,N_9980,N_9937);
and UO_775 (O_775,N_9974,N_9943);
or UO_776 (O_776,N_9939,N_9960);
or UO_777 (O_777,N_9939,N_9915);
and UO_778 (O_778,N_9990,N_9997);
or UO_779 (O_779,N_9933,N_9907);
nand UO_780 (O_780,N_9915,N_9989);
and UO_781 (O_781,N_9987,N_9970);
or UO_782 (O_782,N_9951,N_9937);
and UO_783 (O_783,N_9917,N_9909);
and UO_784 (O_784,N_9917,N_9974);
xor UO_785 (O_785,N_9968,N_9961);
or UO_786 (O_786,N_9935,N_9966);
and UO_787 (O_787,N_9942,N_9987);
nand UO_788 (O_788,N_9994,N_9925);
nand UO_789 (O_789,N_9935,N_9995);
nand UO_790 (O_790,N_9900,N_9929);
and UO_791 (O_791,N_9995,N_9953);
nand UO_792 (O_792,N_9930,N_9973);
nor UO_793 (O_793,N_9975,N_9998);
nand UO_794 (O_794,N_9955,N_9995);
and UO_795 (O_795,N_9906,N_9955);
nand UO_796 (O_796,N_9966,N_9997);
nor UO_797 (O_797,N_9993,N_9940);
nand UO_798 (O_798,N_9932,N_9963);
and UO_799 (O_799,N_9994,N_9909);
nand UO_800 (O_800,N_9910,N_9975);
nor UO_801 (O_801,N_9960,N_9935);
nor UO_802 (O_802,N_9976,N_9962);
nand UO_803 (O_803,N_9971,N_9936);
nor UO_804 (O_804,N_9915,N_9967);
and UO_805 (O_805,N_9952,N_9937);
nand UO_806 (O_806,N_9985,N_9932);
nand UO_807 (O_807,N_9970,N_9919);
nor UO_808 (O_808,N_9931,N_9991);
or UO_809 (O_809,N_9980,N_9985);
or UO_810 (O_810,N_9921,N_9964);
or UO_811 (O_811,N_9992,N_9985);
or UO_812 (O_812,N_9958,N_9955);
or UO_813 (O_813,N_9968,N_9925);
and UO_814 (O_814,N_9945,N_9928);
xnor UO_815 (O_815,N_9906,N_9914);
or UO_816 (O_816,N_9990,N_9970);
or UO_817 (O_817,N_9952,N_9960);
nor UO_818 (O_818,N_9970,N_9923);
or UO_819 (O_819,N_9900,N_9999);
and UO_820 (O_820,N_9907,N_9903);
nor UO_821 (O_821,N_9907,N_9909);
and UO_822 (O_822,N_9951,N_9958);
nor UO_823 (O_823,N_9909,N_9960);
xor UO_824 (O_824,N_9928,N_9979);
nor UO_825 (O_825,N_9938,N_9941);
nand UO_826 (O_826,N_9962,N_9927);
and UO_827 (O_827,N_9968,N_9910);
and UO_828 (O_828,N_9987,N_9985);
xor UO_829 (O_829,N_9942,N_9978);
nor UO_830 (O_830,N_9924,N_9964);
xor UO_831 (O_831,N_9983,N_9957);
or UO_832 (O_832,N_9936,N_9982);
and UO_833 (O_833,N_9949,N_9933);
or UO_834 (O_834,N_9995,N_9942);
or UO_835 (O_835,N_9938,N_9957);
xor UO_836 (O_836,N_9922,N_9938);
or UO_837 (O_837,N_9995,N_9918);
or UO_838 (O_838,N_9911,N_9968);
or UO_839 (O_839,N_9964,N_9916);
or UO_840 (O_840,N_9941,N_9908);
xor UO_841 (O_841,N_9912,N_9909);
nor UO_842 (O_842,N_9902,N_9957);
nand UO_843 (O_843,N_9900,N_9941);
nor UO_844 (O_844,N_9922,N_9987);
or UO_845 (O_845,N_9904,N_9960);
nor UO_846 (O_846,N_9952,N_9924);
nor UO_847 (O_847,N_9906,N_9920);
nor UO_848 (O_848,N_9952,N_9966);
nand UO_849 (O_849,N_9971,N_9942);
or UO_850 (O_850,N_9988,N_9950);
or UO_851 (O_851,N_9995,N_9940);
nand UO_852 (O_852,N_9954,N_9996);
or UO_853 (O_853,N_9991,N_9907);
nor UO_854 (O_854,N_9940,N_9918);
nor UO_855 (O_855,N_9998,N_9955);
and UO_856 (O_856,N_9979,N_9943);
and UO_857 (O_857,N_9992,N_9938);
or UO_858 (O_858,N_9920,N_9921);
or UO_859 (O_859,N_9943,N_9936);
xnor UO_860 (O_860,N_9905,N_9992);
nor UO_861 (O_861,N_9962,N_9900);
nand UO_862 (O_862,N_9985,N_9947);
nor UO_863 (O_863,N_9920,N_9951);
nand UO_864 (O_864,N_9912,N_9922);
nand UO_865 (O_865,N_9951,N_9959);
or UO_866 (O_866,N_9972,N_9978);
nand UO_867 (O_867,N_9906,N_9902);
nor UO_868 (O_868,N_9953,N_9998);
nor UO_869 (O_869,N_9952,N_9997);
nor UO_870 (O_870,N_9935,N_9902);
or UO_871 (O_871,N_9929,N_9974);
xor UO_872 (O_872,N_9971,N_9916);
nor UO_873 (O_873,N_9968,N_9959);
and UO_874 (O_874,N_9933,N_9928);
nor UO_875 (O_875,N_9942,N_9914);
nand UO_876 (O_876,N_9950,N_9911);
or UO_877 (O_877,N_9993,N_9999);
nand UO_878 (O_878,N_9973,N_9916);
nand UO_879 (O_879,N_9980,N_9959);
nor UO_880 (O_880,N_9976,N_9940);
nor UO_881 (O_881,N_9906,N_9925);
nand UO_882 (O_882,N_9949,N_9921);
and UO_883 (O_883,N_9972,N_9976);
and UO_884 (O_884,N_9900,N_9948);
or UO_885 (O_885,N_9998,N_9915);
nor UO_886 (O_886,N_9929,N_9955);
xnor UO_887 (O_887,N_9960,N_9950);
and UO_888 (O_888,N_9940,N_9986);
nand UO_889 (O_889,N_9933,N_9940);
or UO_890 (O_890,N_9999,N_9965);
or UO_891 (O_891,N_9983,N_9987);
and UO_892 (O_892,N_9988,N_9982);
xnor UO_893 (O_893,N_9932,N_9943);
or UO_894 (O_894,N_9914,N_9962);
nor UO_895 (O_895,N_9938,N_9916);
xnor UO_896 (O_896,N_9999,N_9953);
or UO_897 (O_897,N_9917,N_9956);
or UO_898 (O_898,N_9937,N_9939);
nand UO_899 (O_899,N_9973,N_9985);
nor UO_900 (O_900,N_9969,N_9988);
or UO_901 (O_901,N_9952,N_9942);
and UO_902 (O_902,N_9907,N_9986);
nand UO_903 (O_903,N_9915,N_9972);
or UO_904 (O_904,N_9917,N_9951);
nor UO_905 (O_905,N_9976,N_9952);
xnor UO_906 (O_906,N_9976,N_9950);
nand UO_907 (O_907,N_9931,N_9902);
nor UO_908 (O_908,N_9958,N_9917);
or UO_909 (O_909,N_9991,N_9970);
and UO_910 (O_910,N_9996,N_9906);
nand UO_911 (O_911,N_9926,N_9916);
or UO_912 (O_912,N_9951,N_9945);
nor UO_913 (O_913,N_9991,N_9924);
nor UO_914 (O_914,N_9967,N_9968);
nor UO_915 (O_915,N_9960,N_9967);
or UO_916 (O_916,N_9947,N_9942);
or UO_917 (O_917,N_9972,N_9952);
or UO_918 (O_918,N_9955,N_9975);
or UO_919 (O_919,N_9926,N_9902);
or UO_920 (O_920,N_9971,N_9943);
xor UO_921 (O_921,N_9913,N_9900);
and UO_922 (O_922,N_9901,N_9947);
or UO_923 (O_923,N_9981,N_9956);
or UO_924 (O_924,N_9950,N_9903);
and UO_925 (O_925,N_9961,N_9921);
nand UO_926 (O_926,N_9967,N_9918);
xnor UO_927 (O_927,N_9967,N_9942);
and UO_928 (O_928,N_9953,N_9907);
xor UO_929 (O_929,N_9948,N_9901);
and UO_930 (O_930,N_9921,N_9932);
xnor UO_931 (O_931,N_9921,N_9906);
or UO_932 (O_932,N_9943,N_9944);
nor UO_933 (O_933,N_9983,N_9937);
and UO_934 (O_934,N_9954,N_9909);
and UO_935 (O_935,N_9932,N_9930);
and UO_936 (O_936,N_9925,N_9980);
or UO_937 (O_937,N_9919,N_9944);
nand UO_938 (O_938,N_9960,N_9957);
or UO_939 (O_939,N_9989,N_9980);
nand UO_940 (O_940,N_9994,N_9961);
nor UO_941 (O_941,N_9951,N_9934);
or UO_942 (O_942,N_9998,N_9958);
and UO_943 (O_943,N_9902,N_9914);
nor UO_944 (O_944,N_9966,N_9919);
and UO_945 (O_945,N_9911,N_9970);
nand UO_946 (O_946,N_9993,N_9908);
or UO_947 (O_947,N_9956,N_9929);
nand UO_948 (O_948,N_9996,N_9941);
or UO_949 (O_949,N_9963,N_9993);
nand UO_950 (O_950,N_9930,N_9903);
nor UO_951 (O_951,N_9960,N_9948);
nand UO_952 (O_952,N_9954,N_9997);
xor UO_953 (O_953,N_9923,N_9932);
nor UO_954 (O_954,N_9985,N_9914);
and UO_955 (O_955,N_9959,N_9928);
nand UO_956 (O_956,N_9998,N_9916);
or UO_957 (O_957,N_9935,N_9968);
nand UO_958 (O_958,N_9942,N_9911);
nor UO_959 (O_959,N_9934,N_9999);
xor UO_960 (O_960,N_9986,N_9935);
xor UO_961 (O_961,N_9983,N_9981);
nand UO_962 (O_962,N_9902,N_9912);
and UO_963 (O_963,N_9918,N_9904);
nand UO_964 (O_964,N_9978,N_9906);
nor UO_965 (O_965,N_9930,N_9998);
or UO_966 (O_966,N_9930,N_9906);
or UO_967 (O_967,N_9956,N_9972);
and UO_968 (O_968,N_9947,N_9967);
and UO_969 (O_969,N_9970,N_9980);
or UO_970 (O_970,N_9948,N_9978);
or UO_971 (O_971,N_9977,N_9922);
or UO_972 (O_972,N_9968,N_9944);
nand UO_973 (O_973,N_9977,N_9961);
and UO_974 (O_974,N_9913,N_9902);
or UO_975 (O_975,N_9988,N_9922);
and UO_976 (O_976,N_9989,N_9975);
nor UO_977 (O_977,N_9904,N_9915);
nor UO_978 (O_978,N_9912,N_9979);
nand UO_979 (O_979,N_9904,N_9958);
or UO_980 (O_980,N_9913,N_9993);
nand UO_981 (O_981,N_9921,N_9901);
or UO_982 (O_982,N_9929,N_9983);
nor UO_983 (O_983,N_9982,N_9984);
nor UO_984 (O_984,N_9904,N_9933);
nand UO_985 (O_985,N_9923,N_9922);
nor UO_986 (O_986,N_9967,N_9982);
xor UO_987 (O_987,N_9908,N_9954);
nand UO_988 (O_988,N_9911,N_9953);
or UO_989 (O_989,N_9928,N_9916);
nor UO_990 (O_990,N_9926,N_9974);
nand UO_991 (O_991,N_9926,N_9918);
or UO_992 (O_992,N_9967,N_9945);
or UO_993 (O_993,N_9950,N_9999);
and UO_994 (O_994,N_9920,N_9929);
nor UO_995 (O_995,N_9970,N_9999);
nand UO_996 (O_996,N_9983,N_9926);
or UO_997 (O_997,N_9964,N_9938);
nand UO_998 (O_998,N_9987,N_9928);
or UO_999 (O_999,N_9921,N_9981);
nor UO_1000 (O_1000,N_9908,N_9988);
and UO_1001 (O_1001,N_9966,N_9998);
and UO_1002 (O_1002,N_9958,N_9970);
xnor UO_1003 (O_1003,N_9906,N_9980);
and UO_1004 (O_1004,N_9971,N_9995);
xnor UO_1005 (O_1005,N_9935,N_9921);
nor UO_1006 (O_1006,N_9981,N_9985);
nor UO_1007 (O_1007,N_9999,N_9978);
xor UO_1008 (O_1008,N_9996,N_9945);
xnor UO_1009 (O_1009,N_9998,N_9947);
nor UO_1010 (O_1010,N_9944,N_9949);
nor UO_1011 (O_1011,N_9934,N_9916);
nand UO_1012 (O_1012,N_9953,N_9967);
or UO_1013 (O_1013,N_9907,N_9919);
or UO_1014 (O_1014,N_9970,N_9936);
and UO_1015 (O_1015,N_9914,N_9923);
nand UO_1016 (O_1016,N_9967,N_9944);
or UO_1017 (O_1017,N_9983,N_9984);
or UO_1018 (O_1018,N_9928,N_9939);
nand UO_1019 (O_1019,N_9985,N_9997);
or UO_1020 (O_1020,N_9907,N_9982);
nor UO_1021 (O_1021,N_9959,N_9936);
nor UO_1022 (O_1022,N_9982,N_9953);
or UO_1023 (O_1023,N_9999,N_9939);
nand UO_1024 (O_1024,N_9947,N_9903);
nand UO_1025 (O_1025,N_9927,N_9932);
nor UO_1026 (O_1026,N_9935,N_9949);
or UO_1027 (O_1027,N_9918,N_9931);
xnor UO_1028 (O_1028,N_9987,N_9962);
or UO_1029 (O_1029,N_9946,N_9956);
xor UO_1030 (O_1030,N_9931,N_9963);
nand UO_1031 (O_1031,N_9964,N_9928);
nand UO_1032 (O_1032,N_9949,N_9983);
nor UO_1033 (O_1033,N_9971,N_9994);
xnor UO_1034 (O_1034,N_9958,N_9936);
and UO_1035 (O_1035,N_9907,N_9915);
xor UO_1036 (O_1036,N_9992,N_9963);
and UO_1037 (O_1037,N_9956,N_9995);
and UO_1038 (O_1038,N_9923,N_9943);
and UO_1039 (O_1039,N_9923,N_9946);
or UO_1040 (O_1040,N_9902,N_9964);
or UO_1041 (O_1041,N_9950,N_9958);
and UO_1042 (O_1042,N_9971,N_9986);
nor UO_1043 (O_1043,N_9932,N_9970);
nor UO_1044 (O_1044,N_9917,N_9929);
and UO_1045 (O_1045,N_9972,N_9997);
and UO_1046 (O_1046,N_9954,N_9945);
nand UO_1047 (O_1047,N_9918,N_9996);
nand UO_1048 (O_1048,N_9968,N_9901);
nor UO_1049 (O_1049,N_9904,N_9917);
nand UO_1050 (O_1050,N_9933,N_9913);
nor UO_1051 (O_1051,N_9982,N_9915);
nand UO_1052 (O_1052,N_9946,N_9980);
xor UO_1053 (O_1053,N_9972,N_9987);
or UO_1054 (O_1054,N_9994,N_9931);
xor UO_1055 (O_1055,N_9921,N_9985);
nand UO_1056 (O_1056,N_9946,N_9931);
nor UO_1057 (O_1057,N_9977,N_9991);
nand UO_1058 (O_1058,N_9916,N_9902);
nor UO_1059 (O_1059,N_9920,N_9923);
or UO_1060 (O_1060,N_9928,N_9914);
nor UO_1061 (O_1061,N_9918,N_9988);
or UO_1062 (O_1062,N_9937,N_9921);
and UO_1063 (O_1063,N_9960,N_9976);
xor UO_1064 (O_1064,N_9950,N_9972);
and UO_1065 (O_1065,N_9969,N_9938);
nor UO_1066 (O_1066,N_9936,N_9989);
nand UO_1067 (O_1067,N_9939,N_9989);
xnor UO_1068 (O_1068,N_9913,N_9904);
nor UO_1069 (O_1069,N_9946,N_9924);
nand UO_1070 (O_1070,N_9953,N_9933);
nor UO_1071 (O_1071,N_9918,N_9960);
nand UO_1072 (O_1072,N_9951,N_9993);
nor UO_1073 (O_1073,N_9989,N_9963);
and UO_1074 (O_1074,N_9951,N_9901);
nand UO_1075 (O_1075,N_9972,N_9990);
or UO_1076 (O_1076,N_9976,N_9931);
or UO_1077 (O_1077,N_9939,N_9985);
and UO_1078 (O_1078,N_9938,N_9945);
nand UO_1079 (O_1079,N_9957,N_9941);
nand UO_1080 (O_1080,N_9936,N_9956);
nand UO_1081 (O_1081,N_9986,N_9996);
or UO_1082 (O_1082,N_9950,N_9930);
and UO_1083 (O_1083,N_9969,N_9909);
xnor UO_1084 (O_1084,N_9959,N_9912);
and UO_1085 (O_1085,N_9976,N_9955);
and UO_1086 (O_1086,N_9958,N_9956);
nor UO_1087 (O_1087,N_9999,N_9920);
and UO_1088 (O_1088,N_9930,N_9935);
nand UO_1089 (O_1089,N_9951,N_9949);
nand UO_1090 (O_1090,N_9979,N_9987);
and UO_1091 (O_1091,N_9911,N_9903);
nand UO_1092 (O_1092,N_9909,N_9981);
or UO_1093 (O_1093,N_9914,N_9938);
xnor UO_1094 (O_1094,N_9940,N_9984);
nor UO_1095 (O_1095,N_9997,N_9920);
nand UO_1096 (O_1096,N_9939,N_9941);
nand UO_1097 (O_1097,N_9949,N_9966);
or UO_1098 (O_1098,N_9972,N_9939);
or UO_1099 (O_1099,N_9991,N_9916);
and UO_1100 (O_1100,N_9916,N_9989);
nand UO_1101 (O_1101,N_9953,N_9955);
or UO_1102 (O_1102,N_9931,N_9983);
xnor UO_1103 (O_1103,N_9977,N_9988);
or UO_1104 (O_1104,N_9927,N_9936);
nor UO_1105 (O_1105,N_9968,N_9954);
nand UO_1106 (O_1106,N_9956,N_9918);
nand UO_1107 (O_1107,N_9909,N_9930);
and UO_1108 (O_1108,N_9994,N_9927);
or UO_1109 (O_1109,N_9989,N_9943);
or UO_1110 (O_1110,N_9922,N_9940);
nor UO_1111 (O_1111,N_9923,N_9978);
nand UO_1112 (O_1112,N_9921,N_9954);
nor UO_1113 (O_1113,N_9922,N_9952);
xor UO_1114 (O_1114,N_9954,N_9979);
or UO_1115 (O_1115,N_9995,N_9926);
or UO_1116 (O_1116,N_9936,N_9910);
or UO_1117 (O_1117,N_9922,N_9948);
and UO_1118 (O_1118,N_9961,N_9982);
xnor UO_1119 (O_1119,N_9974,N_9907);
nand UO_1120 (O_1120,N_9919,N_9942);
nand UO_1121 (O_1121,N_9964,N_9962);
or UO_1122 (O_1122,N_9953,N_9963);
and UO_1123 (O_1123,N_9985,N_9900);
or UO_1124 (O_1124,N_9925,N_9938);
nand UO_1125 (O_1125,N_9987,N_9917);
or UO_1126 (O_1126,N_9999,N_9990);
xor UO_1127 (O_1127,N_9986,N_9910);
nand UO_1128 (O_1128,N_9955,N_9983);
nand UO_1129 (O_1129,N_9922,N_9959);
xor UO_1130 (O_1130,N_9987,N_9954);
nor UO_1131 (O_1131,N_9932,N_9974);
or UO_1132 (O_1132,N_9950,N_9974);
or UO_1133 (O_1133,N_9926,N_9961);
and UO_1134 (O_1134,N_9929,N_9975);
or UO_1135 (O_1135,N_9967,N_9950);
nand UO_1136 (O_1136,N_9902,N_9974);
nor UO_1137 (O_1137,N_9992,N_9965);
and UO_1138 (O_1138,N_9943,N_9964);
and UO_1139 (O_1139,N_9926,N_9985);
nand UO_1140 (O_1140,N_9954,N_9957);
and UO_1141 (O_1141,N_9926,N_9955);
or UO_1142 (O_1142,N_9966,N_9959);
and UO_1143 (O_1143,N_9963,N_9969);
nor UO_1144 (O_1144,N_9949,N_9950);
or UO_1145 (O_1145,N_9925,N_9996);
or UO_1146 (O_1146,N_9960,N_9930);
nor UO_1147 (O_1147,N_9969,N_9940);
nor UO_1148 (O_1148,N_9940,N_9980);
and UO_1149 (O_1149,N_9967,N_9911);
or UO_1150 (O_1150,N_9905,N_9929);
nor UO_1151 (O_1151,N_9944,N_9988);
and UO_1152 (O_1152,N_9936,N_9984);
and UO_1153 (O_1153,N_9944,N_9987);
and UO_1154 (O_1154,N_9907,N_9973);
nand UO_1155 (O_1155,N_9932,N_9904);
and UO_1156 (O_1156,N_9949,N_9991);
nor UO_1157 (O_1157,N_9996,N_9946);
xor UO_1158 (O_1158,N_9923,N_9944);
and UO_1159 (O_1159,N_9953,N_9939);
or UO_1160 (O_1160,N_9948,N_9934);
nand UO_1161 (O_1161,N_9910,N_9993);
xor UO_1162 (O_1162,N_9948,N_9950);
or UO_1163 (O_1163,N_9961,N_9980);
and UO_1164 (O_1164,N_9962,N_9958);
or UO_1165 (O_1165,N_9919,N_9905);
and UO_1166 (O_1166,N_9970,N_9964);
xnor UO_1167 (O_1167,N_9941,N_9967);
nand UO_1168 (O_1168,N_9974,N_9904);
nor UO_1169 (O_1169,N_9929,N_9985);
nor UO_1170 (O_1170,N_9966,N_9938);
nand UO_1171 (O_1171,N_9966,N_9956);
xnor UO_1172 (O_1172,N_9900,N_9946);
or UO_1173 (O_1173,N_9980,N_9986);
nor UO_1174 (O_1174,N_9991,N_9939);
nor UO_1175 (O_1175,N_9965,N_9972);
nor UO_1176 (O_1176,N_9924,N_9949);
nand UO_1177 (O_1177,N_9912,N_9933);
xnor UO_1178 (O_1178,N_9947,N_9936);
nor UO_1179 (O_1179,N_9915,N_9988);
or UO_1180 (O_1180,N_9974,N_9913);
and UO_1181 (O_1181,N_9943,N_9966);
nand UO_1182 (O_1182,N_9940,N_9968);
or UO_1183 (O_1183,N_9938,N_9973);
nor UO_1184 (O_1184,N_9994,N_9947);
nor UO_1185 (O_1185,N_9924,N_9957);
nand UO_1186 (O_1186,N_9947,N_9931);
and UO_1187 (O_1187,N_9950,N_9922);
or UO_1188 (O_1188,N_9924,N_9921);
xor UO_1189 (O_1189,N_9966,N_9910);
and UO_1190 (O_1190,N_9996,N_9917);
nor UO_1191 (O_1191,N_9936,N_9960);
nand UO_1192 (O_1192,N_9919,N_9921);
nor UO_1193 (O_1193,N_9920,N_9955);
nand UO_1194 (O_1194,N_9945,N_9911);
nand UO_1195 (O_1195,N_9954,N_9986);
xor UO_1196 (O_1196,N_9996,N_9931);
and UO_1197 (O_1197,N_9936,N_9924);
nor UO_1198 (O_1198,N_9910,N_9917);
and UO_1199 (O_1199,N_9903,N_9935);
and UO_1200 (O_1200,N_9918,N_9954);
or UO_1201 (O_1201,N_9995,N_9907);
or UO_1202 (O_1202,N_9918,N_9909);
nand UO_1203 (O_1203,N_9985,N_9905);
and UO_1204 (O_1204,N_9918,N_9983);
or UO_1205 (O_1205,N_9901,N_9993);
nand UO_1206 (O_1206,N_9936,N_9976);
or UO_1207 (O_1207,N_9901,N_9991);
and UO_1208 (O_1208,N_9951,N_9941);
nor UO_1209 (O_1209,N_9916,N_9923);
nand UO_1210 (O_1210,N_9946,N_9937);
nand UO_1211 (O_1211,N_9905,N_9960);
xnor UO_1212 (O_1212,N_9949,N_9988);
and UO_1213 (O_1213,N_9930,N_9995);
and UO_1214 (O_1214,N_9978,N_9967);
nor UO_1215 (O_1215,N_9930,N_9942);
nor UO_1216 (O_1216,N_9923,N_9918);
or UO_1217 (O_1217,N_9913,N_9946);
and UO_1218 (O_1218,N_9937,N_9928);
or UO_1219 (O_1219,N_9915,N_9935);
or UO_1220 (O_1220,N_9982,N_9970);
and UO_1221 (O_1221,N_9928,N_9972);
nand UO_1222 (O_1222,N_9938,N_9963);
nand UO_1223 (O_1223,N_9908,N_9956);
nand UO_1224 (O_1224,N_9927,N_9955);
xnor UO_1225 (O_1225,N_9912,N_9906);
and UO_1226 (O_1226,N_9935,N_9961);
or UO_1227 (O_1227,N_9923,N_9976);
nor UO_1228 (O_1228,N_9955,N_9900);
or UO_1229 (O_1229,N_9909,N_9922);
or UO_1230 (O_1230,N_9941,N_9933);
nor UO_1231 (O_1231,N_9967,N_9902);
and UO_1232 (O_1232,N_9954,N_9926);
or UO_1233 (O_1233,N_9976,N_9954);
xnor UO_1234 (O_1234,N_9958,N_9971);
and UO_1235 (O_1235,N_9907,N_9993);
nor UO_1236 (O_1236,N_9909,N_9977);
or UO_1237 (O_1237,N_9965,N_9935);
xor UO_1238 (O_1238,N_9943,N_9914);
or UO_1239 (O_1239,N_9912,N_9983);
and UO_1240 (O_1240,N_9975,N_9916);
nor UO_1241 (O_1241,N_9926,N_9978);
and UO_1242 (O_1242,N_9999,N_9914);
or UO_1243 (O_1243,N_9951,N_9971);
xor UO_1244 (O_1244,N_9970,N_9939);
xor UO_1245 (O_1245,N_9911,N_9983);
or UO_1246 (O_1246,N_9920,N_9936);
nand UO_1247 (O_1247,N_9945,N_9919);
nand UO_1248 (O_1248,N_9950,N_9921);
nor UO_1249 (O_1249,N_9911,N_9965);
nand UO_1250 (O_1250,N_9992,N_9926);
nand UO_1251 (O_1251,N_9992,N_9931);
nor UO_1252 (O_1252,N_9997,N_9993);
and UO_1253 (O_1253,N_9936,N_9922);
or UO_1254 (O_1254,N_9933,N_9984);
or UO_1255 (O_1255,N_9942,N_9990);
nor UO_1256 (O_1256,N_9996,N_9912);
or UO_1257 (O_1257,N_9964,N_9901);
nand UO_1258 (O_1258,N_9960,N_9958);
nand UO_1259 (O_1259,N_9912,N_9915);
or UO_1260 (O_1260,N_9963,N_9901);
nand UO_1261 (O_1261,N_9906,N_9960);
xor UO_1262 (O_1262,N_9993,N_9980);
or UO_1263 (O_1263,N_9960,N_9962);
nor UO_1264 (O_1264,N_9970,N_9930);
xnor UO_1265 (O_1265,N_9955,N_9961);
or UO_1266 (O_1266,N_9986,N_9950);
nor UO_1267 (O_1267,N_9974,N_9948);
and UO_1268 (O_1268,N_9958,N_9909);
nor UO_1269 (O_1269,N_9976,N_9991);
xor UO_1270 (O_1270,N_9903,N_9979);
or UO_1271 (O_1271,N_9925,N_9989);
or UO_1272 (O_1272,N_9907,N_9976);
or UO_1273 (O_1273,N_9968,N_9974);
nor UO_1274 (O_1274,N_9920,N_9967);
or UO_1275 (O_1275,N_9995,N_9948);
nor UO_1276 (O_1276,N_9963,N_9919);
and UO_1277 (O_1277,N_9910,N_9960);
nand UO_1278 (O_1278,N_9982,N_9990);
and UO_1279 (O_1279,N_9905,N_9920);
or UO_1280 (O_1280,N_9973,N_9936);
and UO_1281 (O_1281,N_9982,N_9994);
nor UO_1282 (O_1282,N_9923,N_9905);
and UO_1283 (O_1283,N_9910,N_9985);
or UO_1284 (O_1284,N_9975,N_9931);
nand UO_1285 (O_1285,N_9907,N_9942);
nor UO_1286 (O_1286,N_9902,N_9991);
nand UO_1287 (O_1287,N_9946,N_9938);
and UO_1288 (O_1288,N_9951,N_9957);
and UO_1289 (O_1289,N_9932,N_9926);
nand UO_1290 (O_1290,N_9965,N_9909);
and UO_1291 (O_1291,N_9906,N_9965);
nand UO_1292 (O_1292,N_9928,N_9951);
and UO_1293 (O_1293,N_9965,N_9973);
xnor UO_1294 (O_1294,N_9943,N_9939);
or UO_1295 (O_1295,N_9937,N_9911);
nand UO_1296 (O_1296,N_9953,N_9935);
nand UO_1297 (O_1297,N_9922,N_9960);
and UO_1298 (O_1298,N_9931,N_9929);
nor UO_1299 (O_1299,N_9939,N_9966);
nor UO_1300 (O_1300,N_9948,N_9911);
xor UO_1301 (O_1301,N_9900,N_9914);
nand UO_1302 (O_1302,N_9951,N_9908);
or UO_1303 (O_1303,N_9988,N_9968);
nand UO_1304 (O_1304,N_9958,N_9911);
or UO_1305 (O_1305,N_9999,N_9924);
nand UO_1306 (O_1306,N_9996,N_9937);
nand UO_1307 (O_1307,N_9936,N_9916);
and UO_1308 (O_1308,N_9984,N_9951);
nor UO_1309 (O_1309,N_9926,N_9946);
nor UO_1310 (O_1310,N_9930,N_9912);
nand UO_1311 (O_1311,N_9910,N_9904);
and UO_1312 (O_1312,N_9961,N_9927);
and UO_1313 (O_1313,N_9921,N_9914);
nand UO_1314 (O_1314,N_9989,N_9982);
nor UO_1315 (O_1315,N_9913,N_9923);
nand UO_1316 (O_1316,N_9915,N_9946);
nor UO_1317 (O_1317,N_9984,N_9969);
and UO_1318 (O_1318,N_9983,N_9996);
nor UO_1319 (O_1319,N_9948,N_9986);
and UO_1320 (O_1320,N_9979,N_9967);
nor UO_1321 (O_1321,N_9951,N_9956);
and UO_1322 (O_1322,N_9954,N_9930);
or UO_1323 (O_1323,N_9947,N_9959);
and UO_1324 (O_1324,N_9991,N_9982);
xnor UO_1325 (O_1325,N_9939,N_9902);
or UO_1326 (O_1326,N_9974,N_9997);
or UO_1327 (O_1327,N_9934,N_9975);
xor UO_1328 (O_1328,N_9963,N_9994);
or UO_1329 (O_1329,N_9950,N_9961);
nor UO_1330 (O_1330,N_9979,N_9910);
nand UO_1331 (O_1331,N_9967,N_9925);
and UO_1332 (O_1332,N_9965,N_9977);
xnor UO_1333 (O_1333,N_9994,N_9998);
nand UO_1334 (O_1334,N_9941,N_9959);
or UO_1335 (O_1335,N_9923,N_9924);
or UO_1336 (O_1336,N_9941,N_9910);
and UO_1337 (O_1337,N_9908,N_9957);
nor UO_1338 (O_1338,N_9980,N_9948);
and UO_1339 (O_1339,N_9965,N_9960);
or UO_1340 (O_1340,N_9998,N_9985);
and UO_1341 (O_1341,N_9919,N_9965);
nor UO_1342 (O_1342,N_9942,N_9937);
nand UO_1343 (O_1343,N_9976,N_9929);
nand UO_1344 (O_1344,N_9982,N_9942);
nand UO_1345 (O_1345,N_9995,N_9993);
nor UO_1346 (O_1346,N_9968,N_9930);
nand UO_1347 (O_1347,N_9930,N_9996);
nand UO_1348 (O_1348,N_9988,N_9954);
nor UO_1349 (O_1349,N_9970,N_9983);
and UO_1350 (O_1350,N_9978,N_9965);
nand UO_1351 (O_1351,N_9917,N_9992);
and UO_1352 (O_1352,N_9905,N_9934);
nor UO_1353 (O_1353,N_9989,N_9908);
or UO_1354 (O_1354,N_9900,N_9903);
xor UO_1355 (O_1355,N_9918,N_9973);
and UO_1356 (O_1356,N_9970,N_9957);
nor UO_1357 (O_1357,N_9975,N_9984);
nand UO_1358 (O_1358,N_9945,N_9922);
xor UO_1359 (O_1359,N_9911,N_9986);
or UO_1360 (O_1360,N_9923,N_9952);
xnor UO_1361 (O_1361,N_9916,N_9909);
and UO_1362 (O_1362,N_9933,N_9969);
xor UO_1363 (O_1363,N_9963,N_9942);
nor UO_1364 (O_1364,N_9924,N_9926);
and UO_1365 (O_1365,N_9913,N_9998);
or UO_1366 (O_1366,N_9912,N_9934);
and UO_1367 (O_1367,N_9947,N_9941);
nand UO_1368 (O_1368,N_9943,N_9907);
nor UO_1369 (O_1369,N_9981,N_9967);
or UO_1370 (O_1370,N_9969,N_9966);
or UO_1371 (O_1371,N_9986,N_9943);
or UO_1372 (O_1372,N_9928,N_9935);
nor UO_1373 (O_1373,N_9970,N_9906);
xor UO_1374 (O_1374,N_9973,N_9952);
and UO_1375 (O_1375,N_9930,N_9976);
nand UO_1376 (O_1376,N_9932,N_9950);
nor UO_1377 (O_1377,N_9906,N_9999);
xor UO_1378 (O_1378,N_9952,N_9946);
or UO_1379 (O_1379,N_9989,N_9991);
nor UO_1380 (O_1380,N_9978,N_9920);
and UO_1381 (O_1381,N_9951,N_9992);
or UO_1382 (O_1382,N_9966,N_9971);
nand UO_1383 (O_1383,N_9922,N_9932);
nor UO_1384 (O_1384,N_9973,N_9994);
xnor UO_1385 (O_1385,N_9937,N_9984);
nand UO_1386 (O_1386,N_9973,N_9967);
or UO_1387 (O_1387,N_9948,N_9936);
or UO_1388 (O_1388,N_9997,N_9902);
and UO_1389 (O_1389,N_9980,N_9916);
nor UO_1390 (O_1390,N_9922,N_9964);
nor UO_1391 (O_1391,N_9999,N_9905);
nor UO_1392 (O_1392,N_9995,N_9987);
nand UO_1393 (O_1393,N_9975,N_9965);
nand UO_1394 (O_1394,N_9960,N_9983);
nand UO_1395 (O_1395,N_9974,N_9985);
nand UO_1396 (O_1396,N_9988,N_9991);
or UO_1397 (O_1397,N_9911,N_9990);
and UO_1398 (O_1398,N_9922,N_9976);
nor UO_1399 (O_1399,N_9919,N_9973);
xor UO_1400 (O_1400,N_9912,N_9980);
nor UO_1401 (O_1401,N_9970,N_9934);
nand UO_1402 (O_1402,N_9944,N_9907);
xnor UO_1403 (O_1403,N_9982,N_9969);
and UO_1404 (O_1404,N_9929,N_9987);
xnor UO_1405 (O_1405,N_9963,N_9958);
or UO_1406 (O_1406,N_9976,N_9938);
xor UO_1407 (O_1407,N_9969,N_9912);
or UO_1408 (O_1408,N_9974,N_9937);
and UO_1409 (O_1409,N_9996,N_9935);
and UO_1410 (O_1410,N_9973,N_9928);
and UO_1411 (O_1411,N_9948,N_9999);
nand UO_1412 (O_1412,N_9921,N_9912);
nand UO_1413 (O_1413,N_9947,N_9933);
xor UO_1414 (O_1414,N_9951,N_9998);
nand UO_1415 (O_1415,N_9953,N_9946);
or UO_1416 (O_1416,N_9978,N_9936);
nand UO_1417 (O_1417,N_9986,N_9953);
and UO_1418 (O_1418,N_9916,N_9986);
and UO_1419 (O_1419,N_9912,N_9943);
nor UO_1420 (O_1420,N_9942,N_9979);
or UO_1421 (O_1421,N_9935,N_9982);
and UO_1422 (O_1422,N_9920,N_9987);
nor UO_1423 (O_1423,N_9943,N_9902);
and UO_1424 (O_1424,N_9966,N_9987);
and UO_1425 (O_1425,N_9947,N_9966);
nor UO_1426 (O_1426,N_9969,N_9951);
nor UO_1427 (O_1427,N_9990,N_9907);
and UO_1428 (O_1428,N_9918,N_9930);
nand UO_1429 (O_1429,N_9972,N_9911);
nand UO_1430 (O_1430,N_9980,N_9987);
nand UO_1431 (O_1431,N_9946,N_9935);
or UO_1432 (O_1432,N_9902,N_9959);
and UO_1433 (O_1433,N_9911,N_9966);
xnor UO_1434 (O_1434,N_9918,N_9970);
or UO_1435 (O_1435,N_9991,N_9972);
nand UO_1436 (O_1436,N_9987,N_9959);
nand UO_1437 (O_1437,N_9933,N_9918);
nand UO_1438 (O_1438,N_9900,N_9930);
nor UO_1439 (O_1439,N_9923,N_9926);
and UO_1440 (O_1440,N_9932,N_9987);
or UO_1441 (O_1441,N_9986,N_9909);
nor UO_1442 (O_1442,N_9942,N_9981);
nor UO_1443 (O_1443,N_9937,N_9923);
nand UO_1444 (O_1444,N_9956,N_9994);
nand UO_1445 (O_1445,N_9993,N_9937);
nand UO_1446 (O_1446,N_9925,N_9992);
or UO_1447 (O_1447,N_9955,N_9944);
nand UO_1448 (O_1448,N_9978,N_9992);
nor UO_1449 (O_1449,N_9933,N_9906);
nand UO_1450 (O_1450,N_9958,N_9968);
and UO_1451 (O_1451,N_9948,N_9959);
nand UO_1452 (O_1452,N_9950,N_9913);
xor UO_1453 (O_1453,N_9966,N_9975);
and UO_1454 (O_1454,N_9917,N_9946);
nand UO_1455 (O_1455,N_9920,N_9991);
xnor UO_1456 (O_1456,N_9928,N_9941);
and UO_1457 (O_1457,N_9947,N_9915);
nand UO_1458 (O_1458,N_9903,N_9924);
and UO_1459 (O_1459,N_9903,N_9964);
nand UO_1460 (O_1460,N_9936,N_9912);
and UO_1461 (O_1461,N_9960,N_9902);
nor UO_1462 (O_1462,N_9980,N_9952);
or UO_1463 (O_1463,N_9944,N_9936);
or UO_1464 (O_1464,N_9984,N_9902);
nor UO_1465 (O_1465,N_9961,N_9918);
and UO_1466 (O_1466,N_9969,N_9968);
xor UO_1467 (O_1467,N_9975,N_9959);
xnor UO_1468 (O_1468,N_9916,N_9960);
or UO_1469 (O_1469,N_9908,N_9929);
or UO_1470 (O_1470,N_9906,N_9916);
xnor UO_1471 (O_1471,N_9948,N_9981);
nand UO_1472 (O_1472,N_9946,N_9990);
and UO_1473 (O_1473,N_9996,N_9955);
and UO_1474 (O_1474,N_9964,N_9920);
xnor UO_1475 (O_1475,N_9954,N_9959);
nor UO_1476 (O_1476,N_9920,N_9968);
nor UO_1477 (O_1477,N_9952,N_9909);
nor UO_1478 (O_1478,N_9911,N_9923);
nor UO_1479 (O_1479,N_9944,N_9909);
nand UO_1480 (O_1480,N_9953,N_9922);
or UO_1481 (O_1481,N_9901,N_9944);
nor UO_1482 (O_1482,N_9994,N_9913);
or UO_1483 (O_1483,N_9913,N_9912);
and UO_1484 (O_1484,N_9933,N_9986);
nand UO_1485 (O_1485,N_9969,N_9962);
or UO_1486 (O_1486,N_9971,N_9960);
nor UO_1487 (O_1487,N_9939,N_9995);
nor UO_1488 (O_1488,N_9924,N_9976);
and UO_1489 (O_1489,N_9915,N_9924);
nor UO_1490 (O_1490,N_9950,N_9991);
and UO_1491 (O_1491,N_9960,N_9986);
or UO_1492 (O_1492,N_9988,N_9935);
nand UO_1493 (O_1493,N_9989,N_9954);
nor UO_1494 (O_1494,N_9912,N_9952);
xnor UO_1495 (O_1495,N_9994,N_9950);
and UO_1496 (O_1496,N_9960,N_9931);
xor UO_1497 (O_1497,N_9940,N_9961);
nand UO_1498 (O_1498,N_9940,N_9925);
or UO_1499 (O_1499,N_9918,N_9924);
endmodule