module basic_1000_10000_1500_100_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_95,In_844);
xnor U1 (N_1,In_563,In_222);
nor U2 (N_2,In_182,In_990);
nand U3 (N_3,In_368,In_531);
nand U4 (N_4,In_426,In_1);
nand U5 (N_5,In_338,In_456);
or U6 (N_6,In_639,In_462);
nor U7 (N_7,In_975,In_232);
or U8 (N_8,In_79,In_525);
nand U9 (N_9,In_300,In_641);
nor U10 (N_10,In_546,In_739);
nand U11 (N_11,In_475,In_996);
or U12 (N_12,In_199,In_309);
nand U13 (N_13,In_480,In_882);
nor U14 (N_14,In_784,In_942);
nand U15 (N_15,In_589,In_828);
nor U16 (N_16,In_434,In_941);
and U17 (N_17,In_241,In_961);
nand U18 (N_18,In_306,In_22);
nand U19 (N_19,In_412,In_217);
xnor U20 (N_20,In_819,In_792);
nor U21 (N_21,In_134,In_335);
xor U22 (N_22,In_176,In_155);
or U23 (N_23,In_69,In_109);
nand U24 (N_24,In_735,In_320);
nor U25 (N_25,In_912,In_272);
and U26 (N_26,In_315,In_48);
nand U27 (N_27,In_999,In_84);
nor U28 (N_28,In_219,In_183);
and U29 (N_29,In_373,In_610);
nor U30 (N_30,In_859,In_181);
or U31 (N_31,In_788,In_213);
nor U32 (N_32,In_408,In_653);
xnor U33 (N_33,In_611,In_27);
or U34 (N_34,In_119,In_956);
nand U35 (N_35,In_842,In_801);
or U36 (N_36,In_311,In_738);
and U37 (N_37,In_264,In_670);
or U38 (N_38,In_561,In_42);
nor U39 (N_39,In_419,In_188);
nand U40 (N_40,In_694,In_489);
xor U41 (N_41,In_866,In_274);
or U42 (N_42,In_152,In_949);
or U43 (N_43,In_687,In_130);
nand U44 (N_44,In_700,In_364);
and U45 (N_45,In_575,In_767);
nand U46 (N_46,In_877,In_562);
nand U47 (N_47,In_33,In_619);
nor U48 (N_48,In_785,In_365);
nor U49 (N_49,In_973,In_609);
and U50 (N_50,In_371,In_601);
nor U51 (N_51,In_400,In_112);
xor U52 (N_52,In_35,In_151);
and U53 (N_53,In_539,In_2);
nand U54 (N_54,In_814,In_359);
nand U55 (N_55,In_225,In_482);
or U56 (N_56,In_711,In_908);
nand U57 (N_57,In_495,In_939);
or U58 (N_58,In_926,In_816);
nand U59 (N_59,In_922,In_790);
nor U60 (N_60,In_30,In_136);
nand U61 (N_61,In_848,In_195);
and U62 (N_62,In_75,In_659);
nor U63 (N_63,In_871,In_421);
nor U64 (N_64,In_576,In_341);
or U65 (N_65,In_645,In_672);
nor U66 (N_66,In_409,In_962);
or U67 (N_67,In_715,In_542);
nand U68 (N_68,In_321,In_584);
nand U69 (N_69,In_564,In_86);
or U70 (N_70,In_757,In_487);
and U71 (N_71,In_148,In_253);
nand U72 (N_72,In_682,In_497);
and U73 (N_73,In_924,In_395);
nand U74 (N_74,In_324,In_781);
nor U75 (N_75,In_102,In_630);
or U76 (N_76,In_722,In_529);
or U77 (N_77,In_839,In_108);
or U78 (N_78,In_932,In_760);
or U79 (N_79,In_793,In_530);
xnor U80 (N_80,In_255,In_286);
nand U81 (N_81,In_501,In_454);
or U82 (N_82,In_350,In_778);
nor U83 (N_83,In_125,In_964);
and U84 (N_84,In_66,In_296);
nand U85 (N_85,In_879,In_725);
nor U86 (N_86,In_65,In_15);
nand U87 (N_87,In_934,In_890);
nor U88 (N_88,In_308,In_696);
or U89 (N_89,In_720,In_634);
nor U90 (N_90,In_804,In_997);
and U91 (N_91,In_673,In_297);
and U92 (N_92,In_588,In_993);
and U93 (N_93,In_796,In_325);
nand U94 (N_94,In_477,In_226);
nand U95 (N_95,In_783,In_508);
or U96 (N_96,In_175,In_343);
or U97 (N_97,In_852,In_913);
nand U98 (N_98,In_940,In_637);
nor U99 (N_99,In_357,In_345);
and U100 (N_100,N_78,In_360);
nand U101 (N_101,In_730,In_969);
nand U102 (N_102,In_276,In_632);
and U103 (N_103,In_745,In_453);
nor U104 (N_104,In_282,In_96);
nand U105 (N_105,In_698,In_332);
nor U106 (N_106,In_773,In_124);
and U107 (N_107,In_719,In_505);
or U108 (N_108,In_688,In_455);
nand U109 (N_109,In_536,In_23);
nand U110 (N_110,In_885,In_958);
nor U111 (N_111,In_499,In_517);
nor U112 (N_112,In_620,In_847);
nand U113 (N_113,In_492,In_41);
nand U114 (N_114,In_731,In_909);
nand U115 (N_115,In_585,In_714);
nand U116 (N_116,In_571,In_976);
nand U117 (N_117,In_503,In_312);
or U118 (N_118,In_423,In_513);
and U119 (N_119,N_64,In_936);
nor U120 (N_120,In_521,In_867);
nand U121 (N_121,In_117,In_31);
or U122 (N_122,In_168,In_957);
nor U123 (N_123,In_110,In_840);
nand U124 (N_124,In_953,In_663);
or U125 (N_125,In_543,In_161);
or U126 (N_126,In_984,In_980);
and U127 (N_127,In_83,In_438);
and U128 (N_128,In_301,In_728);
and U129 (N_129,In_449,In_459);
nor U130 (N_130,In_191,In_390);
nand U131 (N_131,In_707,In_206);
or U132 (N_132,In_774,In_636);
nand U133 (N_133,N_11,In_534);
and U134 (N_134,In_535,In_945);
xor U135 (N_135,In_85,In_293);
nor U136 (N_136,In_411,In_894);
nor U137 (N_137,In_154,In_407);
and U138 (N_138,In_103,In_813);
and U139 (N_139,In_742,In_678);
and U140 (N_140,In_77,In_603);
nor U141 (N_141,In_818,N_93);
and U142 (N_142,In_727,In_834);
nor U143 (N_143,In_260,In_471);
nand U144 (N_144,In_73,In_549);
or U145 (N_145,In_322,N_33);
nor U146 (N_146,N_6,In_149);
and U147 (N_147,In_244,In_709);
or U148 (N_148,N_0,In_938);
or U149 (N_149,In_602,In_986);
and U150 (N_150,In_101,In_662);
or U151 (N_151,In_795,In_7);
and U152 (N_152,N_44,In_855);
and U153 (N_153,In_915,In_626);
and U154 (N_154,In_873,In_458);
or U155 (N_155,In_105,In_968);
nor U156 (N_156,In_811,N_54);
xor U157 (N_157,In_384,In_464);
nand U158 (N_158,In_744,N_26);
nand U159 (N_159,N_12,In_229);
nand U160 (N_160,In_887,In_970);
and U161 (N_161,N_62,In_724);
nand U162 (N_162,In_12,In_649);
or U163 (N_163,In_615,In_669);
nor U164 (N_164,In_808,In_835);
nand U165 (N_165,In_436,In_820);
nand U166 (N_166,In_63,In_88);
or U167 (N_167,In_729,In_930);
or U168 (N_168,In_982,In_246);
nand U169 (N_169,N_4,In_261);
nand U170 (N_170,In_937,In_880);
and U171 (N_171,In_215,In_763);
or U172 (N_172,In_540,In_833);
or U173 (N_173,N_59,N_53);
and U174 (N_174,In_388,N_49);
and U175 (N_175,In_254,In_568);
or U176 (N_176,In_946,In_935);
and U177 (N_177,In_850,In_404);
and U178 (N_178,In_237,In_648);
and U179 (N_179,In_627,In_516);
nor U180 (N_180,In_889,In_120);
or U181 (N_181,In_862,In_18);
or U182 (N_182,In_146,In_787);
or U183 (N_183,In_797,In_494);
xor U184 (N_184,In_876,In_697);
nor U185 (N_185,In_340,In_192);
nand U186 (N_186,In_349,In_666);
and U187 (N_187,In_34,In_207);
xnor U188 (N_188,In_856,In_26);
and U189 (N_189,In_581,In_954);
nand U190 (N_190,In_606,In_824);
or U191 (N_191,In_597,In_342);
or U192 (N_192,In_180,In_914);
nor U193 (N_193,In_317,In_288);
or U194 (N_194,In_44,N_73);
nand U195 (N_195,In_803,In_221);
xnor U196 (N_196,In_905,In_169);
or U197 (N_197,N_57,In_81);
nand U198 (N_198,N_42,In_762);
and U199 (N_199,In_706,N_84);
nand U200 (N_200,In_262,In_732);
nor U201 (N_201,In_684,In_479);
xor U202 (N_202,In_150,In_594);
nor U203 (N_203,In_115,N_95);
nand U204 (N_204,In_690,In_592);
nand U205 (N_205,In_19,In_193);
nand U206 (N_206,In_822,N_110);
or U207 (N_207,N_145,In_40);
nand U208 (N_208,In_772,N_35);
nor U209 (N_209,In_89,In_427);
xnor U210 (N_210,In_116,In_507);
nand U211 (N_211,N_188,In_486);
or U212 (N_212,N_109,In_159);
or U213 (N_213,In_799,In_921);
nor U214 (N_214,In_271,In_553);
and U215 (N_215,In_750,In_328);
nand U216 (N_216,In_46,In_323);
nand U217 (N_217,N_107,N_199);
or U218 (N_218,In_375,In_202);
and U219 (N_219,In_717,In_20);
nor U220 (N_220,In_268,In_614);
nor U221 (N_221,In_74,N_82);
nor U222 (N_222,In_439,N_10);
nor U223 (N_223,In_467,In_337);
nor U224 (N_224,In_650,In_829);
or U225 (N_225,N_124,In_269);
or U226 (N_226,N_134,In_911);
and U227 (N_227,N_142,In_823);
or U228 (N_228,In_316,N_52);
or U229 (N_229,In_474,In_141);
nor U230 (N_230,In_519,In_830);
nand U231 (N_231,In_680,In_548);
and U232 (N_232,In_258,In_263);
or U233 (N_233,In_955,In_979);
nand U234 (N_234,In_171,In_281);
and U235 (N_235,In_794,In_386);
nand U236 (N_236,In_416,In_393);
or U237 (N_237,In_481,In_243);
nand U238 (N_238,N_123,In_743);
or U239 (N_239,N_191,In_613);
nand U240 (N_240,In_617,In_566);
nand U241 (N_241,In_417,In_273);
nand U242 (N_242,In_118,In_607);
and U243 (N_243,In_963,In_703);
nand U244 (N_244,In_3,N_88);
and U245 (N_245,In_425,N_2);
and U246 (N_246,In_651,In_868);
or U247 (N_247,In_230,In_502);
nor U248 (N_248,In_798,In_280);
or U249 (N_249,In_863,In_923);
and U250 (N_250,In_777,N_192);
or U251 (N_251,In_247,In_466);
nand U252 (N_252,In_54,N_36);
and U253 (N_253,In_896,In_392);
nor U254 (N_254,N_151,N_146);
nand U255 (N_255,In_533,In_228);
nand U256 (N_256,In_965,In_29);
nand U257 (N_257,In_410,N_137);
nor U258 (N_258,In_129,In_346);
nor U259 (N_259,In_177,In_864);
nand U260 (N_260,In_644,In_752);
or U261 (N_261,In_71,N_43);
nor U262 (N_262,In_212,In_190);
nor U263 (N_263,In_433,In_555);
and U264 (N_264,In_326,In_741);
nor U265 (N_265,In_749,N_83);
and U266 (N_266,In_422,In_522);
xnor U267 (N_267,In_302,In_216);
or U268 (N_268,N_121,In_577);
or U269 (N_269,In_898,In_370);
or U270 (N_270,In_881,In_205);
nand U271 (N_271,N_47,N_87);
or U272 (N_272,In_259,In_14);
and U273 (N_273,N_60,N_96);
nand U274 (N_274,In_992,N_158);
and U275 (N_275,In_420,In_959);
or U276 (N_276,In_853,In_147);
xnor U277 (N_277,In_559,In_387);
nand U278 (N_278,In_313,In_314);
or U279 (N_279,In_469,In_305);
xnor U280 (N_280,In_872,N_74);
or U281 (N_281,In_10,In_327);
nor U282 (N_282,In_139,In_145);
or U283 (N_283,In_558,In_121);
nand U284 (N_284,N_149,In_726);
and U285 (N_285,N_172,In_172);
and U286 (N_286,N_176,In_189);
nand U287 (N_287,In_39,N_139);
or U288 (N_288,In_201,In_490);
or U289 (N_289,In_802,In_821);
or U290 (N_290,In_99,In_463);
nand U291 (N_291,In_506,In_361);
nor U292 (N_292,N_119,N_5);
or U293 (N_293,In_476,In_838);
nor U294 (N_294,In_210,In_339);
xor U295 (N_295,In_628,In_567);
and U296 (N_296,In_837,In_367);
and U297 (N_297,N_8,In_674);
or U298 (N_298,In_488,N_79);
and U299 (N_299,N_91,In_899);
nor U300 (N_300,In_870,N_167);
nand U301 (N_301,In_330,N_269);
and U302 (N_302,N_92,In_143);
and U303 (N_303,N_287,In_616);
nand U304 (N_304,N_279,In_240);
nand U305 (N_305,N_32,In_208);
nor U306 (N_306,N_173,N_286);
and U307 (N_307,In_658,In_251);
and U308 (N_308,N_218,In_951);
and U309 (N_309,In_618,In_574);
nand U310 (N_310,In_403,N_258);
nand U311 (N_311,In_389,In_443);
or U312 (N_312,In_646,In_713);
and U313 (N_313,In_113,N_174);
and U314 (N_314,In_874,N_185);
nand U315 (N_315,N_246,In_58);
nand U316 (N_316,In_765,In_93);
nor U317 (N_317,N_253,In_319);
nand U318 (N_318,In_557,N_126);
nor U319 (N_319,N_241,N_231);
nand U320 (N_320,In_692,N_162);
and U321 (N_321,In_334,In_608);
or U322 (N_322,In_538,In_196);
nand U323 (N_323,In_366,In_810);
nor U324 (N_324,N_235,N_111);
and U325 (N_325,In_625,In_307);
or U326 (N_326,N_89,N_61);
or U327 (N_327,In_565,In_218);
or U328 (N_328,N_177,In_580);
nand U329 (N_329,N_180,In_396);
or U330 (N_330,In_587,In_836);
or U331 (N_331,N_157,In_705);
or U332 (N_332,In_754,N_228);
and U333 (N_333,In_142,N_99);
xor U334 (N_334,In_194,N_229);
nor U335 (N_335,In_892,N_205);
nor U336 (N_336,In_82,In_446);
nand U337 (N_337,In_655,In_756);
or U338 (N_338,N_166,N_125);
nor U339 (N_339,In_686,In_24);
nand U340 (N_340,In_299,In_138);
or U341 (N_341,In_710,In_483);
nor U342 (N_342,In_352,N_206);
or U343 (N_343,In_805,In_578);
and U344 (N_344,In_746,In_132);
nor U345 (N_345,In_394,In_667);
or U346 (N_346,In_551,In_220);
and U347 (N_347,N_150,In_928);
nor U348 (N_348,In_675,In_527);
and U349 (N_349,N_273,In_51);
and U350 (N_350,In_298,N_224);
or U351 (N_351,In_845,In_764);
nand U352 (N_352,In_812,In_514);
nand U353 (N_353,N_144,In_239);
or U354 (N_354,N_22,N_3);
or U355 (N_355,N_165,In_333);
or U356 (N_356,In_664,N_136);
and U357 (N_357,N_202,N_251);
or U358 (N_358,In_515,In_111);
nand U359 (N_359,N_238,In_76);
nand U360 (N_360,In_524,N_65);
nor U361 (N_361,In_72,In_640);
and U362 (N_362,N_239,In_901);
or U363 (N_363,N_71,In_123);
and U364 (N_364,In_776,In_347);
and U365 (N_365,N_100,In_401);
nor U366 (N_366,In_591,In_657);
nand U367 (N_367,In_579,In_331);
or U368 (N_368,In_989,In_988);
nor U369 (N_369,In_832,N_220);
or U370 (N_370,In_747,In_382);
nor U371 (N_371,In_493,N_230);
or U372 (N_372,N_187,In_283);
nor U373 (N_373,In_943,In_605);
nand U374 (N_374,In_511,In_888);
nor U375 (N_375,In_78,In_496);
nor U376 (N_376,In_902,N_143);
and U377 (N_377,In_817,In_950);
nand U378 (N_378,In_295,In_140);
nor U379 (N_379,In_362,N_23);
nand U380 (N_380,N_50,N_236);
or U381 (N_381,In_621,In_80);
or U382 (N_382,In_920,N_203);
nor U383 (N_383,In_356,In_782);
and U384 (N_384,In_952,In_695);
or U385 (N_385,In_158,N_276);
or U386 (N_386,In_595,N_244);
nor U387 (N_387,N_1,In_424);
nor U388 (N_388,In_484,In_701);
nor U389 (N_389,N_247,In_815);
xnor U390 (N_390,N_221,In_485);
nor U391 (N_391,In_131,In_238);
nand U392 (N_392,In_447,N_18);
xnor U393 (N_393,N_272,In_891);
nor U394 (N_394,N_296,In_917);
and U395 (N_395,N_289,In_846);
or U396 (N_396,N_265,In_849);
or U397 (N_397,In_596,In_509);
or U398 (N_398,In_414,In_59);
nand U399 (N_399,In_442,In_162);
and U400 (N_400,In_60,N_34);
nor U401 (N_401,N_295,In_203);
or U402 (N_402,N_135,N_306);
xor U403 (N_403,N_371,N_9);
nand U404 (N_404,In_380,N_257);
nand U405 (N_405,N_375,In_759);
nor U406 (N_406,N_216,In_668);
nor U407 (N_407,In_600,In_399);
nand U408 (N_408,In_55,N_320);
nor U409 (N_409,In_886,In_21);
or U410 (N_410,N_69,In_265);
or U411 (N_411,In_413,In_133);
nand U412 (N_412,N_102,In_184);
nor U413 (N_413,In_769,N_31);
nand U414 (N_414,N_291,In_478);
and U415 (N_415,N_154,In_869);
or U416 (N_416,N_256,In_789);
and U417 (N_417,N_277,In_170);
and U418 (N_418,N_242,N_94);
and U419 (N_419,In_186,N_360);
or U420 (N_420,In_884,In_294);
or U421 (N_421,In_857,N_171);
and U422 (N_422,N_329,In_523);
nand U423 (N_423,N_350,In_893);
nor U424 (N_424,In_28,N_213);
nand U425 (N_425,N_387,N_370);
or U426 (N_426,In_768,In_385);
and U427 (N_427,N_264,In_284);
or U428 (N_428,In_256,N_232);
nor U429 (N_429,N_13,N_318);
or U430 (N_430,In_437,In_68);
and U431 (N_431,In_174,In_236);
nor U432 (N_432,N_396,N_372);
nand U433 (N_433,N_342,N_313);
nand U434 (N_434,N_30,In_398);
or U435 (N_435,In_363,In_106);
nor U436 (N_436,In_624,N_367);
nand U437 (N_437,N_303,In_165);
nand U438 (N_438,N_20,In_9);
nand U439 (N_439,N_326,In_157);
nor U440 (N_440,N_63,In_791);
xnor U441 (N_441,In_622,N_161);
and U442 (N_442,N_270,N_314);
or U443 (N_443,In_304,In_289);
nor U444 (N_444,In_374,N_308);
and U445 (N_445,In_656,In_683);
and U446 (N_446,In_895,In_878);
nand U447 (N_447,In_586,In_6);
nor U448 (N_448,In_647,N_356);
and U449 (N_449,N_140,N_86);
nor U450 (N_450,In_702,In_925);
or U451 (N_451,N_46,In_661);
and U452 (N_452,In_17,N_357);
nand U453 (N_453,N_267,N_271);
nand U454 (N_454,N_68,N_340);
and U455 (N_455,In_97,In_128);
and U456 (N_456,N_352,In_185);
nor U457 (N_457,N_104,In_665);
xor U458 (N_458,In_178,In_987);
nor U459 (N_459,N_389,In_43);
or U460 (N_460,In_593,In_285);
nand U461 (N_461,N_17,In_329);
nand U462 (N_462,N_333,In_250);
or U463 (N_463,In_751,In_11);
and U464 (N_464,N_132,N_281);
and U465 (N_465,In_461,In_998);
nand U466 (N_466,N_122,N_207);
or U467 (N_467,In_883,N_193);
nor U468 (N_468,N_19,In_13);
and U469 (N_469,N_397,N_331);
nor U470 (N_470,N_153,In_526);
and U471 (N_471,N_29,N_250);
or U472 (N_472,In_635,N_384);
and U473 (N_473,N_399,In_204);
nand U474 (N_474,In_358,In_270);
and U475 (N_475,In_67,N_181);
or U476 (N_476,In_38,In_252);
nor U477 (N_477,In_532,N_332);
nand U478 (N_478,In_126,N_266);
and U479 (N_479,N_245,In_135);
nor U480 (N_480,N_365,N_301);
or U481 (N_481,N_103,N_338);
nand U482 (N_482,In_933,In_100);
nor U483 (N_483,N_97,N_15);
nor U484 (N_484,N_225,N_341);
and U485 (N_485,In_57,N_114);
nand U486 (N_486,In_843,N_152);
or U487 (N_487,In_137,In_224);
nand U488 (N_488,In_61,N_77);
or U489 (N_489,N_385,N_182);
nor U490 (N_490,In_604,In_92);
or U491 (N_491,N_113,In_642);
nand U492 (N_492,N_168,N_398);
nor U493 (N_493,N_310,N_368);
nand U494 (N_494,In_153,N_226);
or U495 (N_495,In_994,In_629);
nand U496 (N_496,In_451,N_278);
nor U497 (N_497,N_322,In_267);
or U498 (N_498,In_107,In_104);
nor U499 (N_499,In_354,In_344);
or U500 (N_500,In_468,In_500);
and U501 (N_501,N_309,N_70);
nor U502 (N_502,In_948,In_179);
and U503 (N_503,In_918,In_740);
or U504 (N_504,N_170,N_175);
and U505 (N_505,N_478,In_991);
nor U506 (N_506,N_381,N_285);
and U507 (N_507,N_319,N_156);
nand U508 (N_508,N_305,N_294);
and U509 (N_509,N_106,N_155);
xnor U510 (N_510,In_248,N_401);
nand U511 (N_511,In_214,N_390);
and U512 (N_512,In_242,N_90);
and U513 (N_513,N_392,N_48);
nor U514 (N_514,In_780,N_485);
xor U515 (N_515,In_291,N_315);
or U516 (N_516,In_173,In_758);
nand U517 (N_517,In_491,In_693);
and U518 (N_518,N_388,In_550);
and U519 (N_519,N_355,In_544);
nand U520 (N_520,N_184,N_444);
nor U521 (N_521,N_456,N_330);
or U522 (N_522,N_25,In_5);
or U523 (N_523,In_573,N_432);
nor U524 (N_524,N_423,N_470);
nor U525 (N_525,N_377,N_237);
xor U526 (N_526,In_405,In_114);
or U527 (N_527,N_56,N_445);
nand U528 (N_528,In_460,In_90);
and U529 (N_529,In_336,N_484);
and U530 (N_530,In_234,N_450);
nor U531 (N_531,N_85,N_349);
nor U532 (N_532,N_492,In_465);
nor U533 (N_533,N_452,N_327);
nand U534 (N_534,In_807,In_676);
nand U535 (N_535,N_449,N_302);
nor U536 (N_536,In_699,N_353);
nor U537 (N_537,In_572,In_860);
nand U538 (N_538,In_748,N_196);
or U539 (N_539,N_481,In_800);
or U540 (N_540,In_978,In_851);
nand U541 (N_541,N_24,In_512);
and U542 (N_542,In_737,N_217);
and U543 (N_543,N_298,N_234);
or U544 (N_544,N_208,N_416);
nor U545 (N_545,In_87,In_854);
or U546 (N_546,N_300,N_204);
and U547 (N_547,In_518,N_299);
nand U548 (N_548,N_465,N_76);
nor U549 (N_549,In_211,N_282);
nand U550 (N_550,N_382,N_406);
and U551 (N_551,N_200,In_355);
or U552 (N_552,N_160,N_422);
or U553 (N_553,In_755,N_263);
and U554 (N_554,N_127,N_28);
nand U555 (N_555,N_210,N_446);
and U556 (N_556,N_128,N_379);
nor U557 (N_557,In_62,In_435);
nand U558 (N_558,N_488,N_227);
nor U559 (N_559,N_497,In_633);
or U560 (N_560,In_841,N_480);
or U561 (N_561,N_366,N_409);
nand U562 (N_562,In_415,N_466);
or U563 (N_563,In_547,N_495);
or U564 (N_564,In_448,In_0);
nand U565 (N_565,In_927,N_441);
and U566 (N_566,N_402,N_437);
or U567 (N_567,N_197,In_197);
or U568 (N_568,N_81,N_101);
and U569 (N_569,In_718,N_316);
and U570 (N_570,In_809,N_189);
nand U571 (N_571,N_255,In_166);
nand U572 (N_572,In_432,In_249);
or U573 (N_573,In_733,N_460);
nand U574 (N_574,N_411,N_487);
nand U575 (N_575,N_404,N_451);
nand U576 (N_576,N_283,N_412);
and U577 (N_577,In_638,N_249);
or U578 (N_578,In_223,N_16);
and U579 (N_579,In_266,N_363);
or U580 (N_580,In_906,In_569);
nand U581 (N_581,In_278,N_211);
or U582 (N_582,N_307,In_56);
or U583 (N_583,N_288,In_287);
nand U584 (N_584,N_259,N_45);
and U585 (N_585,N_130,In_47);
nand U586 (N_586,In_972,N_474);
nand U587 (N_587,N_415,In_983);
nand U588 (N_588,N_413,In_826);
and U589 (N_589,In_406,N_66);
nand U590 (N_590,In_32,In_974);
nor U591 (N_591,N_429,N_483);
nor U592 (N_592,N_240,In_919);
and U593 (N_593,In_277,N_383);
nand U594 (N_594,N_410,In_8);
nor U595 (N_595,N_105,In_560);
or U596 (N_596,In_429,In_910);
or U597 (N_597,In_498,In_723);
and U598 (N_598,N_447,N_98);
nor U599 (N_599,N_420,In_631);
or U600 (N_600,In_430,N_587);
nand U601 (N_601,N_506,In_598);
nor U602 (N_602,N_190,N_569);
and U603 (N_603,N_347,In_582);
and U604 (N_604,In_457,N_201);
or U605 (N_605,In_372,In_827);
nor U606 (N_606,N_120,N_403);
and U607 (N_607,In_831,N_588);
and U608 (N_608,In_233,In_428);
or U609 (N_609,In_770,N_594);
or U610 (N_610,N_219,N_378);
and U611 (N_611,N_476,N_529);
or U612 (N_612,In_378,N_408);
nand U613 (N_613,In_450,In_685);
nand U614 (N_614,In_708,In_198);
or U615 (N_615,In_947,N_562);
and U616 (N_616,N_386,N_583);
nand U617 (N_617,N_115,N_464);
xor U618 (N_618,N_575,N_433);
nand U619 (N_619,N_405,In_127);
or U620 (N_620,N_526,In_520);
nand U621 (N_621,In_318,In_167);
nor U622 (N_622,N_557,N_440);
and U623 (N_623,In_379,N_214);
nand U624 (N_624,N_261,In_227);
nand U625 (N_625,N_418,In_689);
nor U626 (N_626,N_148,In_36);
nand U627 (N_627,N_290,In_510);
and U628 (N_628,N_468,N_354);
or U629 (N_629,N_581,In_402);
nand U630 (N_630,In_583,In_391);
and U631 (N_631,N_500,N_501);
and U632 (N_632,N_520,N_548);
or U633 (N_633,In_552,N_194);
nor U634 (N_634,In_144,N_467);
and U635 (N_635,N_552,N_543);
nor U636 (N_636,N_260,In_554);
and U637 (N_637,N_530,In_671);
or U638 (N_638,In_156,In_45);
nand U639 (N_639,In_652,In_431);
nand U640 (N_640,In_310,N_540);
nor U641 (N_641,N_274,N_38);
nor U642 (N_642,In_977,In_865);
and U643 (N_643,In_966,In_52);
and U644 (N_644,N_510,N_517);
nor U645 (N_645,N_596,N_421);
xnor U646 (N_646,N_335,N_537);
or U647 (N_647,N_293,N_195);
and U648 (N_648,In_25,In_70);
or U649 (N_649,In_94,N_515);
or U650 (N_650,In_995,N_534);
nand U651 (N_651,N_284,N_435);
nor U652 (N_652,In_16,N_523);
nand U653 (N_653,In_444,N_364);
nor U654 (N_654,N_317,N_438);
or U655 (N_655,N_491,N_339);
nor U656 (N_656,In_292,In_771);
or U657 (N_657,In_904,In_556);
nand U658 (N_658,N_58,N_542);
nand U659 (N_659,N_584,In_290);
nand U660 (N_660,N_589,N_544);
nand U661 (N_661,N_461,N_490);
nand U662 (N_662,N_586,N_118);
nand U663 (N_663,N_443,In_691);
or U664 (N_664,In_164,N_545);
or U665 (N_665,In_916,N_431);
and U666 (N_666,N_531,N_494);
or U667 (N_667,N_325,N_328);
or U668 (N_668,In_786,In_504);
nor U669 (N_669,N_505,N_524);
and U670 (N_670,N_112,N_463);
nor U671 (N_671,N_222,N_514);
xor U672 (N_672,In_37,N_380);
nor U673 (N_673,N_164,In_681);
nand U674 (N_674,N_527,N_448);
nand U675 (N_675,N_223,N_578);
nor U676 (N_676,N_457,N_503);
xnor U677 (N_677,N_373,N_519);
nor U678 (N_678,In_861,N_599);
nand U679 (N_679,N_343,N_344);
nand U680 (N_680,In_981,N_233);
nand U681 (N_681,N_564,N_138);
and U682 (N_682,N_55,In_704);
and U683 (N_683,N_324,In_545);
or U684 (N_684,N_376,In_231);
nand U685 (N_685,N_141,In_716);
or U686 (N_686,N_163,In_163);
nor U687 (N_687,N_248,N_212);
and U688 (N_688,N_475,N_254);
or U689 (N_689,N_275,In_541);
xor U690 (N_690,N_7,N_521);
nand U691 (N_691,In_303,N_498);
nand U692 (N_692,In_590,In_736);
nor U693 (N_693,In_712,In_903);
nor U694 (N_694,N_336,In_472);
and U695 (N_695,N_252,N_522);
or U696 (N_696,N_131,In_612);
and U697 (N_697,N_186,N_21);
and U698 (N_698,N_504,N_566);
nor U699 (N_699,N_243,N_183);
and U700 (N_700,N_585,N_558);
nand U701 (N_701,N_159,N_601);
nor U702 (N_702,In_677,N_297);
or U703 (N_703,N_661,N_304);
and U704 (N_704,N_407,N_643);
nand U705 (N_705,N_591,N_27);
nand U706 (N_706,N_623,N_80);
or U707 (N_707,N_550,In_49);
nor U708 (N_708,In_64,N_653);
and U709 (N_709,In_929,N_108);
and U710 (N_710,N_361,N_630);
and U711 (N_711,In_779,In_931);
nand U712 (N_712,N_629,N_369);
xnor U713 (N_713,N_496,N_292);
and U714 (N_714,In_91,N_664);
nor U715 (N_715,N_280,In_907);
or U716 (N_716,In_806,N_618);
nor U717 (N_717,N_439,N_477);
nand U718 (N_718,N_536,N_502);
nand U719 (N_719,N_609,In_279);
or U720 (N_720,In_944,N_268);
nand U721 (N_721,N_605,N_311);
nand U722 (N_722,N_147,N_682);
nand U723 (N_723,N_516,N_462);
or U724 (N_724,N_676,N_428);
and U725 (N_725,N_455,N_613);
nand U726 (N_726,N_359,N_627);
nand U727 (N_727,N_471,N_436);
nor U728 (N_728,N_493,In_160);
nor U729 (N_729,N_14,N_607);
and U730 (N_730,N_486,N_612);
or U731 (N_731,N_669,N_553);
or U732 (N_732,N_400,N_647);
nand U733 (N_733,N_129,N_499);
nand U734 (N_734,In_440,N_632);
or U735 (N_735,N_549,N_323);
and U736 (N_736,N_628,N_116);
nand U737 (N_737,N_674,N_473);
or U738 (N_738,N_641,In_245);
nor U739 (N_739,N_209,N_673);
and U740 (N_740,N_570,In_643);
nor U741 (N_741,In_875,N_568);
and U742 (N_742,N_667,In_351);
or U743 (N_743,N_513,In_900);
and U744 (N_744,N_633,N_658);
nor U745 (N_745,N_178,N_665);
and U746 (N_746,N_620,N_508);
or U747 (N_747,N_602,N_563);
nand U748 (N_748,N_430,N_39);
or U749 (N_749,N_663,N_666);
nor U750 (N_750,N_696,N_453);
nor U751 (N_751,N_512,N_551);
nor U752 (N_752,N_459,In_473);
or U753 (N_753,N_592,In_967);
and U754 (N_754,In_623,N_595);
nor U755 (N_755,N_637,N_321);
and U756 (N_756,In_766,N_656);
and U757 (N_757,In_376,In_200);
and U758 (N_758,N_644,In_470);
nand U759 (N_759,N_604,N_417);
nor U760 (N_760,N_626,N_657);
xor U761 (N_761,N_672,In_187);
and U762 (N_762,N_37,N_611);
nand U763 (N_763,N_391,N_555);
nor U764 (N_764,In_353,N_577);
or U765 (N_765,In_971,In_960);
and U766 (N_766,N_635,N_670);
or U767 (N_767,N_482,N_651);
and U768 (N_768,N_692,N_652);
nor U769 (N_769,N_624,N_619);
xor U770 (N_770,N_688,In_985);
or U771 (N_771,N_358,N_533);
and U772 (N_772,N_631,N_133);
and U773 (N_773,N_511,N_179);
or U774 (N_774,N_489,In_753);
nand U775 (N_775,N_414,In_275);
or U776 (N_776,In_654,N_693);
nand U777 (N_777,In_98,N_579);
nand U778 (N_778,N_434,N_574);
nor U779 (N_779,N_636,N_678);
nor U780 (N_780,N_362,In_418);
nand U781 (N_781,N_655,N_374);
nor U782 (N_782,N_603,In_537);
or U783 (N_783,In_775,N_650);
nor U784 (N_784,N_691,N_262);
nand U785 (N_785,N_677,N_668);
or U786 (N_786,N_606,N_424);
and U787 (N_787,N_598,N_215);
or U788 (N_788,N_642,N_648);
and U789 (N_789,N_597,In_761);
xnor U790 (N_790,N_425,N_469);
nor U791 (N_791,N_695,N_395);
nor U792 (N_792,N_687,N_638);
or U793 (N_793,In_209,N_572);
nand U794 (N_794,In_257,N_671);
nor U795 (N_795,In_452,N_689);
or U796 (N_796,N_617,N_690);
nor U797 (N_797,N_582,N_507);
or U798 (N_798,N_580,In_4);
or U799 (N_799,N_472,N_694);
nand U800 (N_800,N_763,N_739);
nand U801 (N_801,N_756,N_600);
nand U802 (N_802,N_754,In_825);
and U803 (N_803,N_198,In_377);
or U804 (N_804,N_616,N_560);
xor U805 (N_805,N_712,N_442);
nor U806 (N_806,N_702,N_725);
nor U807 (N_807,N_72,In_50);
xnor U808 (N_808,N_608,In_660);
xor U809 (N_809,N_610,N_761);
nor U810 (N_810,N_479,N_726);
and U811 (N_811,N_685,N_744);
and U812 (N_812,In_122,N_758);
nor U813 (N_813,N_684,N_770);
nor U814 (N_814,In_445,In_383);
nor U815 (N_815,N_749,N_41);
or U816 (N_816,In_570,N_535);
nor U817 (N_817,N_732,In_381);
nand U818 (N_818,N_747,N_334);
nand U819 (N_819,N_720,N_715);
nor U820 (N_820,N_778,N_698);
nand U821 (N_821,N_654,N_426);
nand U822 (N_822,N_565,N_788);
nor U823 (N_823,N_762,N_393);
nor U824 (N_824,N_662,N_686);
and U825 (N_825,N_733,N_567);
nor U826 (N_826,N_351,N_752);
and U827 (N_827,N_753,N_659);
nor U828 (N_828,N_615,N_734);
nand U829 (N_829,N_794,N_622);
or U830 (N_830,N_660,N_774);
or U831 (N_831,N_621,N_337);
or U832 (N_832,N_169,N_757);
nand U833 (N_833,N_532,N_760);
and U834 (N_834,N_740,N_716);
or U835 (N_835,N_703,N_556);
and U836 (N_836,In_897,N_719);
or U837 (N_837,N_571,N_427);
and U838 (N_838,N_593,N_764);
nand U839 (N_839,N_769,N_554);
nand U840 (N_840,N_751,N_697);
or U841 (N_841,N_722,N_117);
nand U842 (N_842,N_683,N_708);
or U843 (N_843,N_798,N_528);
and U844 (N_844,N_547,N_675);
nor U845 (N_845,In_721,N_711);
nand U846 (N_846,N_700,N_743);
or U847 (N_847,N_746,N_458);
nor U848 (N_848,N_765,N_748);
nand U849 (N_849,N_51,In_235);
or U850 (N_850,N_646,N_538);
and U851 (N_851,N_729,N_766);
and U852 (N_852,N_782,N_546);
and U853 (N_853,N_727,N_797);
or U854 (N_854,N_783,N_771);
nor U855 (N_855,N_742,N_795);
and U856 (N_856,In_441,N_539);
and U857 (N_857,N_750,N_614);
nor U858 (N_858,N_625,N_312);
nand U859 (N_859,N_710,N_759);
and U860 (N_860,N_346,N_773);
and U861 (N_861,N_728,N_775);
or U862 (N_862,N_714,In_679);
and U863 (N_863,In_528,N_706);
nand U864 (N_864,N_791,In_53);
or U865 (N_865,N_768,N_735);
nor U866 (N_866,N_576,N_779);
or U867 (N_867,N_509,N_590);
nor U868 (N_868,N_796,N_67);
and U869 (N_869,N_731,N_573);
and U870 (N_870,N_772,N_518);
nor U871 (N_871,N_741,N_721);
nor U872 (N_872,N_40,N_634);
nor U873 (N_873,N_348,N_707);
or U874 (N_874,N_559,N_640);
and U875 (N_875,N_790,N_745);
and U876 (N_876,In_734,N_730);
or U877 (N_877,N_789,N_561);
or U878 (N_878,N_785,N_799);
and U879 (N_879,N_704,N_525);
nor U880 (N_880,N_781,N_394);
nand U881 (N_881,N_784,N_724);
or U882 (N_882,N_738,N_767);
nor U883 (N_883,N_345,N_649);
nor U884 (N_884,N_780,N_717);
nand U885 (N_885,N_776,N_680);
nand U886 (N_886,N_701,In_369);
or U887 (N_887,N_681,N_792);
or U888 (N_888,N_787,N_755);
xnor U889 (N_889,N_639,N_713);
or U890 (N_890,N_723,N_679);
or U891 (N_891,In_397,N_75);
nand U892 (N_892,N_645,N_736);
nand U893 (N_893,N_718,N_793);
xnor U894 (N_894,N_737,In_858);
nand U895 (N_895,In_599,N_709);
and U896 (N_896,N_419,N_786);
nand U897 (N_897,N_699,N_541);
or U898 (N_898,N_777,N_454);
nand U899 (N_899,In_348,N_705);
nor U900 (N_900,N_817,N_813);
nor U901 (N_901,N_831,N_895);
nor U902 (N_902,N_841,N_865);
nand U903 (N_903,N_881,N_814);
or U904 (N_904,N_896,N_809);
nand U905 (N_905,N_882,N_869);
and U906 (N_906,N_816,N_825);
and U907 (N_907,N_892,N_802);
nand U908 (N_908,N_880,N_815);
xnor U909 (N_909,N_856,N_861);
or U910 (N_910,N_877,N_886);
nand U911 (N_911,N_822,N_842);
nand U912 (N_912,N_889,N_807);
nand U913 (N_913,N_828,N_875);
or U914 (N_914,N_862,N_832);
nor U915 (N_915,N_887,N_885);
nand U916 (N_916,N_894,N_805);
nor U917 (N_917,N_810,N_834);
nand U918 (N_918,N_888,N_849);
and U919 (N_919,N_863,N_883);
or U920 (N_920,N_812,N_843);
and U921 (N_921,N_873,N_840);
nor U922 (N_922,N_851,N_833);
and U923 (N_923,N_852,N_866);
and U924 (N_924,N_835,N_854);
or U925 (N_925,N_804,N_860);
nand U926 (N_926,N_820,N_848);
or U927 (N_927,N_872,N_879);
and U928 (N_928,N_824,N_839);
nand U929 (N_929,N_800,N_836);
or U930 (N_930,N_837,N_899);
nand U931 (N_931,N_857,N_827);
nand U932 (N_932,N_847,N_846);
or U933 (N_933,N_808,N_801);
and U934 (N_934,N_874,N_819);
nand U935 (N_935,N_890,N_878);
nor U936 (N_936,N_829,N_884);
nor U937 (N_937,N_870,N_898);
or U938 (N_938,N_844,N_803);
and U939 (N_939,N_838,N_876);
nor U940 (N_940,N_867,N_858);
and U941 (N_941,N_821,N_868);
nor U942 (N_942,N_864,N_859);
nor U943 (N_943,N_823,N_897);
or U944 (N_944,N_891,N_871);
nor U945 (N_945,N_893,N_811);
nand U946 (N_946,N_818,N_830);
nor U947 (N_947,N_855,N_826);
or U948 (N_948,N_845,N_853);
nor U949 (N_949,N_806,N_850);
nor U950 (N_950,N_803,N_823);
nor U951 (N_951,N_898,N_825);
and U952 (N_952,N_801,N_879);
and U953 (N_953,N_824,N_815);
nand U954 (N_954,N_886,N_896);
xor U955 (N_955,N_861,N_816);
nor U956 (N_956,N_894,N_885);
and U957 (N_957,N_832,N_872);
nor U958 (N_958,N_818,N_857);
and U959 (N_959,N_813,N_850);
and U960 (N_960,N_880,N_890);
or U961 (N_961,N_859,N_800);
nor U962 (N_962,N_837,N_821);
and U963 (N_963,N_815,N_854);
and U964 (N_964,N_844,N_878);
nand U965 (N_965,N_809,N_850);
or U966 (N_966,N_817,N_805);
and U967 (N_967,N_824,N_833);
or U968 (N_968,N_801,N_890);
nor U969 (N_969,N_824,N_814);
nor U970 (N_970,N_826,N_870);
nor U971 (N_971,N_834,N_800);
or U972 (N_972,N_805,N_898);
and U973 (N_973,N_898,N_822);
or U974 (N_974,N_853,N_837);
nor U975 (N_975,N_831,N_807);
nor U976 (N_976,N_871,N_850);
nor U977 (N_977,N_855,N_876);
nand U978 (N_978,N_832,N_817);
or U979 (N_979,N_863,N_888);
and U980 (N_980,N_888,N_806);
or U981 (N_981,N_899,N_836);
nor U982 (N_982,N_857,N_865);
and U983 (N_983,N_816,N_868);
nor U984 (N_984,N_830,N_890);
xor U985 (N_985,N_870,N_882);
nor U986 (N_986,N_899,N_848);
nor U987 (N_987,N_895,N_852);
or U988 (N_988,N_813,N_865);
or U989 (N_989,N_830,N_873);
or U990 (N_990,N_860,N_862);
or U991 (N_991,N_863,N_800);
nor U992 (N_992,N_897,N_804);
nor U993 (N_993,N_811,N_890);
or U994 (N_994,N_823,N_819);
or U995 (N_995,N_817,N_862);
and U996 (N_996,N_824,N_882);
or U997 (N_997,N_862,N_838);
nor U998 (N_998,N_807,N_858);
nand U999 (N_999,N_863,N_836);
and U1000 (N_1000,N_985,N_936);
or U1001 (N_1001,N_924,N_946);
or U1002 (N_1002,N_918,N_904);
or U1003 (N_1003,N_916,N_986);
and U1004 (N_1004,N_984,N_937);
and U1005 (N_1005,N_962,N_942);
nand U1006 (N_1006,N_954,N_959);
and U1007 (N_1007,N_909,N_975);
nor U1008 (N_1008,N_919,N_935);
nand U1009 (N_1009,N_926,N_928);
and U1010 (N_1010,N_901,N_950);
nor U1011 (N_1011,N_987,N_998);
and U1012 (N_1012,N_991,N_968);
nor U1013 (N_1013,N_972,N_903);
nand U1014 (N_1014,N_915,N_976);
nand U1015 (N_1015,N_902,N_995);
nor U1016 (N_1016,N_980,N_961);
and U1017 (N_1017,N_949,N_905);
or U1018 (N_1018,N_957,N_941);
nand U1019 (N_1019,N_993,N_933);
or U1020 (N_1020,N_944,N_953);
nand U1021 (N_1021,N_999,N_900);
and U1022 (N_1022,N_910,N_920);
or U1023 (N_1023,N_978,N_952);
nor U1024 (N_1024,N_965,N_955);
xnor U1025 (N_1025,N_994,N_948);
or U1026 (N_1026,N_982,N_956);
nor U1027 (N_1027,N_929,N_974);
and U1028 (N_1028,N_932,N_917);
and U1029 (N_1029,N_971,N_913);
or U1030 (N_1030,N_939,N_908);
nand U1031 (N_1031,N_911,N_964);
and U1032 (N_1032,N_973,N_990);
nand U1033 (N_1033,N_947,N_963);
or U1034 (N_1034,N_927,N_922);
or U1035 (N_1035,N_979,N_943);
or U1036 (N_1036,N_988,N_925);
and U1037 (N_1037,N_945,N_907);
or U1038 (N_1038,N_930,N_938);
nor U1039 (N_1039,N_923,N_921);
and U1040 (N_1040,N_983,N_960);
nand U1041 (N_1041,N_931,N_958);
nand U1042 (N_1042,N_906,N_981);
and U1043 (N_1043,N_914,N_970);
or U1044 (N_1044,N_934,N_992);
nand U1045 (N_1045,N_940,N_997);
or U1046 (N_1046,N_912,N_989);
nand U1047 (N_1047,N_977,N_951);
nand U1048 (N_1048,N_967,N_966);
or U1049 (N_1049,N_996,N_969);
or U1050 (N_1050,N_988,N_955);
nor U1051 (N_1051,N_906,N_927);
and U1052 (N_1052,N_956,N_957);
or U1053 (N_1053,N_918,N_944);
and U1054 (N_1054,N_926,N_978);
nand U1055 (N_1055,N_985,N_906);
nand U1056 (N_1056,N_912,N_984);
nor U1057 (N_1057,N_969,N_952);
and U1058 (N_1058,N_918,N_981);
or U1059 (N_1059,N_939,N_904);
or U1060 (N_1060,N_952,N_905);
or U1061 (N_1061,N_996,N_907);
nand U1062 (N_1062,N_978,N_982);
nand U1063 (N_1063,N_955,N_972);
nor U1064 (N_1064,N_970,N_910);
and U1065 (N_1065,N_979,N_946);
and U1066 (N_1066,N_957,N_962);
and U1067 (N_1067,N_981,N_950);
or U1068 (N_1068,N_907,N_905);
and U1069 (N_1069,N_911,N_955);
and U1070 (N_1070,N_952,N_946);
and U1071 (N_1071,N_925,N_924);
and U1072 (N_1072,N_934,N_942);
xnor U1073 (N_1073,N_933,N_929);
and U1074 (N_1074,N_991,N_979);
nand U1075 (N_1075,N_942,N_922);
and U1076 (N_1076,N_940,N_999);
nor U1077 (N_1077,N_937,N_990);
and U1078 (N_1078,N_944,N_972);
nand U1079 (N_1079,N_936,N_923);
xor U1080 (N_1080,N_929,N_951);
nand U1081 (N_1081,N_990,N_980);
nor U1082 (N_1082,N_971,N_923);
nor U1083 (N_1083,N_949,N_927);
nand U1084 (N_1084,N_989,N_959);
and U1085 (N_1085,N_936,N_946);
and U1086 (N_1086,N_906,N_902);
or U1087 (N_1087,N_907,N_952);
and U1088 (N_1088,N_929,N_948);
or U1089 (N_1089,N_904,N_980);
and U1090 (N_1090,N_924,N_993);
or U1091 (N_1091,N_973,N_998);
nor U1092 (N_1092,N_989,N_968);
nand U1093 (N_1093,N_992,N_911);
nand U1094 (N_1094,N_945,N_940);
nor U1095 (N_1095,N_982,N_901);
and U1096 (N_1096,N_970,N_917);
nor U1097 (N_1097,N_984,N_971);
and U1098 (N_1098,N_906,N_946);
nor U1099 (N_1099,N_952,N_989);
nand U1100 (N_1100,N_1041,N_1017);
and U1101 (N_1101,N_1030,N_1035);
and U1102 (N_1102,N_1077,N_1056);
nor U1103 (N_1103,N_1095,N_1043);
nor U1104 (N_1104,N_1065,N_1054);
nand U1105 (N_1105,N_1093,N_1085);
xor U1106 (N_1106,N_1063,N_1071);
nand U1107 (N_1107,N_1066,N_1004);
or U1108 (N_1108,N_1094,N_1036);
nand U1109 (N_1109,N_1020,N_1046);
nand U1110 (N_1110,N_1038,N_1087);
xnor U1111 (N_1111,N_1075,N_1044);
or U1112 (N_1112,N_1076,N_1096);
nand U1113 (N_1113,N_1073,N_1069);
and U1114 (N_1114,N_1008,N_1061);
nor U1115 (N_1115,N_1002,N_1082);
nor U1116 (N_1116,N_1012,N_1029);
nor U1117 (N_1117,N_1049,N_1070);
and U1118 (N_1118,N_1055,N_1081);
or U1119 (N_1119,N_1018,N_1089);
or U1120 (N_1120,N_1051,N_1007);
nand U1121 (N_1121,N_1060,N_1084);
or U1122 (N_1122,N_1067,N_1023);
nor U1123 (N_1123,N_1097,N_1003);
nand U1124 (N_1124,N_1011,N_1005);
and U1125 (N_1125,N_1016,N_1015);
nand U1126 (N_1126,N_1039,N_1025);
nand U1127 (N_1127,N_1074,N_1034);
and U1128 (N_1128,N_1006,N_1014);
nor U1129 (N_1129,N_1033,N_1042);
and U1130 (N_1130,N_1047,N_1083);
nand U1131 (N_1131,N_1013,N_1032);
nand U1132 (N_1132,N_1009,N_1080);
nand U1133 (N_1133,N_1068,N_1021);
nor U1134 (N_1134,N_1031,N_1057);
and U1135 (N_1135,N_1001,N_1079);
nor U1136 (N_1136,N_1010,N_1019);
nor U1137 (N_1137,N_1091,N_1072);
nand U1138 (N_1138,N_1000,N_1098);
or U1139 (N_1139,N_1027,N_1086);
nand U1140 (N_1140,N_1024,N_1062);
or U1141 (N_1141,N_1058,N_1092);
nand U1142 (N_1142,N_1045,N_1090);
nand U1143 (N_1143,N_1028,N_1022);
or U1144 (N_1144,N_1088,N_1064);
nor U1145 (N_1145,N_1040,N_1048);
and U1146 (N_1146,N_1078,N_1026);
nand U1147 (N_1147,N_1050,N_1053);
nor U1148 (N_1148,N_1037,N_1099);
nor U1149 (N_1149,N_1059,N_1052);
nor U1150 (N_1150,N_1010,N_1076);
nor U1151 (N_1151,N_1092,N_1045);
or U1152 (N_1152,N_1087,N_1068);
or U1153 (N_1153,N_1015,N_1017);
nand U1154 (N_1154,N_1016,N_1024);
xor U1155 (N_1155,N_1093,N_1055);
or U1156 (N_1156,N_1036,N_1026);
nor U1157 (N_1157,N_1075,N_1086);
nor U1158 (N_1158,N_1031,N_1078);
nor U1159 (N_1159,N_1029,N_1074);
and U1160 (N_1160,N_1059,N_1043);
nand U1161 (N_1161,N_1007,N_1064);
nand U1162 (N_1162,N_1047,N_1021);
nor U1163 (N_1163,N_1071,N_1043);
or U1164 (N_1164,N_1066,N_1029);
nand U1165 (N_1165,N_1049,N_1003);
nand U1166 (N_1166,N_1035,N_1012);
or U1167 (N_1167,N_1096,N_1089);
nor U1168 (N_1168,N_1083,N_1034);
nand U1169 (N_1169,N_1043,N_1081);
xnor U1170 (N_1170,N_1024,N_1025);
and U1171 (N_1171,N_1047,N_1099);
and U1172 (N_1172,N_1027,N_1059);
nand U1173 (N_1173,N_1021,N_1057);
and U1174 (N_1174,N_1069,N_1040);
nor U1175 (N_1175,N_1053,N_1094);
nor U1176 (N_1176,N_1027,N_1087);
and U1177 (N_1177,N_1069,N_1074);
or U1178 (N_1178,N_1002,N_1040);
nand U1179 (N_1179,N_1060,N_1088);
or U1180 (N_1180,N_1089,N_1054);
or U1181 (N_1181,N_1090,N_1058);
nand U1182 (N_1182,N_1023,N_1093);
nand U1183 (N_1183,N_1069,N_1081);
nor U1184 (N_1184,N_1000,N_1001);
xnor U1185 (N_1185,N_1051,N_1069);
nand U1186 (N_1186,N_1017,N_1092);
and U1187 (N_1187,N_1028,N_1025);
and U1188 (N_1188,N_1051,N_1084);
and U1189 (N_1189,N_1078,N_1049);
nor U1190 (N_1190,N_1036,N_1000);
nand U1191 (N_1191,N_1092,N_1085);
nor U1192 (N_1192,N_1096,N_1095);
and U1193 (N_1193,N_1088,N_1012);
and U1194 (N_1194,N_1099,N_1090);
and U1195 (N_1195,N_1093,N_1003);
nor U1196 (N_1196,N_1026,N_1097);
nor U1197 (N_1197,N_1057,N_1070);
nand U1198 (N_1198,N_1059,N_1080);
or U1199 (N_1199,N_1014,N_1023);
nor U1200 (N_1200,N_1199,N_1144);
and U1201 (N_1201,N_1106,N_1129);
nor U1202 (N_1202,N_1186,N_1125);
nor U1203 (N_1203,N_1198,N_1140);
xnor U1204 (N_1204,N_1176,N_1194);
nand U1205 (N_1205,N_1131,N_1151);
nand U1206 (N_1206,N_1178,N_1175);
and U1207 (N_1207,N_1180,N_1182);
or U1208 (N_1208,N_1128,N_1132);
nand U1209 (N_1209,N_1156,N_1184);
or U1210 (N_1210,N_1110,N_1142);
or U1211 (N_1211,N_1162,N_1164);
nand U1212 (N_1212,N_1113,N_1112);
nand U1213 (N_1213,N_1147,N_1121);
and U1214 (N_1214,N_1168,N_1173);
or U1215 (N_1215,N_1179,N_1152);
or U1216 (N_1216,N_1135,N_1123);
nor U1217 (N_1217,N_1104,N_1108);
nand U1218 (N_1218,N_1117,N_1133);
nor U1219 (N_1219,N_1185,N_1109);
or U1220 (N_1220,N_1195,N_1136);
or U1221 (N_1221,N_1177,N_1124);
and U1222 (N_1222,N_1158,N_1115);
nand U1223 (N_1223,N_1167,N_1174);
nand U1224 (N_1224,N_1100,N_1189);
and U1225 (N_1225,N_1134,N_1103);
nor U1226 (N_1226,N_1118,N_1146);
nand U1227 (N_1227,N_1171,N_1193);
nand U1228 (N_1228,N_1141,N_1165);
nor U1229 (N_1229,N_1122,N_1192);
nor U1230 (N_1230,N_1107,N_1150);
nand U1231 (N_1231,N_1196,N_1138);
and U1232 (N_1232,N_1130,N_1114);
or U1233 (N_1233,N_1127,N_1191);
and U1234 (N_1234,N_1161,N_1172);
and U1235 (N_1235,N_1197,N_1153);
nand U1236 (N_1236,N_1169,N_1120);
nor U1237 (N_1237,N_1159,N_1166);
nand U1238 (N_1238,N_1157,N_1190);
and U1239 (N_1239,N_1183,N_1163);
and U1240 (N_1240,N_1170,N_1137);
and U1241 (N_1241,N_1154,N_1143);
or U1242 (N_1242,N_1126,N_1101);
or U1243 (N_1243,N_1181,N_1119);
or U1244 (N_1244,N_1187,N_1139);
nand U1245 (N_1245,N_1105,N_1116);
and U1246 (N_1246,N_1102,N_1188);
or U1247 (N_1247,N_1149,N_1145);
or U1248 (N_1248,N_1111,N_1160);
xnor U1249 (N_1249,N_1155,N_1148);
and U1250 (N_1250,N_1149,N_1178);
nor U1251 (N_1251,N_1136,N_1115);
nor U1252 (N_1252,N_1153,N_1163);
nor U1253 (N_1253,N_1122,N_1152);
nor U1254 (N_1254,N_1128,N_1125);
and U1255 (N_1255,N_1115,N_1188);
and U1256 (N_1256,N_1177,N_1151);
or U1257 (N_1257,N_1174,N_1181);
and U1258 (N_1258,N_1160,N_1138);
and U1259 (N_1259,N_1195,N_1155);
and U1260 (N_1260,N_1120,N_1111);
and U1261 (N_1261,N_1147,N_1103);
nor U1262 (N_1262,N_1189,N_1176);
and U1263 (N_1263,N_1133,N_1145);
and U1264 (N_1264,N_1125,N_1179);
nand U1265 (N_1265,N_1157,N_1128);
or U1266 (N_1266,N_1192,N_1172);
nor U1267 (N_1267,N_1148,N_1193);
or U1268 (N_1268,N_1182,N_1194);
and U1269 (N_1269,N_1141,N_1146);
nor U1270 (N_1270,N_1163,N_1106);
nor U1271 (N_1271,N_1117,N_1100);
nand U1272 (N_1272,N_1183,N_1143);
and U1273 (N_1273,N_1179,N_1102);
and U1274 (N_1274,N_1151,N_1147);
or U1275 (N_1275,N_1113,N_1133);
or U1276 (N_1276,N_1166,N_1139);
and U1277 (N_1277,N_1143,N_1110);
nand U1278 (N_1278,N_1129,N_1186);
nor U1279 (N_1279,N_1173,N_1147);
and U1280 (N_1280,N_1164,N_1105);
or U1281 (N_1281,N_1156,N_1198);
and U1282 (N_1282,N_1171,N_1138);
or U1283 (N_1283,N_1154,N_1102);
nor U1284 (N_1284,N_1152,N_1153);
and U1285 (N_1285,N_1116,N_1152);
nor U1286 (N_1286,N_1137,N_1190);
nor U1287 (N_1287,N_1110,N_1138);
nand U1288 (N_1288,N_1115,N_1123);
nand U1289 (N_1289,N_1198,N_1130);
and U1290 (N_1290,N_1103,N_1116);
and U1291 (N_1291,N_1106,N_1122);
nor U1292 (N_1292,N_1128,N_1101);
and U1293 (N_1293,N_1146,N_1125);
nand U1294 (N_1294,N_1154,N_1155);
and U1295 (N_1295,N_1103,N_1179);
or U1296 (N_1296,N_1197,N_1169);
and U1297 (N_1297,N_1190,N_1152);
and U1298 (N_1298,N_1122,N_1116);
nor U1299 (N_1299,N_1150,N_1121);
nor U1300 (N_1300,N_1244,N_1288);
nor U1301 (N_1301,N_1215,N_1296);
or U1302 (N_1302,N_1269,N_1243);
nand U1303 (N_1303,N_1209,N_1247);
nor U1304 (N_1304,N_1241,N_1264);
and U1305 (N_1305,N_1218,N_1292);
and U1306 (N_1306,N_1285,N_1289);
or U1307 (N_1307,N_1283,N_1200);
nand U1308 (N_1308,N_1260,N_1256);
nor U1309 (N_1309,N_1263,N_1217);
and U1310 (N_1310,N_1298,N_1266);
nand U1311 (N_1311,N_1268,N_1282);
nor U1312 (N_1312,N_1223,N_1272);
nand U1313 (N_1313,N_1290,N_1253);
nand U1314 (N_1314,N_1291,N_1280);
nand U1315 (N_1315,N_1211,N_1220);
nor U1316 (N_1316,N_1208,N_1238);
and U1317 (N_1317,N_1229,N_1216);
xor U1318 (N_1318,N_1213,N_1237);
nand U1319 (N_1319,N_1259,N_1255);
nand U1320 (N_1320,N_1257,N_1245);
or U1321 (N_1321,N_1240,N_1284);
or U1322 (N_1322,N_1207,N_1203);
nand U1323 (N_1323,N_1222,N_1265);
or U1324 (N_1324,N_1230,N_1277);
or U1325 (N_1325,N_1239,N_1281);
and U1326 (N_1326,N_1219,N_1276);
nand U1327 (N_1327,N_1250,N_1231);
or U1328 (N_1328,N_1261,N_1214);
or U1329 (N_1329,N_1251,N_1294);
and U1330 (N_1330,N_1242,N_1299);
xnor U1331 (N_1331,N_1248,N_1297);
and U1332 (N_1332,N_1225,N_1236);
nand U1333 (N_1333,N_1267,N_1295);
nand U1334 (N_1334,N_1262,N_1202);
nor U1335 (N_1335,N_1226,N_1246);
and U1336 (N_1336,N_1293,N_1221);
and U1337 (N_1337,N_1287,N_1249);
or U1338 (N_1338,N_1279,N_1201);
nand U1339 (N_1339,N_1252,N_1270);
and U1340 (N_1340,N_1275,N_1271);
nor U1341 (N_1341,N_1286,N_1206);
or U1342 (N_1342,N_1228,N_1235);
nand U1343 (N_1343,N_1274,N_1234);
nor U1344 (N_1344,N_1254,N_1233);
nand U1345 (N_1345,N_1212,N_1205);
nand U1346 (N_1346,N_1232,N_1204);
or U1347 (N_1347,N_1273,N_1258);
and U1348 (N_1348,N_1210,N_1224);
nor U1349 (N_1349,N_1227,N_1278);
nor U1350 (N_1350,N_1263,N_1236);
nor U1351 (N_1351,N_1262,N_1228);
and U1352 (N_1352,N_1254,N_1202);
nand U1353 (N_1353,N_1253,N_1209);
and U1354 (N_1354,N_1220,N_1217);
nor U1355 (N_1355,N_1275,N_1280);
or U1356 (N_1356,N_1236,N_1282);
or U1357 (N_1357,N_1210,N_1234);
or U1358 (N_1358,N_1214,N_1217);
nand U1359 (N_1359,N_1234,N_1249);
and U1360 (N_1360,N_1254,N_1289);
or U1361 (N_1361,N_1295,N_1291);
nand U1362 (N_1362,N_1251,N_1237);
and U1363 (N_1363,N_1283,N_1263);
nor U1364 (N_1364,N_1259,N_1290);
and U1365 (N_1365,N_1237,N_1200);
and U1366 (N_1366,N_1283,N_1281);
or U1367 (N_1367,N_1275,N_1200);
nor U1368 (N_1368,N_1293,N_1246);
and U1369 (N_1369,N_1258,N_1248);
and U1370 (N_1370,N_1261,N_1242);
or U1371 (N_1371,N_1274,N_1264);
or U1372 (N_1372,N_1297,N_1227);
nor U1373 (N_1373,N_1226,N_1288);
nand U1374 (N_1374,N_1236,N_1270);
or U1375 (N_1375,N_1280,N_1233);
nand U1376 (N_1376,N_1294,N_1224);
nor U1377 (N_1377,N_1289,N_1216);
nor U1378 (N_1378,N_1284,N_1248);
and U1379 (N_1379,N_1299,N_1290);
nor U1380 (N_1380,N_1236,N_1227);
nand U1381 (N_1381,N_1295,N_1278);
nor U1382 (N_1382,N_1288,N_1225);
nand U1383 (N_1383,N_1286,N_1240);
or U1384 (N_1384,N_1257,N_1288);
and U1385 (N_1385,N_1240,N_1293);
and U1386 (N_1386,N_1237,N_1268);
and U1387 (N_1387,N_1214,N_1225);
or U1388 (N_1388,N_1293,N_1282);
nor U1389 (N_1389,N_1271,N_1262);
nand U1390 (N_1390,N_1219,N_1202);
nand U1391 (N_1391,N_1256,N_1291);
or U1392 (N_1392,N_1236,N_1261);
and U1393 (N_1393,N_1294,N_1220);
nand U1394 (N_1394,N_1273,N_1260);
or U1395 (N_1395,N_1236,N_1228);
nand U1396 (N_1396,N_1204,N_1280);
or U1397 (N_1397,N_1255,N_1238);
and U1398 (N_1398,N_1214,N_1245);
xnor U1399 (N_1399,N_1215,N_1283);
or U1400 (N_1400,N_1356,N_1331);
and U1401 (N_1401,N_1388,N_1307);
xor U1402 (N_1402,N_1363,N_1389);
and U1403 (N_1403,N_1302,N_1327);
or U1404 (N_1404,N_1304,N_1313);
or U1405 (N_1405,N_1306,N_1314);
nor U1406 (N_1406,N_1353,N_1396);
and U1407 (N_1407,N_1319,N_1318);
nand U1408 (N_1408,N_1374,N_1333);
and U1409 (N_1409,N_1394,N_1316);
and U1410 (N_1410,N_1383,N_1322);
nor U1411 (N_1411,N_1326,N_1395);
and U1412 (N_1412,N_1392,N_1336);
and U1413 (N_1413,N_1348,N_1323);
nand U1414 (N_1414,N_1352,N_1397);
or U1415 (N_1415,N_1376,N_1377);
nor U1416 (N_1416,N_1391,N_1305);
and U1417 (N_1417,N_1372,N_1347);
and U1418 (N_1418,N_1334,N_1330);
and U1419 (N_1419,N_1358,N_1345);
xnor U1420 (N_1420,N_1390,N_1384);
or U1421 (N_1421,N_1311,N_1328);
and U1422 (N_1422,N_1351,N_1310);
and U1423 (N_1423,N_1320,N_1321);
xor U1424 (N_1424,N_1369,N_1332);
nand U1425 (N_1425,N_1342,N_1338);
nand U1426 (N_1426,N_1367,N_1387);
and U1427 (N_1427,N_1381,N_1371);
and U1428 (N_1428,N_1300,N_1309);
and U1429 (N_1429,N_1350,N_1382);
nand U1430 (N_1430,N_1301,N_1341);
nand U1431 (N_1431,N_1379,N_1360);
nand U1432 (N_1432,N_1344,N_1315);
and U1433 (N_1433,N_1398,N_1349);
nor U1434 (N_1434,N_1308,N_1325);
nand U1435 (N_1435,N_1329,N_1386);
and U1436 (N_1436,N_1362,N_1312);
nor U1437 (N_1437,N_1368,N_1343);
nor U1438 (N_1438,N_1380,N_1339);
nand U1439 (N_1439,N_1340,N_1378);
nand U1440 (N_1440,N_1399,N_1365);
nor U1441 (N_1441,N_1355,N_1324);
nand U1442 (N_1442,N_1354,N_1335);
nand U1443 (N_1443,N_1393,N_1359);
nand U1444 (N_1444,N_1366,N_1370);
nor U1445 (N_1445,N_1303,N_1373);
and U1446 (N_1446,N_1364,N_1346);
nand U1447 (N_1447,N_1357,N_1337);
and U1448 (N_1448,N_1361,N_1317);
nand U1449 (N_1449,N_1385,N_1375);
nand U1450 (N_1450,N_1351,N_1390);
and U1451 (N_1451,N_1359,N_1370);
nor U1452 (N_1452,N_1367,N_1398);
nand U1453 (N_1453,N_1375,N_1384);
nand U1454 (N_1454,N_1308,N_1335);
or U1455 (N_1455,N_1369,N_1335);
and U1456 (N_1456,N_1318,N_1391);
nor U1457 (N_1457,N_1378,N_1335);
nand U1458 (N_1458,N_1301,N_1345);
or U1459 (N_1459,N_1357,N_1370);
nor U1460 (N_1460,N_1344,N_1332);
or U1461 (N_1461,N_1390,N_1348);
or U1462 (N_1462,N_1347,N_1323);
and U1463 (N_1463,N_1382,N_1344);
nand U1464 (N_1464,N_1369,N_1384);
nor U1465 (N_1465,N_1383,N_1396);
and U1466 (N_1466,N_1383,N_1366);
nand U1467 (N_1467,N_1342,N_1395);
nand U1468 (N_1468,N_1337,N_1304);
nand U1469 (N_1469,N_1324,N_1389);
and U1470 (N_1470,N_1312,N_1353);
nor U1471 (N_1471,N_1377,N_1319);
nor U1472 (N_1472,N_1384,N_1303);
and U1473 (N_1473,N_1348,N_1306);
and U1474 (N_1474,N_1349,N_1370);
and U1475 (N_1475,N_1323,N_1398);
xor U1476 (N_1476,N_1309,N_1310);
and U1477 (N_1477,N_1337,N_1321);
nor U1478 (N_1478,N_1336,N_1300);
nand U1479 (N_1479,N_1379,N_1312);
nand U1480 (N_1480,N_1382,N_1328);
nor U1481 (N_1481,N_1379,N_1307);
and U1482 (N_1482,N_1384,N_1372);
and U1483 (N_1483,N_1341,N_1330);
nand U1484 (N_1484,N_1367,N_1386);
or U1485 (N_1485,N_1350,N_1327);
or U1486 (N_1486,N_1378,N_1341);
or U1487 (N_1487,N_1333,N_1390);
and U1488 (N_1488,N_1362,N_1381);
xor U1489 (N_1489,N_1388,N_1351);
xor U1490 (N_1490,N_1345,N_1336);
nor U1491 (N_1491,N_1384,N_1332);
and U1492 (N_1492,N_1349,N_1315);
nor U1493 (N_1493,N_1370,N_1395);
nor U1494 (N_1494,N_1314,N_1373);
or U1495 (N_1495,N_1388,N_1304);
or U1496 (N_1496,N_1370,N_1345);
and U1497 (N_1497,N_1382,N_1341);
nor U1498 (N_1498,N_1311,N_1344);
nand U1499 (N_1499,N_1356,N_1306);
nand U1500 (N_1500,N_1406,N_1435);
nand U1501 (N_1501,N_1449,N_1465);
nor U1502 (N_1502,N_1453,N_1440);
or U1503 (N_1503,N_1450,N_1490);
and U1504 (N_1504,N_1411,N_1427);
nand U1505 (N_1505,N_1459,N_1455);
nor U1506 (N_1506,N_1495,N_1452);
nor U1507 (N_1507,N_1470,N_1423);
and U1508 (N_1508,N_1429,N_1408);
and U1509 (N_1509,N_1414,N_1428);
and U1510 (N_1510,N_1467,N_1448);
xor U1511 (N_1511,N_1461,N_1472);
and U1512 (N_1512,N_1463,N_1426);
or U1513 (N_1513,N_1476,N_1409);
and U1514 (N_1514,N_1473,N_1454);
and U1515 (N_1515,N_1415,N_1457);
or U1516 (N_1516,N_1486,N_1443);
nor U1517 (N_1517,N_1481,N_1488);
xor U1518 (N_1518,N_1474,N_1484);
and U1519 (N_1519,N_1422,N_1458);
or U1520 (N_1520,N_1413,N_1441);
and U1521 (N_1521,N_1492,N_1477);
nor U1522 (N_1522,N_1498,N_1404);
xnor U1523 (N_1523,N_1478,N_1410);
and U1524 (N_1524,N_1419,N_1451);
nor U1525 (N_1525,N_1479,N_1420);
and U1526 (N_1526,N_1487,N_1462);
and U1527 (N_1527,N_1497,N_1482);
or U1528 (N_1528,N_1436,N_1468);
nand U1529 (N_1529,N_1432,N_1433);
nor U1530 (N_1530,N_1489,N_1456);
nor U1531 (N_1531,N_1421,N_1412);
nor U1532 (N_1532,N_1400,N_1496);
or U1533 (N_1533,N_1445,N_1439);
and U1534 (N_1534,N_1447,N_1464);
xnor U1535 (N_1535,N_1469,N_1460);
or U1536 (N_1536,N_1437,N_1444);
nor U1537 (N_1537,N_1494,N_1446);
or U1538 (N_1538,N_1493,N_1475);
nand U1539 (N_1539,N_1424,N_1402);
nand U1540 (N_1540,N_1438,N_1418);
and U1541 (N_1541,N_1431,N_1407);
nand U1542 (N_1542,N_1483,N_1434);
or U1543 (N_1543,N_1416,N_1485);
nand U1544 (N_1544,N_1405,N_1425);
and U1545 (N_1545,N_1401,N_1442);
and U1546 (N_1546,N_1417,N_1403);
nand U1547 (N_1547,N_1471,N_1466);
nand U1548 (N_1548,N_1499,N_1480);
nand U1549 (N_1549,N_1491,N_1430);
nand U1550 (N_1550,N_1480,N_1441);
nor U1551 (N_1551,N_1429,N_1417);
and U1552 (N_1552,N_1410,N_1418);
and U1553 (N_1553,N_1423,N_1416);
or U1554 (N_1554,N_1492,N_1443);
and U1555 (N_1555,N_1432,N_1417);
nor U1556 (N_1556,N_1454,N_1453);
or U1557 (N_1557,N_1437,N_1415);
nand U1558 (N_1558,N_1410,N_1464);
or U1559 (N_1559,N_1421,N_1420);
and U1560 (N_1560,N_1420,N_1442);
nor U1561 (N_1561,N_1494,N_1403);
nand U1562 (N_1562,N_1470,N_1457);
nand U1563 (N_1563,N_1420,N_1453);
or U1564 (N_1564,N_1444,N_1422);
or U1565 (N_1565,N_1457,N_1405);
and U1566 (N_1566,N_1435,N_1458);
nor U1567 (N_1567,N_1447,N_1432);
or U1568 (N_1568,N_1489,N_1424);
or U1569 (N_1569,N_1406,N_1480);
and U1570 (N_1570,N_1403,N_1496);
and U1571 (N_1571,N_1452,N_1474);
or U1572 (N_1572,N_1448,N_1426);
and U1573 (N_1573,N_1484,N_1469);
xnor U1574 (N_1574,N_1485,N_1479);
nor U1575 (N_1575,N_1406,N_1492);
or U1576 (N_1576,N_1468,N_1477);
or U1577 (N_1577,N_1407,N_1452);
or U1578 (N_1578,N_1461,N_1487);
xnor U1579 (N_1579,N_1412,N_1492);
or U1580 (N_1580,N_1449,N_1479);
or U1581 (N_1581,N_1423,N_1499);
and U1582 (N_1582,N_1421,N_1443);
nor U1583 (N_1583,N_1410,N_1433);
nand U1584 (N_1584,N_1474,N_1465);
nor U1585 (N_1585,N_1498,N_1466);
nand U1586 (N_1586,N_1420,N_1474);
nor U1587 (N_1587,N_1439,N_1424);
nand U1588 (N_1588,N_1413,N_1475);
nor U1589 (N_1589,N_1481,N_1441);
nor U1590 (N_1590,N_1438,N_1406);
and U1591 (N_1591,N_1467,N_1476);
and U1592 (N_1592,N_1451,N_1403);
nand U1593 (N_1593,N_1460,N_1483);
nor U1594 (N_1594,N_1418,N_1478);
and U1595 (N_1595,N_1401,N_1495);
or U1596 (N_1596,N_1443,N_1480);
nand U1597 (N_1597,N_1470,N_1492);
xnor U1598 (N_1598,N_1459,N_1475);
nand U1599 (N_1599,N_1428,N_1465);
and U1600 (N_1600,N_1558,N_1565);
or U1601 (N_1601,N_1572,N_1567);
nor U1602 (N_1602,N_1546,N_1516);
or U1603 (N_1603,N_1573,N_1592);
and U1604 (N_1604,N_1511,N_1559);
or U1605 (N_1605,N_1543,N_1579);
nand U1606 (N_1606,N_1535,N_1522);
and U1607 (N_1607,N_1588,N_1533);
nor U1608 (N_1608,N_1518,N_1561);
nor U1609 (N_1609,N_1508,N_1564);
or U1610 (N_1610,N_1523,N_1506);
and U1611 (N_1611,N_1589,N_1540);
nand U1612 (N_1612,N_1525,N_1545);
and U1613 (N_1613,N_1570,N_1531);
nand U1614 (N_1614,N_1555,N_1552);
and U1615 (N_1615,N_1590,N_1503);
or U1616 (N_1616,N_1593,N_1514);
or U1617 (N_1617,N_1556,N_1594);
and U1618 (N_1618,N_1560,N_1526);
nor U1619 (N_1619,N_1544,N_1517);
and U1620 (N_1620,N_1513,N_1549);
nand U1621 (N_1621,N_1521,N_1574);
nand U1622 (N_1622,N_1548,N_1571);
nand U1623 (N_1623,N_1586,N_1537);
nor U1624 (N_1624,N_1524,N_1542);
nand U1625 (N_1625,N_1566,N_1541);
or U1626 (N_1626,N_1585,N_1597);
nor U1627 (N_1627,N_1528,N_1504);
or U1628 (N_1628,N_1500,N_1539);
and U1629 (N_1629,N_1582,N_1512);
or U1630 (N_1630,N_1563,N_1534);
and U1631 (N_1631,N_1554,N_1562);
nand U1632 (N_1632,N_1584,N_1507);
nand U1633 (N_1633,N_1532,N_1595);
and U1634 (N_1634,N_1520,N_1553);
or U1635 (N_1635,N_1596,N_1530);
nand U1636 (N_1636,N_1578,N_1501);
nor U1637 (N_1637,N_1527,N_1529);
and U1638 (N_1638,N_1568,N_1575);
and U1639 (N_1639,N_1557,N_1505);
nor U1640 (N_1640,N_1550,N_1519);
nor U1641 (N_1641,N_1538,N_1599);
nand U1642 (N_1642,N_1583,N_1576);
nor U1643 (N_1643,N_1551,N_1569);
and U1644 (N_1644,N_1580,N_1598);
nor U1645 (N_1645,N_1502,N_1587);
nand U1646 (N_1646,N_1591,N_1510);
nor U1647 (N_1647,N_1515,N_1581);
nand U1648 (N_1648,N_1509,N_1577);
or U1649 (N_1649,N_1536,N_1547);
nand U1650 (N_1650,N_1537,N_1551);
nand U1651 (N_1651,N_1521,N_1544);
or U1652 (N_1652,N_1591,N_1541);
nor U1653 (N_1653,N_1556,N_1571);
or U1654 (N_1654,N_1592,N_1588);
or U1655 (N_1655,N_1565,N_1514);
or U1656 (N_1656,N_1539,N_1531);
nor U1657 (N_1657,N_1598,N_1514);
xnor U1658 (N_1658,N_1504,N_1580);
or U1659 (N_1659,N_1536,N_1527);
nand U1660 (N_1660,N_1581,N_1595);
or U1661 (N_1661,N_1554,N_1565);
xor U1662 (N_1662,N_1593,N_1542);
or U1663 (N_1663,N_1535,N_1548);
or U1664 (N_1664,N_1529,N_1509);
and U1665 (N_1665,N_1582,N_1589);
nand U1666 (N_1666,N_1528,N_1594);
or U1667 (N_1667,N_1559,N_1502);
and U1668 (N_1668,N_1538,N_1522);
xor U1669 (N_1669,N_1515,N_1578);
nand U1670 (N_1670,N_1536,N_1590);
and U1671 (N_1671,N_1571,N_1578);
and U1672 (N_1672,N_1531,N_1576);
nor U1673 (N_1673,N_1586,N_1569);
nand U1674 (N_1674,N_1561,N_1556);
nand U1675 (N_1675,N_1511,N_1595);
nor U1676 (N_1676,N_1539,N_1529);
or U1677 (N_1677,N_1507,N_1564);
and U1678 (N_1678,N_1541,N_1585);
nand U1679 (N_1679,N_1595,N_1531);
or U1680 (N_1680,N_1503,N_1575);
nand U1681 (N_1681,N_1543,N_1549);
nor U1682 (N_1682,N_1580,N_1511);
nand U1683 (N_1683,N_1598,N_1510);
and U1684 (N_1684,N_1537,N_1592);
or U1685 (N_1685,N_1548,N_1552);
nand U1686 (N_1686,N_1583,N_1575);
nor U1687 (N_1687,N_1532,N_1551);
nand U1688 (N_1688,N_1537,N_1506);
nand U1689 (N_1689,N_1507,N_1574);
or U1690 (N_1690,N_1561,N_1538);
nor U1691 (N_1691,N_1599,N_1578);
nor U1692 (N_1692,N_1568,N_1500);
and U1693 (N_1693,N_1519,N_1564);
nor U1694 (N_1694,N_1593,N_1573);
nand U1695 (N_1695,N_1500,N_1529);
or U1696 (N_1696,N_1559,N_1545);
nor U1697 (N_1697,N_1509,N_1512);
and U1698 (N_1698,N_1507,N_1573);
nand U1699 (N_1699,N_1527,N_1514);
and U1700 (N_1700,N_1680,N_1614);
or U1701 (N_1701,N_1675,N_1636);
nor U1702 (N_1702,N_1628,N_1606);
nand U1703 (N_1703,N_1655,N_1687);
nand U1704 (N_1704,N_1663,N_1641);
nand U1705 (N_1705,N_1623,N_1604);
or U1706 (N_1706,N_1624,N_1658);
nand U1707 (N_1707,N_1661,N_1686);
nor U1708 (N_1708,N_1677,N_1601);
nand U1709 (N_1709,N_1692,N_1647);
xnor U1710 (N_1710,N_1691,N_1632);
nor U1711 (N_1711,N_1670,N_1625);
or U1712 (N_1712,N_1668,N_1613);
xnor U1713 (N_1713,N_1630,N_1695);
or U1714 (N_1714,N_1683,N_1649);
nand U1715 (N_1715,N_1685,N_1689);
nand U1716 (N_1716,N_1694,N_1699);
nand U1717 (N_1717,N_1669,N_1671);
or U1718 (N_1718,N_1605,N_1678);
and U1719 (N_1719,N_1667,N_1611);
nor U1720 (N_1720,N_1642,N_1618);
or U1721 (N_1721,N_1620,N_1674);
nor U1722 (N_1722,N_1634,N_1697);
nand U1723 (N_1723,N_1646,N_1629);
nor U1724 (N_1724,N_1653,N_1603);
nand U1725 (N_1725,N_1682,N_1673);
nor U1726 (N_1726,N_1631,N_1676);
nand U1727 (N_1727,N_1638,N_1600);
nor U1728 (N_1728,N_1688,N_1693);
or U1729 (N_1729,N_1608,N_1684);
nor U1730 (N_1730,N_1652,N_1657);
and U1731 (N_1731,N_1660,N_1609);
nand U1732 (N_1732,N_1626,N_1654);
nor U1733 (N_1733,N_1698,N_1635);
nor U1734 (N_1734,N_1664,N_1662);
or U1735 (N_1735,N_1643,N_1679);
and U1736 (N_1736,N_1659,N_1621);
nand U1737 (N_1737,N_1619,N_1645);
nand U1738 (N_1738,N_1672,N_1650);
or U1739 (N_1739,N_1651,N_1612);
or U1740 (N_1740,N_1627,N_1696);
or U1741 (N_1741,N_1656,N_1666);
nand U1742 (N_1742,N_1639,N_1622);
and U1743 (N_1743,N_1644,N_1690);
or U1744 (N_1744,N_1648,N_1640);
nand U1745 (N_1745,N_1615,N_1637);
nor U1746 (N_1746,N_1633,N_1607);
and U1747 (N_1747,N_1617,N_1602);
and U1748 (N_1748,N_1616,N_1665);
nor U1749 (N_1749,N_1610,N_1681);
or U1750 (N_1750,N_1604,N_1651);
nor U1751 (N_1751,N_1627,N_1622);
nand U1752 (N_1752,N_1667,N_1640);
xnor U1753 (N_1753,N_1698,N_1661);
nor U1754 (N_1754,N_1638,N_1672);
nor U1755 (N_1755,N_1634,N_1685);
nor U1756 (N_1756,N_1633,N_1650);
xor U1757 (N_1757,N_1625,N_1675);
nand U1758 (N_1758,N_1693,N_1669);
nand U1759 (N_1759,N_1608,N_1607);
xnor U1760 (N_1760,N_1692,N_1603);
and U1761 (N_1761,N_1605,N_1624);
nand U1762 (N_1762,N_1678,N_1667);
xnor U1763 (N_1763,N_1643,N_1622);
nand U1764 (N_1764,N_1687,N_1646);
nor U1765 (N_1765,N_1665,N_1690);
nor U1766 (N_1766,N_1645,N_1666);
and U1767 (N_1767,N_1689,N_1633);
nand U1768 (N_1768,N_1627,N_1632);
and U1769 (N_1769,N_1609,N_1654);
nand U1770 (N_1770,N_1635,N_1641);
xor U1771 (N_1771,N_1635,N_1666);
or U1772 (N_1772,N_1693,N_1668);
nor U1773 (N_1773,N_1688,N_1670);
or U1774 (N_1774,N_1634,N_1614);
and U1775 (N_1775,N_1685,N_1614);
and U1776 (N_1776,N_1608,N_1616);
nor U1777 (N_1777,N_1684,N_1647);
nand U1778 (N_1778,N_1616,N_1684);
and U1779 (N_1779,N_1697,N_1686);
nor U1780 (N_1780,N_1649,N_1621);
or U1781 (N_1781,N_1643,N_1616);
nand U1782 (N_1782,N_1605,N_1630);
nor U1783 (N_1783,N_1616,N_1654);
xor U1784 (N_1784,N_1641,N_1604);
nand U1785 (N_1785,N_1614,N_1648);
or U1786 (N_1786,N_1678,N_1612);
or U1787 (N_1787,N_1659,N_1694);
or U1788 (N_1788,N_1632,N_1651);
nor U1789 (N_1789,N_1684,N_1665);
nand U1790 (N_1790,N_1624,N_1639);
nand U1791 (N_1791,N_1673,N_1638);
or U1792 (N_1792,N_1658,N_1625);
nor U1793 (N_1793,N_1632,N_1679);
nand U1794 (N_1794,N_1609,N_1617);
and U1795 (N_1795,N_1653,N_1654);
and U1796 (N_1796,N_1668,N_1681);
nand U1797 (N_1797,N_1644,N_1632);
nor U1798 (N_1798,N_1697,N_1613);
nand U1799 (N_1799,N_1622,N_1646);
nor U1800 (N_1800,N_1703,N_1766);
nor U1801 (N_1801,N_1758,N_1734);
or U1802 (N_1802,N_1738,N_1781);
or U1803 (N_1803,N_1792,N_1719);
nor U1804 (N_1804,N_1716,N_1749);
and U1805 (N_1805,N_1713,N_1731);
nor U1806 (N_1806,N_1722,N_1712);
nand U1807 (N_1807,N_1753,N_1701);
xor U1808 (N_1808,N_1770,N_1721);
or U1809 (N_1809,N_1797,N_1736);
or U1810 (N_1810,N_1710,N_1752);
or U1811 (N_1811,N_1704,N_1735);
nand U1812 (N_1812,N_1720,N_1709);
nand U1813 (N_1813,N_1795,N_1785);
nand U1814 (N_1814,N_1706,N_1774);
nor U1815 (N_1815,N_1776,N_1725);
and U1816 (N_1816,N_1786,N_1724);
nand U1817 (N_1817,N_1760,N_1796);
nor U1818 (N_1818,N_1778,N_1788);
and U1819 (N_1819,N_1787,N_1764);
xnor U1820 (N_1820,N_1798,N_1775);
or U1821 (N_1821,N_1723,N_1777);
nand U1822 (N_1822,N_1747,N_1705);
nand U1823 (N_1823,N_1744,N_1780);
or U1824 (N_1824,N_1793,N_1732);
nor U1825 (N_1825,N_1779,N_1757);
and U1826 (N_1826,N_1761,N_1729);
and U1827 (N_1827,N_1771,N_1754);
nor U1828 (N_1828,N_1790,N_1737);
or U1829 (N_1829,N_1794,N_1750);
nor U1830 (N_1830,N_1784,N_1759);
nor U1831 (N_1831,N_1772,N_1783);
nor U1832 (N_1832,N_1782,N_1700);
xnor U1833 (N_1833,N_1773,N_1741);
and U1834 (N_1834,N_1799,N_1730);
nor U1835 (N_1835,N_1718,N_1791);
and U1836 (N_1836,N_1768,N_1742);
and U1837 (N_1837,N_1746,N_1748);
or U1838 (N_1838,N_1756,N_1733);
nor U1839 (N_1839,N_1739,N_1726);
and U1840 (N_1840,N_1715,N_1711);
nor U1841 (N_1841,N_1707,N_1743);
nor U1842 (N_1842,N_1763,N_1767);
nand U1843 (N_1843,N_1765,N_1769);
or U1844 (N_1844,N_1755,N_1702);
xor U1845 (N_1845,N_1751,N_1762);
nor U1846 (N_1846,N_1714,N_1717);
or U1847 (N_1847,N_1789,N_1727);
or U1848 (N_1848,N_1745,N_1708);
or U1849 (N_1849,N_1740,N_1728);
nand U1850 (N_1850,N_1707,N_1741);
and U1851 (N_1851,N_1783,N_1770);
or U1852 (N_1852,N_1795,N_1772);
or U1853 (N_1853,N_1781,N_1715);
or U1854 (N_1854,N_1778,N_1789);
nand U1855 (N_1855,N_1747,N_1736);
or U1856 (N_1856,N_1765,N_1733);
nor U1857 (N_1857,N_1794,N_1766);
nand U1858 (N_1858,N_1790,N_1726);
xor U1859 (N_1859,N_1796,N_1737);
and U1860 (N_1860,N_1771,N_1741);
nand U1861 (N_1861,N_1730,N_1779);
nand U1862 (N_1862,N_1739,N_1799);
or U1863 (N_1863,N_1770,N_1792);
or U1864 (N_1864,N_1706,N_1714);
or U1865 (N_1865,N_1735,N_1788);
nor U1866 (N_1866,N_1707,N_1727);
and U1867 (N_1867,N_1734,N_1727);
nand U1868 (N_1868,N_1784,N_1771);
nand U1869 (N_1869,N_1709,N_1797);
nor U1870 (N_1870,N_1708,N_1794);
nand U1871 (N_1871,N_1720,N_1727);
nand U1872 (N_1872,N_1749,N_1700);
or U1873 (N_1873,N_1780,N_1726);
nand U1874 (N_1874,N_1759,N_1701);
and U1875 (N_1875,N_1708,N_1795);
nor U1876 (N_1876,N_1770,N_1729);
and U1877 (N_1877,N_1720,N_1724);
nand U1878 (N_1878,N_1762,N_1754);
and U1879 (N_1879,N_1775,N_1746);
or U1880 (N_1880,N_1761,N_1723);
and U1881 (N_1881,N_1770,N_1745);
and U1882 (N_1882,N_1726,N_1743);
xor U1883 (N_1883,N_1732,N_1768);
nand U1884 (N_1884,N_1797,N_1741);
nor U1885 (N_1885,N_1716,N_1724);
nor U1886 (N_1886,N_1767,N_1703);
xnor U1887 (N_1887,N_1749,N_1720);
and U1888 (N_1888,N_1702,N_1719);
nand U1889 (N_1889,N_1794,N_1733);
and U1890 (N_1890,N_1723,N_1709);
or U1891 (N_1891,N_1761,N_1763);
nand U1892 (N_1892,N_1754,N_1782);
xor U1893 (N_1893,N_1759,N_1715);
and U1894 (N_1894,N_1736,N_1787);
nor U1895 (N_1895,N_1736,N_1714);
or U1896 (N_1896,N_1797,N_1778);
nor U1897 (N_1897,N_1754,N_1700);
or U1898 (N_1898,N_1739,N_1704);
or U1899 (N_1899,N_1785,N_1787);
or U1900 (N_1900,N_1818,N_1834);
nand U1901 (N_1901,N_1893,N_1832);
or U1902 (N_1902,N_1807,N_1876);
nand U1903 (N_1903,N_1825,N_1864);
nand U1904 (N_1904,N_1803,N_1846);
nand U1905 (N_1905,N_1894,N_1851);
and U1906 (N_1906,N_1840,N_1830);
or U1907 (N_1907,N_1854,N_1861);
and U1908 (N_1908,N_1859,N_1812);
nand U1909 (N_1909,N_1889,N_1801);
or U1910 (N_1910,N_1831,N_1858);
and U1911 (N_1911,N_1815,N_1848);
nand U1912 (N_1912,N_1808,N_1880);
nor U1913 (N_1913,N_1870,N_1881);
nand U1914 (N_1914,N_1836,N_1860);
and U1915 (N_1915,N_1865,N_1823);
nand U1916 (N_1916,N_1822,N_1849);
and U1917 (N_1917,N_1891,N_1814);
or U1918 (N_1918,N_1843,N_1852);
and U1919 (N_1919,N_1820,N_1857);
xnor U1920 (N_1920,N_1885,N_1863);
nand U1921 (N_1921,N_1816,N_1838);
and U1922 (N_1922,N_1833,N_1883);
and U1923 (N_1923,N_1887,N_1827);
and U1924 (N_1924,N_1829,N_1804);
nor U1925 (N_1925,N_1895,N_1844);
nand U1926 (N_1926,N_1810,N_1875);
or U1927 (N_1927,N_1826,N_1839);
or U1928 (N_1928,N_1837,N_1888);
and U1929 (N_1929,N_1805,N_1811);
or U1930 (N_1930,N_1853,N_1882);
or U1931 (N_1931,N_1845,N_1897);
nand U1932 (N_1932,N_1856,N_1842);
or U1933 (N_1933,N_1873,N_1877);
nand U1934 (N_1934,N_1819,N_1813);
and U1935 (N_1935,N_1872,N_1874);
nand U1936 (N_1936,N_1828,N_1806);
or U1937 (N_1937,N_1886,N_1824);
or U1938 (N_1938,N_1817,N_1871);
and U1939 (N_1939,N_1800,N_1868);
and U1940 (N_1940,N_1890,N_1878);
nand U1941 (N_1941,N_1869,N_1809);
or U1942 (N_1942,N_1850,N_1847);
nor U1943 (N_1943,N_1835,N_1892);
or U1944 (N_1944,N_1866,N_1896);
nand U1945 (N_1945,N_1899,N_1884);
and U1946 (N_1946,N_1879,N_1898);
and U1947 (N_1947,N_1862,N_1841);
nand U1948 (N_1948,N_1867,N_1855);
or U1949 (N_1949,N_1821,N_1802);
and U1950 (N_1950,N_1828,N_1823);
and U1951 (N_1951,N_1833,N_1857);
and U1952 (N_1952,N_1849,N_1861);
or U1953 (N_1953,N_1811,N_1859);
nand U1954 (N_1954,N_1893,N_1862);
nor U1955 (N_1955,N_1888,N_1847);
or U1956 (N_1956,N_1807,N_1866);
or U1957 (N_1957,N_1834,N_1814);
and U1958 (N_1958,N_1840,N_1815);
or U1959 (N_1959,N_1826,N_1892);
and U1960 (N_1960,N_1894,N_1891);
or U1961 (N_1961,N_1813,N_1824);
or U1962 (N_1962,N_1882,N_1831);
or U1963 (N_1963,N_1831,N_1826);
and U1964 (N_1964,N_1897,N_1894);
and U1965 (N_1965,N_1843,N_1872);
or U1966 (N_1966,N_1824,N_1838);
or U1967 (N_1967,N_1864,N_1888);
nor U1968 (N_1968,N_1839,N_1824);
nor U1969 (N_1969,N_1861,N_1865);
or U1970 (N_1970,N_1864,N_1814);
nand U1971 (N_1971,N_1837,N_1816);
or U1972 (N_1972,N_1814,N_1805);
nand U1973 (N_1973,N_1827,N_1893);
nand U1974 (N_1974,N_1816,N_1889);
nand U1975 (N_1975,N_1875,N_1866);
or U1976 (N_1976,N_1848,N_1887);
nor U1977 (N_1977,N_1834,N_1835);
and U1978 (N_1978,N_1867,N_1854);
and U1979 (N_1979,N_1835,N_1866);
or U1980 (N_1980,N_1883,N_1840);
or U1981 (N_1981,N_1839,N_1811);
nand U1982 (N_1982,N_1871,N_1814);
nand U1983 (N_1983,N_1893,N_1836);
nor U1984 (N_1984,N_1822,N_1830);
nor U1985 (N_1985,N_1801,N_1808);
nand U1986 (N_1986,N_1851,N_1845);
nand U1987 (N_1987,N_1874,N_1885);
nand U1988 (N_1988,N_1853,N_1811);
and U1989 (N_1989,N_1829,N_1858);
or U1990 (N_1990,N_1889,N_1891);
xnor U1991 (N_1991,N_1869,N_1860);
or U1992 (N_1992,N_1844,N_1894);
and U1993 (N_1993,N_1871,N_1838);
nor U1994 (N_1994,N_1836,N_1822);
or U1995 (N_1995,N_1858,N_1836);
nand U1996 (N_1996,N_1854,N_1884);
nand U1997 (N_1997,N_1837,N_1851);
nor U1998 (N_1998,N_1877,N_1818);
nor U1999 (N_1999,N_1853,N_1849);
and U2000 (N_2000,N_1924,N_1977);
and U2001 (N_2001,N_1964,N_1984);
nor U2002 (N_2002,N_1969,N_1986);
or U2003 (N_2003,N_1908,N_1985);
or U2004 (N_2004,N_1975,N_1988);
nor U2005 (N_2005,N_1935,N_1947);
nand U2006 (N_2006,N_1958,N_1913);
or U2007 (N_2007,N_1952,N_1925);
and U2008 (N_2008,N_1941,N_1966);
or U2009 (N_2009,N_1983,N_1906);
and U2010 (N_2010,N_1973,N_1938);
and U2011 (N_2011,N_1903,N_1981);
nand U2012 (N_2012,N_1956,N_1979);
or U2013 (N_2013,N_1960,N_1946);
nand U2014 (N_2014,N_1959,N_1912);
nor U2015 (N_2015,N_1997,N_1901);
and U2016 (N_2016,N_1921,N_1950);
or U2017 (N_2017,N_1982,N_1992);
nand U2018 (N_2018,N_1954,N_1961);
and U2019 (N_2019,N_1926,N_1914);
and U2020 (N_2020,N_1905,N_1920);
or U2021 (N_2021,N_1939,N_1917);
nor U2022 (N_2022,N_1937,N_1970);
nor U2023 (N_2023,N_1934,N_1991);
nand U2024 (N_2024,N_1929,N_1972);
and U2025 (N_2025,N_1907,N_1930);
nand U2026 (N_2026,N_1900,N_1932);
nor U2027 (N_2027,N_1927,N_1944);
or U2028 (N_2028,N_1918,N_1990);
or U2029 (N_2029,N_1989,N_1994);
xor U2030 (N_2030,N_1936,N_1957);
and U2031 (N_2031,N_1922,N_1987);
and U2032 (N_2032,N_1971,N_1909);
nor U2033 (N_2033,N_1902,N_1996);
or U2034 (N_2034,N_1948,N_1923);
nor U2035 (N_2035,N_1962,N_1963);
nand U2036 (N_2036,N_1998,N_1945);
and U2037 (N_2037,N_1978,N_1955);
nor U2038 (N_2038,N_1940,N_1931);
nor U2039 (N_2039,N_1974,N_1953);
and U2040 (N_2040,N_1949,N_1993);
nor U2041 (N_2041,N_1968,N_1999);
and U2042 (N_2042,N_1928,N_1995);
nand U2043 (N_2043,N_1980,N_1967);
nor U2044 (N_2044,N_1919,N_1904);
or U2045 (N_2045,N_1910,N_1951);
or U2046 (N_2046,N_1943,N_1911);
or U2047 (N_2047,N_1916,N_1965);
nand U2048 (N_2048,N_1942,N_1976);
nand U2049 (N_2049,N_1915,N_1933);
xnor U2050 (N_2050,N_1996,N_1948);
nand U2051 (N_2051,N_1940,N_1936);
and U2052 (N_2052,N_1989,N_1991);
and U2053 (N_2053,N_1908,N_1963);
nor U2054 (N_2054,N_1971,N_1946);
and U2055 (N_2055,N_1939,N_1936);
or U2056 (N_2056,N_1965,N_1914);
nor U2057 (N_2057,N_1920,N_1993);
and U2058 (N_2058,N_1976,N_1999);
nor U2059 (N_2059,N_1932,N_1951);
and U2060 (N_2060,N_1918,N_1970);
nor U2061 (N_2061,N_1963,N_1967);
or U2062 (N_2062,N_1998,N_1973);
and U2063 (N_2063,N_1985,N_1992);
and U2064 (N_2064,N_1954,N_1930);
or U2065 (N_2065,N_1948,N_1922);
and U2066 (N_2066,N_1900,N_1924);
or U2067 (N_2067,N_1947,N_1985);
or U2068 (N_2068,N_1998,N_1924);
xnor U2069 (N_2069,N_1947,N_1975);
nor U2070 (N_2070,N_1972,N_1977);
nor U2071 (N_2071,N_1977,N_1921);
or U2072 (N_2072,N_1946,N_1915);
nor U2073 (N_2073,N_1908,N_1918);
xnor U2074 (N_2074,N_1970,N_1950);
nor U2075 (N_2075,N_1924,N_1995);
or U2076 (N_2076,N_1943,N_1976);
nand U2077 (N_2077,N_1969,N_1923);
or U2078 (N_2078,N_1933,N_1998);
or U2079 (N_2079,N_1955,N_1988);
and U2080 (N_2080,N_1967,N_1971);
xor U2081 (N_2081,N_1934,N_1924);
nand U2082 (N_2082,N_1911,N_1982);
or U2083 (N_2083,N_1977,N_1938);
and U2084 (N_2084,N_1961,N_1975);
and U2085 (N_2085,N_1983,N_1937);
nor U2086 (N_2086,N_1929,N_1997);
or U2087 (N_2087,N_1930,N_1932);
and U2088 (N_2088,N_1944,N_1946);
nand U2089 (N_2089,N_1977,N_1982);
or U2090 (N_2090,N_1906,N_1931);
nand U2091 (N_2091,N_1937,N_1901);
or U2092 (N_2092,N_1925,N_1923);
and U2093 (N_2093,N_1994,N_1946);
xor U2094 (N_2094,N_1911,N_1994);
or U2095 (N_2095,N_1950,N_1986);
and U2096 (N_2096,N_1914,N_1923);
nor U2097 (N_2097,N_1972,N_1975);
or U2098 (N_2098,N_1923,N_1929);
and U2099 (N_2099,N_1905,N_1974);
xnor U2100 (N_2100,N_2077,N_2089);
and U2101 (N_2101,N_2030,N_2063);
nor U2102 (N_2102,N_2084,N_2068);
nand U2103 (N_2103,N_2016,N_2074);
nand U2104 (N_2104,N_2007,N_2019);
or U2105 (N_2105,N_2027,N_2057);
and U2106 (N_2106,N_2051,N_2040);
nor U2107 (N_2107,N_2060,N_2043);
xnor U2108 (N_2108,N_2013,N_2058);
and U2109 (N_2109,N_2092,N_2093);
nor U2110 (N_2110,N_2090,N_2082);
or U2111 (N_2111,N_2050,N_2034);
nand U2112 (N_2112,N_2046,N_2009);
nand U2113 (N_2113,N_2044,N_2080);
and U2114 (N_2114,N_2099,N_2075);
and U2115 (N_2115,N_2083,N_2096);
nand U2116 (N_2116,N_2098,N_2036);
nor U2117 (N_2117,N_2011,N_2038);
nand U2118 (N_2118,N_2047,N_2079);
nor U2119 (N_2119,N_2070,N_2069);
or U2120 (N_2120,N_2031,N_2012);
or U2121 (N_2121,N_2067,N_2032);
nor U2122 (N_2122,N_2025,N_2010);
nor U2123 (N_2123,N_2037,N_2086);
and U2124 (N_2124,N_2055,N_2020);
and U2125 (N_2125,N_2087,N_2042);
nor U2126 (N_2126,N_2035,N_2029);
nor U2127 (N_2127,N_2064,N_2000);
nand U2128 (N_2128,N_2053,N_2081);
and U2129 (N_2129,N_2097,N_2018);
nand U2130 (N_2130,N_2061,N_2073);
and U2131 (N_2131,N_2006,N_2076);
nor U2132 (N_2132,N_2021,N_2008);
nor U2133 (N_2133,N_2033,N_2001);
and U2134 (N_2134,N_2014,N_2065);
nor U2135 (N_2135,N_2023,N_2049);
nand U2136 (N_2136,N_2024,N_2004);
or U2137 (N_2137,N_2041,N_2066);
or U2138 (N_2138,N_2002,N_2078);
nor U2139 (N_2139,N_2003,N_2072);
nand U2140 (N_2140,N_2039,N_2015);
nor U2141 (N_2141,N_2022,N_2071);
nor U2142 (N_2142,N_2062,N_2095);
nor U2143 (N_2143,N_2005,N_2045);
nor U2144 (N_2144,N_2052,N_2088);
or U2145 (N_2145,N_2017,N_2056);
nor U2146 (N_2146,N_2059,N_2048);
and U2147 (N_2147,N_2026,N_2054);
nand U2148 (N_2148,N_2091,N_2094);
nor U2149 (N_2149,N_2028,N_2085);
or U2150 (N_2150,N_2095,N_2002);
or U2151 (N_2151,N_2088,N_2029);
or U2152 (N_2152,N_2006,N_2074);
nor U2153 (N_2153,N_2034,N_2066);
nand U2154 (N_2154,N_2060,N_2012);
nand U2155 (N_2155,N_2035,N_2089);
xor U2156 (N_2156,N_2083,N_2080);
or U2157 (N_2157,N_2008,N_2031);
nand U2158 (N_2158,N_2016,N_2028);
or U2159 (N_2159,N_2071,N_2053);
and U2160 (N_2160,N_2042,N_2001);
and U2161 (N_2161,N_2055,N_2066);
nand U2162 (N_2162,N_2009,N_2021);
or U2163 (N_2163,N_2086,N_2060);
and U2164 (N_2164,N_2058,N_2005);
nand U2165 (N_2165,N_2099,N_2022);
nand U2166 (N_2166,N_2083,N_2090);
nand U2167 (N_2167,N_2095,N_2067);
nand U2168 (N_2168,N_2049,N_2038);
nor U2169 (N_2169,N_2078,N_2076);
or U2170 (N_2170,N_2060,N_2089);
nand U2171 (N_2171,N_2069,N_2092);
or U2172 (N_2172,N_2099,N_2042);
and U2173 (N_2173,N_2034,N_2025);
and U2174 (N_2174,N_2038,N_2073);
and U2175 (N_2175,N_2063,N_2057);
or U2176 (N_2176,N_2030,N_2077);
or U2177 (N_2177,N_2077,N_2024);
or U2178 (N_2178,N_2082,N_2040);
or U2179 (N_2179,N_2058,N_2033);
nor U2180 (N_2180,N_2043,N_2002);
nor U2181 (N_2181,N_2045,N_2017);
nor U2182 (N_2182,N_2091,N_2016);
nand U2183 (N_2183,N_2017,N_2039);
and U2184 (N_2184,N_2006,N_2032);
and U2185 (N_2185,N_2079,N_2053);
nand U2186 (N_2186,N_2059,N_2061);
and U2187 (N_2187,N_2041,N_2040);
or U2188 (N_2188,N_2050,N_2024);
nor U2189 (N_2189,N_2035,N_2052);
or U2190 (N_2190,N_2066,N_2026);
and U2191 (N_2191,N_2092,N_2008);
or U2192 (N_2192,N_2030,N_2082);
nand U2193 (N_2193,N_2031,N_2072);
and U2194 (N_2194,N_2057,N_2049);
nor U2195 (N_2195,N_2070,N_2090);
or U2196 (N_2196,N_2066,N_2005);
or U2197 (N_2197,N_2051,N_2035);
nand U2198 (N_2198,N_2074,N_2061);
and U2199 (N_2199,N_2093,N_2052);
nor U2200 (N_2200,N_2164,N_2187);
and U2201 (N_2201,N_2125,N_2158);
nor U2202 (N_2202,N_2132,N_2162);
or U2203 (N_2203,N_2102,N_2111);
nor U2204 (N_2204,N_2106,N_2100);
and U2205 (N_2205,N_2155,N_2101);
and U2206 (N_2206,N_2139,N_2113);
or U2207 (N_2207,N_2146,N_2154);
and U2208 (N_2208,N_2138,N_2185);
or U2209 (N_2209,N_2152,N_2120);
or U2210 (N_2210,N_2104,N_2151);
nand U2211 (N_2211,N_2148,N_2191);
and U2212 (N_2212,N_2161,N_2149);
nand U2213 (N_2213,N_2181,N_2112);
nor U2214 (N_2214,N_2173,N_2179);
or U2215 (N_2215,N_2168,N_2189);
nand U2216 (N_2216,N_2192,N_2186);
or U2217 (N_2217,N_2166,N_2128);
nor U2218 (N_2218,N_2188,N_2180);
and U2219 (N_2219,N_2143,N_2170);
and U2220 (N_2220,N_2114,N_2177);
or U2221 (N_2221,N_2135,N_2178);
nor U2222 (N_2222,N_2197,N_2107);
nor U2223 (N_2223,N_2142,N_2110);
nand U2224 (N_2224,N_2122,N_2190);
nor U2225 (N_2225,N_2163,N_2171);
and U2226 (N_2226,N_2116,N_2150);
and U2227 (N_2227,N_2199,N_2137);
nand U2228 (N_2228,N_2167,N_2176);
and U2229 (N_2229,N_2123,N_2108);
or U2230 (N_2230,N_2153,N_2145);
nand U2231 (N_2231,N_2121,N_2156);
nor U2232 (N_2232,N_2127,N_2196);
nand U2233 (N_2233,N_2133,N_2117);
and U2234 (N_2234,N_2140,N_2147);
or U2235 (N_2235,N_2105,N_2160);
nor U2236 (N_2236,N_2198,N_2159);
or U2237 (N_2237,N_2129,N_2109);
or U2238 (N_2238,N_2157,N_2172);
and U2239 (N_2239,N_2183,N_2144);
and U2240 (N_2240,N_2141,N_2130);
nor U2241 (N_2241,N_2118,N_2103);
and U2242 (N_2242,N_2184,N_2131);
nor U2243 (N_2243,N_2134,N_2194);
nor U2244 (N_2244,N_2124,N_2126);
and U2245 (N_2245,N_2193,N_2119);
or U2246 (N_2246,N_2136,N_2165);
or U2247 (N_2247,N_2169,N_2182);
nor U2248 (N_2248,N_2195,N_2115);
or U2249 (N_2249,N_2174,N_2175);
nand U2250 (N_2250,N_2138,N_2157);
or U2251 (N_2251,N_2168,N_2109);
nand U2252 (N_2252,N_2109,N_2160);
and U2253 (N_2253,N_2173,N_2144);
and U2254 (N_2254,N_2143,N_2113);
nand U2255 (N_2255,N_2120,N_2182);
or U2256 (N_2256,N_2193,N_2142);
or U2257 (N_2257,N_2163,N_2136);
nand U2258 (N_2258,N_2158,N_2130);
and U2259 (N_2259,N_2191,N_2151);
or U2260 (N_2260,N_2138,N_2128);
xor U2261 (N_2261,N_2135,N_2189);
nand U2262 (N_2262,N_2133,N_2142);
and U2263 (N_2263,N_2100,N_2159);
xor U2264 (N_2264,N_2138,N_2170);
and U2265 (N_2265,N_2102,N_2157);
nand U2266 (N_2266,N_2144,N_2135);
or U2267 (N_2267,N_2127,N_2188);
and U2268 (N_2268,N_2156,N_2152);
and U2269 (N_2269,N_2157,N_2128);
nand U2270 (N_2270,N_2122,N_2124);
nor U2271 (N_2271,N_2151,N_2117);
and U2272 (N_2272,N_2183,N_2151);
or U2273 (N_2273,N_2198,N_2158);
nand U2274 (N_2274,N_2182,N_2115);
nand U2275 (N_2275,N_2154,N_2195);
or U2276 (N_2276,N_2168,N_2120);
and U2277 (N_2277,N_2196,N_2106);
nor U2278 (N_2278,N_2124,N_2181);
nand U2279 (N_2279,N_2189,N_2165);
nor U2280 (N_2280,N_2109,N_2145);
or U2281 (N_2281,N_2112,N_2174);
nand U2282 (N_2282,N_2199,N_2143);
nand U2283 (N_2283,N_2177,N_2129);
nand U2284 (N_2284,N_2113,N_2176);
and U2285 (N_2285,N_2141,N_2117);
nand U2286 (N_2286,N_2118,N_2191);
nand U2287 (N_2287,N_2150,N_2172);
and U2288 (N_2288,N_2149,N_2164);
nand U2289 (N_2289,N_2107,N_2192);
or U2290 (N_2290,N_2196,N_2101);
or U2291 (N_2291,N_2136,N_2116);
or U2292 (N_2292,N_2186,N_2161);
nand U2293 (N_2293,N_2162,N_2102);
nand U2294 (N_2294,N_2165,N_2139);
nor U2295 (N_2295,N_2191,N_2112);
or U2296 (N_2296,N_2194,N_2196);
and U2297 (N_2297,N_2187,N_2165);
and U2298 (N_2298,N_2107,N_2176);
or U2299 (N_2299,N_2135,N_2183);
and U2300 (N_2300,N_2298,N_2265);
and U2301 (N_2301,N_2297,N_2278);
nand U2302 (N_2302,N_2225,N_2202);
nand U2303 (N_2303,N_2215,N_2299);
nand U2304 (N_2304,N_2214,N_2235);
or U2305 (N_2305,N_2261,N_2210);
and U2306 (N_2306,N_2291,N_2288);
or U2307 (N_2307,N_2227,N_2285);
nand U2308 (N_2308,N_2224,N_2242);
xnor U2309 (N_2309,N_2211,N_2233);
or U2310 (N_2310,N_2248,N_2240);
nand U2311 (N_2311,N_2289,N_2203);
nand U2312 (N_2312,N_2251,N_2260);
nand U2313 (N_2313,N_2284,N_2287);
nor U2314 (N_2314,N_2219,N_2252);
nand U2315 (N_2315,N_2246,N_2216);
or U2316 (N_2316,N_2237,N_2217);
or U2317 (N_2317,N_2279,N_2241);
and U2318 (N_2318,N_2212,N_2286);
nand U2319 (N_2319,N_2218,N_2295);
xor U2320 (N_2320,N_2209,N_2253);
nand U2321 (N_2321,N_2282,N_2213);
nand U2322 (N_2322,N_2266,N_2271);
nand U2323 (N_2323,N_2239,N_2231);
and U2324 (N_2324,N_2275,N_2268);
nor U2325 (N_2325,N_2277,N_2222);
and U2326 (N_2326,N_2236,N_2206);
or U2327 (N_2327,N_2230,N_2244);
nand U2328 (N_2328,N_2272,N_2280);
and U2329 (N_2329,N_2256,N_2259);
and U2330 (N_2330,N_2255,N_2267);
or U2331 (N_2331,N_2207,N_2293);
nor U2332 (N_2332,N_2249,N_2296);
nand U2333 (N_2333,N_2247,N_2245);
and U2334 (N_2334,N_2264,N_2229);
nand U2335 (N_2335,N_2232,N_2208);
and U2336 (N_2336,N_2276,N_2223);
nand U2337 (N_2337,N_2201,N_2228);
nand U2338 (N_2338,N_2294,N_2220);
xnor U2339 (N_2339,N_2281,N_2258);
and U2340 (N_2340,N_2234,N_2250);
nor U2341 (N_2341,N_2200,N_2254);
nor U2342 (N_2342,N_2226,N_2263);
or U2343 (N_2343,N_2262,N_2273);
and U2344 (N_2344,N_2269,N_2221);
or U2345 (N_2345,N_2274,N_2243);
nand U2346 (N_2346,N_2270,N_2292);
nand U2347 (N_2347,N_2257,N_2290);
nor U2348 (N_2348,N_2283,N_2238);
and U2349 (N_2349,N_2204,N_2205);
xnor U2350 (N_2350,N_2246,N_2247);
nand U2351 (N_2351,N_2226,N_2234);
nand U2352 (N_2352,N_2269,N_2212);
and U2353 (N_2353,N_2253,N_2252);
nand U2354 (N_2354,N_2298,N_2280);
nand U2355 (N_2355,N_2232,N_2217);
nand U2356 (N_2356,N_2225,N_2252);
nand U2357 (N_2357,N_2273,N_2222);
and U2358 (N_2358,N_2277,N_2237);
nand U2359 (N_2359,N_2235,N_2221);
nor U2360 (N_2360,N_2251,N_2266);
nand U2361 (N_2361,N_2206,N_2278);
xor U2362 (N_2362,N_2286,N_2207);
nor U2363 (N_2363,N_2213,N_2223);
nor U2364 (N_2364,N_2228,N_2224);
nand U2365 (N_2365,N_2278,N_2289);
or U2366 (N_2366,N_2231,N_2275);
or U2367 (N_2367,N_2296,N_2212);
or U2368 (N_2368,N_2247,N_2215);
nand U2369 (N_2369,N_2299,N_2297);
nor U2370 (N_2370,N_2260,N_2277);
or U2371 (N_2371,N_2287,N_2204);
nand U2372 (N_2372,N_2227,N_2238);
nand U2373 (N_2373,N_2277,N_2265);
or U2374 (N_2374,N_2259,N_2289);
or U2375 (N_2375,N_2258,N_2285);
nor U2376 (N_2376,N_2211,N_2258);
nor U2377 (N_2377,N_2299,N_2210);
or U2378 (N_2378,N_2290,N_2227);
nor U2379 (N_2379,N_2211,N_2246);
or U2380 (N_2380,N_2258,N_2234);
nand U2381 (N_2381,N_2251,N_2232);
and U2382 (N_2382,N_2238,N_2212);
and U2383 (N_2383,N_2213,N_2248);
xor U2384 (N_2384,N_2216,N_2245);
or U2385 (N_2385,N_2246,N_2228);
nand U2386 (N_2386,N_2207,N_2223);
nor U2387 (N_2387,N_2263,N_2250);
xnor U2388 (N_2388,N_2290,N_2295);
and U2389 (N_2389,N_2206,N_2299);
nand U2390 (N_2390,N_2212,N_2294);
nor U2391 (N_2391,N_2203,N_2200);
nor U2392 (N_2392,N_2285,N_2231);
nand U2393 (N_2393,N_2228,N_2210);
or U2394 (N_2394,N_2209,N_2206);
or U2395 (N_2395,N_2247,N_2290);
nor U2396 (N_2396,N_2207,N_2203);
nand U2397 (N_2397,N_2297,N_2204);
nand U2398 (N_2398,N_2205,N_2295);
and U2399 (N_2399,N_2239,N_2206);
nor U2400 (N_2400,N_2345,N_2343);
or U2401 (N_2401,N_2354,N_2367);
nor U2402 (N_2402,N_2319,N_2337);
xor U2403 (N_2403,N_2379,N_2305);
nor U2404 (N_2404,N_2308,N_2380);
and U2405 (N_2405,N_2330,N_2383);
nor U2406 (N_2406,N_2346,N_2387);
nor U2407 (N_2407,N_2369,N_2398);
nor U2408 (N_2408,N_2378,N_2338);
nor U2409 (N_2409,N_2312,N_2364);
and U2410 (N_2410,N_2348,N_2322);
or U2411 (N_2411,N_2324,N_2344);
and U2412 (N_2412,N_2363,N_2356);
nor U2413 (N_2413,N_2392,N_2329);
nor U2414 (N_2414,N_2373,N_2384);
nand U2415 (N_2415,N_2311,N_2323);
nor U2416 (N_2416,N_2339,N_2303);
or U2417 (N_2417,N_2351,N_2389);
nor U2418 (N_2418,N_2349,N_2310);
and U2419 (N_2419,N_2353,N_2393);
nand U2420 (N_2420,N_2300,N_2366);
nand U2421 (N_2421,N_2315,N_2385);
and U2422 (N_2422,N_2302,N_2314);
nor U2423 (N_2423,N_2371,N_2395);
and U2424 (N_2424,N_2331,N_2301);
nor U2425 (N_2425,N_2336,N_2399);
xor U2426 (N_2426,N_2382,N_2307);
nand U2427 (N_2427,N_2352,N_2334);
and U2428 (N_2428,N_2332,N_2316);
xor U2429 (N_2429,N_2340,N_2318);
nand U2430 (N_2430,N_2362,N_2342);
or U2431 (N_2431,N_2321,N_2306);
nor U2432 (N_2432,N_2397,N_2309);
nor U2433 (N_2433,N_2320,N_2313);
nand U2434 (N_2434,N_2374,N_2396);
xor U2435 (N_2435,N_2368,N_2341);
or U2436 (N_2436,N_2377,N_2370);
or U2437 (N_2437,N_2365,N_2391);
nand U2438 (N_2438,N_2359,N_2347);
nand U2439 (N_2439,N_2325,N_2386);
and U2440 (N_2440,N_2328,N_2317);
and U2441 (N_2441,N_2355,N_2372);
or U2442 (N_2442,N_2335,N_2388);
nand U2443 (N_2443,N_2390,N_2357);
nor U2444 (N_2444,N_2350,N_2360);
nand U2445 (N_2445,N_2375,N_2304);
and U2446 (N_2446,N_2358,N_2327);
or U2447 (N_2447,N_2361,N_2326);
and U2448 (N_2448,N_2376,N_2394);
nand U2449 (N_2449,N_2333,N_2381);
xor U2450 (N_2450,N_2350,N_2372);
nor U2451 (N_2451,N_2375,N_2320);
or U2452 (N_2452,N_2397,N_2303);
and U2453 (N_2453,N_2378,N_2312);
nand U2454 (N_2454,N_2391,N_2359);
or U2455 (N_2455,N_2389,N_2384);
and U2456 (N_2456,N_2357,N_2314);
or U2457 (N_2457,N_2385,N_2312);
or U2458 (N_2458,N_2307,N_2384);
nand U2459 (N_2459,N_2374,N_2369);
nand U2460 (N_2460,N_2341,N_2336);
nor U2461 (N_2461,N_2390,N_2348);
and U2462 (N_2462,N_2392,N_2373);
or U2463 (N_2463,N_2306,N_2389);
and U2464 (N_2464,N_2306,N_2385);
and U2465 (N_2465,N_2397,N_2350);
or U2466 (N_2466,N_2396,N_2373);
nand U2467 (N_2467,N_2399,N_2350);
nand U2468 (N_2468,N_2308,N_2307);
nand U2469 (N_2469,N_2355,N_2323);
nand U2470 (N_2470,N_2379,N_2301);
and U2471 (N_2471,N_2396,N_2348);
and U2472 (N_2472,N_2342,N_2311);
nor U2473 (N_2473,N_2315,N_2366);
nand U2474 (N_2474,N_2380,N_2327);
or U2475 (N_2475,N_2384,N_2347);
nor U2476 (N_2476,N_2357,N_2327);
nand U2477 (N_2477,N_2342,N_2379);
nand U2478 (N_2478,N_2397,N_2355);
or U2479 (N_2479,N_2375,N_2321);
nand U2480 (N_2480,N_2374,N_2388);
and U2481 (N_2481,N_2365,N_2359);
nor U2482 (N_2482,N_2351,N_2396);
nand U2483 (N_2483,N_2373,N_2335);
and U2484 (N_2484,N_2341,N_2360);
nand U2485 (N_2485,N_2315,N_2358);
nand U2486 (N_2486,N_2341,N_2397);
nand U2487 (N_2487,N_2382,N_2313);
and U2488 (N_2488,N_2377,N_2319);
or U2489 (N_2489,N_2391,N_2309);
nor U2490 (N_2490,N_2371,N_2304);
nor U2491 (N_2491,N_2358,N_2318);
nand U2492 (N_2492,N_2385,N_2326);
xnor U2493 (N_2493,N_2333,N_2326);
and U2494 (N_2494,N_2347,N_2340);
or U2495 (N_2495,N_2330,N_2313);
nor U2496 (N_2496,N_2365,N_2358);
nand U2497 (N_2497,N_2389,N_2381);
and U2498 (N_2498,N_2368,N_2352);
nor U2499 (N_2499,N_2327,N_2313);
nor U2500 (N_2500,N_2456,N_2452);
nor U2501 (N_2501,N_2445,N_2480);
nand U2502 (N_2502,N_2408,N_2442);
nand U2503 (N_2503,N_2431,N_2404);
xor U2504 (N_2504,N_2468,N_2423);
nor U2505 (N_2505,N_2449,N_2414);
or U2506 (N_2506,N_2441,N_2479);
nand U2507 (N_2507,N_2484,N_2426);
and U2508 (N_2508,N_2466,N_2432);
or U2509 (N_2509,N_2467,N_2438);
nor U2510 (N_2510,N_2487,N_2443);
or U2511 (N_2511,N_2413,N_2410);
nand U2512 (N_2512,N_2478,N_2406);
nor U2513 (N_2513,N_2488,N_2473);
or U2514 (N_2514,N_2494,N_2498);
and U2515 (N_2515,N_2440,N_2495);
nand U2516 (N_2516,N_2481,N_2428);
and U2517 (N_2517,N_2475,N_2430);
or U2518 (N_2518,N_2477,N_2412);
nand U2519 (N_2519,N_2482,N_2435);
and U2520 (N_2520,N_2489,N_2454);
or U2521 (N_2521,N_2419,N_2459);
nor U2522 (N_2522,N_2493,N_2463);
and U2523 (N_2523,N_2417,N_2465);
nand U2524 (N_2524,N_2451,N_2499);
or U2525 (N_2525,N_2434,N_2415);
or U2526 (N_2526,N_2433,N_2421);
nor U2527 (N_2527,N_2469,N_2458);
nand U2528 (N_2528,N_2422,N_2483);
nand U2529 (N_2529,N_2471,N_2446);
nand U2530 (N_2530,N_2491,N_2472);
or U2531 (N_2531,N_2457,N_2485);
and U2532 (N_2532,N_2407,N_2409);
nor U2533 (N_2533,N_2492,N_2453);
nand U2534 (N_2534,N_2420,N_2418);
xnor U2535 (N_2535,N_2402,N_2450);
nor U2536 (N_2536,N_2448,N_2425);
and U2537 (N_2537,N_2405,N_2464);
nand U2538 (N_2538,N_2447,N_2429);
nand U2539 (N_2539,N_2416,N_2460);
or U2540 (N_2540,N_2436,N_2462);
nand U2541 (N_2541,N_2411,N_2427);
or U2542 (N_2542,N_2461,N_2497);
or U2543 (N_2543,N_2400,N_2401);
nor U2544 (N_2544,N_2486,N_2474);
nor U2545 (N_2545,N_2470,N_2444);
or U2546 (N_2546,N_2424,N_2455);
nand U2547 (N_2547,N_2476,N_2403);
nand U2548 (N_2548,N_2496,N_2439);
or U2549 (N_2549,N_2437,N_2490);
or U2550 (N_2550,N_2454,N_2453);
and U2551 (N_2551,N_2406,N_2480);
nor U2552 (N_2552,N_2487,N_2451);
nand U2553 (N_2553,N_2401,N_2447);
nor U2554 (N_2554,N_2407,N_2405);
and U2555 (N_2555,N_2423,N_2403);
xnor U2556 (N_2556,N_2409,N_2424);
or U2557 (N_2557,N_2422,N_2494);
and U2558 (N_2558,N_2462,N_2490);
and U2559 (N_2559,N_2425,N_2468);
and U2560 (N_2560,N_2473,N_2420);
or U2561 (N_2561,N_2444,N_2436);
and U2562 (N_2562,N_2496,N_2457);
nor U2563 (N_2563,N_2492,N_2405);
or U2564 (N_2564,N_2464,N_2440);
and U2565 (N_2565,N_2444,N_2478);
or U2566 (N_2566,N_2453,N_2418);
or U2567 (N_2567,N_2474,N_2487);
nand U2568 (N_2568,N_2474,N_2430);
or U2569 (N_2569,N_2402,N_2428);
and U2570 (N_2570,N_2463,N_2424);
or U2571 (N_2571,N_2496,N_2485);
nand U2572 (N_2572,N_2476,N_2423);
nand U2573 (N_2573,N_2459,N_2432);
or U2574 (N_2574,N_2404,N_2401);
or U2575 (N_2575,N_2440,N_2489);
and U2576 (N_2576,N_2482,N_2472);
or U2577 (N_2577,N_2430,N_2419);
or U2578 (N_2578,N_2492,N_2433);
or U2579 (N_2579,N_2435,N_2416);
nand U2580 (N_2580,N_2445,N_2429);
and U2581 (N_2581,N_2495,N_2468);
and U2582 (N_2582,N_2476,N_2440);
or U2583 (N_2583,N_2427,N_2498);
xnor U2584 (N_2584,N_2455,N_2496);
nand U2585 (N_2585,N_2492,N_2484);
or U2586 (N_2586,N_2464,N_2400);
and U2587 (N_2587,N_2467,N_2426);
nand U2588 (N_2588,N_2432,N_2460);
xor U2589 (N_2589,N_2455,N_2489);
or U2590 (N_2590,N_2436,N_2479);
and U2591 (N_2591,N_2479,N_2498);
nor U2592 (N_2592,N_2439,N_2433);
nor U2593 (N_2593,N_2456,N_2446);
nor U2594 (N_2594,N_2499,N_2444);
nor U2595 (N_2595,N_2447,N_2457);
nand U2596 (N_2596,N_2450,N_2404);
and U2597 (N_2597,N_2445,N_2441);
or U2598 (N_2598,N_2484,N_2443);
or U2599 (N_2599,N_2488,N_2412);
nand U2600 (N_2600,N_2522,N_2547);
nand U2601 (N_2601,N_2576,N_2539);
and U2602 (N_2602,N_2511,N_2530);
nor U2603 (N_2603,N_2537,N_2598);
nor U2604 (N_2604,N_2579,N_2552);
nor U2605 (N_2605,N_2523,N_2536);
nor U2606 (N_2606,N_2514,N_2500);
or U2607 (N_2607,N_2548,N_2585);
nor U2608 (N_2608,N_2554,N_2589);
nor U2609 (N_2609,N_2542,N_2533);
nor U2610 (N_2610,N_2508,N_2582);
nand U2611 (N_2611,N_2509,N_2557);
nand U2612 (N_2612,N_2592,N_2587);
nor U2613 (N_2613,N_2549,N_2574);
nor U2614 (N_2614,N_2546,N_2563);
nand U2615 (N_2615,N_2507,N_2553);
or U2616 (N_2616,N_2515,N_2512);
or U2617 (N_2617,N_2575,N_2513);
nand U2618 (N_2618,N_2588,N_2538);
nand U2619 (N_2619,N_2551,N_2518);
and U2620 (N_2620,N_2525,N_2529);
and U2621 (N_2621,N_2544,N_2555);
and U2622 (N_2622,N_2519,N_2581);
nor U2623 (N_2623,N_2567,N_2502);
nor U2624 (N_2624,N_2535,N_2594);
nor U2625 (N_2625,N_2590,N_2532);
and U2626 (N_2626,N_2597,N_2503);
or U2627 (N_2627,N_2564,N_2568);
nor U2628 (N_2628,N_2531,N_2534);
and U2629 (N_2629,N_2571,N_2566);
or U2630 (N_2630,N_2545,N_2516);
nand U2631 (N_2631,N_2550,N_2505);
nand U2632 (N_2632,N_2565,N_2593);
nand U2633 (N_2633,N_2524,N_2543);
nand U2634 (N_2634,N_2586,N_2583);
nor U2635 (N_2635,N_2596,N_2595);
nand U2636 (N_2636,N_2541,N_2572);
nor U2637 (N_2637,N_2570,N_2584);
nand U2638 (N_2638,N_2558,N_2504);
and U2639 (N_2639,N_2501,N_2526);
nand U2640 (N_2640,N_2562,N_2510);
or U2641 (N_2641,N_2560,N_2517);
nor U2642 (N_2642,N_2591,N_2528);
or U2643 (N_2643,N_2573,N_2540);
nand U2644 (N_2644,N_2578,N_2556);
or U2645 (N_2645,N_2520,N_2521);
nand U2646 (N_2646,N_2561,N_2577);
nor U2647 (N_2647,N_2527,N_2506);
and U2648 (N_2648,N_2599,N_2559);
or U2649 (N_2649,N_2580,N_2569);
nor U2650 (N_2650,N_2523,N_2513);
and U2651 (N_2651,N_2526,N_2502);
or U2652 (N_2652,N_2559,N_2514);
nand U2653 (N_2653,N_2532,N_2578);
and U2654 (N_2654,N_2558,N_2516);
nand U2655 (N_2655,N_2566,N_2551);
and U2656 (N_2656,N_2533,N_2528);
and U2657 (N_2657,N_2541,N_2569);
nor U2658 (N_2658,N_2581,N_2518);
nor U2659 (N_2659,N_2513,N_2566);
or U2660 (N_2660,N_2575,N_2521);
or U2661 (N_2661,N_2510,N_2555);
and U2662 (N_2662,N_2566,N_2534);
and U2663 (N_2663,N_2592,N_2589);
nand U2664 (N_2664,N_2528,N_2588);
nor U2665 (N_2665,N_2598,N_2568);
and U2666 (N_2666,N_2550,N_2573);
or U2667 (N_2667,N_2507,N_2592);
nand U2668 (N_2668,N_2557,N_2553);
nor U2669 (N_2669,N_2528,N_2553);
nor U2670 (N_2670,N_2518,N_2528);
nand U2671 (N_2671,N_2525,N_2598);
nor U2672 (N_2672,N_2580,N_2532);
nor U2673 (N_2673,N_2547,N_2500);
and U2674 (N_2674,N_2520,N_2553);
nor U2675 (N_2675,N_2502,N_2573);
and U2676 (N_2676,N_2592,N_2530);
nor U2677 (N_2677,N_2541,N_2594);
or U2678 (N_2678,N_2599,N_2555);
nand U2679 (N_2679,N_2521,N_2569);
nor U2680 (N_2680,N_2522,N_2550);
nand U2681 (N_2681,N_2593,N_2544);
and U2682 (N_2682,N_2552,N_2567);
and U2683 (N_2683,N_2563,N_2593);
nor U2684 (N_2684,N_2556,N_2566);
or U2685 (N_2685,N_2500,N_2526);
and U2686 (N_2686,N_2563,N_2542);
nand U2687 (N_2687,N_2585,N_2509);
or U2688 (N_2688,N_2543,N_2547);
nand U2689 (N_2689,N_2586,N_2556);
and U2690 (N_2690,N_2546,N_2594);
and U2691 (N_2691,N_2597,N_2513);
and U2692 (N_2692,N_2578,N_2591);
or U2693 (N_2693,N_2505,N_2513);
or U2694 (N_2694,N_2590,N_2534);
nor U2695 (N_2695,N_2582,N_2572);
nor U2696 (N_2696,N_2501,N_2565);
and U2697 (N_2697,N_2518,N_2579);
nor U2698 (N_2698,N_2551,N_2516);
nand U2699 (N_2699,N_2532,N_2531);
and U2700 (N_2700,N_2634,N_2616);
nor U2701 (N_2701,N_2649,N_2614);
nand U2702 (N_2702,N_2625,N_2656);
and U2703 (N_2703,N_2695,N_2653);
and U2704 (N_2704,N_2631,N_2619);
nor U2705 (N_2705,N_2691,N_2650);
and U2706 (N_2706,N_2682,N_2605);
nand U2707 (N_2707,N_2699,N_2617);
or U2708 (N_2708,N_2697,N_2673);
nor U2709 (N_2709,N_2669,N_2678);
or U2710 (N_2710,N_2688,N_2621);
or U2711 (N_2711,N_2643,N_2610);
nand U2712 (N_2712,N_2659,N_2684);
nand U2713 (N_2713,N_2612,N_2615);
nor U2714 (N_2714,N_2651,N_2632);
xnor U2715 (N_2715,N_2655,N_2694);
and U2716 (N_2716,N_2604,N_2609);
xor U2717 (N_2717,N_2628,N_2667);
or U2718 (N_2718,N_2674,N_2601);
nor U2719 (N_2719,N_2663,N_2644);
nand U2720 (N_2720,N_2629,N_2677);
or U2721 (N_2721,N_2608,N_2661);
and U2722 (N_2722,N_2624,N_2645);
nor U2723 (N_2723,N_2635,N_2672);
and U2724 (N_2724,N_2662,N_2637);
or U2725 (N_2725,N_2696,N_2692);
nor U2726 (N_2726,N_2689,N_2620);
or U2727 (N_2727,N_2654,N_2642);
or U2728 (N_2728,N_2646,N_2686);
and U2729 (N_2729,N_2641,N_2687);
or U2730 (N_2730,N_2600,N_2664);
or U2731 (N_2731,N_2613,N_2665);
nand U2732 (N_2732,N_2630,N_2648);
or U2733 (N_2733,N_2640,N_2622);
nand U2734 (N_2734,N_2607,N_2679);
and U2735 (N_2735,N_2670,N_2618);
or U2736 (N_2736,N_2685,N_2668);
or U2737 (N_2737,N_2636,N_2603);
and U2738 (N_2738,N_2633,N_2657);
nor U2739 (N_2739,N_2681,N_2683);
xnor U2740 (N_2740,N_2638,N_2652);
or U2741 (N_2741,N_2626,N_2602);
or U2742 (N_2742,N_2647,N_2623);
and U2743 (N_2743,N_2671,N_2611);
or U2744 (N_2744,N_2606,N_2639);
nand U2745 (N_2745,N_2627,N_2675);
or U2746 (N_2746,N_2676,N_2658);
xnor U2747 (N_2747,N_2666,N_2680);
nand U2748 (N_2748,N_2693,N_2698);
and U2749 (N_2749,N_2660,N_2690);
nor U2750 (N_2750,N_2675,N_2647);
and U2751 (N_2751,N_2637,N_2622);
nor U2752 (N_2752,N_2676,N_2648);
and U2753 (N_2753,N_2630,N_2624);
or U2754 (N_2754,N_2618,N_2679);
nor U2755 (N_2755,N_2620,N_2698);
nor U2756 (N_2756,N_2613,N_2694);
and U2757 (N_2757,N_2636,N_2654);
nor U2758 (N_2758,N_2669,N_2695);
nor U2759 (N_2759,N_2647,N_2671);
and U2760 (N_2760,N_2602,N_2648);
or U2761 (N_2761,N_2683,N_2673);
nor U2762 (N_2762,N_2607,N_2660);
nand U2763 (N_2763,N_2691,N_2676);
xor U2764 (N_2764,N_2641,N_2683);
nand U2765 (N_2765,N_2649,N_2628);
nand U2766 (N_2766,N_2697,N_2605);
nand U2767 (N_2767,N_2610,N_2654);
or U2768 (N_2768,N_2658,N_2606);
or U2769 (N_2769,N_2697,N_2643);
nor U2770 (N_2770,N_2627,N_2612);
or U2771 (N_2771,N_2616,N_2636);
and U2772 (N_2772,N_2666,N_2658);
nor U2773 (N_2773,N_2682,N_2696);
and U2774 (N_2774,N_2663,N_2615);
nand U2775 (N_2775,N_2650,N_2601);
and U2776 (N_2776,N_2655,N_2682);
nor U2777 (N_2777,N_2675,N_2625);
and U2778 (N_2778,N_2645,N_2600);
or U2779 (N_2779,N_2620,N_2640);
or U2780 (N_2780,N_2693,N_2649);
or U2781 (N_2781,N_2653,N_2696);
or U2782 (N_2782,N_2654,N_2699);
or U2783 (N_2783,N_2685,N_2630);
nand U2784 (N_2784,N_2621,N_2613);
xnor U2785 (N_2785,N_2678,N_2696);
nand U2786 (N_2786,N_2664,N_2630);
nand U2787 (N_2787,N_2669,N_2655);
or U2788 (N_2788,N_2696,N_2636);
or U2789 (N_2789,N_2604,N_2636);
nor U2790 (N_2790,N_2606,N_2691);
and U2791 (N_2791,N_2637,N_2617);
xor U2792 (N_2792,N_2652,N_2689);
nor U2793 (N_2793,N_2610,N_2639);
nand U2794 (N_2794,N_2671,N_2667);
or U2795 (N_2795,N_2635,N_2659);
or U2796 (N_2796,N_2600,N_2650);
or U2797 (N_2797,N_2613,N_2670);
or U2798 (N_2798,N_2622,N_2633);
nand U2799 (N_2799,N_2614,N_2624);
or U2800 (N_2800,N_2736,N_2768);
nand U2801 (N_2801,N_2778,N_2750);
or U2802 (N_2802,N_2793,N_2713);
nor U2803 (N_2803,N_2786,N_2798);
and U2804 (N_2804,N_2767,N_2728);
and U2805 (N_2805,N_2724,N_2764);
and U2806 (N_2806,N_2791,N_2729);
xnor U2807 (N_2807,N_2766,N_2796);
xnor U2808 (N_2808,N_2745,N_2732);
and U2809 (N_2809,N_2759,N_2742);
xnor U2810 (N_2810,N_2747,N_2757);
nor U2811 (N_2811,N_2702,N_2721);
nand U2812 (N_2812,N_2752,N_2744);
nand U2813 (N_2813,N_2787,N_2754);
nor U2814 (N_2814,N_2769,N_2700);
or U2815 (N_2815,N_2782,N_2781);
and U2816 (N_2816,N_2771,N_2741);
nand U2817 (N_2817,N_2704,N_2714);
nand U2818 (N_2818,N_2719,N_2709);
or U2819 (N_2819,N_2784,N_2780);
or U2820 (N_2820,N_2773,N_2774);
and U2821 (N_2821,N_2723,N_2733);
and U2822 (N_2822,N_2790,N_2753);
nor U2823 (N_2823,N_2727,N_2716);
or U2824 (N_2824,N_2726,N_2722);
and U2825 (N_2825,N_2749,N_2755);
nand U2826 (N_2826,N_2708,N_2776);
nor U2827 (N_2827,N_2739,N_2788);
or U2828 (N_2828,N_2779,N_2707);
and U2829 (N_2829,N_2763,N_2775);
and U2830 (N_2830,N_2795,N_2751);
or U2831 (N_2831,N_2758,N_2734);
or U2832 (N_2832,N_2765,N_2799);
nor U2833 (N_2833,N_2760,N_2738);
nor U2834 (N_2834,N_2705,N_2746);
nand U2835 (N_2835,N_2743,N_2740);
and U2836 (N_2836,N_2785,N_2715);
and U2837 (N_2837,N_2783,N_2735);
or U2838 (N_2838,N_2770,N_2731);
and U2839 (N_2839,N_2725,N_2792);
nor U2840 (N_2840,N_2712,N_2701);
and U2841 (N_2841,N_2789,N_2710);
nand U2842 (N_2842,N_2748,N_2794);
or U2843 (N_2843,N_2761,N_2703);
nand U2844 (N_2844,N_2711,N_2756);
nor U2845 (N_2845,N_2718,N_2762);
and U2846 (N_2846,N_2772,N_2717);
or U2847 (N_2847,N_2720,N_2737);
or U2848 (N_2848,N_2706,N_2730);
or U2849 (N_2849,N_2777,N_2797);
nor U2850 (N_2850,N_2762,N_2701);
and U2851 (N_2851,N_2785,N_2796);
nand U2852 (N_2852,N_2751,N_2757);
or U2853 (N_2853,N_2744,N_2750);
nor U2854 (N_2854,N_2722,N_2788);
nand U2855 (N_2855,N_2732,N_2734);
nand U2856 (N_2856,N_2736,N_2719);
nor U2857 (N_2857,N_2701,N_2760);
and U2858 (N_2858,N_2758,N_2715);
or U2859 (N_2859,N_2764,N_2779);
or U2860 (N_2860,N_2706,N_2737);
nand U2861 (N_2861,N_2756,N_2704);
nand U2862 (N_2862,N_2779,N_2741);
nor U2863 (N_2863,N_2773,N_2785);
or U2864 (N_2864,N_2780,N_2726);
nor U2865 (N_2865,N_2742,N_2792);
xnor U2866 (N_2866,N_2783,N_2754);
nor U2867 (N_2867,N_2774,N_2743);
and U2868 (N_2868,N_2794,N_2753);
or U2869 (N_2869,N_2727,N_2778);
nor U2870 (N_2870,N_2727,N_2702);
nand U2871 (N_2871,N_2788,N_2765);
or U2872 (N_2872,N_2765,N_2778);
nand U2873 (N_2873,N_2744,N_2764);
nand U2874 (N_2874,N_2736,N_2785);
or U2875 (N_2875,N_2722,N_2787);
nand U2876 (N_2876,N_2747,N_2754);
nand U2877 (N_2877,N_2778,N_2760);
nand U2878 (N_2878,N_2753,N_2727);
or U2879 (N_2879,N_2793,N_2790);
and U2880 (N_2880,N_2799,N_2758);
or U2881 (N_2881,N_2778,N_2790);
xnor U2882 (N_2882,N_2791,N_2706);
and U2883 (N_2883,N_2774,N_2715);
and U2884 (N_2884,N_2713,N_2751);
and U2885 (N_2885,N_2737,N_2755);
nand U2886 (N_2886,N_2792,N_2782);
and U2887 (N_2887,N_2708,N_2737);
nor U2888 (N_2888,N_2719,N_2734);
nor U2889 (N_2889,N_2701,N_2770);
nand U2890 (N_2890,N_2710,N_2701);
nor U2891 (N_2891,N_2747,N_2715);
nand U2892 (N_2892,N_2761,N_2779);
and U2893 (N_2893,N_2709,N_2750);
nor U2894 (N_2894,N_2753,N_2719);
or U2895 (N_2895,N_2758,N_2726);
nand U2896 (N_2896,N_2768,N_2794);
nand U2897 (N_2897,N_2732,N_2779);
nand U2898 (N_2898,N_2761,N_2749);
or U2899 (N_2899,N_2774,N_2704);
and U2900 (N_2900,N_2840,N_2859);
and U2901 (N_2901,N_2847,N_2814);
or U2902 (N_2902,N_2881,N_2861);
and U2903 (N_2903,N_2819,N_2851);
nor U2904 (N_2904,N_2879,N_2816);
and U2905 (N_2905,N_2873,N_2871);
nor U2906 (N_2906,N_2817,N_2858);
and U2907 (N_2907,N_2857,N_2807);
nor U2908 (N_2908,N_2835,N_2842);
nand U2909 (N_2909,N_2862,N_2888);
nor U2910 (N_2910,N_2867,N_2827);
and U2911 (N_2911,N_2854,N_2866);
or U2912 (N_2912,N_2885,N_2828);
nand U2913 (N_2913,N_2845,N_2824);
nand U2914 (N_2914,N_2826,N_2836);
and U2915 (N_2915,N_2850,N_2822);
and U2916 (N_2916,N_2860,N_2891);
nor U2917 (N_2917,N_2877,N_2812);
nor U2918 (N_2918,N_2874,N_2844);
nor U2919 (N_2919,N_2876,N_2892);
or U2920 (N_2920,N_2880,N_2823);
or U2921 (N_2921,N_2849,N_2800);
nor U2922 (N_2922,N_2897,N_2875);
xnor U2923 (N_2923,N_2820,N_2869);
and U2924 (N_2924,N_2853,N_2834);
nor U2925 (N_2925,N_2868,N_2898);
and U2926 (N_2926,N_2886,N_2831);
nor U2927 (N_2927,N_2833,N_2878);
and U2928 (N_2928,N_2809,N_2803);
nor U2929 (N_2929,N_2806,N_2818);
nor U2930 (N_2930,N_2884,N_2864);
and U2931 (N_2931,N_2843,N_2852);
and U2932 (N_2932,N_2838,N_2804);
nand U2933 (N_2933,N_2813,N_2832);
nor U2934 (N_2934,N_2825,N_2872);
nor U2935 (N_2935,N_2837,N_2821);
xor U2936 (N_2936,N_2887,N_2895);
nor U2937 (N_2937,N_2870,N_2865);
xor U2938 (N_2938,N_2830,N_2894);
nand U2939 (N_2939,N_2839,N_2802);
nor U2940 (N_2940,N_2855,N_2890);
xnor U2941 (N_2941,N_2883,N_2889);
or U2942 (N_2942,N_2829,N_2811);
and U2943 (N_2943,N_2882,N_2801);
nor U2944 (N_2944,N_2863,N_2808);
nand U2945 (N_2945,N_2846,N_2810);
nor U2946 (N_2946,N_2848,N_2815);
or U2947 (N_2947,N_2841,N_2899);
nand U2948 (N_2948,N_2896,N_2893);
and U2949 (N_2949,N_2805,N_2856);
or U2950 (N_2950,N_2887,N_2801);
and U2951 (N_2951,N_2821,N_2819);
nor U2952 (N_2952,N_2807,N_2891);
and U2953 (N_2953,N_2816,N_2823);
nand U2954 (N_2954,N_2858,N_2866);
nand U2955 (N_2955,N_2840,N_2863);
nand U2956 (N_2956,N_2833,N_2832);
and U2957 (N_2957,N_2860,N_2885);
xnor U2958 (N_2958,N_2807,N_2862);
nand U2959 (N_2959,N_2861,N_2848);
nand U2960 (N_2960,N_2865,N_2882);
nand U2961 (N_2961,N_2821,N_2810);
nand U2962 (N_2962,N_2834,N_2835);
nor U2963 (N_2963,N_2852,N_2835);
and U2964 (N_2964,N_2881,N_2887);
nor U2965 (N_2965,N_2829,N_2861);
xor U2966 (N_2966,N_2875,N_2861);
nor U2967 (N_2967,N_2802,N_2896);
nor U2968 (N_2968,N_2821,N_2888);
nand U2969 (N_2969,N_2867,N_2840);
nor U2970 (N_2970,N_2817,N_2889);
and U2971 (N_2971,N_2875,N_2847);
nor U2972 (N_2972,N_2861,N_2838);
nor U2973 (N_2973,N_2838,N_2845);
and U2974 (N_2974,N_2858,N_2894);
nor U2975 (N_2975,N_2832,N_2862);
or U2976 (N_2976,N_2811,N_2819);
nor U2977 (N_2977,N_2840,N_2800);
and U2978 (N_2978,N_2826,N_2854);
nor U2979 (N_2979,N_2801,N_2830);
nand U2980 (N_2980,N_2883,N_2822);
nor U2981 (N_2981,N_2842,N_2863);
nor U2982 (N_2982,N_2883,N_2854);
nor U2983 (N_2983,N_2853,N_2846);
or U2984 (N_2984,N_2831,N_2888);
nor U2985 (N_2985,N_2865,N_2838);
xnor U2986 (N_2986,N_2867,N_2896);
nor U2987 (N_2987,N_2820,N_2892);
and U2988 (N_2988,N_2892,N_2832);
nand U2989 (N_2989,N_2850,N_2801);
nand U2990 (N_2990,N_2849,N_2886);
nor U2991 (N_2991,N_2850,N_2807);
or U2992 (N_2992,N_2824,N_2838);
and U2993 (N_2993,N_2808,N_2811);
and U2994 (N_2994,N_2889,N_2818);
nor U2995 (N_2995,N_2822,N_2832);
and U2996 (N_2996,N_2839,N_2849);
nor U2997 (N_2997,N_2812,N_2857);
xnor U2998 (N_2998,N_2837,N_2880);
and U2999 (N_2999,N_2879,N_2840);
or U3000 (N_3000,N_2923,N_2978);
nor U3001 (N_3001,N_2912,N_2919);
nor U3002 (N_3002,N_2939,N_2930);
or U3003 (N_3003,N_2997,N_2949);
nand U3004 (N_3004,N_2987,N_2943);
or U3005 (N_3005,N_2973,N_2979);
nor U3006 (N_3006,N_2906,N_2913);
or U3007 (N_3007,N_2904,N_2975);
nand U3008 (N_3008,N_2903,N_2989);
and U3009 (N_3009,N_2993,N_2931);
or U3010 (N_3010,N_2991,N_2907);
and U3011 (N_3011,N_2924,N_2940);
or U3012 (N_3012,N_2974,N_2938);
nor U3013 (N_3013,N_2980,N_2925);
and U3014 (N_3014,N_2954,N_2901);
or U3015 (N_3015,N_2936,N_2995);
and U3016 (N_3016,N_2988,N_2928);
or U3017 (N_3017,N_2985,N_2964);
or U3018 (N_3018,N_2962,N_2920);
or U3019 (N_3019,N_2915,N_2937);
and U3020 (N_3020,N_2958,N_2982);
or U3021 (N_3021,N_2959,N_2900);
nor U3022 (N_3022,N_2934,N_2957);
nor U3023 (N_3023,N_2908,N_2999);
and U3024 (N_3024,N_2956,N_2971);
nand U3025 (N_3025,N_2953,N_2967);
nor U3026 (N_3026,N_2914,N_2910);
and U3027 (N_3027,N_2972,N_2921);
nand U3028 (N_3028,N_2909,N_2994);
or U3029 (N_3029,N_2917,N_2998);
nor U3030 (N_3030,N_2952,N_2902);
or U3031 (N_3031,N_2966,N_2922);
nand U3032 (N_3032,N_2947,N_2942);
or U3033 (N_3033,N_2927,N_2929);
nor U3034 (N_3034,N_2926,N_2944);
or U3035 (N_3035,N_2945,N_2983);
nand U3036 (N_3036,N_2911,N_2965);
and U3037 (N_3037,N_2941,N_2970);
xnor U3038 (N_3038,N_2984,N_2932);
or U3039 (N_3039,N_2946,N_2950);
and U3040 (N_3040,N_2996,N_2948);
nand U3041 (N_3041,N_2963,N_2918);
or U3042 (N_3042,N_2977,N_2981);
nor U3043 (N_3043,N_2955,N_2916);
and U3044 (N_3044,N_2986,N_2935);
and U3045 (N_3045,N_2976,N_2968);
or U3046 (N_3046,N_2992,N_2969);
xor U3047 (N_3047,N_2951,N_2960);
or U3048 (N_3048,N_2990,N_2961);
or U3049 (N_3049,N_2933,N_2905);
nor U3050 (N_3050,N_2937,N_2990);
nand U3051 (N_3051,N_2902,N_2995);
nor U3052 (N_3052,N_2985,N_2927);
and U3053 (N_3053,N_2964,N_2963);
and U3054 (N_3054,N_2903,N_2986);
nand U3055 (N_3055,N_2959,N_2927);
nor U3056 (N_3056,N_2936,N_2923);
nand U3057 (N_3057,N_2990,N_2999);
nor U3058 (N_3058,N_2984,N_2928);
nor U3059 (N_3059,N_2972,N_2904);
nor U3060 (N_3060,N_2989,N_2944);
or U3061 (N_3061,N_2934,N_2990);
nor U3062 (N_3062,N_2961,N_2913);
or U3063 (N_3063,N_2912,N_2924);
and U3064 (N_3064,N_2942,N_2902);
nor U3065 (N_3065,N_2932,N_2921);
and U3066 (N_3066,N_2908,N_2996);
nor U3067 (N_3067,N_2985,N_2921);
and U3068 (N_3068,N_2921,N_2957);
or U3069 (N_3069,N_2917,N_2968);
nand U3070 (N_3070,N_2979,N_2984);
or U3071 (N_3071,N_2937,N_2903);
and U3072 (N_3072,N_2944,N_2970);
or U3073 (N_3073,N_2908,N_2932);
nor U3074 (N_3074,N_2959,N_2952);
nand U3075 (N_3075,N_2901,N_2990);
or U3076 (N_3076,N_2996,N_2962);
or U3077 (N_3077,N_2981,N_2928);
nand U3078 (N_3078,N_2919,N_2905);
and U3079 (N_3079,N_2901,N_2920);
nand U3080 (N_3080,N_2948,N_2979);
or U3081 (N_3081,N_2953,N_2949);
nand U3082 (N_3082,N_2958,N_2946);
xor U3083 (N_3083,N_2964,N_2987);
nand U3084 (N_3084,N_2946,N_2997);
and U3085 (N_3085,N_2927,N_2940);
nand U3086 (N_3086,N_2995,N_2967);
or U3087 (N_3087,N_2980,N_2996);
nand U3088 (N_3088,N_2908,N_2961);
or U3089 (N_3089,N_2991,N_2970);
nand U3090 (N_3090,N_2962,N_2993);
nor U3091 (N_3091,N_2980,N_2973);
or U3092 (N_3092,N_2909,N_2970);
and U3093 (N_3093,N_2968,N_2999);
nand U3094 (N_3094,N_2939,N_2984);
nand U3095 (N_3095,N_2968,N_2946);
nand U3096 (N_3096,N_2955,N_2989);
nor U3097 (N_3097,N_2945,N_2993);
or U3098 (N_3098,N_2930,N_2982);
or U3099 (N_3099,N_2973,N_2921);
nand U3100 (N_3100,N_3032,N_3038);
nand U3101 (N_3101,N_3088,N_3061);
nand U3102 (N_3102,N_3025,N_3017);
xor U3103 (N_3103,N_3076,N_3085);
xor U3104 (N_3104,N_3027,N_3018);
nand U3105 (N_3105,N_3051,N_3029);
and U3106 (N_3106,N_3054,N_3042);
or U3107 (N_3107,N_3055,N_3048);
or U3108 (N_3108,N_3007,N_3014);
or U3109 (N_3109,N_3053,N_3010);
nand U3110 (N_3110,N_3033,N_3099);
nor U3111 (N_3111,N_3068,N_3003);
nor U3112 (N_3112,N_3049,N_3050);
and U3113 (N_3113,N_3031,N_3034);
nor U3114 (N_3114,N_3071,N_3060);
nor U3115 (N_3115,N_3078,N_3091);
nand U3116 (N_3116,N_3075,N_3044);
or U3117 (N_3117,N_3011,N_3022);
nand U3118 (N_3118,N_3024,N_3095);
nand U3119 (N_3119,N_3016,N_3040);
nand U3120 (N_3120,N_3063,N_3065);
nand U3121 (N_3121,N_3004,N_3058);
xor U3122 (N_3122,N_3039,N_3072);
and U3123 (N_3123,N_3002,N_3020);
or U3124 (N_3124,N_3006,N_3036);
or U3125 (N_3125,N_3023,N_3087);
nand U3126 (N_3126,N_3047,N_3043);
xor U3127 (N_3127,N_3093,N_3056);
nor U3128 (N_3128,N_3096,N_3090);
nand U3129 (N_3129,N_3041,N_3086);
or U3130 (N_3130,N_3080,N_3045);
nor U3131 (N_3131,N_3001,N_3092);
nand U3132 (N_3132,N_3057,N_3013);
or U3133 (N_3133,N_3052,N_3035);
nor U3134 (N_3134,N_3081,N_3064);
or U3135 (N_3135,N_3015,N_3069);
or U3136 (N_3136,N_3009,N_3079);
nand U3137 (N_3137,N_3059,N_3097);
nor U3138 (N_3138,N_3084,N_3067);
nand U3139 (N_3139,N_3021,N_3012);
or U3140 (N_3140,N_3083,N_3030);
nor U3141 (N_3141,N_3028,N_3005);
and U3142 (N_3142,N_3098,N_3077);
and U3143 (N_3143,N_3037,N_3062);
or U3144 (N_3144,N_3026,N_3046);
or U3145 (N_3145,N_3070,N_3089);
or U3146 (N_3146,N_3073,N_3074);
and U3147 (N_3147,N_3000,N_3094);
nand U3148 (N_3148,N_3019,N_3066);
and U3149 (N_3149,N_3008,N_3082);
and U3150 (N_3150,N_3070,N_3055);
or U3151 (N_3151,N_3011,N_3004);
nand U3152 (N_3152,N_3016,N_3074);
or U3153 (N_3153,N_3049,N_3013);
and U3154 (N_3154,N_3005,N_3089);
and U3155 (N_3155,N_3011,N_3099);
or U3156 (N_3156,N_3078,N_3072);
or U3157 (N_3157,N_3009,N_3035);
and U3158 (N_3158,N_3055,N_3035);
nand U3159 (N_3159,N_3035,N_3042);
nor U3160 (N_3160,N_3099,N_3022);
nor U3161 (N_3161,N_3019,N_3018);
and U3162 (N_3162,N_3013,N_3097);
and U3163 (N_3163,N_3096,N_3082);
nor U3164 (N_3164,N_3066,N_3016);
nand U3165 (N_3165,N_3032,N_3084);
and U3166 (N_3166,N_3073,N_3058);
and U3167 (N_3167,N_3097,N_3075);
or U3168 (N_3168,N_3041,N_3022);
nor U3169 (N_3169,N_3085,N_3041);
nor U3170 (N_3170,N_3046,N_3022);
nor U3171 (N_3171,N_3070,N_3075);
and U3172 (N_3172,N_3074,N_3078);
and U3173 (N_3173,N_3014,N_3051);
or U3174 (N_3174,N_3001,N_3073);
nand U3175 (N_3175,N_3084,N_3093);
xor U3176 (N_3176,N_3027,N_3032);
nor U3177 (N_3177,N_3048,N_3034);
nor U3178 (N_3178,N_3099,N_3023);
and U3179 (N_3179,N_3005,N_3001);
and U3180 (N_3180,N_3017,N_3071);
nor U3181 (N_3181,N_3050,N_3079);
nor U3182 (N_3182,N_3047,N_3079);
or U3183 (N_3183,N_3085,N_3004);
xor U3184 (N_3184,N_3066,N_3040);
and U3185 (N_3185,N_3084,N_3059);
or U3186 (N_3186,N_3025,N_3077);
xnor U3187 (N_3187,N_3002,N_3053);
and U3188 (N_3188,N_3097,N_3077);
nor U3189 (N_3189,N_3005,N_3046);
or U3190 (N_3190,N_3026,N_3034);
or U3191 (N_3191,N_3047,N_3074);
nand U3192 (N_3192,N_3002,N_3090);
or U3193 (N_3193,N_3077,N_3004);
and U3194 (N_3194,N_3061,N_3071);
nand U3195 (N_3195,N_3071,N_3002);
nor U3196 (N_3196,N_3034,N_3043);
nor U3197 (N_3197,N_3000,N_3073);
and U3198 (N_3198,N_3001,N_3098);
or U3199 (N_3199,N_3054,N_3086);
nand U3200 (N_3200,N_3196,N_3133);
and U3201 (N_3201,N_3100,N_3157);
or U3202 (N_3202,N_3122,N_3142);
and U3203 (N_3203,N_3155,N_3120);
and U3204 (N_3204,N_3147,N_3126);
nand U3205 (N_3205,N_3182,N_3162);
nor U3206 (N_3206,N_3101,N_3130);
and U3207 (N_3207,N_3174,N_3105);
and U3208 (N_3208,N_3188,N_3173);
nor U3209 (N_3209,N_3197,N_3123);
nand U3210 (N_3210,N_3154,N_3134);
or U3211 (N_3211,N_3136,N_3168);
nand U3212 (N_3212,N_3107,N_3160);
nand U3213 (N_3213,N_3193,N_3113);
nor U3214 (N_3214,N_3180,N_3138);
and U3215 (N_3215,N_3170,N_3111);
or U3216 (N_3216,N_3141,N_3108);
nor U3217 (N_3217,N_3139,N_3125);
and U3218 (N_3218,N_3159,N_3128);
nand U3219 (N_3219,N_3143,N_3177);
nand U3220 (N_3220,N_3109,N_3103);
nand U3221 (N_3221,N_3186,N_3117);
or U3222 (N_3222,N_3119,N_3129);
or U3223 (N_3223,N_3184,N_3112);
nand U3224 (N_3224,N_3169,N_3151);
and U3225 (N_3225,N_3163,N_3140);
or U3226 (N_3226,N_3185,N_3172);
nand U3227 (N_3227,N_3115,N_3132);
nand U3228 (N_3228,N_3198,N_3148);
and U3229 (N_3229,N_3191,N_3127);
nand U3230 (N_3230,N_3124,N_3145);
xnor U3231 (N_3231,N_3149,N_3195);
and U3232 (N_3232,N_3152,N_3102);
nand U3233 (N_3233,N_3118,N_3110);
or U3234 (N_3234,N_3137,N_3167);
and U3235 (N_3235,N_3153,N_3165);
nand U3236 (N_3236,N_3146,N_3187);
nand U3237 (N_3237,N_3189,N_3116);
nor U3238 (N_3238,N_3178,N_3158);
nand U3239 (N_3239,N_3183,N_3150);
nand U3240 (N_3240,N_3156,N_3194);
nand U3241 (N_3241,N_3179,N_3181);
or U3242 (N_3242,N_3104,N_3106);
nand U3243 (N_3243,N_3166,N_3190);
nand U3244 (N_3244,N_3171,N_3135);
nand U3245 (N_3245,N_3114,N_3121);
or U3246 (N_3246,N_3164,N_3161);
nand U3247 (N_3247,N_3199,N_3192);
nand U3248 (N_3248,N_3176,N_3175);
and U3249 (N_3249,N_3144,N_3131);
nor U3250 (N_3250,N_3148,N_3100);
nor U3251 (N_3251,N_3145,N_3168);
or U3252 (N_3252,N_3188,N_3198);
and U3253 (N_3253,N_3106,N_3161);
or U3254 (N_3254,N_3122,N_3100);
or U3255 (N_3255,N_3136,N_3137);
or U3256 (N_3256,N_3194,N_3190);
nor U3257 (N_3257,N_3125,N_3184);
xnor U3258 (N_3258,N_3199,N_3124);
or U3259 (N_3259,N_3174,N_3156);
and U3260 (N_3260,N_3161,N_3141);
and U3261 (N_3261,N_3157,N_3174);
or U3262 (N_3262,N_3142,N_3150);
nand U3263 (N_3263,N_3118,N_3158);
nor U3264 (N_3264,N_3185,N_3177);
nor U3265 (N_3265,N_3125,N_3137);
nor U3266 (N_3266,N_3102,N_3170);
nand U3267 (N_3267,N_3104,N_3105);
or U3268 (N_3268,N_3192,N_3141);
nor U3269 (N_3269,N_3193,N_3196);
nand U3270 (N_3270,N_3137,N_3108);
or U3271 (N_3271,N_3111,N_3196);
nor U3272 (N_3272,N_3169,N_3155);
nand U3273 (N_3273,N_3190,N_3155);
nand U3274 (N_3274,N_3123,N_3114);
or U3275 (N_3275,N_3167,N_3198);
or U3276 (N_3276,N_3161,N_3159);
nor U3277 (N_3277,N_3178,N_3116);
nand U3278 (N_3278,N_3143,N_3176);
or U3279 (N_3279,N_3111,N_3178);
or U3280 (N_3280,N_3158,N_3121);
and U3281 (N_3281,N_3134,N_3139);
xnor U3282 (N_3282,N_3157,N_3138);
and U3283 (N_3283,N_3107,N_3102);
or U3284 (N_3284,N_3118,N_3121);
xor U3285 (N_3285,N_3139,N_3107);
or U3286 (N_3286,N_3120,N_3130);
and U3287 (N_3287,N_3183,N_3167);
nand U3288 (N_3288,N_3113,N_3134);
nor U3289 (N_3289,N_3150,N_3180);
and U3290 (N_3290,N_3129,N_3102);
nor U3291 (N_3291,N_3159,N_3174);
nand U3292 (N_3292,N_3173,N_3126);
or U3293 (N_3293,N_3181,N_3142);
nand U3294 (N_3294,N_3172,N_3126);
or U3295 (N_3295,N_3189,N_3138);
nor U3296 (N_3296,N_3168,N_3159);
or U3297 (N_3297,N_3138,N_3100);
nand U3298 (N_3298,N_3148,N_3116);
nand U3299 (N_3299,N_3167,N_3170);
nor U3300 (N_3300,N_3208,N_3286);
nor U3301 (N_3301,N_3247,N_3265);
nand U3302 (N_3302,N_3299,N_3230);
and U3303 (N_3303,N_3238,N_3224);
or U3304 (N_3304,N_3200,N_3267);
or U3305 (N_3305,N_3268,N_3233);
and U3306 (N_3306,N_3262,N_3205);
or U3307 (N_3307,N_3217,N_3220);
nor U3308 (N_3308,N_3250,N_3234);
nor U3309 (N_3309,N_3207,N_3219);
and U3310 (N_3310,N_3275,N_3229);
nor U3311 (N_3311,N_3239,N_3295);
nor U3312 (N_3312,N_3251,N_3289);
nand U3313 (N_3313,N_3288,N_3227);
or U3314 (N_3314,N_3270,N_3298);
or U3315 (N_3315,N_3257,N_3246);
or U3316 (N_3316,N_3294,N_3218);
nor U3317 (N_3317,N_3261,N_3241);
or U3318 (N_3318,N_3221,N_3282);
and U3319 (N_3319,N_3287,N_3263);
xnor U3320 (N_3320,N_3209,N_3201);
or U3321 (N_3321,N_3280,N_3264);
nor U3322 (N_3322,N_3253,N_3248);
or U3323 (N_3323,N_3215,N_3240);
nand U3324 (N_3324,N_3276,N_3204);
nand U3325 (N_3325,N_3271,N_3285);
nor U3326 (N_3326,N_3252,N_3293);
nor U3327 (N_3327,N_3242,N_3256);
nand U3328 (N_3328,N_3206,N_3272);
nand U3329 (N_3329,N_3266,N_3213);
or U3330 (N_3330,N_3243,N_3260);
nand U3331 (N_3331,N_3296,N_3212);
nor U3332 (N_3332,N_3258,N_3223);
and U3333 (N_3333,N_3297,N_3274);
nand U3334 (N_3334,N_3203,N_3225);
nor U3335 (N_3335,N_3292,N_3259);
or U3336 (N_3336,N_3231,N_3254);
and U3337 (N_3337,N_3236,N_3273);
nand U3338 (N_3338,N_3255,N_3269);
nor U3339 (N_3339,N_3278,N_3210);
nor U3340 (N_3340,N_3235,N_3202);
nand U3341 (N_3341,N_3279,N_3216);
nor U3342 (N_3342,N_3249,N_3284);
nand U3343 (N_3343,N_3222,N_3226);
nor U3344 (N_3344,N_3291,N_3211);
nor U3345 (N_3345,N_3237,N_3281);
nor U3346 (N_3346,N_3214,N_3277);
nor U3347 (N_3347,N_3283,N_3228);
nor U3348 (N_3348,N_3232,N_3244);
nand U3349 (N_3349,N_3245,N_3290);
nor U3350 (N_3350,N_3233,N_3205);
nor U3351 (N_3351,N_3263,N_3278);
or U3352 (N_3352,N_3209,N_3287);
nand U3353 (N_3353,N_3257,N_3293);
nand U3354 (N_3354,N_3251,N_3216);
nor U3355 (N_3355,N_3280,N_3286);
nand U3356 (N_3356,N_3290,N_3204);
or U3357 (N_3357,N_3209,N_3203);
or U3358 (N_3358,N_3205,N_3226);
nor U3359 (N_3359,N_3227,N_3259);
nor U3360 (N_3360,N_3269,N_3202);
or U3361 (N_3361,N_3261,N_3227);
and U3362 (N_3362,N_3207,N_3273);
or U3363 (N_3363,N_3238,N_3279);
and U3364 (N_3364,N_3296,N_3255);
and U3365 (N_3365,N_3282,N_3229);
nand U3366 (N_3366,N_3246,N_3262);
and U3367 (N_3367,N_3208,N_3230);
nor U3368 (N_3368,N_3268,N_3267);
or U3369 (N_3369,N_3263,N_3208);
nand U3370 (N_3370,N_3252,N_3241);
nor U3371 (N_3371,N_3249,N_3221);
or U3372 (N_3372,N_3287,N_3202);
nand U3373 (N_3373,N_3281,N_3257);
or U3374 (N_3374,N_3228,N_3252);
nor U3375 (N_3375,N_3282,N_3218);
nor U3376 (N_3376,N_3257,N_3274);
and U3377 (N_3377,N_3269,N_3284);
nand U3378 (N_3378,N_3238,N_3298);
or U3379 (N_3379,N_3210,N_3220);
nand U3380 (N_3380,N_3252,N_3226);
and U3381 (N_3381,N_3252,N_3250);
nand U3382 (N_3382,N_3270,N_3248);
and U3383 (N_3383,N_3203,N_3235);
or U3384 (N_3384,N_3222,N_3225);
nor U3385 (N_3385,N_3224,N_3285);
xnor U3386 (N_3386,N_3205,N_3219);
and U3387 (N_3387,N_3247,N_3269);
or U3388 (N_3388,N_3291,N_3272);
nand U3389 (N_3389,N_3254,N_3243);
nor U3390 (N_3390,N_3205,N_3238);
and U3391 (N_3391,N_3231,N_3220);
and U3392 (N_3392,N_3298,N_3222);
and U3393 (N_3393,N_3258,N_3209);
or U3394 (N_3394,N_3269,N_3270);
nor U3395 (N_3395,N_3271,N_3217);
nand U3396 (N_3396,N_3245,N_3222);
and U3397 (N_3397,N_3238,N_3248);
nor U3398 (N_3398,N_3203,N_3210);
nor U3399 (N_3399,N_3243,N_3265);
nand U3400 (N_3400,N_3343,N_3302);
nor U3401 (N_3401,N_3308,N_3321);
nand U3402 (N_3402,N_3378,N_3337);
or U3403 (N_3403,N_3358,N_3327);
and U3404 (N_3404,N_3355,N_3380);
or U3405 (N_3405,N_3399,N_3373);
nor U3406 (N_3406,N_3395,N_3352);
nand U3407 (N_3407,N_3375,N_3379);
or U3408 (N_3408,N_3388,N_3336);
and U3409 (N_3409,N_3349,N_3338);
nand U3410 (N_3410,N_3329,N_3344);
and U3411 (N_3411,N_3312,N_3357);
and U3412 (N_3412,N_3384,N_3350);
and U3413 (N_3413,N_3319,N_3383);
and U3414 (N_3414,N_3332,N_3323);
nor U3415 (N_3415,N_3301,N_3348);
or U3416 (N_3416,N_3305,N_3307);
or U3417 (N_3417,N_3389,N_3333);
and U3418 (N_3418,N_3371,N_3341);
nand U3419 (N_3419,N_3342,N_3316);
nand U3420 (N_3420,N_3306,N_3372);
nand U3421 (N_3421,N_3325,N_3377);
or U3422 (N_3422,N_3346,N_3311);
xnor U3423 (N_3423,N_3366,N_3351);
or U3424 (N_3424,N_3387,N_3328);
nor U3425 (N_3425,N_3361,N_3376);
nor U3426 (N_3426,N_3360,N_3340);
nand U3427 (N_3427,N_3310,N_3397);
nor U3428 (N_3428,N_3370,N_3368);
nand U3429 (N_3429,N_3369,N_3304);
and U3430 (N_3430,N_3322,N_3335);
or U3431 (N_3431,N_3393,N_3309);
nand U3432 (N_3432,N_3330,N_3318);
or U3433 (N_3433,N_3356,N_3359);
and U3434 (N_3434,N_3364,N_3334);
nor U3435 (N_3435,N_3363,N_3391);
nor U3436 (N_3436,N_3324,N_3354);
nor U3437 (N_3437,N_3386,N_3315);
nor U3438 (N_3438,N_3314,N_3317);
and U3439 (N_3439,N_3392,N_3353);
nor U3440 (N_3440,N_3300,N_3374);
and U3441 (N_3441,N_3381,N_3331);
nor U3442 (N_3442,N_3367,N_3320);
nand U3443 (N_3443,N_3390,N_3303);
nor U3444 (N_3444,N_3396,N_3394);
or U3445 (N_3445,N_3398,N_3339);
or U3446 (N_3446,N_3326,N_3345);
nor U3447 (N_3447,N_3365,N_3382);
or U3448 (N_3448,N_3313,N_3347);
and U3449 (N_3449,N_3362,N_3385);
nor U3450 (N_3450,N_3368,N_3388);
nor U3451 (N_3451,N_3386,N_3366);
nand U3452 (N_3452,N_3340,N_3381);
nand U3453 (N_3453,N_3399,N_3390);
and U3454 (N_3454,N_3368,N_3320);
nor U3455 (N_3455,N_3370,N_3396);
nand U3456 (N_3456,N_3323,N_3311);
xor U3457 (N_3457,N_3386,N_3304);
nand U3458 (N_3458,N_3381,N_3374);
or U3459 (N_3459,N_3330,N_3368);
or U3460 (N_3460,N_3316,N_3326);
or U3461 (N_3461,N_3343,N_3375);
nor U3462 (N_3462,N_3317,N_3300);
nand U3463 (N_3463,N_3358,N_3314);
or U3464 (N_3464,N_3372,N_3339);
and U3465 (N_3465,N_3382,N_3357);
nor U3466 (N_3466,N_3350,N_3324);
nor U3467 (N_3467,N_3364,N_3391);
and U3468 (N_3468,N_3384,N_3363);
and U3469 (N_3469,N_3304,N_3318);
nor U3470 (N_3470,N_3321,N_3387);
or U3471 (N_3471,N_3316,N_3379);
nor U3472 (N_3472,N_3393,N_3324);
nor U3473 (N_3473,N_3327,N_3360);
or U3474 (N_3474,N_3310,N_3347);
xnor U3475 (N_3475,N_3391,N_3323);
nor U3476 (N_3476,N_3333,N_3376);
nor U3477 (N_3477,N_3389,N_3359);
and U3478 (N_3478,N_3348,N_3383);
and U3479 (N_3479,N_3344,N_3306);
or U3480 (N_3480,N_3308,N_3399);
or U3481 (N_3481,N_3327,N_3312);
nand U3482 (N_3482,N_3373,N_3344);
nand U3483 (N_3483,N_3357,N_3343);
or U3484 (N_3484,N_3329,N_3377);
nor U3485 (N_3485,N_3394,N_3351);
nor U3486 (N_3486,N_3301,N_3303);
nor U3487 (N_3487,N_3398,N_3356);
or U3488 (N_3488,N_3398,N_3300);
and U3489 (N_3489,N_3392,N_3366);
and U3490 (N_3490,N_3310,N_3365);
nand U3491 (N_3491,N_3316,N_3303);
nor U3492 (N_3492,N_3328,N_3350);
nor U3493 (N_3493,N_3330,N_3341);
and U3494 (N_3494,N_3302,N_3317);
nor U3495 (N_3495,N_3357,N_3316);
or U3496 (N_3496,N_3387,N_3318);
or U3497 (N_3497,N_3388,N_3335);
nor U3498 (N_3498,N_3370,N_3378);
nand U3499 (N_3499,N_3364,N_3388);
and U3500 (N_3500,N_3485,N_3463);
and U3501 (N_3501,N_3411,N_3429);
or U3502 (N_3502,N_3400,N_3490);
nor U3503 (N_3503,N_3407,N_3468);
nand U3504 (N_3504,N_3440,N_3423);
and U3505 (N_3505,N_3433,N_3439);
nor U3506 (N_3506,N_3450,N_3415);
nand U3507 (N_3507,N_3462,N_3442);
and U3508 (N_3508,N_3457,N_3483);
nor U3509 (N_3509,N_3458,N_3441);
nand U3510 (N_3510,N_3437,N_3491);
xnor U3511 (N_3511,N_3425,N_3413);
and U3512 (N_3512,N_3424,N_3477);
nor U3513 (N_3513,N_3469,N_3416);
nand U3514 (N_3514,N_3480,N_3452);
and U3515 (N_3515,N_3461,N_3474);
and U3516 (N_3516,N_3481,N_3436);
nand U3517 (N_3517,N_3476,N_3430);
nand U3518 (N_3518,N_3448,N_3451);
nor U3519 (N_3519,N_3486,N_3492);
nor U3520 (N_3520,N_3446,N_3418);
nor U3521 (N_3521,N_3421,N_3406);
or U3522 (N_3522,N_3464,N_3489);
and U3523 (N_3523,N_3449,N_3470);
nor U3524 (N_3524,N_3495,N_3459);
or U3525 (N_3525,N_3478,N_3498);
nor U3526 (N_3526,N_3456,N_3401);
or U3527 (N_3527,N_3405,N_3460);
nand U3528 (N_3528,N_3472,N_3465);
or U3529 (N_3529,N_3496,N_3494);
nand U3530 (N_3530,N_3482,N_3475);
xor U3531 (N_3531,N_3403,N_3427);
or U3532 (N_3532,N_3466,N_3454);
and U3533 (N_3533,N_3473,N_3420);
or U3534 (N_3534,N_3443,N_3493);
nor U3535 (N_3535,N_3414,N_3497);
or U3536 (N_3536,N_3431,N_3408);
nor U3537 (N_3537,N_3410,N_3471);
nand U3538 (N_3538,N_3467,N_3487);
xnor U3539 (N_3539,N_3404,N_3445);
or U3540 (N_3540,N_3453,N_3435);
and U3541 (N_3541,N_3402,N_3428);
and U3542 (N_3542,N_3444,N_3419);
nand U3543 (N_3543,N_3455,N_3412);
and U3544 (N_3544,N_3488,N_3438);
nor U3545 (N_3545,N_3499,N_3417);
nand U3546 (N_3546,N_3432,N_3426);
or U3547 (N_3547,N_3447,N_3409);
and U3548 (N_3548,N_3422,N_3434);
and U3549 (N_3549,N_3484,N_3479);
and U3550 (N_3550,N_3437,N_3463);
nor U3551 (N_3551,N_3430,N_3492);
and U3552 (N_3552,N_3462,N_3463);
and U3553 (N_3553,N_3496,N_3429);
and U3554 (N_3554,N_3432,N_3480);
or U3555 (N_3555,N_3439,N_3413);
and U3556 (N_3556,N_3499,N_3452);
or U3557 (N_3557,N_3417,N_3426);
nand U3558 (N_3558,N_3484,N_3423);
nand U3559 (N_3559,N_3482,N_3478);
nor U3560 (N_3560,N_3403,N_3441);
xor U3561 (N_3561,N_3444,N_3472);
and U3562 (N_3562,N_3492,N_3431);
or U3563 (N_3563,N_3463,N_3421);
nor U3564 (N_3564,N_3404,N_3495);
nor U3565 (N_3565,N_3433,N_3458);
nand U3566 (N_3566,N_3413,N_3415);
and U3567 (N_3567,N_3408,N_3446);
or U3568 (N_3568,N_3425,N_3458);
nor U3569 (N_3569,N_3445,N_3449);
xnor U3570 (N_3570,N_3443,N_3401);
nand U3571 (N_3571,N_3466,N_3449);
and U3572 (N_3572,N_3437,N_3405);
nor U3573 (N_3573,N_3414,N_3465);
nand U3574 (N_3574,N_3444,N_3434);
nand U3575 (N_3575,N_3466,N_3490);
or U3576 (N_3576,N_3409,N_3465);
nand U3577 (N_3577,N_3406,N_3489);
xnor U3578 (N_3578,N_3405,N_3402);
nor U3579 (N_3579,N_3434,N_3418);
and U3580 (N_3580,N_3460,N_3471);
and U3581 (N_3581,N_3439,N_3405);
nor U3582 (N_3582,N_3401,N_3486);
or U3583 (N_3583,N_3435,N_3406);
nor U3584 (N_3584,N_3488,N_3407);
or U3585 (N_3585,N_3485,N_3441);
nor U3586 (N_3586,N_3450,N_3473);
nand U3587 (N_3587,N_3410,N_3463);
nor U3588 (N_3588,N_3453,N_3492);
xor U3589 (N_3589,N_3466,N_3404);
or U3590 (N_3590,N_3409,N_3492);
nor U3591 (N_3591,N_3411,N_3439);
and U3592 (N_3592,N_3406,N_3459);
or U3593 (N_3593,N_3417,N_3498);
nand U3594 (N_3594,N_3400,N_3421);
and U3595 (N_3595,N_3419,N_3416);
nand U3596 (N_3596,N_3467,N_3415);
nor U3597 (N_3597,N_3485,N_3408);
or U3598 (N_3598,N_3499,N_3483);
or U3599 (N_3599,N_3439,N_3424);
and U3600 (N_3600,N_3546,N_3553);
or U3601 (N_3601,N_3590,N_3501);
and U3602 (N_3602,N_3532,N_3548);
or U3603 (N_3603,N_3574,N_3543);
and U3604 (N_3604,N_3514,N_3504);
and U3605 (N_3605,N_3584,N_3593);
or U3606 (N_3606,N_3579,N_3551);
or U3607 (N_3607,N_3500,N_3536);
or U3608 (N_3608,N_3559,N_3525);
and U3609 (N_3609,N_3518,N_3545);
nand U3610 (N_3610,N_3506,N_3552);
and U3611 (N_3611,N_3520,N_3503);
nor U3612 (N_3612,N_3519,N_3547);
and U3613 (N_3613,N_3516,N_3567);
or U3614 (N_3614,N_3595,N_3563);
nor U3615 (N_3615,N_3570,N_3573);
nor U3616 (N_3616,N_3527,N_3569);
or U3617 (N_3617,N_3588,N_3556);
or U3618 (N_3618,N_3538,N_3507);
nand U3619 (N_3619,N_3597,N_3526);
nor U3620 (N_3620,N_3565,N_3508);
nor U3621 (N_3621,N_3522,N_3576);
and U3622 (N_3622,N_3596,N_3557);
or U3623 (N_3623,N_3578,N_3564);
nand U3624 (N_3624,N_3542,N_3537);
or U3625 (N_3625,N_3550,N_3528);
and U3626 (N_3626,N_3530,N_3577);
and U3627 (N_3627,N_3587,N_3580);
nand U3628 (N_3628,N_3575,N_3592);
and U3629 (N_3629,N_3523,N_3572);
or U3630 (N_3630,N_3598,N_3502);
nor U3631 (N_3631,N_3586,N_3581);
and U3632 (N_3632,N_3599,N_3509);
or U3633 (N_3633,N_3539,N_3591);
and U3634 (N_3634,N_3585,N_3513);
nor U3635 (N_3635,N_3583,N_3534);
and U3636 (N_3636,N_3571,N_3589);
or U3637 (N_3637,N_3560,N_3594);
nor U3638 (N_3638,N_3540,N_3582);
nor U3639 (N_3639,N_3521,N_3529);
or U3640 (N_3640,N_3511,N_3562);
or U3641 (N_3641,N_3549,N_3555);
xnor U3642 (N_3642,N_3512,N_3554);
and U3643 (N_3643,N_3568,N_3541);
nor U3644 (N_3644,N_3535,N_3566);
nor U3645 (N_3645,N_3544,N_3561);
nor U3646 (N_3646,N_3517,N_3558);
and U3647 (N_3647,N_3510,N_3515);
or U3648 (N_3648,N_3531,N_3524);
nor U3649 (N_3649,N_3533,N_3505);
nor U3650 (N_3650,N_3558,N_3593);
and U3651 (N_3651,N_3507,N_3519);
or U3652 (N_3652,N_3523,N_3511);
or U3653 (N_3653,N_3507,N_3500);
or U3654 (N_3654,N_3588,N_3540);
or U3655 (N_3655,N_3592,N_3540);
nand U3656 (N_3656,N_3519,N_3549);
nor U3657 (N_3657,N_3502,N_3570);
nor U3658 (N_3658,N_3505,N_3585);
or U3659 (N_3659,N_3514,N_3586);
xnor U3660 (N_3660,N_3581,N_3544);
nand U3661 (N_3661,N_3566,N_3577);
or U3662 (N_3662,N_3569,N_3545);
and U3663 (N_3663,N_3598,N_3568);
and U3664 (N_3664,N_3526,N_3500);
and U3665 (N_3665,N_3582,N_3534);
nor U3666 (N_3666,N_3550,N_3576);
and U3667 (N_3667,N_3578,N_3530);
nand U3668 (N_3668,N_3597,N_3565);
nor U3669 (N_3669,N_3520,N_3570);
and U3670 (N_3670,N_3503,N_3529);
nand U3671 (N_3671,N_3544,N_3594);
nand U3672 (N_3672,N_3593,N_3594);
or U3673 (N_3673,N_3586,N_3521);
nand U3674 (N_3674,N_3553,N_3556);
or U3675 (N_3675,N_3586,N_3599);
xor U3676 (N_3676,N_3585,N_3533);
nor U3677 (N_3677,N_3555,N_3520);
nand U3678 (N_3678,N_3536,N_3522);
nand U3679 (N_3679,N_3568,N_3502);
nor U3680 (N_3680,N_3565,N_3593);
and U3681 (N_3681,N_3527,N_3557);
nor U3682 (N_3682,N_3549,N_3556);
nor U3683 (N_3683,N_3514,N_3530);
or U3684 (N_3684,N_3595,N_3569);
or U3685 (N_3685,N_3509,N_3585);
and U3686 (N_3686,N_3551,N_3595);
nand U3687 (N_3687,N_3557,N_3562);
nor U3688 (N_3688,N_3561,N_3598);
and U3689 (N_3689,N_3501,N_3560);
nor U3690 (N_3690,N_3506,N_3518);
or U3691 (N_3691,N_3595,N_3509);
and U3692 (N_3692,N_3526,N_3564);
or U3693 (N_3693,N_3579,N_3537);
or U3694 (N_3694,N_3513,N_3559);
nand U3695 (N_3695,N_3526,N_3531);
xnor U3696 (N_3696,N_3533,N_3508);
nand U3697 (N_3697,N_3503,N_3580);
nor U3698 (N_3698,N_3517,N_3553);
or U3699 (N_3699,N_3548,N_3583);
or U3700 (N_3700,N_3665,N_3672);
nor U3701 (N_3701,N_3644,N_3611);
and U3702 (N_3702,N_3691,N_3688);
or U3703 (N_3703,N_3694,N_3660);
nor U3704 (N_3704,N_3600,N_3696);
and U3705 (N_3705,N_3654,N_3662);
and U3706 (N_3706,N_3655,N_3626);
nor U3707 (N_3707,N_3682,N_3687);
nor U3708 (N_3708,N_3619,N_3678);
and U3709 (N_3709,N_3621,N_3604);
nor U3710 (N_3710,N_3658,N_3620);
nand U3711 (N_3711,N_3679,N_3638);
or U3712 (N_3712,N_3641,N_3607);
nand U3713 (N_3713,N_3601,N_3693);
nand U3714 (N_3714,N_3629,N_3645);
nand U3715 (N_3715,N_3615,N_3648);
and U3716 (N_3716,N_3657,N_3636);
nand U3717 (N_3717,N_3627,N_3622);
nand U3718 (N_3718,N_3639,N_3617);
nor U3719 (N_3719,N_3631,N_3612);
and U3720 (N_3720,N_3647,N_3668);
or U3721 (N_3721,N_3646,N_3669);
and U3722 (N_3722,N_3602,N_3603);
or U3723 (N_3723,N_3640,N_3699);
and U3724 (N_3724,N_3642,N_3616);
nor U3725 (N_3725,N_3606,N_3625);
nand U3726 (N_3726,N_3697,N_3661);
nand U3727 (N_3727,N_3650,N_3698);
nand U3728 (N_3728,N_3608,N_3695);
or U3729 (N_3729,N_3690,N_3663);
nor U3730 (N_3730,N_3651,N_3675);
nor U3731 (N_3731,N_3605,N_3609);
nand U3732 (N_3732,N_3674,N_3637);
and U3733 (N_3733,N_3613,N_3681);
and U3734 (N_3734,N_3680,N_3692);
or U3735 (N_3735,N_3683,N_3649);
and U3736 (N_3736,N_3659,N_3630);
or U3737 (N_3737,N_3623,N_3673);
nor U3738 (N_3738,N_3684,N_3634);
and U3739 (N_3739,N_3633,N_3667);
nand U3740 (N_3740,N_3664,N_3635);
xnor U3741 (N_3741,N_3677,N_3685);
or U3742 (N_3742,N_3689,N_3628);
and U3743 (N_3743,N_3656,N_3676);
xnor U3744 (N_3744,N_3614,N_3671);
nor U3745 (N_3745,N_3652,N_3686);
or U3746 (N_3746,N_3653,N_3618);
or U3747 (N_3747,N_3624,N_3643);
and U3748 (N_3748,N_3670,N_3632);
nor U3749 (N_3749,N_3666,N_3610);
nand U3750 (N_3750,N_3692,N_3667);
nand U3751 (N_3751,N_3660,N_3653);
or U3752 (N_3752,N_3637,N_3639);
or U3753 (N_3753,N_3693,N_3667);
or U3754 (N_3754,N_3622,N_3628);
and U3755 (N_3755,N_3635,N_3686);
nor U3756 (N_3756,N_3610,N_3605);
and U3757 (N_3757,N_3618,N_3691);
nand U3758 (N_3758,N_3671,N_3667);
xnor U3759 (N_3759,N_3633,N_3662);
and U3760 (N_3760,N_3674,N_3691);
nor U3761 (N_3761,N_3688,N_3632);
or U3762 (N_3762,N_3636,N_3621);
or U3763 (N_3763,N_3613,N_3657);
or U3764 (N_3764,N_3679,N_3641);
and U3765 (N_3765,N_3637,N_3609);
and U3766 (N_3766,N_3689,N_3648);
nand U3767 (N_3767,N_3688,N_3623);
nand U3768 (N_3768,N_3612,N_3632);
nor U3769 (N_3769,N_3696,N_3618);
nand U3770 (N_3770,N_3649,N_3612);
or U3771 (N_3771,N_3633,N_3682);
nor U3772 (N_3772,N_3636,N_3698);
nand U3773 (N_3773,N_3649,N_3621);
and U3774 (N_3774,N_3672,N_3650);
or U3775 (N_3775,N_3612,N_3671);
or U3776 (N_3776,N_3612,N_3640);
or U3777 (N_3777,N_3666,N_3637);
nand U3778 (N_3778,N_3660,N_3691);
nand U3779 (N_3779,N_3643,N_3661);
and U3780 (N_3780,N_3640,N_3603);
or U3781 (N_3781,N_3656,N_3679);
nand U3782 (N_3782,N_3629,N_3612);
or U3783 (N_3783,N_3660,N_3662);
and U3784 (N_3784,N_3640,N_3608);
nor U3785 (N_3785,N_3670,N_3613);
or U3786 (N_3786,N_3650,N_3611);
nor U3787 (N_3787,N_3611,N_3668);
and U3788 (N_3788,N_3651,N_3670);
nor U3789 (N_3789,N_3646,N_3601);
nand U3790 (N_3790,N_3675,N_3672);
and U3791 (N_3791,N_3614,N_3662);
nor U3792 (N_3792,N_3691,N_3695);
nor U3793 (N_3793,N_3648,N_3640);
or U3794 (N_3794,N_3690,N_3643);
and U3795 (N_3795,N_3690,N_3648);
and U3796 (N_3796,N_3611,N_3608);
nand U3797 (N_3797,N_3657,N_3616);
and U3798 (N_3798,N_3658,N_3600);
and U3799 (N_3799,N_3614,N_3653);
and U3800 (N_3800,N_3775,N_3746);
nor U3801 (N_3801,N_3785,N_3714);
or U3802 (N_3802,N_3712,N_3707);
and U3803 (N_3803,N_3735,N_3781);
nor U3804 (N_3804,N_3722,N_3737);
or U3805 (N_3805,N_3784,N_3742);
or U3806 (N_3806,N_3710,N_3749);
nand U3807 (N_3807,N_3769,N_3789);
nor U3808 (N_3808,N_3728,N_3726);
and U3809 (N_3809,N_3753,N_3734);
nor U3810 (N_3810,N_3773,N_3791);
and U3811 (N_3811,N_3709,N_3760);
nand U3812 (N_3812,N_3718,N_3771);
and U3813 (N_3813,N_3748,N_3732);
or U3814 (N_3814,N_3711,N_3750);
nor U3815 (N_3815,N_3717,N_3761);
nor U3816 (N_3816,N_3796,N_3754);
nor U3817 (N_3817,N_3758,N_3721);
nor U3818 (N_3818,N_3776,N_3700);
or U3819 (N_3819,N_3778,N_3763);
nand U3820 (N_3820,N_3768,N_3767);
and U3821 (N_3821,N_3715,N_3724);
and U3822 (N_3822,N_3731,N_3759);
nor U3823 (N_3823,N_3702,N_3727);
nor U3824 (N_3824,N_3747,N_3783);
nor U3825 (N_3825,N_3739,N_3762);
or U3826 (N_3826,N_3741,N_3770);
and U3827 (N_3827,N_3740,N_3713);
nand U3828 (N_3828,N_3798,N_3729);
nand U3829 (N_3829,N_3780,N_3751);
and U3830 (N_3830,N_3705,N_3792);
or U3831 (N_3831,N_3782,N_3706);
or U3832 (N_3832,N_3755,N_3797);
or U3833 (N_3833,N_3793,N_3766);
nor U3834 (N_3834,N_3720,N_3703);
xnor U3835 (N_3835,N_3790,N_3788);
nor U3836 (N_3836,N_3733,N_3765);
nor U3837 (N_3837,N_3701,N_3786);
and U3838 (N_3838,N_3774,N_3723);
nand U3839 (N_3839,N_3704,N_3744);
xor U3840 (N_3840,N_3756,N_3738);
and U3841 (N_3841,N_3779,N_3772);
nand U3842 (N_3842,N_3730,N_3799);
and U3843 (N_3843,N_3777,N_3745);
or U3844 (N_3844,N_3757,N_3795);
and U3845 (N_3845,N_3725,N_3743);
nand U3846 (N_3846,N_3752,N_3708);
and U3847 (N_3847,N_3794,N_3719);
or U3848 (N_3848,N_3716,N_3764);
and U3849 (N_3849,N_3736,N_3787);
nand U3850 (N_3850,N_3791,N_3781);
and U3851 (N_3851,N_3716,N_3714);
or U3852 (N_3852,N_3706,N_3770);
nor U3853 (N_3853,N_3704,N_3771);
nor U3854 (N_3854,N_3774,N_3794);
or U3855 (N_3855,N_3740,N_3793);
nor U3856 (N_3856,N_3731,N_3785);
nand U3857 (N_3857,N_3708,N_3773);
xnor U3858 (N_3858,N_3714,N_3713);
nor U3859 (N_3859,N_3785,N_3726);
and U3860 (N_3860,N_3790,N_3721);
nand U3861 (N_3861,N_3781,N_3782);
or U3862 (N_3862,N_3731,N_3771);
or U3863 (N_3863,N_3788,N_3756);
nor U3864 (N_3864,N_3775,N_3709);
nor U3865 (N_3865,N_3768,N_3765);
or U3866 (N_3866,N_3743,N_3753);
and U3867 (N_3867,N_3741,N_3783);
and U3868 (N_3868,N_3716,N_3752);
and U3869 (N_3869,N_3746,N_3710);
or U3870 (N_3870,N_3772,N_3794);
and U3871 (N_3871,N_3788,N_3791);
or U3872 (N_3872,N_3781,N_3724);
or U3873 (N_3873,N_3764,N_3746);
or U3874 (N_3874,N_3760,N_3722);
or U3875 (N_3875,N_3720,N_3757);
nor U3876 (N_3876,N_3721,N_3786);
nor U3877 (N_3877,N_3795,N_3749);
and U3878 (N_3878,N_3787,N_3781);
and U3879 (N_3879,N_3764,N_3790);
or U3880 (N_3880,N_3715,N_3708);
and U3881 (N_3881,N_3729,N_3733);
nand U3882 (N_3882,N_3718,N_3747);
nand U3883 (N_3883,N_3796,N_3762);
nand U3884 (N_3884,N_3796,N_3778);
nand U3885 (N_3885,N_3726,N_3700);
or U3886 (N_3886,N_3741,N_3796);
nor U3887 (N_3887,N_3772,N_3701);
or U3888 (N_3888,N_3789,N_3745);
nor U3889 (N_3889,N_3737,N_3728);
or U3890 (N_3890,N_3762,N_3715);
or U3891 (N_3891,N_3740,N_3792);
or U3892 (N_3892,N_3700,N_3793);
nor U3893 (N_3893,N_3756,N_3784);
or U3894 (N_3894,N_3782,N_3765);
and U3895 (N_3895,N_3728,N_3723);
or U3896 (N_3896,N_3795,N_3743);
nor U3897 (N_3897,N_3772,N_3769);
nand U3898 (N_3898,N_3793,N_3714);
nor U3899 (N_3899,N_3701,N_3741);
or U3900 (N_3900,N_3804,N_3814);
nor U3901 (N_3901,N_3899,N_3834);
nand U3902 (N_3902,N_3890,N_3851);
or U3903 (N_3903,N_3853,N_3865);
and U3904 (N_3904,N_3837,N_3871);
and U3905 (N_3905,N_3884,N_3832);
nor U3906 (N_3906,N_3801,N_3891);
nor U3907 (N_3907,N_3828,N_3898);
nor U3908 (N_3908,N_3840,N_3803);
nor U3909 (N_3909,N_3805,N_3836);
and U3910 (N_3910,N_3835,N_3819);
nand U3911 (N_3911,N_3876,N_3867);
nor U3912 (N_3912,N_3806,N_3823);
and U3913 (N_3913,N_3882,N_3892);
and U3914 (N_3914,N_3815,N_3813);
and U3915 (N_3915,N_3846,N_3820);
nand U3916 (N_3916,N_3856,N_3855);
nand U3917 (N_3917,N_3843,N_3872);
nand U3918 (N_3918,N_3879,N_3829);
nand U3919 (N_3919,N_3866,N_3838);
or U3920 (N_3920,N_3849,N_3818);
or U3921 (N_3921,N_3824,N_3850);
nand U3922 (N_3922,N_3878,N_3848);
and U3923 (N_3923,N_3864,N_3881);
nor U3924 (N_3924,N_3852,N_3817);
or U3925 (N_3925,N_3897,N_3880);
nand U3926 (N_3926,N_3812,N_3810);
or U3927 (N_3927,N_3886,N_3845);
nand U3928 (N_3928,N_3889,N_3883);
nand U3929 (N_3929,N_3862,N_3807);
nor U3930 (N_3930,N_3802,N_3844);
xnor U3931 (N_3931,N_3861,N_3859);
or U3932 (N_3932,N_3842,N_3833);
and U3933 (N_3933,N_3860,N_3857);
or U3934 (N_3934,N_3874,N_3863);
and U3935 (N_3935,N_3858,N_3822);
nor U3936 (N_3936,N_3825,N_3887);
nand U3937 (N_3937,N_3831,N_3809);
or U3938 (N_3938,N_3875,N_3873);
or U3939 (N_3939,N_3869,N_3800);
nand U3940 (N_3940,N_3821,N_3847);
and U3941 (N_3941,N_3854,N_3877);
nand U3942 (N_3942,N_3893,N_3841);
nand U3943 (N_3943,N_3870,N_3888);
and U3944 (N_3944,N_3896,N_3894);
nor U3945 (N_3945,N_3868,N_3826);
nor U3946 (N_3946,N_3808,N_3885);
or U3947 (N_3947,N_3830,N_3816);
nand U3948 (N_3948,N_3839,N_3827);
nand U3949 (N_3949,N_3811,N_3895);
nor U3950 (N_3950,N_3841,N_3865);
or U3951 (N_3951,N_3829,N_3883);
or U3952 (N_3952,N_3853,N_3898);
or U3953 (N_3953,N_3846,N_3876);
and U3954 (N_3954,N_3819,N_3881);
nor U3955 (N_3955,N_3824,N_3864);
or U3956 (N_3956,N_3862,N_3884);
or U3957 (N_3957,N_3826,N_3832);
nor U3958 (N_3958,N_3875,N_3832);
and U3959 (N_3959,N_3842,N_3854);
or U3960 (N_3960,N_3890,N_3874);
nand U3961 (N_3961,N_3844,N_3895);
nor U3962 (N_3962,N_3817,N_3865);
and U3963 (N_3963,N_3878,N_3814);
and U3964 (N_3964,N_3883,N_3817);
nor U3965 (N_3965,N_3864,N_3890);
nor U3966 (N_3966,N_3893,N_3898);
nand U3967 (N_3967,N_3803,N_3823);
nand U3968 (N_3968,N_3821,N_3826);
nand U3969 (N_3969,N_3808,N_3866);
and U3970 (N_3970,N_3897,N_3854);
nand U3971 (N_3971,N_3884,N_3838);
nand U3972 (N_3972,N_3863,N_3839);
nor U3973 (N_3973,N_3866,N_3864);
or U3974 (N_3974,N_3897,N_3881);
and U3975 (N_3975,N_3801,N_3847);
nand U3976 (N_3976,N_3847,N_3898);
and U3977 (N_3977,N_3805,N_3824);
and U3978 (N_3978,N_3878,N_3811);
nand U3979 (N_3979,N_3879,N_3840);
nor U3980 (N_3980,N_3836,N_3820);
nand U3981 (N_3981,N_3861,N_3863);
nand U3982 (N_3982,N_3858,N_3842);
or U3983 (N_3983,N_3825,N_3839);
nor U3984 (N_3984,N_3810,N_3841);
nand U3985 (N_3985,N_3824,N_3825);
or U3986 (N_3986,N_3852,N_3892);
and U3987 (N_3987,N_3825,N_3808);
or U3988 (N_3988,N_3883,N_3881);
nand U3989 (N_3989,N_3876,N_3899);
nor U3990 (N_3990,N_3872,N_3883);
and U3991 (N_3991,N_3867,N_3890);
nor U3992 (N_3992,N_3883,N_3862);
and U3993 (N_3993,N_3888,N_3860);
nand U3994 (N_3994,N_3823,N_3870);
nand U3995 (N_3995,N_3873,N_3824);
or U3996 (N_3996,N_3813,N_3845);
nand U3997 (N_3997,N_3805,N_3841);
and U3998 (N_3998,N_3848,N_3829);
nand U3999 (N_3999,N_3838,N_3840);
nand U4000 (N_4000,N_3971,N_3976);
and U4001 (N_4001,N_3996,N_3931);
nand U4002 (N_4002,N_3912,N_3919);
nor U4003 (N_4003,N_3917,N_3972);
nand U4004 (N_4004,N_3960,N_3982);
nor U4005 (N_4005,N_3997,N_3907);
nor U4006 (N_4006,N_3995,N_3928);
nand U4007 (N_4007,N_3905,N_3944);
and U4008 (N_4008,N_3989,N_3908);
nor U4009 (N_4009,N_3923,N_3925);
or U4010 (N_4010,N_3965,N_3947);
nor U4011 (N_4011,N_3929,N_3934);
and U4012 (N_4012,N_3924,N_3926);
xnor U4013 (N_4013,N_3951,N_3910);
nand U4014 (N_4014,N_3988,N_3903);
nand U4015 (N_4015,N_3954,N_3969);
nor U4016 (N_4016,N_3973,N_3978);
and U4017 (N_4017,N_3932,N_3992);
or U4018 (N_4018,N_3958,N_3911);
and U4019 (N_4019,N_3940,N_3999);
nand U4020 (N_4020,N_3987,N_3914);
or U4021 (N_4021,N_3990,N_3955);
nor U4022 (N_4022,N_3985,N_3902);
nand U4023 (N_4023,N_3922,N_3977);
nor U4024 (N_4024,N_3964,N_3906);
nor U4025 (N_4025,N_3937,N_3980);
nand U4026 (N_4026,N_3963,N_3946);
nand U4027 (N_4027,N_3949,N_3975);
nand U4028 (N_4028,N_3984,N_3901);
and U4029 (N_4029,N_3938,N_3933);
or U4030 (N_4030,N_3900,N_3916);
nor U4031 (N_4031,N_3956,N_3974);
xor U4032 (N_4032,N_3993,N_3909);
xnor U4033 (N_4033,N_3998,N_3913);
or U4034 (N_4034,N_3939,N_3921);
nor U4035 (N_4035,N_3915,N_3953);
and U4036 (N_4036,N_3983,N_3961);
nand U4037 (N_4037,N_3904,N_3966);
or U4038 (N_4038,N_3935,N_3981);
or U4039 (N_4039,N_3920,N_3991);
nand U4040 (N_4040,N_3986,N_3936);
nor U4041 (N_4041,N_3967,N_3962);
nor U4042 (N_4042,N_3970,N_3957);
xor U4043 (N_4043,N_3979,N_3950);
nand U4044 (N_4044,N_3945,N_3948);
nor U4045 (N_4045,N_3943,N_3952);
xnor U4046 (N_4046,N_3941,N_3918);
and U4047 (N_4047,N_3942,N_3994);
xor U4048 (N_4048,N_3959,N_3927);
or U4049 (N_4049,N_3930,N_3968);
nand U4050 (N_4050,N_3904,N_3902);
nand U4051 (N_4051,N_3959,N_3955);
nand U4052 (N_4052,N_3947,N_3960);
nor U4053 (N_4053,N_3983,N_3927);
nand U4054 (N_4054,N_3966,N_3928);
nand U4055 (N_4055,N_3990,N_3923);
or U4056 (N_4056,N_3926,N_3996);
or U4057 (N_4057,N_3901,N_3972);
or U4058 (N_4058,N_3986,N_3929);
or U4059 (N_4059,N_3960,N_3968);
nand U4060 (N_4060,N_3941,N_3956);
nand U4061 (N_4061,N_3938,N_3956);
nand U4062 (N_4062,N_3930,N_3925);
nand U4063 (N_4063,N_3938,N_3916);
or U4064 (N_4064,N_3910,N_3994);
nand U4065 (N_4065,N_3923,N_3961);
and U4066 (N_4066,N_3952,N_3996);
nor U4067 (N_4067,N_3974,N_3976);
nand U4068 (N_4068,N_3963,N_3987);
or U4069 (N_4069,N_3952,N_3926);
and U4070 (N_4070,N_3930,N_3935);
nor U4071 (N_4071,N_3930,N_3967);
xor U4072 (N_4072,N_3969,N_3943);
nand U4073 (N_4073,N_3924,N_3939);
or U4074 (N_4074,N_3982,N_3925);
or U4075 (N_4075,N_3932,N_3959);
or U4076 (N_4076,N_3954,N_3927);
and U4077 (N_4077,N_3930,N_3950);
or U4078 (N_4078,N_3911,N_3989);
or U4079 (N_4079,N_3942,N_3984);
nand U4080 (N_4080,N_3910,N_3903);
nand U4081 (N_4081,N_3972,N_3980);
and U4082 (N_4082,N_3916,N_3905);
nor U4083 (N_4083,N_3931,N_3912);
or U4084 (N_4084,N_3991,N_3961);
and U4085 (N_4085,N_3935,N_3990);
nand U4086 (N_4086,N_3925,N_3918);
nand U4087 (N_4087,N_3937,N_3905);
and U4088 (N_4088,N_3943,N_3985);
and U4089 (N_4089,N_3901,N_3940);
nand U4090 (N_4090,N_3931,N_3954);
or U4091 (N_4091,N_3953,N_3951);
or U4092 (N_4092,N_3951,N_3961);
and U4093 (N_4093,N_3975,N_3938);
nand U4094 (N_4094,N_3960,N_3931);
or U4095 (N_4095,N_3961,N_3939);
or U4096 (N_4096,N_3970,N_3947);
xnor U4097 (N_4097,N_3951,N_3997);
nor U4098 (N_4098,N_3975,N_3953);
nor U4099 (N_4099,N_3934,N_3962);
and U4100 (N_4100,N_4089,N_4032);
xnor U4101 (N_4101,N_4004,N_4040);
nor U4102 (N_4102,N_4061,N_4085);
xor U4103 (N_4103,N_4025,N_4022);
and U4104 (N_4104,N_4028,N_4046);
and U4105 (N_4105,N_4002,N_4067);
nand U4106 (N_4106,N_4091,N_4095);
or U4107 (N_4107,N_4055,N_4053);
nand U4108 (N_4108,N_4012,N_4069);
nand U4109 (N_4109,N_4072,N_4020);
or U4110 (N_4110,N_4011,N_4001);
and U4111 (N_4111,N_4041,N_4000);
or U4112 (N_4112,N_4026,N_4052);
nor U4113 (N_4113,N_4008,N_4080);
and U4114 (N_4114,N_4083,N_4050);
and U4115 (N_4115,N_4010,N_4078);
and U4116 (N_4116,N_4079,N_4084);
nand U4117 (N_4117,N_4098,N_4019);
nand U4118 (N_4118,N_4054,N_4034);
xnor U4119 (N_4119,N_4070,N_4013);
and U4120 (N_4120,N_4039,N_4092);
and U4121 (N_4121,N_4087,N_4076);
and U4122 (N_4122,N_4037,N_4062);
or U4123 (N_4123,N_4017,N_4096);
and U4124 (N_4124,N_4093,N_4063);
or U4125 (N_4125,N_4097,N_4042);
nor U4126 (N_4126,N_4048,N_4099);
nand U4127 (N_4127,N_4086,N_4033);
nor U4128 (N_4128,N_4060,N_4049);
nand U4129 (N_4129,N_4024,N_4059);
and U4130 (N_4130,N_4075,N_4029);
nand U4131 (N_4131,N_4030,N_4051);
nor U4132 (N_4132,N_4043,N_4066);
or U4133 (N_4133,N_4009,N_4007);
nor U4134 (N_4134,N_4014,N_4044);
or U4135 (N_4135,N_4077,N_4003);
or U4136 (N_4136,N_4045,N_4023);
or U4137 (N_4137,N_4056,N_4073);
or U4138 (N_4138,N_4068,N_4082);
xnor U4139 (N_4139,N_4005,N_4018);
nor U4140 (N_4140,N_4006,N_4071);
or U4141 (N_4141,N_4031,N_4038);
or U4142 (N_4142,N_4064,N_4015);
or U4143 (N_4143,N_4081,N_4047);
nor U4144 (N_4144,N_4090,N_4088);
nor U4145 (N_4145,N_4057,N_4027);
nor U4146 (N_4146,N_4094,N_4065);
or U4147 (N_4147,N_4036,N_4074);
xnor U4148 (N_4148,N_4016,N_4035);
nor U4149 (N_4149,N_4058,N_4021);
nor U4150 (N_4150,N_4018,N_4096);
nand U4151 (N_4151,N_4023,N_4005);
nor U4152 (N_4152,N_4083,N_4097);
or U4153 (N_4153,N_4069,N_4030);
nor U4154 (N_4154,N_4091,N_4083);
or U4155 (N_4155,N_4098,N_4022);
and U4156 (N_4156,N_4059,N_4038);
nor U4157 (N_4157,N_4063,N_4038);
nor U4158 (N_4158,N_4011,N_4025);
or U4159 (N_4159,N_4096,N_4000);
xnor U4160 (N_4160,N_4049,N_4013);
or U4161 (N_4161,N_4026,N_4094);
or U4162 (N_4162,N_4044,N_4049);
and U4163 (N_4163,N_4026,N_4038);
and U4164 (N_4164,N_4036,N_4076);
nand U4165 (N_4165,N_4095,N_4006);
nand U4166 (N_4166,N_4034,N_4062);
nand U4167 (N_4167,N_4086,N_4081);
and U4168 (N_4168,N_4067,N_4057);
or U4169 (N_4169,N_4003,N_4049);
nor U4170 (N_4170,N_4070,N_4098);
nand U4171 (N_4171,N_4008,N_4012);
nor U4172 (N_4172,N_4078,N_4009);
and U4173 (N_4173,N_4055,N_4071);
or U4174 (N_4174,N_4027,N_4036);
or U4175 (N_4175,N_4090,N_4021);
xor U4176 (N_4176,N_4021,N_4000);
nand U4177 (N_4177,N_4067,N_4081);
nor U4178 (N_4178,N_4098,N_4023);
and U4179 (N_4179,N_4096,N_4062);
nand U4180 (N_4180,N_4024,N_4069);
and U4181 (N_4181,N_4082,N_4033);
nand U4182 (N_4182,N_4041,N_4003);
nand U4183 (N_4183,N_4088,N_4085);
or U4184 (N_4184,N_4011,N_4009);
or U4185 (N_4185,N_4046,N_4027);
or U4186 (N_4186,N_4060,N_4016);
nand U4187 (N_4187,N_4030,N_4039);
nor U4188 (N_4188,N_4083,N_4092);
nand U4189 (N_4189,N_4090,N_4081);
or U4190 (N_4190,N_4015,N_4078);
nor U4191 (N_4191,N_4001,N_4079);
and U4192 (N_4192,N_4032,N_4093);
nor U4193 (N_4193,N_4013,N_4067);
and U4194 (N_4194,N_4040,N_4082);
nand U4195 (N_4195,N_4071,N_4012);
xnor U4196 (N_4196,N_4064,N_4018);
and U4197 (N_4197,N_4039,N_4049);
and U4198 (N_4198,N_4049,N_4002);
or U4199 (N_4199,N_4054,N_4060);
or U4200 (N_4200,N_4131,N_4172);
and U4201 (N_4201,N_4135,N_4149);
or U4202 (N_4202,N_4185,N_4164);
and U4203 (N_4203,N_4167,N_4171);
nor U4204 (N_4204,N_4196,N_4190);
and U4205 (N_4205,N_4143,N_4138);
or U4206 (N_4206,N_4125,N_4189);
nand U4207 (N_4207,N_4174,N_4126);
and U4208 (N_4208,N_4106,N_4194);
or U4209 (N_4209,N_4173,N_4184);
or U4210 (N_4210,N_4179,N_4152);
or U4211 (N_4211,N_4137,N_4163);
and U4212 (N_4212,N_4151,N_4108);
nand U4213 (N_4213,N_4105,N_4109);
nor U4214 (N_4214,N_4146,N_4117);
or U4215 (N_4215,N_4100,N_4150);
or U4216 (N_4216,N_4168,N_4161);
and U4217 (N_4217,N_4195,N_4188);
and U4218 (N_4218,N_4160,N_4129);
or U4219 (N_4219,N_4165,N_4155);
nand U4220 (N_4220,N_4133,N_4118);
nor U4221 (N_4221,N_4186,N_4198);
nor U4222 (N_4222,N_4193,N_4158);
and U4223 (N_4223,N_4128,N_4148);
or U4224 (N_4224,N_4191,N_4166);
or U4225 (N_4225,N_4124,N_4182);
nand U4226 (N_4226,N_4136,N_4144);
nand U4227 (N_4227,N_4147,N_4177);
and U4228 (N_4228,N_4122,N_4159);
and U4229 (N_4229,N_4101,N_4175);
or U4230 (N_4230,N_4112,N_4192);
nor U4231 (N_4231,N_4107,N_4176);
and U4232 (N_4232,N_4111,N_4140);
or U4233 (N_4233,N_4114,N_4120);
nand U4234 (N_4234,N_4169,N_4116);
nand U4235 (N_4235,N_4102,N_4145);
nand U4236 (N_4236,N_4141,N_4121);
and U4237 (N_4237,N_4156,N_4199);
nor U4238 (N_4238,N_4197,N_4183);
or U4239 (N_4239,N_4142,N_4110);
and U4240 (N_4240,N_4162,N_4132);
nor U4241 (N_4241,N_4119,N_4139);
or U4242 (N_4242,N_4178,N_4181);
and U4243 (N_4243,N_4130,N_4154);
nand U4244 (N_4244,N_4170,N_4157);
nand U4245 (N_4245,N_4115,N_4127);
and U4246 (N_4246,N_4134,N_4180);
nand U4247 (N_4247,N_4153,N_4123);
nor U4248 (N_4248,N_4103,N_4187);
nor U4249 (N_4249,N_4113,N_4104);
nand U4250 (N_4250,N_4174,N_4185);
nor U4251 (N_4251,N_4118,N_4136);
and U4252 (N_4252,N_4140,N_4174);
nand U4253 (N_4253,N_4160,N_4164);
and U4254 (N_4254,N_4139,N_4183);
nand U4255 (N_4255,N_4186,N_4123);
nor U4256 (N_4256,N_4107,N_4126);
or U4257 (N_4257,N_4122,N_4147);
nand U4258 (N_4258,N_4151,N_4105);
nand U4259 (N_4259,N_4190,N_4156);
or U4260 (N_4260,N_4191,N_4140);
or U4261 (N_4261,N_4195,N_4114);
or U4262 (N_4262,N_4142,N_4179);
nor U4263 (N_4263,N_4183,N_4147);
and U4264 (N_4264,N_4149,N_4116);
and U4265 (N_4265,N_4147,N_4101);
and U4266 (N_4266,N_4136,N_4197);
xnor U4267 (N_4267,N_4120,N_4112);
or U4268 (N_4268,N_4181,N_4110);
nand U4269 (N_4269,N_4129,N_4187);
and U4270 (N_4270,N_4197,N_4146);
and U4271 (N_4271,N_4135,N_4108);
or U4272 (N_4272,N_4173,N_4111);
and U4273 (N_4273,N_4180,N_4185);
or U4274 (N_4274,N_4125,N_4186);
nor U4275 (N_4275,N_4163,N_4185);
or U4276 (N_4276,N_4178,N_4135);
and U4277 (N_4277,N_4101,N_4130);
nand U4278 (N_4278,N_4157,N_4132);
nand U4279 (N_4279,N_4110,N_4180);
nor U4280 (N_4280,N_4158,N_4110);
nand U4281 (N_4281,N_4147,N_4196);
and U4282 (N_4282,N_4136,N_4135);
or U4283 (N_4283,N_4117,N_4116);
and U4284 (N_4284,N_4121,N_4120);
and U4285 (N_4285,N_4128,N_4100);
and U4286 (N_4286,N_4195,N_4125);
and U4287 (N_4287,N_4152,N_4181);
or U4288 (N_4288,N_4193,N_4159);
nand U4289 (N_4289,N_4187,N_4128);
nand U4290 (N_4290,N_4138,N_4105);
and U4291 (N_4291,N_4108,N_4145);
nor U4292 (N_4292,N_4104,N_4116);
nand U4293 (N_4293,N_4171,N_4127);
nor U4294 (N_4294,N_4128,N_4131);
nand U4295 (N_4295,N_4137,N_4161);
nor U4296 (N_4296,N_4187,N_4197);
nand U4297 (N_4297,N_4114,N_4163);
and U4298 (N_4298,N_4184,N_4159);
or U4299 (N_4299,N_4140,N_4152);
and U4300 (N_4300,N_4295,N_4257);
or U4301 (N_4301,N_4247,N_4283);
nor U4302 (N_4302,N_4228,N_4207);
nor U4303 (N_4303,N_4249,N_4255);
and U4304 (N_4304,N_4284,N_4210);
nand U4305 (N_4305,N_4240,N_4237);
nor U4306 (N_4306,N_4222,N_4264);
or U4307 (N_4307,N_4238,N_4245);
or U4308 (N_4308,N_4250,N_4272);
nand U4309 (N_4309,N_4293,N_4205);
xnor U4310 (N_4310,N_4204,N_4267);
or U4311 (N_4311,N_4273,N_4271);
nor U4312 (N_4312,N_4212,N_4282);
nand U4313 (N_4313,N_4269,N_4258);
nor U4314 (N_4314,N_4242,N_4266);
and U4315 (N_4315,N_4221,N_4248);
nor U4316 (N_4316,N_4291,N_4298);
and U4317 (N_4317,N_4294,N_4254);
nor U4318 (N_4318,N_4288,N_4223);
nand U4319 (N_4319,N_4290,N_4251);
and U4320 (N_4320,N_4217,N_4208);
and U4321 (N_4321,N_4202,N_4234);
or U4322 (N_4322,N_4276,N_4286);
nor U4323 (N_4323,N_4292,N_4299);
nand U4324 (N_4324,N_4233,N_4278);
nand U4325 (N_4325,N_4260,N_4243);
or U4326 (N_4326,N_4268,N_4232);
nor U4327 (N_4327,N_4213,N_4200);
nor U4328 (N_4328,N_4256,N_4201);
and U4329 (N_4329,N_4246,N_4227);
nand U4330 (N_4330,N_4224,N_4279);
and U4331 (N_4331,N_4209,N_4218);
nor U4332 (N_4332,N_4253,N_4297);
nor U4333 (N_4333,N_4262,N_4281);
nor U4334 (N_4334,N_4239,N_4275);
xnor U4335 (N_4335,N_4259,N_4280);
and U4336 (N_4336,N_4206,N_4203);
or U4337 (N_4337,N_4215,N_4244);
nand U4338 (N_4338,N_4261,N_4225);
nand U4339 (N_4339,N_4220,N_4231);
nor U4340 (N_4340,N_4219,N_4252);
and U4341 (N_4341,N_4230,N_4287);
or U4342 (N_4342,N_4214,N_4226);
nor U4343 (N_4343,N_4241,N_4236);
or U4344 (N_4344,N_4229,N_4263);
or U4345 (N_4345,N_4270,N_4216);
or U4346 (N_4346,N_4296,N_4211);
or U4347 (N_4347,N_4285,N_4265);
nor U4348 (N_4348,N_4274,N_4277);
nand U4349 (N_4349,N_4289,N_4235);
nand U4350 (N_4350,N_4296,N_4230);
nor U4351 (N_4351,N_4222,N_4291);
nor U4352 (N_4352,N_4216,N_4277);
or U4353 (N_4353,N_4234,N_4248);
nand U4354 (N_4354,N_4220,N_4276);
and U4355 (N_4355,N_4275,N_4270);
nor U4356 (N_4356,N_4245,N_4282);
or U4357 (N_4357,N_4221,N_4290);
and U4358 (N_4358,N_4255,N_4272);
nand U4359 (N_4359,N_4270,N_4247);
nor U4360 (N_4360,N_4242,N_4212);
nor U4361 (N_4361,N_4245,N_4207);
or U4362 (N_4362,N_4298,N_4210);
nor U4363 (N_4363,N_4269,N_4209);
nor U4364 (N_4364,N_4279,N_4241);
or U4365 (N_4365,N_4294,N_4287);
or U4366 (N_4366,N_4278,N_4241);
nand U4367 (N_4367,N_4231,N_4221);
or U4368 (N_4368,N_4233,N_4293);
and U4369 (N_4369,N_4248,N_4250);
nor U4370 (N_4370,N_4212,N_4245);
or U4371 (N_4371,N_4296,N_4201);
nand U4372 (N_4372,N_4269,N_4247);
nand U4373 (N_4373,N_4234,N_4290);
and U4374 (N_4374,N_4274,N_4283);
or U4375 (N_4375,N_4272,N_4249);
nand U4376 (N_4376,N_4237,N_4286);
nor U4377 (N_4377,N_4212,N_4269);
and U4378 (N_4378,N_4288,N_4244);
and U4379 (N_4379,N_4278,N_4279);
nand U4380 (N_4380,N_4255,N_4280);
nor U4381 (N_4381,N_4290,N_4281);
nor U4382 (N_4382,N_4209,N_4228);
nor U4383 (N_4383,N_4230,N_4248);
nand U4384 (N_4384,N_4280,N_4262);
or U4385 (N_4385,N_4293,N_4292);
nor U4386 (N_4386,N_4262,N_4273);
or U4387 (N_4387,N_4281,N_4237);
nand U4388 (N_4388,N_4217,N_4294);
nand U4389 (N_4389,N_4261,N_4203);
xor U4390 (N_4390,N_4258,N_4205);
nor U4391 (N_4391,N_4247,N_4257);
nor U4392 (N_4392,N_4264,N_4263);
nor U4393 (N_4393,N_4266,N_4223);
nand U4394 (N_4394,N_4241,N_4239);
nand U4395 (N_4395,N_4263,N_4251);
or U4396 (N_4396,N_4278,N_4295);
nor U4397 (N_4397,N_4207,N_4263);
nand U4398 (N_4398,N_4227,N_4221);
nand U4399 (N_4399,N_4249,N_4262);
nand U4400 (N_4400,N_4325,N_4331);
nor U4401 (N_4401,N_4391,N_4324);
or U4402 (N_4402,N_4300,N_4375);
xor U4403 (N_4403,N_4339,N_4322);
or U4404 (N_4404,N_4393,N_4328);
nor U4405 (N_4405,N_4388,N_4395);
nor U4406 (N_4406,N_4316,N_4397);
nor U4407 (N_4407,N_4349,N_4350);
nor U4408 (N_4408,N_4353,N_4392);
or U4409 (N_4409,N_4344,N_4332);
nor U4410 (N_4410,N_4351,N_4382);
nor U4411 (N_4411,N_4365,N_4335);
or U4412 (N_4412,N_4304,N_4317);
or U4413 (N_4413,N_4329,N_4334);
or U4414 (N_4414,N_4326,N_4368);
nand U4415 (N_4415,N_4319,N_4379);
nand U4416 (N_4416,N_4312,N_4363);
nor U4417 (N_4417,N_4333,N_4327);
nand U4418 (N_4418,N_4370,N_4345);
nor U4419 (N_4419,N_4341,N_4348);
or U4420 (N_4420,N_4389,N_4394);
or U4421 (N_4421,N_4367,N_4398);
or U4422 (N_4422,N_4381,N_4302);
or U4423 (N_4423,N_4390,N_4354);
nor U4424 (N_4424,N_4366,N_4373);
nand U4425 (N_4425,N_4355,N_4346);
nor U4426 (N_4426,N_4343,N_4337);
nand U4427 (N_4427,N_4323,N_4396);
nor U4428 (N_4428,N_4357,N_4361);
and U4429 (N_4429,N_4386,N_4362);
nor U4430 (N_4430,N_4380,N_4342);
and U4431 (N_4431,N_4315,N_4347);
or U4432 (N_4432,N_4369,N_4378);
nand U4433 (N_4433,N_4320,N_4309);
or U4434 (N_4434,N_4314,N_4359);
or U4435 (N_4435,N_4306,N_4364);
and U4436 (N_4436,N_4303,N_4371);
nor U4437 (N_4437,N_4305,N_4352);
nand U4438 (N_4438,N_4338,N_4356);
or U4439 (N_4439,N_4340,N_4374);
nor U4440 (N_4440,N_4330,N_4377);
nor U4441 (N_4441,N_4307,N_4321);
nor U4442 (N_4442,N_4301,N_4399);
or U4443 (N_4443,N_4313,N_4384);
and U4444 (N_4444,N_4387,N_4360);
or U4445 (N_4445,N_4318,N_4311);
or U4446 (N_4446,N_4372,N_4358);
nand U4447 (N_4447,N_4383,N_4308);
nor U4448 (N_4448,N_4385,N_4336);
or U4449 (N_4449,N_4310,N_4376);
nand U4450 (N_4450,N_4307,N_4325);
nor U4451 (N_4451,N_4381,N_4372);
or U4452 (N_4452,N_4338,N_4350);
nand U4453 (N_4453,N_4367,N_4392);
nor U4454 (N_4454,N_4367,N_4361);
and U4455 (N_4455,N_4376,N_4336);
nand U4456 (N_4456,N_4359,N_4307);
xor U4457 (N_4457,N_4366,N_4313);
or U4458 (N_4458,N_4396,N_4363);
or U4459 (N_4459,N_4336,N_4322);
nand U4460 (N_4460,N_4324,N_4367);
or U4461 (N_4461,N_4369,N_4335);
and U4462 (N_4462,N_4356,N_4377);
nor U4463 (N_4463,N_4346,N_4358);
and U4464 (N_4464,N_4387,N_4311);
nand U4465 (N_4465,N_4334,N_4395);
nor U4466 (N_4466,N_4325,N_4385);
and U4467 (N_4467,N_4342,N_4353);
or U4468 (N_4468,N_4344,N_4327);
and U4469 (N_4469,N_4333,N_4365);
or U4470 (N_4470,N_4373,N_4337);
or U4471 (N_4471,N_4388,N_4381);
nor U4472 (N_4472,N_4326,N_4380);
and U4473 (N_4473,N_4385,N_4361);
nand U4474 (N_4474,N_4379,N_4351);
nand U4475 (N_4475,N_4353,N_4391);
nor U4476 (N_4476,N_4345,N_4337);
nor U4477 (N_4477,N_4322,N_4369);
nor U4478 (N_4478,N_4373,N_4369);
and U4479 (N_4479,N_4308,N_4380);
nand U4480 (N_4480,N_4394,N_4305);
and U4481 (N_4481,N_4379,N_4353);
nand U4482 (N_4482,N_4383,N_4366);
nand U4483 (N_4483,N_4334,N_4390);
and U4484 (N_4484,N_4348,N_4332);
and U4485 (N_4485,N_4329,N_4366);
nor U4486 (N_4486,N_4336,N_4363);
and U4487 (N_4487,N_4355,N_4320);
xor U4488 (N_4488,N_4363,N_4377);
nand U4489 (N_4489,N_4343,N_4357);
nand U4490 (N_4490,N_4332,N_4323);
and U4491 (N_4491,N_4355,N_4308);
nand U4492 (N_4492,N_4348,N_4351);
nor U4493 (N_4493,N_4319,N_4324);
nor U4494 (N_4494,N_4328,N_4301);
and U4495 (N_4495,N_4398,N_4313);
and U4496 (N_4496,N_4319,N_4342);
nand U4497 (N_4497,N_4341,N_4369);
nand U4498 (N_4498,N_4338,N_4370);
and U4499 (N_4499,N_4316,N_4320);
nor U4500 (N_4500,N_4435,N_4483);
nand U4501 (N_4501,N_4448,N_4481);
and U4502 (N_4502,N_4473,N_4421);
or U4503 (N_4503,N_4408,N_4409);
nor U4504 (N_4504,N_4456,N_4469);
or U4505 (N_4505,N_4498,N_4458);
and U4506 (N_4506,N_4437,N_4466);
and U4507 (N_4507,N_4472,N_4474);
and U4508 (N_4508,N_4470,N_4454);
nor U4509 (N_4509,N_4447,N_4410);
nand U4510 (N_4510,N_4403,N_4453);
nand U4511 (N_4511,N_4427,N_4416);
nor U4512 (N_4512,N_4432,N_4485);
nand U4513 (N_4513,N_4486,N_4495);
and U4514 (N_4514,N_4450,N_4428);
nand U4515 (N_4515,N_4401,N_4440);
nand U4516 (N_4516,N_4436,N_4444);
nand U4517 (N_4517,N_4417,N_4487);
nor U4518 (N_4518,N_4484,N_4492);
nand U4519 (N_4519,N_4455,N_4406);
or U4520 (N_4520,N_4405,N_4461);
and U4521 (N_4521,N_4497,N_4434);
and U4522 (N_4522,N_4419,N_4496);
and U4523 (N_4523,N_4429,N_4423);
nand U4524 (N_4524,N_4442,N_4446);
or U4525 (N_4525,N_4490,N_4424);
and U4526 (N_4526,N_4477,N_4452);
or U4527 (N_4527,N_4499,N_4489);
or U4528 (N_4528,N_4411,N_4475);
xor U4529 (N_4529,N_4459,N_4438);
nand U4530 (N_4530,N_4413,N_4482);
nand U4531 (N_4531,N_4460,N_4478);
nor U4532 (N_4532,N_4493,N_4445);
nor U4533 (N_4533,N_4404,N_4462);
and U4534 (N_4534,N_4491,N_4465);
nor U4535 (N_4535,N_4441,N_4439);
or U4536 (N_4536,N_4443,N_4418);
nand U4537 (N_4537,N_4480,N_4494);
nor U4538 (N_4538,N_4402,N_4479);
and U4539 (N_4539,N_4464,N_4420);
nor U4540 (N_4540,N_4407,N_4471);
and U4541 (N_4541,N_4430,N_4431);
nor U4542 (N_4542,N_4457,N_4426);
nor U4543 (N_4543,N_4467,N_4415);
or U4544 (N_4544,N_4414,N_4468);
nand U4545 (N_4545,N_4400,N_4412);
or U4546 (N_4546,N_4463,N_4476);
nor U4547 (N_4547,N_4488,N_4422);
and U4548 (N_4548,N_4451,N_4425);
nor U4549 (N_4549,N_4449,N_4433);
or U4550 (N_4550,N_4456,N_4422);
and U4551 (N_4551,N_4480,N_4417);
nand U4552 (N_4552,N_4411,N_4470);
nor U4553 (N_4553,N_4418,N_4471);
and U4554 (N_4554,N_4423,N_4443);
or U4555 (N_4555,N_4471,N_4416);
or U4556 (N_4556,N_4462,N_4400);
and U4557 (N_4557,N_4471,N_4408);
nand U4558 (N_4558,N_4404,N_4454);
xnor U4559 (N_4559,N_4474,N_4401);
and U4560 (N_4560,N_4484,N_4445);
and U4561 (N_4561,N_4404,N_4471);
nor U4562 (N_4562,N_4425,N_4435);
nand U4563 (N_4563,N_4403,N_4496);
nor U4564 (N_4564,N_4429,N_4437);
nor U4565 (N_4565,N_4449,N_4455);
nor U4566 (N_4566,N_4428,N_4456);
or U4567 (N_4567,N_4428,N_4449);
nand U4568 (N_4568,N_4452,N_4435);
nand U4569 (N_4569,N_4415,N_4455);
and U4570 (N_4570,N_4413,N_4445);
and U4571 (N_4571,N_4481,N_4438);
nor U4572 (N_4572,N_4427,N_4418);
and U4573 (N_4573,N_4400,N_4461);
and U4574 (N_4574,N_4413,N_4406);
nand U4575 (N_4575,N_4422,N_4458);
nor U4576 (N_4576,N_4442,N_4406);
nor U4577 (N_4577,N_4467,N_4461);
nor U4578 (N_4578,N_4491,N_4432);
or U4579 (N_4579,N_4480,N_4428);
and U4580 (N_4580,N_4422,N_4408);
and U4581 (N_4581,N_4463,N_4490);
nor U4582 (N_4582,N_4416,N_4419);
or U4583 (N_4583,N_4475,N_4403);
or U4584 (N_4584,N_4424,N_4444);
and U4585 (N_4585,N_4481,N_4425);
and U4586 (N_4586,N_4433,N_4413);
nand U4587 (N_4587,N_4428,N_4404);
and U4588 (N_4588,N_4474,N_4453);
or U4589 (N_4589,N_4429,N_4489);
or U4590 (N_4590,N_4456,N_4444);
nand U4591 (N_4591,N_4440,N_4456);
nand U4592 (N_4592,N_4456,N_4496);
and U4593 (N_4593,N_4430,N_4453);
nor U4594 (N_4594,N_4424,N_4461);
and U4595 (N_4595,N_4417,N_4486);
and U4596 (N_4596,N_4444,N_4405);
nand U4597 (N_4597,N_4498,N_4453);
nor U4598 (N_4598,N_4457,N_4498);
or U4599 (N_4599,N_4414,N_4449);
xnor U4600 (N_4600,N_4556,N_4542);
or U4601 (N_4601,N_4586,N_4538);
nor U4602 (N_4602,N_4534,N_4515);
nor U4603 (N_4603,N_4595,N_4593);
nand U4604 (N_4604,N_4544,N_4550);
nor U4605 (N_4605,N_4577,N_4510);
nor U4606 (N_4606,N_4511,N_4520);
or U4607 (N_4607,N_4565,N_4569);
or U4608 (N_4608,N_4561,N_4526);
xor U4609 (N_4609,N_4500,N_4588);
nor U4610 (N_4610,N_4591,N_4560);
and U4611 (N_4611,N_4555,N_4553);
or U4612 (N_4612,N_4585,N_4572);
nor U4613 (N_4613,N_4571,N_4531);
nor U4614 (N_4614,N_4547,N_4583);
and U4615 (N_4615,N_4541,N_4558);
and U4616 (N_4616,N_4570,N_4533);
and U4617 (N_4617,N_4513,N_4543);
nor U4618 (N_4618,N_4527,N_4557);
nor U4619 (N_4619,N_4517,N_4530);
or U4620 (N_4620,N_4532,N_4578);
nor U4621 (N_4621,N_4502,N_4582);
or U4622 (N_4622,N_4599,N_4574);
or U4623 (N_4623,N_4575,N_4594);
nand U4624 (N_4624,N_4592,N_4567);
and U4625 (N_4625,N_4576,N_4554);
and U4626 (N_4626,N_4564,N_4546);
or U4627 (N_4627,N_4590,N_4524);
and U4628 (N_4628,N_4516,N_4584);
nand U4629 (N_4629,N_4508,N_4589);
or U4630 (N_4630,N_4539,N_4514);
nand U4631 (N_4631,N_4537,N_4580);
nor U4632 (N_4632,N_4579,N_4507);
nand U4633 (N_4633,N_4545,N_4598);
nor U4634 (N_4634,N_4559,N_4529);
nor U4635 (N_4635,N_4522,N_4512);
nand U4636 (N_4636,N_4505,N_4521);
or U4637 (N_4637,N_4503,N_4536);
nor U4638 (N_4638,N_4519,N_4581);
nor U4639 (N_4639,N_4597,N_4549);
nand U4640 (N_4640,N_4596,N_4562);
nand U4641 (N_4641,N_4509,N_4540);
nor U4642 (N_4642,N_4587,N_4573);
nand U4643 (N_4643,N_4525,N_4551);
nand U4644 (N_4644,N_4566,N_4563);
nand U4645 (N_4645,N_4528,N_4548);
or U4646 (N_4646,N_4523,N_4568);
or U4647 (N_4647,N_4552,N_4518);
nand U4648 (N_4648,N_4506,N_4504);
nor U4649 (N_4649,N_4535,N_4501);
and U4650 (N_4650,N_4554,N_4502);
xor U4651 (N_4651,N_4599,N_4552);
and U4652 (N_4652,N_4541,N_4585);
xnor U4653 (N_4653,N_4586,N_4565);
nor U4654 (N_4654,N_4581,N_4599);
nand U4655 (N_4655,N_4553,N_4532);
nand U4656 (N_4656,N_4549,N_4581);
or U4657 (N_4657,N_4545,N_4558);
and U4658 (N_4658,N_4583,N_4593);
or U4659 (N_4659,N_4578,N_4540);
nand U4660 (N_4660,N_4509,N_4531);
or U4661 (N_4661,N_4561,N_4538);
nor U4662 (N_4662,N_4527,N_4576);
nor U4663 (N_4663,N_4508,N_4599);
xnor U4664 (N_4664,N_4558,N_4554);
and U4665 (N_4665,N_4597,N_4551);
nand U4666 (N_4666,N_4584,N_4596);
or U4667 (N_4667,N_4554,N_4508);
nor U4668 (N_4668,N_4501,N_4597);
xnor U4669 (N_4669,N_4564,N_4531);
nand U4670 (N_4670,N_4530,N_4588);
and U4671 (N_4671,N_4557,N_4551);
nor U4672 (N_4672,N_4551,N_4549);
and U4673 (N_4673,N_4519,N_4551);
nor U4674 (N_4674,N_4564,N_4589);
nand U4675 (N_4675,N_4575,N_4553);
nand U4676 (N_4676,N_4540,N_4594);
nor U4677 (N_4677,N_4594,N_4572);
nand U4678 (N_4678,N_4593,N_4569);
or U4679 (N_4679,N_4533,N_4535);
nor U4680 (N_4680,N_4581,N_4569);
nand U4681 (N_4681,N_4537,N_4593);
nand U4682 (N_4682,N_4553,N_4581);
nand U4683 (N_4683,N_4570,N_4520);
nand U4684 (N_4684,N_4525,N_4544);
and U4685 (N_4685,N_4552,N_4564);
nand U4686 (N_4686,N_4569,N_4516);
nor U4687 (N_4687,N_4519,N_4513);
nand U4688 (N_4688,N_4508,N_4538);
nor U4689 (N_4689,N_4583,N_4511);
and U4690 (N_4690,N_4526,N_4535);
and U4691 (N_4691,N_4599,N_4515);
or U4692 (N_4692,N_4506,N_4583);
nand U4693 (N_4693,N_4553,N_4501);
or U4694 (N_4694,N_4571,N_4533);
or U4695 (N_4695,N_4529,N_4582);
or U4696 (N_4696,N_4502,N_4547);
and U4697 (N_4697,N_4582,N_4584);
nor U4698 (N_4698,N_4526,N_4595);
nor U4699 (N_4699,N_4564,N_4576);
nand U4700 (N_4700,N_4692,N_4662);
nor U4701 (N_4701,N_4643,N_4657);
and U4702 (N_4702,N_4623,N_4680);
or U4703 (N_4703,N_4619,N_4606);
nor U4704 (N_4704,N_4620,N_4650);
nor U4705 (N_4705,N_4676,N_4649);
or U4706 (N_4706,N_4616,N_4603);
or U4707 (N_4707,N_4673,N_4677);
nand U4708 (N_4708,N_4655,N_4640);
xnor U4709 (N_4709,N_4681,N_4613);
and U4710 (N_4710,N_4685,N_4667);
nor U4711 (N_4711,N_4663,N_4670);
and U4712 (N_4712,N_4630,N_4696);
xor U4713 (N_4713,N_4647,N_4656);
nor U4714 (N_4714,N_4629,N_4635);
or U4715 (N_4715,N_4633,N_4689);
or U4716 (N_4716,N_4637,N_4632);
nand U4717 (N_4717,N_4644,N_4664);
and U4718 (N_4718,N_4634,N_4672);
nand U4719 (N_4719,N_4698,N_4611);
and U4720 (N_4720,N_4694,N_4608);
nand U4721 (N_4721,N_4695,N_4674);
or U4722 (N_4722,N_4665,N_4600);
nor U4723 (N_4723,N_4617,N_4671);
or U4724 (N_4724,N_4621,N_4638);
nand U4725 (N_4725,N_4651,N_4625);
nand U4726 (N_4726,N_4624,N_4602);
and U4727 (N_4727,N_4699,N_4652);
nor U4728 (N_4728,N_4627,N_4607);
and U4729 (N_4729,N_4614,N_4683);
nor U4730 (N_4730,N_4601,N_4605);
and U4731 (N_4731,N_4684,N_4669);
and U4732 (N_4732,N_4691,N_4639);
nor U4733 (N_4733,N_4615,N_4618);
and U4734 (N_4734,N_4641,N_4675);
nor U4735 (N_4735,N_4661,N_4686);
or U4736 (N_4736,N_4660,N_4679);
nor U4737 (N_4737,N_4688,N_4612);
or U4738 (N_4738,N_4609,N_4653);
nand U4739 (N_4739,N_4666,N_4636);
xor U4740 (N_4740,N_4658,N_4622);
nand U4741 (N_4741,N_4648,N_4693);
nand U4742 (N_4742,N_4659,N_4646);
nand U4743 (N_4743,N_4654,N_4631);
and U4744 (N_4744,N_4687,N_4645);
nand U4745 (N_4745,N_4682,N_4642);
nor U4746 (N_4746,N_4697,N_4668);
and U4747 (N_4747,N_4690,N_4604);
nand U4748 (N_4748,N_4628,N_4610);
nand U4749 (N_4749,N_4678,N_4626);
xor U4750 (N_4750,N_4640,N_4610);
nor U4751 (N_4751,N_4664,N_4620);
nor U4752 (N_4752,N_4627,N_4600);
nor U4753 (N_4753,N_4663,N_4675);
nand U4754 (N_4754,N_4643,N_4674);
nand U4755 (N_4755,N_4625,N_4692);
nand U4756 (N_4756,N_4604,N_4642);
or U4757 (N_4757,N_4605,N_4619);
or U4758 (N_4758,N_4662,N_4682);
nand U4759 (N_4759,N_4611,N_4634);
nor U4760 (N_4760,N_4644,N_4636);
and U4761 (N_4761,N_4669,N_4624);
or U4762 (N_4762,N_4634,N_4676);
or U4763 (N_4763,N_4675,N_4633);
xnor U4764 (N_4764,N_4614,N_4664);
nor U4765 (N_4765,N_4693,N_4606);
nor U4766 (N_4766,N_4609,N_4612);
and U4767 (N_4767,N_4686,N_4642);
or U4768 (N_4768,N_4683,N_4660);
xnor U4769 (N_4769,N_4656,N_4661);
and U4770 (N_4770,N_4624,N_4694);
nand U4771 (N_4771,N_4602,N_4629);
and U4772 (N_4772,N_4608,N_4615);
and U4773 (N_4773,N_4638,N_4628);
and U4774 (N_4774,N_4641,N_4651);
nand U4775 (N_4775,N_4653,N_4680);
or U4776 (N_4776,N_4612,N_4629);
nand U4777 (N_4777,N_4671,N_4684);
nor U4778 (N_4778,N_4686,N_4637);
and U4779 (N_4779,N_4688,N_4646);
or U4780 (N_4780,N_4672,N_4620);
and U4781 (N_4781,N_4643,N_4638);
or U4782 (N_4782,N_4668,N_4642);
or U4783 (N_4783,N_4650,N_4652);
and U4784 (N_4784,N_4670,N_4626);
or U4785 (N_4785,N_4618,N_4621);
nand U4786 (N_4786,N_4624,N_4610);
and U4787 (N_4787,N_4691,N_4645);
nor U4788 (N_4788,N_4695,N_4632);
xnor U4789 (N_4789,N_4689,N_4665);
nand U4790 (N_4790,N_4691,N_4649);
xor U4791 (N_4791,N_4641,N_4611);
or U4792 (N_4792,N_4687,N_4686);
nor U4793 (N_4793,N_4689,N_4675);
nor U4794 (N_4794,N_4634,N_4600);
nor U4795 (N_4795,N_4621,N_4609);
nand U4796 (N_4796,N_4672,N_4628);
or U4797 (N_4797,N_4663,N_4607);
nand U4798 (N_4798,N_4665,N_4671);
nand U4799 (N_4799,N_4656,N_4673);
nor U4800 (N_4800,N_4749,N_4795);
nor U4801 (N_4801,N_4793,N_4780);
xor U4802 (N_4802,N_4755,N_4765);
nor U4803 (N_4803,N_4792,N_4783);
nor U4804 (N_4804,N_4727,N_4701);
nor U4805 (N_4805,N_4770,N_4771);
and U4806 (N_4806,N_4725,N_4743);
and U4807 (N_4807,N_4744,N_4742);
and U4808 (N_4808,N_4787,N_4710);
or U4809 (N_4809,N_4704,N_4796);
nor U4810 (N_4810,N_4791,N_4745);
and U4811 (N_4811,N_4726,N_4768);
or U4812 (N_4812,N_4773,N_4733);
nand U4813 (N_4813,N_4724,N_4775);
and U4814 (N_4814,N_4707,N_4794);
nor U4815 (N_4815,N_4736,N_4746);
and U4816 (N_4816,N_4790,N_4714);
or U4817 (N_4817,N_4760,N_4720);
nand U4818 (N_4818,N_4785,N_4767);
nor U4819 (N_4819,N_4731,N_4799);
or U4820 (N_4820,N_4750,N_4729);
and U4821 (N_4821,N_4757,N_4779);
and U4822 (N_4822,N_4711,N_4772);
nand U4823 (N_4823,N_4761,N_4763);
or U4824 (N_4824,N_4748,N_4712);
nor U4825 (N_4825,N_4735,N_4782);
nor U4826 (N_4826,N_4797,N_4713);
nand U4827 (N_4827,N_4719,N_4778);
and U4828 (N_4828,N_4769,N_4798);
and U4829 (N_4829,N_4741,N_4738);
or U4830 (N_4830,N_4789,N_4784);
nand U4831 (N_4831,N_4753,N_4730);
or U4832 (N_4832,N_4766,N_4776);
nand U4833 (N_4833,N_4723,N_4702);
and U4834 (N_4834,N_4747,N_4722);
or U4835 (N_4835,N_4703,N_4751);
and U4836 (N_4836,N_4764,N_4721);
and U4837 (N_4837,N_4705,N_4756);
and U4838 (N_4838,N_4781,N_4728);
nor U4839 (N_4839,N_4759,N_4709);
and U4840 (N_4840,N_4739,N_4754);
and U4841 (N_4841,N_4752,N_4758);
nor U4842 (N_4842,N_4715,N_4716);
nand U4843 (N_4843,N_4717,N_4786);
nor U4844 (N_4844,N_4708,N_4732);
nand U4845 (N_4845,N_4706,N_4777);
xnor U4846 (N_4846,N_4788,N_4740);
and U4847 (N_4847,N_4774,N_4718);
or U4848 (N_4848,N_4762,N_4734);
nor U4849 (N_4849,N_4737,N_4700);
nand U4850 (N_4850,N_4799,N_4744);
or U4851 (N_4851,N_4731,N_4775);
nor U4852 (N_4852,N_4721,N_4775);
or U4853 (N_4853,N_4782,N_4755);
or U4854 (N_4854,N_4757,N_4710);
nor U4855 (N_4855,N_4712,N_4786);
and U4856 (N_4856,N_4744,N_4746);
nand U4857 (N_4857,N_4714,N_4737);
nor U4858 (N_4858,N_4746,N_4763);
or U4859 (N_4859,N_4766,N_4762);
or U4860 (N_4860,N_4795,N_4745);
nand U4861 (N_4861,N_4703,N_4719);
and U4862 (N_4862,N_4710,N_4716);
and U4863 (N_4863,N_4796,N_4719);
nand U4864 (N_4864,N_4774,N_4731);
nand U4865 (N_4865,N_4703,N_4764);
or U4866 (N_4866,N_4780,N_4744);
or U4867 (N_4867,N_4707,N_4749);
and U4868 (N_4868,N_4706,N_4748);
nand U4869 (N_4869,N_4750,N_4703);
nor U4870 (N_4870,N_4731,N_4752);
and U4871 (N_4871,N_4761,N_4744);
nor U4872 (N_4872,N_4756,N_4766);
nand U4873 (N_4873,N_4760,N_4715);
nor U4874 (N_4874,N_4753,N_4704);
or U4875 (N_4875,N_4785,N_4774);
and U4876 (N_4876,N_4762,N_4701);
nor U4877 (N_4877,N_4788,N_4795);
or U4878 (N_4878,N_4733,N_4780);
nand U4879 (N_4879,N_4722,N_4758);
and U4880 (N_4880,N_4741,N_4716);
xor U4881 (N_4881,N_4718,N_4721);
and U4882 (N_4882,N_4759,N_4765);
nor U4883 (N_4883,N_4741,N_4763);
nor U4884 (N_4884,N_4706,N_4702);
xor U4885 (N_4885,N_4744,N_4723);
and U4886 (N_4886,N_4783,N_4733);
nor U4887 (N_4887,N_4718,N_4784);
nand U4888 (N_4888,N_4741,N_4773);
or U4889 (N_4889,N_4706,N_4710);
and U4890 (N_4890,N_4756,N_4787);
or U4891 (N_4891,N_4731,N_4704);
nor U4892 (N_4892,N_4762,N_4732);
or U4893 (N_4893,N_4705,N_4760);
or U4894 (N_4894,N_4704,N_4735);
or U4895 (N_4895,N_4778,N_4717);
nand U4896 (N_4896,N_4731,N_4746);
nand U4897 (N_4897,N_4775,N_4766);
or U4898 (N_4898,N_4789,N_4783);
nor U4899 (N_4899,N_4790,N_4742);
xor U4900 (N_4900,N_4838,N_4820);
or U4901 (N_4901,N_4859,N_4814);
nand U4902 (N_4902,N_4860,N_4898);
or U4903 (N_4903,N_4800,N_4874);
nand U4904 (N_4904,N_4828,N_4849);
nand U4905 (N_4905,N_4845,N_4878);
nor U4906 (N_4906,N_4851,N_4804);
or U4907 (N_4907,N_4810,N_4819);
and U4908 (N_4908,N_4888,N_4867);
or U4909 (N_4909,N_4825,N_4862);
nand U4910 (N_4910,N_4872,N_4895);
nand U4911 (N_4911,N_4890,N_4821);
and U4912 (N_4912,N_4873,N_4892);
and U4913 (N_4913,N_4831,N_4842);
nand U4914 (N_4914,N_4864,N_4854);
and U4915 (N_4915,N_4894,N_4827);
nand U4916 (N_4916,N_4824,N_4869);
or U4917 (N_4917,N_4808,N_4879);
nand U4918 (N_4918,N_4801,N_4863);
and U4919 (N_4919,N_4812,N_4850);
and U4920 (N_4920,N_4881,N_4880);
or U4921 (N_4921,N_4885,N_4858);
nand U4922 (N_4922,N_4855,N_4818);
nand U4923 (N_4923,N_4847,N_4848);
nor U4924 (N_4924,N_4852,N_4805);
nand U4925 (N_4925,N_4891,N_4832);
nor U4926 (N_4926,N_4856,N_4829);
nand U4927 (N_4927,N_4837,N_4840);
nor U4928 (N_4928,N_4817,N_4877);
and U4929 (N_4929,N_4861,N_4834);
nand U4930 (N_4930,N_4802,N_4826);
nand U4931 (N_4931,N_4870,N_4866);
nand U4932 (N_4932,N_4833,N_4897);
nand U4933 (N_4933,N_4807,N_4813);
nand U4934 (N_4934,N_4803,N_4889);
and U4935 (N_4935,N_4811,N_4844);
or U4936 (N_4936,N_4835,N_4887);
nor U4937 (N_4937,N_4843,N_4865);
nand U4938 (N_4938,N_4883,N_4899);
nor U4939 (N_4939,N_4857,N_4853);
nand U4940 (N_4940,N_4815,N_4875);
and U4941 (N_4941,N_4823,N_4896);
or U4942 (N_4942,N_4806,N_4830);
nand U4943 (N_4943,N_4876,N_4836);
or U4944 (N_4944,N_4884,N_4846);
or U4945 (N_4945,N_4839,N_4886);
or U4946 (N_4946,N_4871,N_4893);
and U4947 (N_4947,N_4822,N_4841);
or U4948 (N_4948,N_4816,N_4868);
and U4949 (N_4949,N_4882,N_4809);
nor U4950 (N_4950,N_4870,N_4822);
or U4951 (N_4951,N_4856,N_4889);
and U4952 (N_4952,N_4891,N_4813);
or U4953 (N_4953,N_4871,N_4878);
nand U4954 (N_4954,N_4862,N_4800);
nor U4955 (N_4955,N_4847,N_4862);
nor U4956 (N_4956,N_4861,N_4895);
nor U4957 (N_4957,N_4826,N_4822);
and U4958 (N_4958,N_4875,N_4802);
and U4959 (N_4959,N_4858,N_4842);
and U4960 (N_4960,N_4884,N_4856);
and U4961 (N_4961,N_4812,N_4823);
nor U4962 (N_4962,N_4843,N_4814);
nand U4963 (N_4963,N_4896,N_4872);
nand U4964 (N_4964,N_4849,N_4836);
nand U4965 (N_4965,N_4857,N_4835);
or U4966 (N_4966,N_4867,N_4892);
nor U4967 (N_4967,N_4833,N_4878);
nor U4968 (N_4968,N_4890,N_4859);
nor U4969 (N_4969,N_4890,N_4852);
nor U4970 (N_4970,N_4885,N_4829);
and U4971 (N_4971,N_4811,N_4809);
nor U4972 (N_4972,N_4843,N_4827);
nor U4973 (N_4973,N_4860,N_4817);
nand U4974 (N_4974,N_4864,N_4881);
nand U4975 (N_4975,N_4823,N_4828);
or U4976 (N_4976,N_4838,N_4811);
or U4977 (N_4977,N_4810,N_4876);
and U4978 (N_4978,N_4840,N_4896);
and U4979 (N_4979,N_4842,N_4814);
and U4980 (N_4980,N_4869,N_4851);
or U4981 (N_4981,N_4816,N_4846);
and U4982 (N_4982,N_4861,N_4856);
nand U4983 (N_4983,N_4893,N_4854);
nand U4984 (N_4984,N_4847,N_4885);
nand U4985 (N_4985,N_4824,N_4871);
nand U4986 (N_4986,N_4897,N_4808);
nand U4987 (N_4987,N_4882,N_4827);
or U4988 (N_4988,N_4888,N_4810);
nand U4989 (N_4989,N_4892,N_4875);
and U4990 (N_4990,N_4899,N_4888);
nor U4991 (N_4991,N_4845,N_4814);
nor U4992 (N_4992,N_4866,N_4830);
or U4993 (N_4993,N_4870,N_4886);
nand U4994 (N_4994,N_4845,N_4890);
nand U4995 (N_4995,N_4807,N_4892);
nand U4996 (N_4996,N_4897,N_4848);
or U4997 (N_4997,N_4836,N_4812);
or U4998 (N_4998,N_4807,N_4881);
nor U4999 (N_4999,N_4843,N_4846);
and U5000 (N_5000,N_4965,N_4903);
or U5001 (N_5001,N_4974,N_4966);
nor U5002 (N_5002,N_4917,N_4958);
or U5003 (N_5003,N_4907,N_4915);
or U5004 (N_5004,N_4984,N_4948);
xor U5005 (N_5005,N_4987,N_4947);
nor U5006 (N_5006,N_4921,N_4976);
nand U5007 (N_5007,N_4905,N_4960);
nor U5008 (N_5008,N_4970,N_4981);
or U5009 (N_5009,N_4969,N_4982);
or U5010 (N_5010,N_4953,N_4929);
and U5011 (N_5011,N_4962,N_4926);
or U5012 (N_5012,N_4942,N_4931);
and U5013 (N_5013,N_4983,N_4968);
or U5014 (N_5014,N_4964,N_4944);
nor U5015 (N_5015,N_4913,N_4945);
or U5016 (N_5016,N_4990,N_4918);
nand U5017 (N_5017,N_4975,N_4930);
and U5018 (N_5018,N_4995,N_4928);
nor U5019 (N_5019,N_4985,N_4955);
or U5020 (N_5020,N_4941,N_4925);
and U5021 (N_5021,N_4910,N_4937);
and U5022 (N_5022,N_4933,N_4943);
nor U5023 (N_5023,N_4906,N_4911);
nand U5024 (N_5024,N_4932,N_4939);
nor U5025 (N_5025,N_4998,N_4992);
nand U5026 (N_5026,N_4936,N_4935);
or U5027 (N_5027,N_4954,N_4951);
or U5028 (N_5028,N_4999,N_4963);
or U5029 (N_5029,N_4980,N_4919);
nand U5030 (N_5030,N_4949,N_4934);
nor U5031 (N_5031,N_4916,N_4946);
or U5032 (N_5032,N_4956,N_4938);
and U5033 (N_5033,N_4994,N_4904);
nor U5034 (N_5034,N_4988,N_4961);
nor U5035 (N_5035,N_4940,N_4973);
nand U5036 (N_5036,N_4989,N_4952);
nor U5037 (N_5037,N_4971,N_4993);
nor U5038 (N_5038,N_4986,N_4996);
nor U5039 (N_5039,N_4959,N_4977);
and U5040 (N_5040,N_4909,N_4914);
and U5041 (N_5041,N_4902,N_4922);
nor U5042 (N_5042,N_4950,N_4908);
and U5043 (N_5043,N_4923,N_4967);
nor U5044 (N_5044,N_4972,N_4900);
and U5045 (N_5045,N_4997,N_4978);
and U5046 (N_5046,N_4924,N_4957);
nand U5047 (N_5047,N_4927,N_4920);
or U5048 (N_5048,N_4991,N_4901);
nand U5049 (N_5049,N_4912,N_4979);
nand U5050 (N_5050,N_4975,N_4950);
nor U5051 (N_5051,N_4921,N_4907);
or U5052 (N_5052,N_4971,N_4989);
and U5053 (N_5053,N_4915,N_4901);
or U5054 (N_5054,N_4955,N_4960);
or U5055 (N_5055,N_4933,N_4927);
and U5056 (N_5056,N_4970,N_4925);
or U5057 (N_5057,N_4934,N_4948);
and U5058 (N_5058,N_4992,N_4964);
or U5059 (N_5059,N_4952,N_4929);
and U5060 (N_5060,N_4986,N_4987);
nor U5061 (N_5061,N_4939,N_4945);
or U5062 (N_5062,N_4950,N_4907);
and U5063 (N_5063,N_4964,N_4995);
or U5064 (N_5064,N_4987,N_4914);
and U5065 (N_5065,N_4911,N_4968);
or U5066 (N_5066,N_4905,N_4989);
nand U5067 (N_5067,N_4910,N_4981);
nand U5068 (N_5068,N_4993,N_4913);
nor U5069 (N_5069,N_4953,N_4907);
or U5070 (N_5070,N_4964,N_4913);
nor U5071 (N_5071,N_4907,N_4924);
nor U5072 (N_5072,N_4929,N_4977);
nor U5073 (N_5073,N_4931,N_4935);
nand U5074 (N_5074,N_4935,N_4947);
xor U5075 (N_5075,N_4910,N_4952);
and U5076 (N_5076,N_4932,N_4924);
nor U5077 (N_5077,N_4988,N_4903);
nor U5078 (N_5078,N_4959,N_4908);
and U5079 (N_5079,N_4991,N_4998);
and U5080 (N_5080,N_4938,N_4984);
nor U5081 (N_5081,N_4902,N_4913);
and U5082 (N_5082,N_4957,N_4975);
nand U5083 (N_5083,N_4970,N_4961);
nand U5084 (N_5084,N_4906,N_4925);
nand U5085 (N_5085,N_4937,N_4954);
nor U5086 (N_5086,N_4932,N_4959);
or U5087 (N_5087,N_4963,N_4978);
nor U5088 (N_5088,N_4973,N_4923);
and U5089 (N_5089,N_4914,N_4946);
and U5090 (N_5090,N_4956,N_4950);
or U5091 (N_5091,N_4959,N_4998);
nand U5092 (N_5092,N_4932,N_4900);
nor U5093 (N_5093,N_4946,N_4966);
nand U5094 (N_5094,N_4952,N_4950);
or U5095 (N_5095,N_4982,N_4987);
nand U5096 (N_5096,N_4943,N_4911);
and U5097 (N_5097,N_4973,N_4920);
nor U5098 (N_5098,N_4905,N_4949);
nor U5099 (N_5099,N_4924,N_4992);
xnor U5100 (N_5100,N_5005,N_5032);
xnor U5101 (N_5101,N_5079,N_5091);
and U5102 (N_5102,N_5012,N_5088);
or U5103 (N_5103,N_5014,N_5011);
nor U5104 (N_5104,N_5061,N_5013);
nand U5105 (N_5105,N_5070,N_5053);
or U5106 (N_5106,N_5026,N_5065);
or U5107 (N_5107,N_5010,N_5009);
nor U5108 (N_5108,N_5063,N_5072);
or U5109 (N_5109,N_5069,N_5086);
or U5110 (N_5110,N_5073,N_5033);
and U5111 (N_5111,N_5007,N_5056);
nand U5112 (N_5112,N_5003,N_5092);
or U5113 (N_5113,N_5097,N_5001);
or U5114 (N_5114,N_5058,N_5047);
xnor U5115 (N_5115,N_5084,N_5085);
nand U5116 (N_5116,N_5059,N_5043);
xor U5117 (N_5117,N_5002,N_5095);
and U5118 (N_5118,N_5046,N_5045);
nand U5119 (N_5119,N_5096,N_5048);
nor U5120 (N_5120,N_5075,N_5080);
and U5121 (N_5121,N_5074,N_5083);
and U5122 (N_5122,N_5021,N_5000);
and U5123 (N_5123,N_5022,N_5094);
nand U5124 (N_5124,N_5015,N_5039);
nor U5125 (N_5125,N_5028,N_5041);
or U5126 (N_5126,N_5030,N_5023);
nand U5127 (N_5127,N_5035,N_5060);
nor U5128 (N_5128,N_5027,N_5018);
nor U5129 (N_5129,N_5025,N_5093);
nor U5130 (N_5130,N_5090,N_5036);
or U5131 (N_5131,N_5037,N_5038);
and U5132 (N_5132,N_5019,N_5087);
nor U5133 (N_5133,N_5020,N_5078);
nand U5134 (N_5134,N_5024,N_5052);
nand U5135 (N_5135,N_5004,N_5099);
and U5136 (N_5136,N_5049,N_5071);
or U5137 (N_5137,N_5068,N_5006);
nand U5138 (N_5138,N_5057,N_5066);
or U5139 (N_5139,N_5082,N_5098);
or U5140 (N_5140,N_5044,N_5076);
and U5141 (N_5141,N_5029,N_5081);
or U5142 (N_5142,N_5089,N_5042);
xnor U5143 (N_5143,N_5064,N_5034);
nand U5144 (N_5144,N_5031,N_5067);
nand U5145 (N_5145,N_5050,N_5055);
nor U5146 (N_5146,N_5054,N_5051);
or U5147 (N_5147,N_5062,N_5008);
nand U5148 (N_5148,N_5077,N_5040);
or U5149 (N_5149,N_5016,N_5017);
or U5150 (N_5150,N_5071,N_5013);
nand U5151 (N_5151,N_5010,N_5040);
or U5152 (N_5152,N_5088,N_5062);
and U5153 (N_5153,N_5042,N_5065);
nor U5154 (N_5154,N_5030,N_5048);
or U5155 (N_5155,N_5082,N_5083);
nand U5156 (N_5156,N_5022,N_5059);
nand U5157 (N_5157,N_5038,N_5086);
nand U5158 (N_5158,N_5061,N_5039);
or U5159 (N_5159,N_5031,N_5066);
nor U5160 (N_5160,N_5074,N_5014);
nor U5161 (N_5161,N_5034,N_5051);
nor U5162 (N_5162,N_5016,N_5033);
and U5163 (N_5163,N_5070,N_5081);
nand U5164 (N_5164,N_5036,N_5076);
nor U5165 (N_5165,N_5012,N_5044);
nand U5166 (N_5166,N_5062,N_5051);
or U5167 (N_5167,N_5027,N_5067);
and U5168 (N_5168,N_5046,N_5071);
and U5169 (N_5169,N_5009,N_5066);
nand U5170 (N_5170,N_5019,N_5086);
nor U5171 (N_5171,N_5008,N_5093);
nand U5172 (N_5172,N_5071,N_5010);
or U5173 (N_5173,N_5080,N_5060);
nand U5174 (N_5174,N_5051,N_5078);
xnor U5175 (N_5175,N_5013,N_5048);
nor U5176 (N_5176,N_5016,N_5021);
or U5177 (N_5177,N_5078,N_5062);
and U5178 (N_5178,N_5018,N_5068);
and U5179 (N_5179,N_5035,N_5079);
or U5180 (N_5180,N_5002,N_5007);
nor U5181 (N_5181,N_5070,N_5086);
and U5182 (N_5182,N_5092,N_5067);
nor U5183 (N_5183,N_5043,N_5030);
and U5184 (N_5184,N_5053,N_5027);
nand U5185 (N_5185,N_5023,N_5039);
and U5186 (N_5186,N_5022,N_5056);
xnor U5187 (N_5187,N_5036,N_5017);
nand U5188 (N_5188,N_5096,N_5082);
and U5189 (N_5189,N_5022,N_5088);
nor U5190 (N_5190,N_5077,N_5087);
nor U5191 (N_5191,N_5061,N_5078);
and U5192 (N_5192,N_5043,N_5010);
and U5193 (N_5193,N_5083,N_5050);
and U5194 (N_5194,N_5030,N_5055);
or U5195 (N_5195,N_5094,N_5098);
nand U5196 (N_5196,N_5021,N_5055);
nor U5197 (N_5197,N_5030,N_5014);
nand U5198 (N_5198,N_5065,N_5058);
or U5199 (N_5199,N_5032,N_5074);
and U5200 (N_5200,N_5185,N_5159);
and U5201 (N_5201,N_5166,N_5102);
and U5202 (N_5202,N_5132,N_5148);
and U5203 (N_5203,N_5174,N_5183);
or U5204 (N_5204,N_5105,N_5138);
nand U5205 (N_5205,N_5188,N_5109);
or U5206 (N_5206,N_5103,N_5152);
nor U5207 (N_5207,N_5114,N_5146);
or U5208 (N_5208,N_5111,N_5108);
or U5209 (N_5209,N_5119,N_5190);
nand U5210 (N_5210,N_5182,N_5184);
and U5211 (N_5211,N_5164,N_5112);
or U5212 (N_5212,N_5197,N_5175);
nor U5213 (N_5213,N_5180,N_5123);
or U5214 (N_5214,N_5133,N_5113);
nor U5215 (N_5215,N_5144,N_5172);
xor U5216 (N_5216,N_5155,N_5161);
or U5217 (N_5217,N_5165,N_5179);
or U5218 (N_5218,N_5107,N_5191);
nor U5219 (N_5219,N_5151,N_5117);
or U5220 (N_5220,N_5127,N_5160);
and U5221 (N_5221,N_5142,N_5131);
nand U5222 (N_5222,N_5140,N_5153);
and U5223 (N_5223,N_5139,N_5187);
nor U5224 (N_5224,N_5128,N_5192);
nor U5225 (N_5225,N_5157,N_5150);
and U5226 (N_5226,N_5124,N_5149);
and U5227 (N_5227,N_5121,N_5100);
or U5228 (N_5228,N_5177,N_5163);
nand U5229 (N_5229,N_5125,N_5194);
and U5230 (N_5230,N_5176,N_5143);
nor U5231 (N_5231,N_5178,N_5170);
nand U5232 (N_5232,N_5162,N_5141);
nand U5233 (N_5233,N_5196,N_5158);
nand U5234 (N_5234,N_5101,N_5181);
nand U5235 (N_5235,N_5106,N_5110);
or U5236 (N_5236,N_5198,N_5145);
and U5237 (N_5237,N_5154,N_5134);
nand U5238 (N_5238,N_5136,N_5115);
and U5239 (N_5239,N_5168,N_5167);
nor U5240 (N_5240,N_5195,N_5104);
or U5241 (N_5241,N_5156,N_5169);
nand U5242 (N_5242,N_5147,N_5130);
nor U5243 (N_5243,N_5193,N_5126);
and U5244 (N_5244,N_5171,N_5173);
or U5245 (N_5245,N_5186,N_5199);
and U5246 (N_5246,N_5129,N_5120);
and U5247 (N_5247,N_5189,N_5116);
and U5248 (N_5248,N_5135,N_5118);
xnor U5249 (N_5249,N_5137,N_5122);
nand U5250 (N_5250,N_5145,N_5124);
nand U5251 (N_5251,N_5127,N_5107);
or U5252 (N_5252,N_5109,N_5106);
nor U5253 (N_5253,N_5198,N_5103);
nor U5254 (N_5254,N_5100,N_5115);
nand U5255 (N_5255,N_5166,N_5134);
or U5256 (N_5256,N_5145,N_5189);
and U5257 (N_5257,N_5185,N_5166);
nand U5258 (N_5258,N_5164,N_5104);
xor U5259 (N_5259,N_5113,N_5165);
nor U5260 (N_5260,N_5122,N_5143);
or U5261 (N_5261,N_5151,N_5107);
or U5262 (N_5262,N_5141,N_5155);
nor U5263 (N_5263,N_5133,N_5124);
nand U5264 (N_5264,N_5124,N_5155);
or U5265 (N_5265,N_5186,N_5163);
or U5266 (N_5266,N_5123,N_5127);
or U5267 (N_5267,N_5158,N_5133);
nand U5268 (N_5268,N_5131,N_5146);
and U5269 (N_5269,N_5147,N_5156);
nand U5270 (N_5270,N_5147,N_5153);
and U5271 (N_5271,N_5153,N_5146);
and U5272 (N_5272,N_5188,N_5118);
and U5273 (N_5273,N_5114,N_5129);
xnor U5274 (N_5274,N_5123,N_5119);
and U5275 (N_5275,N_5156,N_5167);
or U5276 (N_5276,N_5158,N_5124);
nand U5277 (N_5277,N_5175,N_5140);
nor U5278 (N_5278,N_5110,N_5135);
or U5279 (N_5279,N_5140,N_5132);
or U5280 (N_5280,N_5181,N_5117);
nor U5281 (N_5281,N_5145,N_5166);
and U5282 (N_5282,N_5198,N_5174);
and U5283 (N_5283,N_5144,N_5119);
nor U5284 (N_5284,N_5158,N_5125);
nor U5285 (N_5285,N_5104,N_5173);
xnor U5286 (N_5286,N_5137,N_5132);
nand U5287 (N_5287,N_5129,N_5187);
and U5288 (N_5288,N_5124,N_5195);
nand U5289 (N_5289,N_5198,N_5156);
nor U5290 (N_5290,N_5167,N_5182);
or U5291 (N_5291,N_5150,N_5124);
and U5292 (N_5292,N_5196,N_5172);
and U5293 (N_5293,N_5128,N_5100);
nor U5294 (N_5294,N_5124,N_5188);
or U5295 (N_5295,N_5107,N_5115);
nor U5296 (N_5296,N_5142,N_5182);
nor U5297 (N_5297,N_5124,N_5197);
nor U5298 (N_5298,N_5177,N_5197);
and U5299 (N_5299,N_5105,N_5117);
and U5300 (N_5300,N_5248,N_5200);
xor U5301 (N_5301,N_5286,N_5279);
nand U5302 (N_5302,N_5272,N_5265);
nor U5303 (N_5303,N_5208,N_5255);
or U5304 (N_5304,N_5261,N_5238);
nand U5305 (N_5305,N_5236,N_5278);
or U5306 (N_5306,N_5268,N_5250);
or U5307 (N_5307,N_5299,N_5258);
and U5308 (N_5308,N_5285,N_5291);
or U5309 (N_5309,N_5204,N_5253);
or U5310 (N_5310,N_5257,N_5287);
nand U5311 (N_5311,N_5232,N_5237);
nor U5312 (N_5312,N_5274,N_5252);
and U5313 (N_5313,N_5240,N_5209);
and U5314 (N_5314,N_5277,N_5275);
and U5315 (N_5315,N_5216,N_5293);
nand U5316 (N_5316,N_5244,N_5276);
nand U5317 (N_5317,N_5266,N_5217);
nand U5318 (N_5318,N_5207,N_5225);
nor U5319 (N_5319,N_5214,N_5201);
nand U5320 (N_5320,N_5215,N_5295);
and U5321 (N_5321,N_5221,N_5227);
nor U5322 (N_5322,N_5219,N_5212);
nor U5323 (N_5323,N_5269,N_5239);
or U5324 (N_5324,N_5273,N_5230);
xnor U5325 (N_5325,N_5292,N_5202);
nor U5326 (N_5326,N_5270,N_5226);
nor U5327 (N_5327,N_5211,N_5262);
and U5328 (N_5328,N_5223,N_5288);
or U5329 (N_5329,N_5254,N_5267);
or U5330 (N_5330,N_5281,N_5247);
nand U5331 (N_5331,N_5206,N_5203);
and U5332 (N_5332,N_5220,N_5284);
nand U5333 (N_5333,N_5228,N_5290);
nor U5334 (N_5334,N_5298,N_5241);
nor U5335 (N_5335,N_5294,N_5245);
xor U5336 (N_5336,N_5229,N_5222);
and U5337 (N_5337,N_5243,N_5282);
nor U5338 (N_5338,N_5283,N_5210);
nand U5339 (N_5339,N_5249,N_5264);
nor U5340 (N_5340,N_5256,N_5280);
or U5341 (N_5341,N_5297,N_5296);
nand U5342 (N_5342,N_5234,N_5260);
and U5343 (N_5343,N_5224,N_5259);
and U5344 (N_5344,N_5271,N_5242);
or U5345 (N_5345,N_5235,N_5233);
nor U5346 (N_5346,N_5213,N_5205);
or U5347 (N_5347,N_5218,N_5263);
nand U5348 (N_5348,N_5231,N_5246);
or U5349 (N_5349,N_5251,N_5289);
and U5350 (N_5350,N_5257,N_5263);
nand U5351 (N_5351,N_5288,N_5254);
nor U5352 (N_5352,N_5261,N_5284);
nand U5353 (N_5353,N_5243,N_5247);
xnor U5354 (N_5354,N_5289,N_5278);
nand U5355 (N_5355,N_5232,N_5275);
nand U5356 (N_5356,N_5252,N_5216);
or U5357 (N_5357,N_5229,N_5207);
or U5358 (N_5358,N_5253,N_5297);
nand U5359 (N_5359,N_5229,N_5221);
or U5360 (N_5360,N_5206,N_5290);
nor U5361 (N_5361,N_5239,N_5293);
nor U5362 (N_5362,N_5200,N_5289);
nand U5363 (N_5363,N_5256,N_5249);
and U5364 (N_5364,N_5220,N_5296);
and U5365 (N_5365,N_5273,N_5225);
and U5366 (N_5366,N_5210,N_5235);
or U5367 (N_5367,N_5241,N_5216);
nor U5368 (N_5368,N_5287,N_5209);
nor U5369 (N_5369,N_5278,N_5246);
nand U5370 (N_5370,N_5249,N_5255);
and U5371 (N_5371,N_5294,N_5219);
and U5372 (N_5372,N_5226,N_5256);
nor U5373 (N_5373,N_5277,N_5254);
or U5374 (N_5374,N_5266,N_5235);
or U5375 (N_5375,N_5272,N_5250);
nand U5376 (N_5376,N_5212,N_5214);
or U5377 (N_5377,N_5285,N_5278);
and U5378 (N_5378,N_5238,N_5239);
nand U5379 (N_5379,N_5243,N_5233);
or U5380 (N_5380,N_5212,N_5224);
and U5381 (N_5381,N_5211,N_5265);
or U5382 (N_5382,N_5200,N_5244);
nor U5383 (N_5383,N_5279,N_5226);
or U5384 (N_5384,N_5210,N_5295);
nand U5385 (N_5385,N_5239,N_5223);
or U5386 (N_5386,N_5295,N_5290);
and U5387 (N_5387,N_5262,N_5215);
nor U5388 (N_5388,N_5236,N_5208);
or U5389 (N_5389,N_5265,N_5291);
nand U5390 (N_5390,N_5280,N_5283);
and U5391 (N_5391,N_5205,N_5295);
nor U5392 (N_5392,N_5234,N_5290);
xnor U5393 (N_5393,N_5272,N_5251);
nand U5394 (N_5394,N_5241,N_5284);
nor U5395 (N_5395,N_5280,N_5275);
nor U5396 (N_5396,N_5253,N_5221);
or U5397 (N_5397,N_5202,N_5200);
or U5398 (N_5398,N_5262,N_5238);
nand U5399 (N_5399,N_5270,N_5217);
nor U5400 (N_5400,N_5376,N_5377);
and U5401 (N_5401,N_5305,N_5354);
nand U5402 (N_5402,N_5303,N_5375);
nand U5403 (N_5403,N_5334,N_5314);
or U5404 (N_5404,N_5384,N_5357);
and U5405 (N_5405,N_5339,N_5343);
and U5406 (N_5406,N_5327,N_5382);
and U5407 (N_5407,N_5390,N_5394);
or U5408 (N_5408,N_5396,N_5368);
or U5409 (N_5409,N_5320,N_5389);
nand U5410 (N_5410,N_5324,N_5367);
or U5411 (N_5411,N_5315,N_5330);
and U5412 (N_5412,N_5301,N_5308);
or U5413 (N_5413,N_5369,N_5326);
nor U5414 (N_5414,N_5363,N_5359);
nor U5415 (N_5415,N_5345,N_5306);
or U5416 (N_5416,N_5352,N_5348);
or U5417 (N_5417,N_5328,N_5333);
and U5418 (N_5418,N_5388,N_5331);
nor U5419 (N_5419,N_5341,N_5349);
and U5420 (N_5420,N_5381,N_5380);
or U5421 (N_5421,N_5304,N_5351);
and U5422 (N_5422,N_5399,N_5329);
nand U5423 (N_5423,N_5332,N_5360);
nor U5424 (N_5424,N_5340,N_5336);
or U5425 (N_5425,N_5361,N_5300);
and U5426 (N_5426,N_5358,N_5313);
and U5427 (N_5427,N_5323,N_5344);
or U5428 (N_5428,N_5317,N_5307);
and U5429 (N_5429,N_5392,N_5325);
nor U5430 (N_5430,N_5373,N_5316);
or U5431 (N_5431,N_5347,N_5385);
nand U5432 (N_5432,N_5310,N_5374);
nor U5433 (N_5433,N_5365,N_5395);
nand U5434 (N_5434,N_5335,N_5371);
nand U5435 (N_5435,N_5321,N_5318);
nand U5436 (N_5436,N_5312,N_5337);
and U5437 (N_5437,N_5398,N_5342);
nand U5438 (N_5438,N_5366,N_5387);
nor U5439 (N_5439,N_5370,N_5356);
and U5440 (N_5440,N_5346,N_5379);
or U5441 (N_5441,N_5386,N_5319);
and U5442 (N_5442,N_5309,N_5350);
nand U5443 (N_5443,N_5338,N_5355);
nand U5444 (N_5444,N_5383,N_5397);
or U5445 (N_5445,N_5378,N_5372);
nand U5446 (N_5446,N_5391,N_5393);
and U5447 (N_5447,N_5302,N_5362);
and U5448 (N_5448,N_5322,N_5311);
or U5449 (N_5449,N_5353,N_5364);
nand U5450 (N_5450,N_5359,N_5369);
or U5451 (N_5451,N_5350,N_5377);
nand U5452 (N_5452,N_5345,N_5355);
nand U5453 (N_5453,N_5344,N_5373);
or U5454 (N_5454,N_5377,N_5338);
and U5455 (N_5455,N_5376,N_5306);
or U5456 (N_5456,N_5304,N_5366);
nor U5457 (N_5457,N_5385,N_5354);
nor U5458 (N_5458,N_5353,N_5379);
and U5459 (N_5459,N_5349,N_5364);
and U5460 (N_5460,N_5371,N_5396);
and U5461 (N_5461,N_5326,N_5389);
or U5462 (N_5462,N_5327,N_5351);
or U5463 (N_5463,N_5329,N_5316);
and U5464 (N_5464,N_5336,N_5379);
nand U5465 (N_5465,N_5368,N_5335);
nor U5466 (N_5466,N_5377,N_5343);
or U5467 (N_5467,N_5335,N_5365);
nand U5468 (N_5468,N_5395,N_5392);
nor U5469 (N_5469,N_5360,N_5389);
and U5470 (N_5470,N_5310,N_5332);
or U5471 (N_5471,N_5330,N_5339);
nand U5472 (N_5472,N_5301,N_5328);
or U5473 (N_5473,N_5334,N_5371);
or U5474 (N_5474,N_5333,N_5376);
or U5475 (N_5475,N_5310,N_5386);
xor U5476 (N_5476,N_5387,N_5344);
or U5477 (N_5477,N_5360,N_5326);
and U5478 (N_5478,N_5301,N_5359);
and U5479 (N_5479,N_5302,N_5310);
and U5480 (N_5480,N_5360,N_5378);
nand U5481 (N_5481,N_5302,N_5340);
or U5482 (N_5482,N_5359,N_5323);
or U5483 (N_5483,N_5349,N_5395);
nand U5484 (N_5484,N_5376,N_5304);
nor U5485 (N_5485,N_5312,N_5340);
or U5486 (N_5486,N_5377,N_5326);
nor U5487 (N_5487,N_5337,N_5357);
nor U5488 (N_5488,N_5328,N_5352);
nand U5489 (N_5489,N_5355,N_5354);
nor U5490 (N_5490,N_5371,N_5328);
and U5491 (N_5491,N_5351,N_5398);
or U5492 (N_5492,N_5344,N_5318);
and U5493 (N_5493,N_5370,N_5380);
and U5494 (N_5494,N_5398,N_5379);
and U5495 (N_5495,N_5395,N_5315);
and U5496 (N_5496,N_5370,N_5363);
nor U5497 (N_5497,N_5302,N_5301);
nor U5498 (N_5498,N_5313,N_5347);
xor U5499 (N_5499,N_5300,N_5369);
nand U5500 (N_5500,N_5443,N_5428);
and U5501 (N_5501,N_5494,N_5418);
nor U5502 (N_5502,N_5478,N_5461);
or U5503 (N_5503,N_5459,N_5458);
and U5504 (N_5504,N_5465,N_5469);
or U5505 (N_5505,N_5407,N_5485);
nand U5506 (N_5506,N_5439,N_5431);
or U5507 (N_5507,N_5432,N_5447);
nor U5508 (N_5508,N_5415,N_5445);
nor U5509 (N_5509,N_5460,N_5436);
nand U5510 (N_5510,N_5466,N_5401);
xnor U5511 (N_5511,N_5400,N_5419);
nand U5512 (N_5512,N_5403,N_5437);
nand U5513 (N_5513,N_5492,N_5425);
nor U5514 (N_5514,N_5471,N_5438);
or U5515 (N_5515,N_5412,N_5481);
xnor U5516 (N_5516,N_5404,N_5430);
and U5517 (N_5517,N_5470,N_5414);
nor U5518 (N_5518,N_5422,N_5450);
and U5519 (N_5519,N_5490,N_5487);
nor U5520 (N_5520,N_5464,N_5402);
nor U5521 (N_5521,N_5496,N_5444);
or U5522 (N_5522,N_5495,N_5486);
nor U5523 (N_5523,N_5480,N_5493);
or U5524 (N_5524,N_5499,N_5498);
nor U5525 (N_5525,N_5449,N_5477);
or U5526 (N_5526,N_5476,N_5475);
nor U5527 (N_5527,N_5497,N_5405);
nor U5528 (N_5528,N_5427,N_5411);
and U5529 (N_5529,N_5462,N_5479);
and U5530 (N_5530,N_5488,N_5456);
and U5531 (N_5531,N_5433,N_5420);
or U5532 (N_5532,N_5463,N_5484);
and U5533 (N_5533,N_5417,N_5491);
and U5534 (N_5534,N_5409,N_5408);
and U5535 (N_5535,N_5446,N_5455);
and U5536 (N_5536,N_5423,N_5467);
nor U5537 (N_5537,N_5472,N_5440);
or U5538 (N_5538,N_5483,N_5482);
nor U5539 (N_5539,N_5473,N_5442);
nor U5540 (N_5540,N_5454,N_5489);
and U5541 (N_5541,N_5448,N_5435);
nand U5542 (N_5542,N_5429,N_5441);
xor U5543 (N_5543,N_5468,N_5453);
nand U5544 (N_5544,N_5434,N_5451);
nand U5545 (N_5545,N_5410,N_5416);
and U5546 (N_5546,N_5452,N_5424);
nor U5547 (N_5547,N_5406,N_5421);
or U5548 (N_5548,N_5457,N_5474);
or U5549 (N_5549,N_5413,N_5426);
or U5550 (N_5550,N_5423,N_5437);
and U5551 (N_5551,N_5458,N_5453);
nand U5552 (N_5552,N_5411,N_5497);
nand U5553 (N_5553,N_5499,N_5491);
nor U5554 (N_5554,N_5433,N_5451);
and U5555 (N_5555,N_5485,N_5440);
xnor U5556 (N_5556,N_5445,N_5457);
nor U5557 (N_5557,N_5474,N_5489);
nand U5558 (N_5558,N_5414,N_5459);
or U5559 (N_5559,N_5406,N_5471);
and U5560 (N_5560,N_5461,N_5484);
nor U5561 (N_5561,N_5486,N_5453);
nand U5562 (N_5562,N_5474,N_5464);
or U5563 (N_5563,N_5459,N_5436);
nor U5564 (N_5564,N_5442,N_5486);
and U5565 (N_5565,N_5468,N_5437);
nand U5566 (N_5566,N_5438,N_5401);
or U5567 (N_5567,N_5406,N_5446);
nor U5568 (N_5568,N_5451,N_5418);
xnor U5569 (N_5569,N_5475,N_5438);
nand U5570 (N_5570,N_5420,N_5401);
nor U5571 (N_5571,N_5477,N_5447);
or U5572 (N_5572,N_5498,N_5460);
nor U5573 (N_5573,N_5452,N_5446);
and U5574 (N_5574,N_5453,N_5494);
nor U5575 (N_5575,N_5427,N_5454);
nand U5576 (N_5576,N_5487,N_5460);
and U5577 (N_5577,N_5456,N_5421);
nor U5578 (N_5578,N_5474,N_5420);
or U5579 (N_5579,N_5476,N_5468);
nor U5580 (N_5580,N_5485,N_5437);
and U5581 (N_5581,N_5459,N_5424);
nand U5582 (N_5582,N_5464,N_5473);
xor U5583 (N_5583,N_5487,N_5483);
and U5584 (N_5584,N_5420,N_5411);
nor U5585 (N_5585,N_5409,N_5459);
or U5586 (N_5586,N_5441,N_5467);
nor U5587 (N_5587,N_5438,N_5452);
and U5588 (N_5588,N_5414,N_5415);
and U5589 (N_5589,N_5428,N_5442);
nand U5590 (N_5590,N_5431,N_5481);
nand U5591 (N_5591,N_5432,N_5426);
nand U5592 (N_5592,N_5497,N_5442);
and U5593 (N_5593,N_5495,N_5438);
and U5594 (N_5594,N_5466,N_5431);
and U5595 (N_5595,N_5499,N_5492);
or U5596 (N_5596,N_5460,N_5493);
or U5597 (N_5597,N_5458,N_5464);
or U5598 (N_5598,N_5474,N_5492);
or U5599 (N_5599,N_5492,N_5409);
and U5600 (N_5600,N_5577,N_5515);
nand U5601 (N_5601,N_5543,N_5594);
and U5602 (N_5602,N_5592,N_5570);
nor U5603 (N_5603,N_5527,N_5588);
and U5604 (N_5604,N_5542,N_5538);
and U5605 (N_5605,N_5533,N_5520);
or U5606 (N_5606,N_5597,N_5503);
or U5607 (N_5607,N_5579,N_5540);
and U5608 (N_5608,N_5510,N_5502);
or U5609 (N_5609,N_5557,N_5555);
xnor U5610 (N_5610,N_5580,N_5563);
nor U5611 (N_5611,N_5585,N_5501);
or U5612 (N_5612,N_5587,N_5530);
or U5613 (N_5613,N_5573,N_5514);
nor U5614 (N_5614,N_5596,N_5508);
nor U5615 (N_5615,N_5551,N_5547);
nor U5616 (N_5616,N_5584,N_5536);
or U5617 (N_5617,N_5518,N_5568);
or U5618 (N_5618,N_5539,N_5589);
nand U5619 (N_5619,N_5553,N_5565);
or U5620 (N_5620,N_5571,N_5564);
nor U5621 (N_5621,N_5545,N_5544);
and U5622 (N_5622,N_5599,N_5521);
nor U5623 (N_5623,N_5525,N_5575);
nand U5624 (N_5624,N_5517,N_5581);
and U5625 (N_5625,N_5528,N_5582);
nor U5626 (N_5626,N_5569,N_5529);
nand U5627 (N_5627,N_5535,N_5583);
and U5628 (N_5628,N_5523,N_5574);
and U5629 (N_5629,N_5559,N_5561);
nor U5630 (N_5630,N_5549,N_5506);
nor U5631 (N_5631,N_5572,N_5519);
and U5632 (N_5632,N_5513,N_5516);
nand U5633 (N_5633,N_5537,N_5598);
nor U5634 (N_5634,N_5586,N_5562);
or U5635 (N_5635,N_5593,N_5554);
nand U5636 (N_5636,N_5550,N_5558);
nor U5637 (N_5637,N_5524,N_5595);
nor U5638 (N_5638,N_5534,N_5556);
and U5639 (N_5639,N_5541,N_5509);
nor U5640 (N_5640,N_5505,N_5566);
nor U5641 (N_5641,N_5590,N_5546);
and U5642 (N_5642,N_5507,N_5511);
and U5643 (N_5643,N_5567,N_5500);
and U5644 (N_5644,N_5531,N_5552);
nand U5645 (N_5645,N_5512,N_5591);
or U5646 (N_5646,N_5526,N_5522);
xor U5647 (N_5647,N_5578,N_5504);
and U5648 (N_5648,N_5548,N_5560);
or U5649 (N_5649,N_5532,N_5576);
or U5650 (N_5650,N_5528,N_5550);
or U5651 (N_5651,N_5500,N_5544);
nand U5652 (N_5652,N_5554,N_5588);
nor U5653 (N_5653,N_5595,N_5506);
or U5654 (N_5654,N_5574,N_5593);
and U5655 (N_5655,N_5542,N_5594);
nand U5656 (N_5656,N_5583,N_5571);
nand U5657 (N_5657,N_5509,N_5544);
and U5658 (N_5658,N_5589,N_5578);
or U5659 (N_5659,N_5535,N_5546);
and U5660 (N_5660,N_5590,N_5504);
nand U5661 (N_5661,N_5556,N_5539);
nand U5662 (N_5662,N_5532,N_5530);
nand U5663 (N_5663,N_5547,N_5574);
nand U5664 (N_5664,N_5524,N_5588);
nand U5665 (N_5665,N_5587,N_5507);
nor U5666 (N_5666,N_5532,N_5508);
nand U5667 (N_5667,N_5502,N_5538);
or U5668 (N_5668,N_5587,N_5529);
or U5669 (N_5669,N_5553,N_5510);
nor U5670 (N_5670,N_5544,N_5560);
or U5671 (N_5671,N_5531,N_5547);
and U5672 (N_5672,N_5507,N_5575);
nor U5673 (N_5673,N_5503,N_5506);
and U5674 (N_5674,N_5517,N_5520);
nand U5675 (N_5675,N_5509,N_5581);
nand U5676 (N_5676,N_5513,N_5570);
and U5677 (N_5677,N_5506,N_5532);
or U5678 (N_5678,N_5534,N_5506);
and U5679 (N_5679,N_5510,N_5546);
nor U5680 (N_5680,N_5544,N_5570);
or U5681 (N_5681,N_5560,N_5567);
and U5682 (N_5682,N_5518,N_5523);
nand U5683 (N_5683,N_5518,N_5556);
nor U5684 (N_5684,N_5542,N_5522);
or U5685 (N_5685,N_5523,N_5562);
nor U5686 (N_5686,N_5570,N_5554);
nor U5687 (N_5687,N_5582,N_5562);
xor U5688 (N_5688,N_5536,N_5549);
nand U5689 (N_5689,N_5588,N_5513);
nor U5690 (N_5690,N_5521,N_5546);
or U5691 (N_5691,N_5543,N_5558);
and U5692 (N_5692,N_5585,N_5541);
and U5693 (N_5693,N_5560,N_5531);
or U5694 (N_5694,N_5538,N_5525);
and U5695 (N_5695,N_5583,N_5596);
nand U5696 (N_5696,N_5529,N_5525);
and U5697 (N_5697,N_5577,N_5535);
nor U5698 (N_5698,N_5577,N_5501);
nand U5699 (N_5699,N_5529,N_5572);
and U5700 (N_5700,N_5658,N_5654);
and U5701 (N_5701,N_5622,N_5600);
nor U5702 (N_5702,N_5620,N_5677);
and U5703 (N_5703,N_5669,N_5684);
and U5704 (N_5704,N_5601,N_5691);
nor U5705 (N_5705,N_5689,N_5695);
or U5706 (N_5706,N_5623,N_5665);
or U5707 (N_5707,N_5698,N_5611);
nor U5708 (N_5708,N_5618,N_5627);
nor U5709 (N_5709,N_5678,N_5639);
nand U5710 (N_5710,N_5625,N_5638);
and U5711 (N_5711,N_5664,N_5679);
nand U5712 (N_5712,N_5632,N_5653);
nor U5713 (N_5713,N_5651,N_5662);
nor U5714 (N_5714,N_5641,N_5631);
nand U5715 (N_5715,N_5692,N_5685);
nand U5716 (N_5716,N_5661,N_5696);
and U5717 (N_5717,N_5630,N_5667);
or U5718 (N_5718,N_5629,N_5633);
xnor U5719 (N_5719,N_5674,N_5682);
nand U5720 (N_5720,N_5604,N_5616);
nand U5721 (N_5721,N_5655,N_5635);
nand U5722 (N_5722,N_5652,N_5602);
or U5723 (N_5723,N_5687,N_5681);
and U5724 (N_5724,N_5636,N_5645);
nand U5725 (N_5725,N_5672,N_5673);
xnor U5726 (N_5726,N_5683,N_5670);
or U5727 (N_5727,N_5608,N_5617);
nor U5728 (N_5728,N_5626,N_5614);
and U5729 (N_5729,N_5647,N_5643);
and U5730 (N_5730,N_5640,N_5668);
nor U5731 (N_5731,N_5609,N_5650);
nand U5732 (N_5732,N_5688,N_5663);
nand U5733 (N_5733,N_5605,N_5657);
nand U5734 (N_5734,N_5680,N_5612);
nand U5735 (N_5735,N_5656,N_5648);
and U5736 (N_5736,N_5697,N_5660);
or U5737 (N_5737,N_5646,N_5610);
nand U5738 (N_5738,N_5606,N_5644);
nor U5739 (N_5739,N_5699,N_5676);
nor U5740 (N_5740,N_5642,N_5613);
nor U5741 (N_5741,N_5607,N_5624);
or U5742 (N_5742,N_5603,N_5628);
or U5743 (N_5743,N_5621,N_5671);
or U5744 (N_5744,N_5686,N_5615);
or U5745 (N_5745,N_5694,N_5659);
or U5746 (N_5746,N_5675,N_5637);
and U5747 (N_5747,N_5649,N_5666);
nand U5748 (N_5748,N_5693,N_5619);
nor U5749 (N_5749,N_5690,N_5634);
nand U5750 (N_5750,N_5673,N_5642);
nor U5751 (N_5751,N_5636,N_5696);
xor U5752 (N_5752,N_5618,N_5638);
or U5753 (N_5753,N_5677,N_5635);
or U5754 (N_5754,N_5657,N_5608);
nand U5755 (N_5755,N_5608,N_5683);
nand U5756 (N_5756,N_5616,N_5652);
nor U5757 (N_5757,N_5638,N_5632);
and U5758 (N_5758,N_5664,N_5638);
or U5759 (N_5759,N_5647,N_5640);
nand U5760 (N_5760,N_5626,N_5676);
nand U5761 (N_5761,N_5600,N_5617);
or U5762 (N_5762,N_5652,N_5638);
nand U5763 (N_5763,N_5663,N_5677);
nand U5764 (N_5764,N_5674,N_5656);
nor U5765 (N_5765,N_5671,N_5659);
nor U5766 (N_5766,N_5654,N_5677);
nand U5767 (N_5767,N_5630,N_5605);
or U5768 (N_5768,N_5693,N_5687);
or U5769 (N_5769,N_5625,N_5603);
or U5770 (N_5770,N_5653,N_5640);
nor U5771 (N_5771,N_5643,N_5613);
nor U5772 (N_5772,N_5684,N_5658);
nand U5773 (N_5773,N_5677,N_5640);
nand U5774 (N_5774,N_5627,N_5616);
and U5775 (N_5775,N_5649,N_5690);
nand U5776 (N_5776,N_5662,N_5682);
and U5777 (N_5777,N_5654,N_5683);
and U5778 (N_5778,N_5624,N_5685);
and U5779 (N_5779,N_5666,N_5626);
nor U5780 (N_5780,N_5655,N_5640);
and U5781 (N_5781,N_5603,N_5672);
and U5782 (N_5782,N_5631,N_5672);
nor U5783 (N_5783,N_5666,N_5682);
xor U5784 (N_5784,N_5646,N_5645);
nand U5785 (N_5785,N_5655,N_5627);
nor U5786 (N_5786,N_5690,N_5615);
nor U5787 (N_5787,N_5617,N_5606);
nor U5788 (N_5788,N_5665,N_5686);
and U5789 (N_5789,N_5622,N_5608);
nand U5790 (N_5790,N_5683,N_5658);
and U5791 (N_5791,N_5687,N_5696);
nand U5792 (N_5792,N_5657,N_5685);
nor U5793 (N_5793,N_5615,N_5653);
and U5794 (N_5794,N_5615,N_5682);
nor U5795 (N_5795,N_5602,N_5642);
xnor U5796 (N_5796,N_5649,N_5607);
or U5797 (N_5797,N_5647,N_5692);
or U5798 (N_5798,N_5676,N_5629);
nor U5799 (N_5799,N_5690,N_5627);
and U5800 (N_5800,N_5727,N_5702);
and U5801 (N_5801,N_5785,N_5770);
or U5802 (N_5802,N_5725,N_5720);
nor U5803 (N_5803,N_5705,N_5763);
nor U5804 (N_5804,N_5703,N_5784);
nand U5805 (N_5805,N_5767,N_5710);
and U5806 (N_5806,N_5789,N_5700);
nor U5807 (N_5807,N_5772,N_5738);
nor U5808 (N_5808,N_5771,N_5708);
or U5809 (N_5809,N_5786,N_5792);
and U5810 (N_5810,N_5764,N_5750);
or U5811 (N_5811,N_5707,N_5709);
nand U5812 (N_5812,N_5740,N_5749);
nor U5813 (N_5813,N_5774,N_5783);
or U5814 (N_5814,N_5712,N_5757);
nand U5815 (N_5815,N_5713,N_5775);
or U5816 (N_5816,N_5747,N_5723);
or U5817 (N_5817,N_5762,N_5797);
or U5818 (N_5818,N_5754,N_5756);
and U5819 (N_5819,N_5746,N_5798);
or U5820 (N_5820,N_5731,N_5794);
or U5821 (N_5821,N_5793,N_5717);
and U5822 (N_5822,N_5758,N_5722);
nand U5823 (N_5823,N_5755,N_5780);
nor U5824 (N_5824,N_5768,N_5799);
or U5825 (N_5825,N_5773,N_5711);
and U5826 (N_5826,N_5721,N_5735);
or U5827 (N_5827,N_5718,N_5704);
nand U5828 (N_5828,N_5732,N_5777);
nor U5829 (N_5829,N_5759,N_5745);
nor U5830 (N_5830,N_5737,N_5726);
nor U5831 (N_5831,N_5715,N_5761);
nand U5832 (N_5832,N_5795,N_5752);
and U5833 (N_5833,N_5743,N_5776);
nor U5834 (N_5834,N_5753,N_5765);
or U5835 (N_5835,N_5734,N_5779);
or U5836 (N_5836,N_5766,N_5790);
nand U5837 (N_5837,N_5787,N_5791);
nor U5838 (N_5838,N_5769,N_5760);
nor U5839 (N_5839,N_5719,N_5788);
or U5840 (N_5840,N_5782,N_5751);
or U5841 (N_5841,N_5736,N_5742);
nor U5842 (N_5842,N_5748,N_5730);
and U5843 (N_5843,N_5728,N_5781);
and U5844 (N_5844,N_5706,N_5724);
and U5845 (N_5845,N_5739,N_5714);
or U5846 (N_5846,N_5741,N_5796);
and U5847 (N_5847,N_5778,N_5701);
nand U5848 (N_5848,N_5744,N_5733);
nor U5849 (N_5849,N_5716,N_5729);
xor U5850 (N_5850,N_5784,N_5773);
or U5851 (N_5851,N_5774,N_5740);
nor U5852 (N_5852,N_5727,N_5757);
nor U5853 (N_5853,N_5774,N_5722);
or U5854 (N_5854,N_5749,N_5772);
nor U5855 (N_5855,N_5742,N_5724);
nand U5856 (N_5856,N_5799,N_5734);
or U5857 (N_5857,N_5706,N_5715);
and U5858 (N_5858,N_5707,N_5779);
or U5859 (N_5859,N_5793,N_5798);
and U5860 (N_5860,N_5708,N_5743);
nand U5861 (N_5861,N_5713,N_5760);
or U5862 (N_5862,N_5728,N_5752);
nand U5863 (N_5863,N_5724,N_5761);
or U5864 (N_5864,N_5767,N_5761);
and U5865 (N_5865,N_5778,N_5736);
xor U5866 (N_5866,N_5778,N_5708);
and U5867 (N_5867,N_5773,N_5765);
nand U5868 (N_5868,N_5748,N_5720);
or U5869 (N_5869,N_5798,N_5732);
nor U5870 (N_5870,N_5739,N_5733);
xor U5871 (N_5871,N_5769,N_5703);
and U5872 (N_5872,N_5747,N_5750);
nand U5873 (N_5873,N_5725,N_5711);
nand U5874 (N_5874,N_5724,N_5765);
or U5875 (N_5875,N_5769,N_5710);
or U5876 (N_5876,N_5704,N_5760);
or U5877 (N_5877,N_5761,N_5780);
nand U5878 (N_5878,N_5712,N_5786);
nand U5879 (N_5879,N_5787,N_5736);
or U5880 (N_5880,N_5712,N_5763);
nand U5881 (N_5881,N_5712,N_5746);
nand U5882 (N_5882,N_5793,N_5787);
nor U5883 (N_5883,N_5737,N_5713);
nand U5884 (N_5884,N_5792,N_5773);
or U5885 (N_5885,N_5736,N_5709);
nor U5886 (N_5886,N_5779,N_5791);
nor U5887 (N_5887,N_5772,N_5739);
nand U5888 (N_5888,N_5764,N_5708);
nand U5889 (N_5889,N_5759,N_5717);
and U5890 (N_5890,N_5758,N_5781);
or U5891 (N_5891,N_5732,N_5742);
nor U5892 (N_5892,N_5714,N_5722);
nor U5893 (N_5893,N_5701,N_5733);
nor U5894 (N_5894,N_5704,N_5705);
nand U5895 (N_5895,N_5738,N_5759);
nor U5896 (N_5896,N_5710,N_5723);
nand U5897 (N_5897,N_5712,N_5700);
nand U5898 (N_5898,N_5755,N_5712);
and U5899 (N_5899,N_5787,N_5732);
and U5900 (N_5900,N_5821,N_5813);
and U5901 (N_5901,N_5846,N_5831);
or U5902 (N_5902,N_5857,N_5801);
or U5903 (N_5903,N_5899,N_5882);
nor U5904 (N_5904,N_5858,N_5866);
and U5905 (N_5905,N_5872,N_5803);
nor U5906 (N_5906,N_5815,N_5829);
nor U5907 (N_5907,N_5845,N_5863);
nor U5908 (N_5908,N_5868,N_5825);
nand U5909 (N_5909,N_5808,N_5834);
and U5910 (N_5910,N_5887,N_5880);
nand U5911 (N_5911,N_5886,N_5893);
nand U5912 (N_5912,N_5802,N_5824);
nor U5913 (N_5913,N_5850,N_5874);
nor U5914 (N_5914,N_5873,N_5853);
or U5915 (N_5915,N_5804,N_5851);
nand U5916 (N_5916,N_5871,N_5827);
or U5917 (N_5917,N_5830,N_5826);
and U5918 (N_5918,N_5888,N_5814);
xor U5919 (N_5919,N_5875,N_5895);
and U5920 (N_5920,N_5833,N_5843);
nor U5921 (N_5921,N_5838,N_5807);
nand U5922 (N_5922,N_5856,N_5865);
or U5923 (N_5923,N_5877,N_5864);
nor U5924 (N_5924,N_5869,N_5839);
or U5925 (N_5925,N_5884,N_5867);
nor U5926 (N_5926,N_5870,N_5896);
and U5927 (N_5927,N_5885,N_5894);
nand U5928 (N_5928,N_5892,N_5890);
xnor U5929 (N_5929,N_5847,N_5879);
and U5930 (N_5930,N_5811,N_5820);
and U5931 (N_5931,N_5823,N_5878);
and U5932 (N_5932,N_5844,N_5854);
or U5933 (N_5933,N_5835,N_5809);
and U5934 (N_5934,N_5862,N_5819);
nor U5935 (N_5935,N_5861,N_5883);
and U5936 (N_5936,N_5822,N_5837);
and U5937 (N_5937,N_5898,N_5848);
nand U5938 (N_5938,N_5849,N_5889);
and U5939 (N_5939,N_5842,N_5876);
and U5940 (N_5940,N_5818,N_5855);
nand U5941 (N_5941,N_5812,N_5841);
nor U5942 (N_5942,N_5828,N_5840);
nor U5943 (N_5943,N_5852,N_5832);
nor U5944 (N_5944,N_5806,N_5816);
nand U5945 (N_5945,N_5891,N_5810);
nor U5946 (N_5946,N_5897,N_5881);
and U5947 (N_5947,N_5800,N_5817);
and U5948 (N_5948,N_5836,N_5860);
and U5949 (N_5949,N_5859,N_5805);
nor U5950 (N_5950,N_5849,N_5850);
and U5951 (N_5951,N_5892,N_5865);
or U5952 (N_5952,N_5814,N_5841);
nand U5953 (N_5953,N_5825,N_5858);
nand U5954 (N_5954,N_5838,N_5841);
nand U5955 (N_5955,N_5853,N_5890);
and U5956 (N_5956,N_5826,N_5808);
and U5957 (N_5957,N_5866,N_5841);
nor U5958 (N_5958,N_5874,N_5879);
nor U5959 (N_5959,N_5872,N_5857);
nand U5960 (N_5960,N_5893,N_5833);
nand U5961 (N_5961,N_5892,N_5830);
xnor U5962 (N_5962,N_5811,N_5877);
or U5963 (N_5963,N_5883,N_5839);
nor U5964 (N_5964,N_5885,N_5812);
nor U5965 (N_5965,N_5820,N_5842);
or U5966 (N_5966,N_5884,N_5898);
nor U5967 (N_5967,N_5849,N_5869);
and U5968 (N_5968,N_5897,N_5801);
nand U5969 (N_5969,N_5837,N_5889);
nand U5970 (N_5970,N_5828,N_5831);
nand U5971 (N_5971,N_5857,N_5865);
or U5972 (N_5972,N_5879,N_5803);
or U5973 (N_5973,N_5852,N_5863);
and U5974 (N_5974,N_5866,N_5803);
nand U5975 (N_5975,N_5890,N_5889);
or U5976 (N_5976,N_5802,N_5865);
and U5977 (N_5977,N_5847,N_5857);
or U5978 (N_5978,N_5835,N_5849);
nor U5979 (N_5979,N_5812,N_5832);
nand U5980 (N_5980,N_5850,N_5858);
and U5981 (N_5981,N_5885,N_5875);
and U5982 (N_5982,N_5884,N_5830);
or U5983 (N_5983,N_5844,N_5831);
nand U5984 (N_5984,N_5822,N_5890);
or U5985 (N_5985,N_5885,N_5893);
and U5986 (N_5986,N_5808,N_5849);
or U5987 (N_5987,N_5858,N_5839);
or U5988 (N_5988,N_5864,N_5872);
nor U5989 (N_5989,N_5854,N_5877);
nor U5990 (N_5990,N_5814,N_5853);
or U5991 (N_5991,N_5837,N_5843);
nand U5992 (N_5992,N_5889,N_5858);
nor U5993 (N_5993,N_5831,N_5835);
or U5994 (N_5994,N_5887,N_5812);
or U5995 (N_5995,N_5893,N_5820);
nor U5996 (N_5996,N_5830,N_5878);
nor U5997 (N_5997,N_5881,N_5846);
nand U5998 (N_5998,N_5804,N_5821);
nor U5999 (N_5999,N_5875,N_5887);
nand U6000 (N_6000,N_5917,N_5931);
and U6001 (N_6001,N_5933,N_5941);
and U6002 (N_6002,N_5937,N_5909);
nand U6003 (N_6003,N_5958,N_5963);
or U6004 (N_6004,N_5990,N_5950);
or U6005 (N_6005,N_5905,N_5994);
nand U6006 (N_6006,N_5964,N_5919);
or U6007 (N_6007,N_5962,N_5968);
nor U6008 (N_6008,N_5929,N_5954);
or U6009 (N_6009,N_5913,N_5975);
or U6010 (N_6010,N_5916,N_5902);
or U6011 (N_6011,N_5914,N_5996);
and U6012 (N_6012,N_5921,N_5922);
and U6013 (N_6013,N_5915,N_5903);
nand U6014 (N_6014,N_5928,N_5957);
nor U6015 (N_6015,N_5939,N_5982);
or U6016 (N_6016,N_5995,N_5978);
nand U6017 (N_6017,N_5980,N_5925);
nor U6018 (N_6018,N_5989,N_5945);
and U6019 (N_6019,N_5910,N_5946);
or U6020 (N_6020,N_5951,N_5942);
and U6021 (N_6021,N_5977,N_5960);
and U6022 (N_6022,N_5998,N_5992);
nor U6023 (N_6023,N_5971,N_5967);
xor U6024 (N_6024,N_5983,N_5970);
and U6025 (N_6025,N_5986,N_5927);
and U6026 (N_6026,N_5924,N_5911);
nor U6027 (N_6027,N_5940,N_5938);
or U6028 (N_6028,N_5900,N_5961);
nand U6029 (N_6029,N_5932,N_5974);
and U6030 (N_6030,N_5923,N_5906);
nor U6031 (N_6031,N_5956,N_5979);
nor U6032 (N_6032,N_5935,N_5981);
or U6033 (N_6033,N_5973,N_5984);
and U6034 (N_6034,N_5948,N_5944);
or U6035 (N_6035,N_5987,N_5972);
nor U6036 (N_6036,N_5953,N_5904);
and U6037 (N_6037,N_5943,N_5947);
nand U6038 (N_6038,N_5965,N_5920);
and U6039 (N_6039,N_5955,N_5926);
nand U6040 (N_6040,N_5912,N_5930);
nand U6041 (N_6041,N_5985,N_5993);
nor U6042 (N_6042,N_5997,N_5988);
nand U6043 (N_6043,N_5999,N_5907);
xor U6044 (N_6044,N_5976,N_5908);
nor U6045 (N_6045,N_5934,N_5901);
and U6046 (N_6046,N_5949,N_5936);
nor U6047 (N_6047,N_5952,N_5969);
and U6048 (N_6048,N_5918,N_5959);
and U6049 (N_6049,N_5966,N_5991);
nor U6050 (N_6050,N_5910,N_5925);
or U6051 (N_6051,N_5997,N_5983);
nand U6052 (N_6052,N_5926,N_5923);
and U6053 (N_6053,N_5964,N_5962);
xnor U6054 (N_6054,N_5960,N_5948);
nor U6055 (N_6055,N_5937,N_5950);
or U6056 (N_6056,N_5995,N_5967);
nor U6057 (N_6057,N_5936,N_5958);
nand U6058 (N_6058,N_5905,N_5989);
nor U6059 (N_6059,N_5942,N_5946);
nand U6060 (N_6060,N_5932,N_5920);
nand U6061 (N_6061,N_5952,N_5925);
or U6062 (N_6062,N_5956,N_5959);
and U6063 (N_6063,N_5923,N_5900);
nand U6064 (N_6064,N_5928,N_5915);
and U6065 (N_6065,N_5915,N_5995);
nand U6066 (N_6066,N_5928,N_5982);
and U6067 (N_6067,N_5983,N_5962);
and U6068 (N_6068,N_5979,N_5915);
and U6069 (N_6069,N_5997,N_5979);
xor U6070 (N_6070,N_5945,N_5917);
xnor U6071 (N_6071,N_5993,N_5949);
nor U6072 (N_6072,N_5981,N_5910);
or U6073 (N_6073,N_5981,N_5946);
nand U6074 (N_6074,N_5917,N_5977);
and U6075 (N_6075,N_5941,N_5950);
nor U6076 (N_6076,N_5941,N_5924);
and U6077 (N_6077,N_5990,N_5941);
nor U6078 (N_6078,N_5958,N_5933);
and U6079 (N_6079,N_5950,N_5973);
nand U6080 (N_6080,N_5901,N_5928);
and U6081 (N_6081,N_5976,N_5977);
nor U6082 (N_6082,N_5974,N_5903);
and U6083 (N_6083,N_5956,N_5921);
nor U6084 (N_6084,N_5916,N_5905);
nor U6085 (N_6085,N_5947,N_5914);
nor U6086 (N_6086,N_5938,N_5942);
or U6087 (N_6087,N_5920,N_5951);
nand U6088 (N_6088,N_5985,N_5901);
or U6089 (N_6089,N_5922,N_5985);
and U6090 (N_6090,N_5966,N_5926);
or U6091 (N_6091,N_5924,N_5970);
nor U6092 (N_6092,N_5934,N_5976);
nor U6093 (N_6093,N_5936,N_5961);
nand U6094 (N_6094,N_5956,N_5932);
or U6095 (N_6095,N_5969,N_5911);
nor U6096 (N_6096,N_5964,N_5953);
or U6097 (N_6097,N_5990,N_5909);
and U6098 (N_6098,N_5964,N_5981);
and U6099 (N_6099,N_5902,N_5961);
and U6100 (N_6100,N_6035,N_6012);
nor U6101 (N_6101,N_6052,N_6070);
nand U6102 (N_6102,N_6023,N_6075);
nand U6103 (N_6103,N_6033,N_6004);
or U6104 (N_6104,N_6050,N_6005);
nand U6105 (N_6105,N_6048,N_6022);
or U6106 (N_6106,N_6041,N_6027);
nor U6107 (N_6107,N_6088,N_6055);
and U6108 (N_6108,N_6080,N_6065);
or U6109 (N_6109,N_6029,N_6015);
nor U6110 (N_6110,N_6069,N_6061);
and U6111 (N_6111,N_6021,N_6047);
and U6112 (N_6112,N_6011,N_6000);
and U6113 (N_6113,N_6006,N_6078);
and U6114 (N_6114,N_6073,N_6002);
and U6115 (N_6115,N_6085,N_6090);
and U6116 (N_6116,N_6056,N_6018);
and U6117 (N_6117,N_6042,N_6097);
nor U6118 (N_6118,N_6092,N_6068);
and U6119 (N_6119,N_6045,N_6058);
nor U6120 (N_6120,N_6084,N_6044);
and U6121 (N_6121,N_6019,N_6083);
or U6122 (N_6122,N_6016,N_6057);
or U6123 (N_6123,N_6008,N_6040);
or U6124 (N_6124,N_6098,N_6072);
nor U6125 (N_6125,N_6077,N_6081);
nor U6126 (N_6126,N_6020,N_6099);
and U6127 (N_6127,N_6038,N_6001);
nand U6128 (N_6128,N_6026,N_6049);
nand U6129 (N_6129,N_6043,N_6024);
nand U6130 (N_6130,N_6031,N_6060);
and U6131 (N_6131,N_6067,N_6074);
xnor U6132 (N_6132,N_6091,N_6036);
or U6133 (N_6133,N_6093,N_6096);
and U6134 (N_6134,N_6051,N_6087);
nor U6135 (N_6135,N_6025,N_6046);
or U6136 (N_6136,N_6039,N_6082);
and U6137 (N_6137,N_6095,N_6032);
nand U6138 (N_6138,N_6030,N_6054);
or U6139 (N_6139,N_6010,N_6007);
and U6140 (N_6140,N_6017,N_6064);
nand U6141 (N_6141,N_6037,N_6079);
nand U6142 (N_6142,N_6003,N_6086);
nand U6143 (N_6143,N_6053,N_6063);
nor U6144 (N_6144,N_6066,N_6014);
and U6145 (N_6145,N_6009,N_6062);
and U6146 (N_6146,N_6059,N_6094);
and U6147 (N_6147,N_6034,N_6028);
nor U6148 (N_6148,N_6076,N_6089);
nor U6149 (N_6149,N_6071,N_6013);
nand U6150 (N_6150,N_6097,N_6040);
nor U6151 (N_6151,N_6043,N_6025);
xnor U6152 (N_6152,N_6039,N_6017);
nor U6153 (N_6153,N_6062,N_6040);
nand U6154 (N_6154,N_6000,N_6059);
nand U6155 (N_6155,N_6055,N_6046);
or U6156 (N_6156,N_6075,N_6067);
and U6157 (N_6157,N_6043,N_6045);
nand U6158 (N_6158,N_6000,N_6097);
and U6159 (N_6159,N_6021,N_6058);
nand U6160 (N_6160,N_6003,N_6098);
and U6161 (N_6161,N_6004,N_6072);
nand U6162 (N_6162,N_6009,N_6084);
and U6163 (N_6163,N_6000,N_6033);
nor U6164 (N_6164,N_6012,N_6037);
nor U6165 (N_6165,N_6019,N_6031);
nor U6166 (N_6166,N_6091,N_6016);
or U6167 (N_6167,N_6075,N_6064);
nor U6168 (N_6168,N_6064,N_6000);
nand U6169 (N_6169,N_6090,N_6023);
nand U6170 (N_6170,N_6022,N_6014);
nor U6171 (N_6171,N_6017,N_6080);
nor U6172 (N_6172,N_6035,N_6080);
nand U6173 (N_6173,N_6052,N_6082);
nor U6174 (N_6174,N_6062,N_6000);
nor U6175 (N_6175,N_6054,N_6057);
and U6176 (N_6176,N_6047,N_6088);
nor U6177 (N_6177,N_6002,N_6061);
or U6178 (N_6178,N_6052,N_6059);
and U6179 (N_6179,N_6073,N_6020);
nand U6180 (N_6180,N_6080,N_6014);
and U6181 (N_6181,N_6001,N_6056);
nand U6182 (N_6182,N_6086,N_6028);
nor U6183 (N_6183,N_6052,N_6050);
or U6184 (N_6184,N_6075,N_6055);
or U6185 (N_6185,N_6065,N_6041);
nor U6186 (N_6186,N_6099,N_6014);
nand U6187 (N_6187,N_6083,N_6052);
and U6188 (N_6188,N_6025,N_6023);
and U6189 (N_6189,N_6065,N_6085);
or U6190 (N_6190,N_6032,N_6088);
nand U6191 (N_6191,N_6075,N_6058);
nand U6192 (N_6192,N_6099,N_6088);
nor U6193 (N_6193,N_6041,N_6072);
nor U6194 (N_6194,N_6098,N_6027);
nor U6195 (N_6195,N_6092,N_6031);
or U6196 (N_6196,N_6085,N_6069);
or U6197 (N_6197,N_6032,N_6013);
or U6198 (N_6198,N_6037,N_6083);
and U6199 (N_6199,N_6090,N_6019);
or U6200 (N_6200,N_6177,N_6165);
nor U6201 (N_6201,N_6193,N_6191);
nor U6202 (N_6202,N_6118,N_6157);
nand U6203 (N_6203,N_6102,N_6184);
or U6204 (N_6204,N_6178,N_6176);
nor U6205 (N_6205,N_6147,N_6146);
nand U6206 (N_6206,N_6187,N_6154);
or U6207 (N_6207,N_6106,N_6198);
and U6208 (N_6208,N_6169,N_6197);
or U6209 (N_6209,N_6190,N_6108);
or U6210 (N_6210,N_6181,N_6182);
nor U6211 (N_6211,N_6173,N_6137);
and U6212 (N_6212,N_6166,N_6183);
or U6213 (N_6213,N_6174,N_6172);
and U6214 (N_6214,N_6151,N_6189);
and U6215 (N_6215,N_6104,N_6179);
or U6216 (N_6216,N_6192,N_6180);
xnor U6217 (N_6217,N_6160,N_6164);
nand U6218 (N_6218,N_6116,N_6141);
and U6219 (N_6219,N_6188,N_6123);
or U6220 (N_6220,N_6148,N_6194);
or U6221 (N_6221,N_6139,N_6135);
and U6222 (N_6222,N_6126,N_6170);
nand U6223 (N_6223,N_6149,N_6129);
nor U6224 (N_6224,N_6119,N_6163);
or U6225 (N_6225,N_6175,N_6145);
and U6226 (N_6226,N_6122,N_6195);
and U6227 (N_6227,N_6171,N_6134);
nand U6228 (N_6228,N_6107,N_6131);
nand U6229 (N_6229,N_6150,N_6120);
nor U6230 (N_6230,N_6186,N_6105);
or U6231 (N_6231,N_6113,N_6100);
nor U6232 (N_6232,N_6144,N_6103);
or U6233 (N_6233,N_6138,N_6143);
nand U6234 (N_6234,N_6153,N_6140);
or U6235 (N_6235,N_6124,N_6101);
nor U6236 (N_6236,N_6199,N_6125);
or U6237 (N_6237,N_6168,N_6185);
or U6238 (N_6238,N_6121,N_6155);
nand U6239 (N_6239,N_6152,N_6127);
or U6240 (N_6240,N_6162,N_6161);
or U6241 (N_6241,N_6130,N_6133);
and U6242 (N_6242,N_6132,N_6110);
nand U6243 (N_6243,N_6158,N_6159);
and U6244 (N_6244,N_6196,N_6111);
and U6245 (N_6245,N_6109,N_6136);
nor U6246 (N_6246,N_6142,N_6156);
nand U6247 (N_6247,N_6112,N_6117);
or U6248 (N_6248,N_6115,N_6167);
and U6249 (N_6249,N_6114,N_6128);
nor U6250 (N_6250,N_6117,N_6179);
or U6251 (N_6251,N_6147,N_6168);
or U6252 (N_6252,N_6123,N_6185);
or U6253 (N_6253,N_6178,N_6170);
and U6254 (N_6254,N_6114,N_6178);
and U6255 (N_6255,N_6163,N_6126);
and U6256 (N_6256,N_6193,N_6189);
or U6257 (N_6257,N_6169,N_6158);
or U6258 (N_6258,N_6196,N_6183);
nand U6259 (N_6259,N_6196,N_6182);
or U6260 (N_6260,N_6186,N_6183);
and U6261 (N_6261,N_6129,N_6109);
or U6262 (N_6262,N_6178,N_6116);
nor U6263 (N_6263,N_6189,N_6142);
and U6264 (N_6264,N_6186,N_6156);
nor U6265 (N_6265,N_6176,N_6159);
nor U6266 (N_6266,N_6153,N_6111);
or U6267 (N_6267,N_6129,N_6167);
and U6268 (N_6268,N_6159,N_6135);
or U6269 (N_6269,N_6119,N_6180);
or U6270 (N_6270,N_6190,N_6122);
and U6271 (N_6271,N_6156,N_6164);
or U6272 (N_6272,N_6170,N_6118);
nand U6273 (N_6273,N_6107,N_6165);
and U6274 (N_6274,N_6193,N_6163);
and U6275 (N_6275,N_6103,N_6153);
nand U6276 (N_6276,N_6104,N_6184);
and U6277 (N_6277,N_6137,N_6184);
nor U6278 (N_6278,N_6133,N_6125);
nor U6279 (N_6279,N_6164,N_6109);
nand U6280 (N_6280,N_6159,N_6191);
nor U6281 (N_6281,N_6190,N_6129);
and U6282 (N_6282,N_6143,N_6134);
nand U6283 (N_6283,N_6133,N_6146);
nand U6284 (N_6284,N_6144,N_6133);
nand U6285 (N_6285,N_6182,N_6142);
xor U6286 (N_6286,N_6191,N_6117);
nand U6287 (N_6287,N_6114,N_6155);
or U6288 (N_6288,N_6152,N_6110);
or U6289 (N_6289,N_6143,N_6187);
nor U6290 (N_6290,N_6158,N_6179);
nor U6291 (N_6291,N_6161,N_6168);
nand U6292 (N_6292,N_6175,N_6139);
nor U6293 (N_6293,N_6171,N_6149);
nand U6294 (N_6294,N_6124,N_6187);
nand U6295 (N_6295,N_6130,N_6170);
nor U6296 (N_6296,N_6176,N_6150);
xnor U6297 (N_6297,N_6163,N_6140);
and U6298 (N_6298,N_6117,N_6138);
nand U6299 (N_6299,N_6150,N_6190);
nand U6300 (N_6300,N_6256,N_6245);
or U6301 (N_6301,N_6236,N_6285);
and U6302 (N_6302,N_6206,N_6281);
nor U6303 (N_6303,N_6218,N_6272);
and U6304 (N_6304,N_6292,N_6229);
nor U6305 (N_6305,N_6268,N_6214);
and U6306 (N_6306,N_6259,N_6233);
nor U6307 (N_6307,N_6287,N_6260);
or U6308 (N_6308,N_6277,N_6261);
nand U6309 (N_6309,N_6298,N_6207);
or U6310 (N_6310,N_6297,N_6274);
nand U6311 (N_6311,N_6271,N_6262);
or U6312 (N_6312,N_6263,N_6222);
or U6313 (N_6313,N_6284,N_6205);
and U6314 (N_6314,N_6220,N_6203);
or U6315 (N_6315,N_6293,N_6208);
nand U6316 (N_6316,N_6217,N_6227);
nor U6317 (N_6317,N_6282,N_6212);
nand U6318 (N_6318,N_6238,N_6209);
nand U6319 (N_6319,N_6211,N_6253);
and U6320 (N_6320,N_6279,N_6286);
nand U6321 (N_6321,N_6276,N_6202);
or U6322 (N_6322,N_6249,N_6223);
and U6323 (N_6323,N_6228,N_6235);
nand U6324 (N_6324,N_6204,N_6290);
nor U6325 (N_6325,N_6247,N_6226);
or U6326 (N_6326,N_6225,N_6240);
nand U6327 (N_6327,N_6280,N_6254);
or U6328 (N_6328,N_6295,N_6288);
or U6329 (N_6329,N_6296,N_6270);
or U6330 (N_6330,N_6283,N_6278);
and U6331 (N_6331,N_6231,N_6234);
nor U6332 (N_6332,N_6269,N_6246);
or U6333 (N_6333,N_6232,N_6299);
nand U6334 (N_6334,N_6213,N_6242);
nor U6335 (N_6335,N_6248,N_6258);
nor U6336 (N_6336,N_6243,N_6267);
nor U6337 (N_6337,N_6266,N_6264);
nand U6338 (N_6338,N_6230,N_6252);
nand U6339 (N_6339,N_6257,N_6275);
and U6340 (N_6340,N_6250,N_6239);
nand U6341 (N_6341,N_6200,N_6241);
and U6342 (N_6342,N_6244,N_6273);
or U6343 (N_6343,N_6291,N_6289);
nand U6344 (N_6344,N_6255,N_6251);
or U6345 (N_6345,N_6216,N_6265);
and U6346 (N_6346,N_6237,N_6294);
or U6347 (N_6347,N_6201,N_6210);
nor U6348 (N_6348,N_6219,N_6224);
nand U6349 (N_6349,N_6215,N_6221);
xor U6350 (N_6350,N_6299,N_6297);
nor U6351 (N_6351,N_6249,N_6230);
or U6352 (N_6352,N_6243,N_6222);
nand U6353 (N_6353,N_6203,N_6244);
or U6354 (N_6354,N_6237,N_6200);
nand U6355 (N_6355,N_6269,N_6223);
nand U6356 (N_6356,N_6249,N_6268);
and U6357 (N_6357,N_6202,N_6246);
and U6358 (N_6358,N_6220,N_6277);
nor U6359 (N_6359,N_6251,N_6286);
nor U6360 (N_6360,N_6285,N_6234);
or U6361 (N_6361,N_6274,N_6276);
nor U6362 (N_6362,N_6243,N_6237);
nand U6363 (N_6363,N_6212,N_6285);
nand U6364 (N_6364,N_6257,N_6280);
and U6365 (N_6365,N_6220,N_6283);
and U6366 (N_6366,N_6211,N_6214);
nor U6367 (N_6367,N_6223,N_6236);
nand U6368 (N_6368,N_6246,N_6244);
xnor U6369 (N_6369,N_6285,N_6238);
or U6370 (N_6370,N_6252,N_6232);
nand U6371 (N_6371,N_6259,N_6264);
or U6372 (N_6372,N_6284,N_6276);
or U6373 (N_6373,N_6226,N_6285);
nor U6374 (N_6374,N_6229,N_6277);
nor U6375 (N_6375,N_6229,N_6275);
nor U6376 (N_6376,N_6220,N_6255);
nand U6377 (N_6377,N_6245,N_6200);
or U6378 (N_6378,N_6219,N_6258);
nor U6379 (N_6379,N_6211,N_6225);
or U6380 (N_6380,N_6211,N_6208);
nand U6381 (N_6381,N_6262,N_6211);
nor U6382 (N_6382,N_6257,N_6273);
and U6383 (N_6383,N_6223,N_6240);
and U6384 (N_6384,N_6278,N_6290);
and U6385 (N_6385,N_6281,N_6226);
nor U6386 (N_6386,N_6280,N_6295);
nand U6387 (N_6387,N_6266,N_6265);
or U6388 (N_6388,N_6219,N_6234);
and U6389 (N_6389,N_6268,N_6296);
and U6390 (N_6390,N_6298,N_6235);
nand U6391 (N_6391,N_6262,N_6291);
nand U6392 (N_6392,N_6202,N_6206);
nor U6393 (N_6393,N_6296,N_6211);
nor U6394 (N_6394,N_6223,N_6221);
and U6395 (N_6395,N_6209,N_6266);
or U6396 (N_6396,N_6230,N_6203);
and U6397 (N_6397,N_6267,N_6201);
nand U6398 (N_6398,N_6287,N_6210);
nor U6399 (N_6399,N_6249,N_6293);
or U6400 (N_6400,N_6313,N_6362);
nand U6401 (N_6401,N_6339,N_6347);
nand U6402 (N_6402,N_6329,N_6398);
nor U6403 (N_6403,N_6325,N_6377);
nor U6404 (N_6404,N_6393,N_6376);
nand U6405 (N_6405,N_6315,N_6365);
and U6406 (N_6406,N_6319,N_6389);
nand U6407 (N_6407,N_6316,N_6351);
xor U6408 (N_6408,N_6358,N_6307);
xnor U6409 (N_6409,N_6332,N_6357);
nor U6410 (N_6410,N_6337,N_6363);
or U6411 (N_6411,N_6312,N_6388);
or U6412 (N_6412,N_6333,N_6360);
nor U6413 (N_6413,N_6334,N_6350);
or U6414 (N_6414,N_6349,N_6391);
and U6415 (N_6415,N_6341,N_6385);
nand U6416 (N_6416,N_6306,N_6321);
or U6417 (N_6417,N_6305,N_6322);
or U6418 (N_6418,N_6369,N_6368);
or U6419 (N_6419,N_6320,N_6338);
or U6420 (N_6420,N_6379,N_6317);
or U6421 (N_6421,N_6326,N_6383);
and U6422 (N_6422,N_6375,N_6331);
and U6423 (N_6423,N_6372,N_6395);
or U6424 (N_6424,N_6345,N_6373);
and U6425 (N_6425,N_6354,N_6323);
or U6426 (N_6426,N_6303,N_6302);
nor U6427 (N_6427,N_6394,N_6378);
nand U6428 (N_6428,N_6356,N_6318);
and U6429 (N_6429,N_6361,N_6314);
or U6430 (N_6430,N_6390,N_6364);
nand U6431 (N_6431,N_6324,N_6353);
nand U6432 (N_6432,N_6387,N_6336);
and U6433 (N_6433,N_6359,N_6311);
nor U6434 (N_6434,N_6308,N_6384);
nand U6435 (N_6435,N_6382,N_6301);
nor U6436 (N_6436,N_6327,N_6310);
and U6437 (N_6437,N_6335,N_6346);
or U6438 (N_6438,N_6343,N_6371);
nor U6439 (N_6439,N_6328,N_6344);
nor U6440 (N_6440,N_6397,N_6370);
and U6441 (N_6441,N_6396,N_6300);
or U6442 (N_6442,N_6392,N_6381);
nor U6443 (N_6443,N_6309,N_6330);
nand U6444 (N_6444,N_6342,N_6386);
nor U6445 (N_6445,N_6366,N_6399);
or U6446 (N_6446,N_6374,N_6380);
and U6447 (N_6447,N_6304,N_6355);
and U6448 (N_6448,N_6352,N_6340);
and U6449 (N_6449,N_6367,N_6348);
or U6450 (N_6450,N_6390,N_6387);
nand U6451 (N_6451,N_6362,N_6383);
or U6452 (N_6452,N_6363,N_6396);
nor U6453 (N_6453,N_6334,N_6379);
and U6454 (N_6454,N_6329,N_6316);
or U6455 (N_6455,N_6384,N_6320);
and U6456 (N_6456,N_6398,N_6320);
nand U6457 (N_6457,N_6332,N_6396);
nor U6458 (N_6458,N_6346,N_6389);
nand U6459 (N_6459,N_6313,N_6336);
nand U6460 (N_6460,N_6330,N_6321);
nor U6461 (N_6461,N_6398,N_6395);
nand U6462 (N_6462,N_6319,N_6320);
nor U6463 (N_6463,N_6307,N_6381);
xor U6464 (N_6464,N_6301,N_6343);
or U6465 (N_6465,N_6379,N_6315);
or U6466 (N_6466,N_6344,N_6394);
or U6467 (N_6467,N_6382,N_6316);
nand U6468 (N_6468,N_6336,N_6382);
or U6469 (N_6469,N_6313,N_6380);
xor U6470 (N_6470,N_6319,N_6357);
and U6471 (N_6471,N_6369,N_6342);
and U6472 (N_6472,N_6394,N_6347);
or U6473 (N_6473,N_6333,N_6371);
and U6474 (N_6474,N_6389,N_6363);
and U6475 (N_6475,N_6363,N_6312);
or U6476 (N_6476,N_6349,N_6360);
and U6477 (N_6477,N_6331,N_6308);
or U6478 (N_6478,N_6376,N_6355);
or U6479 (N_6479,N_6303,N_6384);
and U6480 (N_6480,N_6387,N_6370);
nand U6481 (N_6481,N_6330,N_6356);
or U6482 (N_6482,N_6307,N_6329);
or U6483 (N_6483,N_6355,N_6362);
nand U6484 (N_6484,N_6368,N_6340);
xnor U6485 (N_6485,N_6375,N_6300);
and U6486 (N_6486,N_6301,N_6398);
nor U6487 (N_6487,N_6320,N_6349);
xor U6488 (N_6488,N_6327,N_6367);
or U6489 (N_6489,N_6372,N_6333);
and U6490 (N_6490,N_6379,N_6343);
nor U6491 (N_6491,N_6392,N_6352);
or U6492 (N_6492,N_6349,N_6309);
nand U6493 (N_6493,N_6355,N_6329);
nor U6494 (N_6494,N_6335,N_6348);
or U6495 (N_6495,N_6371,N_6337);
nor U6496 (N_6496,N_6355,N_6327);
or U6497 (N_6497,N_6334,N_6398);
nor U6498 (N_6498,N_6354,N_6350);
nand U6499 (N_6499,N_6310,N_6330);
or U6500 (N_6500,N_6489,N_6473);
nor U6501 (N_6501,N_6422,N_6487);
nand U6502 (N_6502,N_6417,N_6433);
and U6503 (N_6503,N_6491,N_6499);
and U6504 (N_6504,N_6447,N_6420);
and U6505 (N_6505,N_6455,N_6477);
nor U6506 (N_6506,N_6468,N_6425);
or U6507 (N_6507,N_6486,N_6481);
or U6508 (N_6508,N_6412,N_6423);
or U6509 (N_6509,N_6450,N_6472);
and U6510 (N_6510,N_6488,N_6495);
and U6511 (N_6511,N_6403,N_6480);
and U6512 (N_6512,N_6419,N_6471);
and U6513 (N_6513,N_6466,N_6458);
and U6514 (N_6514,N_6401,N_6498);
nor U6515 (N_6515,N_6482,N_6470);
nor U6516 (N_6516,N_6406,N_6400);
or U6517 (N_6517,N_6463,N_6494);
nand U6518 (N_6518,N_6496,N_6456);
nand U6519 (N_6519,N_6475,N_6405);
or U6520 (N_6520,N_6459,N_6445);
and U6521 (N_6521,N_6424,N_6490);
or U6522 (N_6522,N_6409,N_6469);
and U6523 (N_6523,N_6436,N_6454);
or U6524 (N_6524,N_6444,N_6438);
nor U6525 (N_6525,N_6408,N_6448);
nor U6526 (N_6526,N_6476,N_6411);
and U6527 (N_6527,N_6442,N_6410);
or U6528 (N_6528,N_6402,N_6439);
and U6529 (N_6529,N_6434,N_6427);
or U6530 (N_6530,N_6432,N_6446);
and U6531 (N_6531,N_6453,N_6413);
and U6532 (N_6532,N_6493,N_6492);
nor U6533 (N_6533,N_6443,N_6435);
nor U6534 (N_6534,N_6462,N_6407);
nor U6535 (N_6535,N_6451,N_6431);
and U6536 (N_6536,N_6464,N_6430);
and U6537 (N_6537,N_6452,N_6441);
nand U6538 (N_6538,N_6479,N_6426);
nand U6539 (N_6539,N_6467,N_6418);
nor U6540 (N_6540,N_6460,N_6497);
nand U6541 (N_6541,N_6414,N_6474);
and U6542 (N_6542,N_6484,N_6440);
and U6543 (N_6543,N_6416,N_6415);
or U6544 (N_6544,N_6465,N_6421);
and U6545 (N_6545,N_6485,N_6429);
or U6546 (N_6546,N_6449,N_6461);
and U6547 (N_6547,N_6457,N_6428);
or U6548 (N_6548,N_6483,N_6404);
and U6549 (N_6549,N_6478,N_6437);
and U6550 (N_6550,N_6405,N_6476);
nor U6551 (N_6551,N_6428,N_6424);
nor U6552 (N_6552,N_6489,N_6494);
or U6553 (N_6553,N_6409,N_6415);
and U6554 (N_6554,N_6422,N_6499);
and U6555 (N_6555,N_6498,N_6473);
or U6556 (N_6556,N_6410,N_6424);
and U6557 (N_6557,N_6490,N_6416);
nor U6558 (N_6558,N_6447,N_6414);
or U6559 (N_6559,N_6424,N_6480);
nand U6560 (N_6560,N_6478,N_6499);
xor U6561 (N_6561,N_6434,N_6493);
nand U6562 (N_6562,N_6493,N_6438);
nand U6563 (N_6563,N_6468,N_6454);
xnor U6564 (N_6564,N_6474,N_6456);
and U6565 (N_6565,N_6444,N_6415);
or U6566 (N_6566,N_6439,N_6411);
nand U6567 (N_6567,N_6495,N_6468);
and U6568 (N_6568,N_6485,N_6422);
and U6569 (N_6569,N_6486,N_6427);
or U6570 (N_6570,N_6465,N_6423);
and U6571 (N_6571,N_6471,N_6490);
nand U6572 (N_6572,N_6416,N_6453);
nand U6573 (N_6573,N_6447,N_6485);
xor U6574 (N_6574,N_6468,N_6410);
or U6575 (N_6575,N_6469,N_6431);
and U6576 (N_6576,N_6485,N_6420);
or U6577 (N_6577,N_6445,N_6455);
or U6578 (N_6578,N_6405,N_6460);
nor U6579 (N_6579,N_6479,N_6438);
or U6580 (N_6580,N_6446,N_6465);
nand U6581 (N_6581,N_6481,N_6447);
or U6582 (N_6582,N_6476,N_6439);
nand U6583 (N_6583,N_6458,N_6430);
nand U6584 (N_6584,N_6424,N_6484);
nor U6585 (N_6585,N_6495,N_6465);
nor U6586 (N_6586,N_6477,N_6406);
xor U6587 (N_6587,N_6457,N_6465);
nand U6588 (N_6588,N_6462,N_6451);
nor U6589 (N_6589,N_6421,N_6481);
xor U6590 (N_6590,N_6418,N_6410);
or U6591 (N_6591,N_6452,N_6442);
nor U6592 (N_6592,N_6450,N_6435);
or U6593 (N_6593,N_6457,N_6495);
nand U6594 (N_6594,N_6457,N_6410);
and U6595 (N_6595,N_6477,N_6413);
or U6596 (N_6596,N_6403,N_6485);
nand U6597 (N_6597,N_6428,N_6406);
or U6598 (N_6598,N_6400,N_6437);
or U6599 (N_6599,N_6499,N_6435);
and U6600 (N_6600,N_6525,N_6506);
and U6601 (N_6601,N_6531,N_6538);
and U6602 (N_6602,N_6524,N_6573);
nand U6603 (N_6603,N_6593,N_6548);
nand U6604 (N_6604,N_6550,N_6546);
nand U6605 (N_6605,N_6503,N_6586);
nand U6606 (N_6606,N_6540,N_6534);
or U6607 (N_6607,N_6590,N_6528);
or U6608 (N_6608,N_6560,N_6507);
nand U6609 (N_6609,N_6535,N_6598);
nor U6610 (N_6610,N_6545,N_6589);
nand U6611 (N_6611,N_6574,N_6597);
nand U6612 (N_6612,N_6588,N_6551);
nand U6613 (N_6613,N_6572,N_6515);
nor U6614 (N_6614,N_6500,N_6579);
or U6615 (N_6615,N_6558,N_6582);
nand U6616 (N_6616,N_6514,N_6508);
nor U6617 (N_6617,N_6585,N_6526);
nand U6618 (N_6618,N_6513,N_6581);
nor U6619 (N_6619,N_6553,N_6596);
nand U6620 (N_6620,N_6544,N_6599);
nor U6621 (N_6621,N_6587,N_6547);
nand U6622 (N_6622,N_6584,N_6504);
nand U6623 (N_6623,N_6527,N_6563);
and U6624 (N_6624,N_6591,N_6561);
and U6625 (N_6625,N_6519,N_6512);
xnor U6626 (N_6626,N_6510,N_6522);
and U6627 (N_6627,N_6568,N_6567);
nor U6628 (N_6628,N_6559,N_6543);
or U6629 (N_6629,N_6530,N_6571);
and U6630 (N_6630,N_6516,N_6583);
and U6631 (N_6631,N_6564,N_6565);
nand U6632 (N_6632,N_6539,N_6502);
or U6633 (N_6633,N_6509,N_6532);
or U6634 (N_6634,N_6517,N_6541);
nand U6635 (N_6635,N_6523,N_6533);
and U6636 (N_6636,N_6562,N_6575);
and U6637 (N_6637,N_6521,N_6549);
or U6638 (N_6638,N_6569,N_6536);
or U6639 (N_6639,N_6557,N_6518);
nor U6640 (N_6640,N_6555,N_6592);
nor U6641 (N_6641,N_6570,N_6542);
nor U6642 (N_6642,N_6566,N_6537);
or U6643 (N_6643,N_6556,N_6505);
and U6644 (N_6644,N_6595,N_6578);
or U6645 (N_6645,N_6511,N_6552);
nor U6646 (N_6646,N_6501,N_6594);
nand U6647 (N_6647,N_6520,N_6577);
nor U6648 (N_6648,N_6580,N_6529);
and U6649 (N_6649,N_6554,N_6576);
nand U6650 (N_6650,N_6577,N_6566);
and U6651 (N_6651,N_6516,N_6542);
xnor U6652 (N_6652,N_6558,N_6557);
nor U6653 (N_6653,N_6519,N_6509);
xor U6654 (N_6654,N_6545,N_6580);
nor U6655 (N_6655,N_6513,N_6599);
nand U6656 (N_6656,N_6542,N_6574);
nor U6657 (N_6657,N_6589,N_6533);
or U6658 (N_6658,N_6581,N_6502);
nand U6659 (N_6659,N_6514,N_6558);
or U6660 (N_6660,N_6573,N_6543);
or U6661 (N_6661,N_6596,N_6569);
and U6662 (N_6662,N_6545,N_6560);
nand U6663 (N_6663,N_6577,N_6578);
nor U6664 (N_6664,N_6550,N_6584);
nor U6665 (N_6665,N_6564,N_6583);
nor U6666 (N_6666,N_6551,N_6501);
and U6667 (N_6667,N_6537,N_6579);
nand U6668 (N_6668,N_6567,N_6535);
nand U6669 (N_6669,N_6519,N_6506);
and U6670 (N_6670,N_6501,N_6564);
nand U6671 (N_6671,N_6528,N_6502);
nand U6672 (N_6672,N_6555,N_6562);
or U6673 (N_6673,N_6524,N_6586);
and U6674 (N_6674,N_6515,N_6545);
or U6675 (N_6675,N_6536,N_6529);
or U6676 (N_6676,N_6500,N_6546);
and U6677 (N_6677,N_6575,N_6507);
xnor U6678 (N_6678,N_6531,N_6556);
and U6679 (N_6679,N_6566,N_6538);
nor U6680 (N_6680,N_6543,N_6507);
or U6681 (N_6681,N_6545,N_6564);
nand U6682 (N_6682,N_6556,N_6519);
or U6683 (N_6683,N_6588,N_6547);
or U6684 (N_6684,N_6519,N_6501);
or U6685 (N_6685,N_6558,N_6578);
nor U6686 (N_6686,N_6533,N_6550);
nor U6687 (N_6687,N_6540,N_6525);
or U6688 (N_6688,N_6584,N_6532);
nand U6689 (N_6689,N_6587,N_6532);
or U6690 (N_6690,N_6595,N_6526);
nand U6691 (N_6691,N_6503,N_6535);
and U6692 (N_6692,N_6509,N_6591);
nand U6693 (N_6693,N_6598,N_6521);
nand U6694 (N_6694,N_6555,N_6537);
nor U6695 (N_6695,N_6589,N_6550);
nor U6696 (N_6696,N_6530,N_6594);
nor U6697 (N_6697,N_6503,N_6530);
nor U6698 (N_6698,N_6538,N_6505);
nor U6699 (N_6699,N_6559,N_6546);
or U6700 (N_6700,N_6690,N_6659);
and U6701 (N_6701,N_6600,N_6680);
or U6702 (N_6702,N_6657,N_6628);
nor U6703 (N_6703,N_6604,N_6688);
xnor U6704 (N_6704,N_6691,N_6679);
nor U6705 (N_6705,N_6641,N_6678);
nor U6706 (N_6706,N_6622,N_6647);
or U6707 (N_6707,N_6638,N_6692);
nor U6708 (N_6708,N_6665,N_6669);
nor U6709 (N_6709,N_6697,N_6618);
nand U6710 (N_6710,N_6671,N_6667);
nand U6711 (N_6711,N_6660,N_6601);
or U6712 (N_6712,N_6617,N_6672);
and U6713 (N_6713,N_6650,N_6602);
nor U6714 (N_6714,N_6674,N_6643);
and U6715 (N_6715,N_6687,N_6615);
or U6716 (N_6716,N_6645,N_6619);
or U6717 (N_6717,N_6636,N_6614);
or U6718 (N_6718,N_6685,N_6610);
nor U6719 (N_6719,N_6620,N_6699);
and U6720 (N_6720,N_6640,N_6648);
or U6721 (N_6721,N_6611,N_6658);
and U6722 (N_6722,N_6662,N_6653);
and U6723 (N_6723,N_6663,N_6666);
nand U6724 (N_6724,N_6609,N_6635);
nand U6725 (N_6725,N_6629,N_6621);
and U6726 (N_6726,N_6695,N_6676);
or U6727 (N_6727,N_6608,N_6644);
or U6728 (N_6728,N_6670,N_6651);
nand U6729 (N_6729,N_6624,N_6642);
and U6730 (N_6730,N_6683,N_6631);
nand U6731 (N_6731,N_6607,N_6693);
nand U6732 (N_6732,N_6633,N_6625);
and U6733 (N_6733,N_6694,N_6652);
nand U6734 (N_6734,N_6677,N_6681);
or U6735 (N_6735,N_6627,N_6630);
nand U6736 (N_6736,N_6612,N_6649);
nand U6737 (N_6737,N_6606,N_6698);
nand U6738 (N_6738,N_6654,N_6684);
nand U6739 (N_6739,N_6686,N_6696);
or U6740 (N_6740,N_6646,N_6632);
nor U6741 (N_6741,N_6637,N_6656);
nand U6742 (N_6742,N_6668,N_6655);
nor U6743 (N_6743,N_6616,N_6682);
or U6744 (N_6744,N_6675,N_6639);
and U6745 (N_6745,N_6613,N_6634);
nor U6746 (N_6746,N_6689,N_6623);
nor U6747 (N_6747,N_6673,N_6603);
or U6748 (N_6748,N_6661,N_6626);
and U6749 (N_6749,N_6605,N_6664);
nor U6750 (N_6750,N_6686,N_6624);
and U6751 (N_6751,N_6601,N_6659);
or U6752 (N_6752,N_6617,N_6685);
nor U6753 (N_6753,N_6654,N_6663);
or U6754 (N_6754,N_6687,N_6644);
nor U6755 (N_6755,N_6681,N_6617);
nor U6756 (N_6756,N_6661,N_6666);
and U6757 (N_6757,N_6633,N_6624);
or U6758 (N_6758,N_6640,N_6677);
nor U6759 (N_6759,N_6672,N_6656);
nor U6760 (N_6760,N_6618,N_6673);
nand U6761 (N_6761,N_6658,N_6687);
or U6762 (N_6762,N_6614,N_6606);
nor U6763 (N_6763,N_6663,N_6665);
nand U6764 (N_6764,N_6661,N_6658);
nand U6765 (N_6765,N_6667,N_6602);
nand U6766 (N_6766,N_6618,N_6653);
and U6767 (N_6767,N_6654,N_6632);
nor U6768 (N_6768,N_6603,N_6694);
nor U6769 (N_6769,N_6637,N_6685);
or U6770 (N_6770,N_6676,N_6671);
nand U6771 (N_6771,N_6627,N_6687);
or U6772 (N_6772,N_6617,N_6660);
or U6773 (N_6773,N_6605,N_6622);
or U6774 (N_6774,N_6627,N_6670);
and U6775 (N_6775,N_6680,N_6678);
nand U6776 (N_6776,N_6640,N_6636);
nor U6777 (N_6777,N_6659,N_6642);
nor U6778 (N_6778,N_6632,N_6671);
nand U6779 (N_6779,N_6607,N_6683);
and U6780 (N_6780,N_6663,N_6682);
or U6781 (N_6781,N_6620,N_6662);
and U6782 (N_6782,N_6619,N_6669);
nand U6783 (N_6783,N_6644,N_6678);
nor U6784 (N_6784,N_6660,N_6662);
and U6785 (N_6785,N_6658,N_6668);
nand U6786 (N_6786,N_6659,N_6649);
nor U6787 (N_6787,N_6696,N_6693);
or U6788 (N_6788,N_6609,N_6607);
nand U6789 (N_6789,N_6659,N_6622);
or U6790 (N_6790,N_6668,N_6657);
or U6791 (N_6791,N_6697,N_6667);
nor U6792 (N_6792,N_6687,N_6656);
nor U6793 (N_6793,N_6665,N_6639);
nor U6794 (N_6794,N_6683,N_6651);
or U6795 (N_6795,N_6686,N_6603);
and U6796 (N_6796,N_6627,N_6669);
and U6797 (N_6797,N_6639,N_6672);
nor U6798 (N_6798,N_6616,N_6679);
and U6799 (N_6799,N_6675,N_6612);
nand U6800 (N_6800,N_6752,N_6729);
or U6801 (N_6801,N_6760,N_6764);
and U6802 (N_6802,N_6767,N_6785);
nand U6803 (N_6803,N_6734,N_6709);
and U6804 (N_6804,N_6750,N_6744);
or U6805 (N_6805,N_6775,N_6722);
nor U6806 (N_6806,N_6706,N_6755);
or U6807 (N_6807,N_6781,N_6795);
nand U6808 (N_6808,N_6704,N_6784);
nand U6809 (N_6809,N_6783,N_6705);
and U6810 (N_6810,N_6717,N_6728);
nand U6811 (N_6811,N_6761,N_6723);
nor U6812 (N_6812,N_6770,N_6799);
nand U6813 (N_6813,N_6745,N_6772);
and U6814 (N_6814,N_6769,N_6777);
or U6815 (N_6815,N_6701,N_6794);
nand U6816 (N_6816,N_6700,N_6763);
and U6817 (N_6817,N_6727,N_6766);
nor U6818 (N_6818,N_6774,N_6707);
nand U6819 (N_6819,N_6797,N_6751);
or U6820 (N_6820,N_6733,N_6792);
xnor U6821 (N_6821,N_6713,N_6786);
xor U6822 (N_6822,N_6748,N_6771);
or U6823 (N_6823,N_6749,N_6716);
or U6824 (N_6824,N_6735,N_6724);
nor U6825 (N_6825,N_6756,N_6773);
or U6826 (N_6826,N_6721,N_6757);
and U6827 (N_6827,N_6793,N_6796);
or U6828 (N_6828,N_6798,N_6718);
nand U6829 (N_6829,N_6703,N_6754);
nor U6830 (N_6830,N_6789,N_6738);
nor U6831 (N_6831,N_6726,N_6708);
and U6832 (N_6832,N_6739,N_6740);
or U6833 (N_6833,N_6737,N_6736);
nand U6834 (N_6834,N_6710,N_6782);
or U6835 (N_6835,N_6743,N_6732);
nor U6836 (N_6836,N_6753,N_6791);
or U6837 (N_6837,N_6742,N_6776);
nor U6838 (N_6838,N_6731,N_6759);
or U6839 (N_6839,N_6712,N_6702);
nand U6840 (N_6840,N_6780,N_6730);
or U6841 (N_6841,N_6768,N_6746);
nor U6842 (N_6842,N_6725,N_6715);
and U6843 (N_6843,N_6711,N_6762);
nand U6844 (N_6844,N_6779,N_6758);
and U6845 (N_6845,N_6765,N_6788);
nand U6846 (N_6846,N_6719,N_6787);
or U6847 (N_6847,N_6741,N_6747);
or U6848 (N_6848,N_6714,N_6790);
and U6849 (N_6849,N_6778,N_6720);
nand U6850 (N_6850,N_6735,N_6789);
or U6851 (N_6851,N_6710,N_6796);
or U6852 (N_6852,N_6732,N_6796);
and U6853 (N_6853,N_6742,N_6785);
xor U6854 (N_6854,N_6739,N_6721);
nand U6855 (N_6855,N_6726,N_6745);
or U6856 (N_6856,N_6754,N_6758);
nor U6857 (N_6857,N_6701,N_6705);
nand U6858 (N_6858,N_6741,N_6792);
or U6859 (N_6859,N_6718,N_6707);
nand U6860 (N_6860,N_6726,N_6757);
xnor U6861 (N_6861,N_6736,N_6742);
nor U6862 (N_6862,N_6762,N_6713);
and U6863 (N_6863,N_6775,N_6730);
nand U6864 (N_6864,N_6782,N_6780);
nand U6865 (N_6865,N_6763,N_6791);
nor U6866 (N_6866,N_6721,N_6703);
nor U6867 (N_6867,N_6775,N_6767);
and U6868 (N_6868,N_6745,N_6736);
nor U6869 (N_6869,N_6715,N_6794);
or U6870 (N_6870,N_6759,N_6752);
or U6871 (N_6871,N_6786,N_6752);
or U6872 (N_6872,N_6748,N_6735);
or U6873 (N_6873,N_6785,N_6727);
or U6874 (N_6874,N_6749,N_6718);
nand U6875 (N_6875,N_6790,N_6728);
xnor U6876 (N_6876,N_6709,N_6726);
nand U6877 (N_6877,N_6736,N_6757);
or U6878 (N_6878,N_6791,N_6768);
nand U6879 (N_6879,N_6763,N_6744);
or U6880 (N_6880,N_6714,N_6766);
and U6881 (N_6881,N_6774,N_6783);
nor U6882 (N_6882,N_6769,N_6701);
nand U6883 (N_6883,N_6724,N_6771);
or U6884 (N_6884,N_6703,N_6782);
or U6885 (N_6885,N_6720,N_6784);
nor U6886 (N_6886,N_6744,N_6798);
and U6887 (N_6887,N_6777,N_6748);
or U6888 (N_6888,N_6742,N_6720);
nor U6889 (N_6889,N_6712,N_6796);
nor U6890 (N_6890,N_6729,N_6773);
nand U6891 (N_6891,N_6792,N_6764);
and U6892 (N_6892,N_6727,N_6784);
or U6893 (N_6893,N_6770,N_6786);
nor U6894 (N_6894,N_6709,N_6751);
xnor U6895 (N_6895,N_6726,N_6736);
nand U6896 (N_6896,N_6793,N_6799);
or U6897 (N_6897,N_6758,N_6714);
nor U6898 (N_6898,N_6758,N_6732);
and U6899 (N_6899,N_6733,N_6781);
and U6900 (N_6900,N_6827,N_6881);
nand U6901 (N_6901,N_6879,N_6825);
nor U6902 (N_6902,N_6818,N_6895);
nor U6903 (N_6903,N_6814,N_6829);
nand U6904 (N_6904,N_6826,N_6846);
and U6905 (N_6905,N_6845,N_6889);
nand U6906 (N_6906,N_6875,N_6809);
nand U6907 (N_6907,N_6897,N_6821);
nand U6908 (N_6908,N_6807,N_6888);
or U6909 (N_6909,N_6850,N_6847);
and U6910 (N_6910,N_6859,N_6887);
nor U6911 (N_6911,N_6898,N_6806);
nand U6912 (N_6912,N_6884,N_6822);
nor U6913 (N_6913,N_6836,N_6865);
nor U6914 (N_6914,N_6800,N_6852);
or U6915 (N_6915,N_6863,N_6801);
nor U6916 (N_6916,N_6853,N_6868);
and U6917 (N_6917,N_6861,N_6802);
nor U6918 (N_6918,N_6860,N_6891);
nand U6919 (N_6919,N_6873,N_6878);
nor U6920 (N_6920,N_6874,N_6851);
and U6921 (N_6921,N_6837,N_6864);
nor U6922 (N_6922,N_6877,N_6838);
and U6923 (N_6923,N_6848,N_6858);
nand U6924 (N_6924,N_6849,N_6870);
nor U6925 (N_6925,N_6819,N_6880);
and U6926 (N_6926,N_6815,N_6842);
nor U6927 (N_6927,N_6841,N_6824);
nand U6928 (N_6928,N_6867,N_6823);
and U6929 (N_6929,N_6803,N_6816);
nand U6930 (N_6930,N_6832,N_6813);
or U6931 (N_6931,N_6840,N_6854);
nor U6932 (N_6932,N_6811,N_6885);
nand U6933 (N_6933,N_6839,N_6871);
nor U6934 (N_6934,N_6833,N_6857);
and U6935 (N_6935,N_6856,N_6820);
and U6936 (N_6936,N_6805,N_6892);
or U6937 (N_6937,N_6866,N_6835);
and U6938 (N_6938,N_6893,N_6843);
nor U6939 (N_6939,N_6844,N_6899);
nand U6940 (N_6940,N_6828,N_6830);
or U6941 (N_6941,N_6817,N_6883);
and U6942 (N_6942,N_6862,N_6872);
or U6943 (N_6943,N_6810,N_6896);
nand U6944 (N_6944,N_6804,N_6834);
and U6945 (N_6945,N_6855,N_6869);
nor U6946 (N_6946,N_6890,N_6894);
nor U6947 (N_6947,N_6876,N_6831);
nor U6948 (N_6948,N_6808,N_6882);
or U6949 (N_6949,N_6886,N_6812);
nor U6950 (N_6950,N_6816,N_6830);
or U6951 (N_6951,N_6894,N_6883);
or U6952 (N_6952,N_6842,N_6897);
xnor U6953 (N_6953,N_6882,N_6897);
and U6954 (N_6954,N_6854,N_6897);
nand U6955 (N_6955,N_6841,N_6861);
and U6956 (N_6956,N_6860,N_6862);
nor U6957 (N_6957,N_6877,N_6878);
or U6958 (N_6958,N_6840,N_6809);
nand U6959 (N_6959,N_6879,N_6899);
nor U6960 (N_6960,N_6871,N_6859);
xnor U6961 (N_6961,N_6823,N_6895);
nand U6962 (N_6962,N_6881,N_6846);
nand U6963 (N_6963,N_6807,N_6850);
or U6964 (N_6964,N_6891,N_6866);
or U6965 (N_6965,N_6812,N_6811);
and U6966 (N_6966,N_6821,N_6837);
and U6967 (N_6967,N_6896,N_6867);
and U6968 (N_6968,N_6816,N_6874);
and U6969 (N_6969,N_6843,N_6889);
nand U6970 (N_6970,N_6814,N_6874);
nand U6971 (N_6971,N_6864,N_6885);
nand U6972 (N_6972,N_6822,N_6872);
and U6973 (N_6973,N_6886,N_6818);
and U6974 (N_6974,N_6803,N_6812);
and U6975 (N_6975,N_6842,N_6855);
nand U6976 (N_6976,N_6897,N_6857);
and U6977 (N_6977,N_6876,N_6888);
nand U6978 (N_6978,N_6821,N_6829);
xnor U6979 (N_6979,N_6810,N_6872);
and U6980 (N_6980,N_6826,N_6841);
nand U6981 (N_6981,N_6802,N_6846);
or U6982 (N_6982,N_6872,N_6825);
nand U6983 (N_6983,N_6869,N_6898);
nand U6984 (N_6984,N_6868,N_6878);
and U6985 (N_6985,N_6804,N_6857);
nor U6986 (N_6986,N_6849,N_6816);
and U6987 (N_6987,N_6821,N_6895);
nand U6988 (N_6988,N_6871,N_6879);
or U6989 (N_6989,N_6895,N_6898);
nor U6990 (N_6990,N_6882,N_6805);
and U6991 (N_6991,N_6816,N_6857);
or U6992 (N_6992,N_6830,N_6802);
and U6993 (N_6993,N_6863,N_6826);
or U6994 (N_6994,N_6830,N_6840);
nor U6995 (N_6995,N_6812,N_6816);
nand U6996 (N_6996,N_6829,N_6878);
and U6997 (N_6997,N_6815,N_6875);
nand U6998 (N_6998,N_6892,N_6825);
or U6999 (N_6999,N_6838,N_6815);
nand U7000 (N_7000,N_6973,N_6991);
nand U7001 (N_7001,N_6924,N_6919);
and U7002 (N_7002,N_6928,N_6918);
nor U7003 (N_7003,N_6982,N_6934);
nand U7004 (N_7004,N_6990,N_6917);
xor U7005 (N_7005,N_6938,N_6941);
or U7006 (N_7006,N_6961,N_6988);
nor U7007 (N_7007,N_6957,N_6909);
and U7008 (N_7008,N_6940,N_6954);
and U7009 (N_7009,N_6996,N_6997);
and U7010 (N_7010,N_6915,N_6955);
and U7011 (N_7011,N_6911,N_6964);
xnor U7012 (N_7012,N_6913,N_6975);
nand U7013 (N_7013,N_6989,N_6974);
and U7014 (N_7014,N_6953,N_6910);
nand U7015 (N_7015,N_6993,N_6921);
or U7016 (N_7016,N_6966,N_6979);
and U7017 (N_7017,N_6976,N_6925);
nand U7018 (N_7018,N_6956,N_6969);
and U7019 (N_7019,N_6999,N_6986);
nand U7020 (N_7020,N_6980,N_6942);
nor U7021 (N_7021,N_6968,N_6922);
nand U7022 (N_7022,N_6994,N_6970);
nand U7023 (N_7023,N_6985,N_6962);
and U7024 (N_7024,N_6903,N_6984);
nand U7025 (N_7025,N_6960,N_6929);
nand U7026 (N_7026,N_6952,N_6939);
nor U7027 (N_7027,N_6987,N_6916);
nand U7028 (N_7028,N_6906,N_6923);
nand U7029 (N_7029,N_6932,N_6902);
nand U7030 (N_7030,N_6943,N_6931);
nand U7031 (N_7031,N_6912,N_6981);
and U7032 (N_7032,N_6958,N_6920);
nor U7033 (N_7033,N_6937,N_6998);
nand U7034 (N_7034,N_6978,N_6901);
or U7035 (N_7035,N_6965,N_6951);
nand U7036 (N_7036,N_6983,N_6905);
or U7037 (N_7037,N_6963,N_6992);
nand U7038 (N_7038,N_6933,N_6936);
or U7039 (N_7039,N_6927,N_6967);
nand U7040 (N_7040,N_6914,N_6945);
nand U7041 (N_7041,N_6946,N_6977);
nand U7042 (N_7042,N_6944,N_6971);
nor U7043 (N_7043,N_6904,N_6950);
nor U7044 (N_7044,N_6935,N_6948);
or U7045 (N_7045,N_6907,N_6930);
and U7046 (N_7046,N_6926,N_6949);
xnor U7047 (N_7047,N_6959,N_6972);
nand U7048 (N_7048,N_6908,N_6947);
or U7049 (N_7049,N_6900,N_6995);
nor U7050 (N_7050,N_6979,N_6930);
and U7051 (N_7051,N_6947,N_6983);
nand U7052 (N_7052,N_6905,N_6908);
and U7053 (N_7053,N_6985,N_6907);
xor U7054 (N_7054,N_6923,N_6958);
or U7055 (N_7055,N_6969,N_6995);
nor U7056 (N_7056,N_6982,N_6989);
and U7057 (N_7057,N_6968,N_6955);
and U7058 (N_7058,N_6990,N_6903);
and U7059 (N_7059,N_6937,N_6919);
and U7060 (N_7060,N_6949,N_6957);
nor U7061 (N_7061,N_6995,N_6953);
nor U7062 (N_7062,N_6984,N_6900);
nor U7063 (N_7063,N_6915,N_6901);
nand U7064 (N_7064,N_6984,N_6961);
nor U7065 (N_7065,N_6997,N_6900);
nor U7066 (N_7066,N_6978,N_6984);
and U7067 (N_7067,N_6912,N_6911);
and U7068 (N_7068,N_6900,N_6917);
nand U7069 (N_7069,N_6906,N_6998);
nand U7070 (N_7070,N_6902,N_6984);
nand U7071 (N_7071,N_6994,N_6967);
nor U7072 (N_7072,N_6907,N_6952);
and U7073 (N_7073,N_6906,N_6937);
or U7074 (N_7074,N_6911,N_6982);
xnor U7075 (N_7075,N_6908,N_6930);
nor U7076 (N_7076,N_6973,N_6917);
and U7077 (N_7077,N_6958,N_6919);
nand U7078 (N_7078,N_6959,N_6928);
nor U7079 (N_7079,N_6913,N_6915);
nand U7080 (N_7080,N_6956,N_6917);
and U7081 (N_7081,N_6923,N_6900);
and U7082 (N_7082,N_6963,N_6967);
and U7083 (N_7083,N_6927,N_6982);
nand U7084 (N_7084,N_6982,N_6904);
nor U7085 (N_7085,N_6925,N_6909);
and U7086 (N_7086,N_6905,N_6961);
nor U7087 (N_7087,N_6998,N_6996);
nand U7088 (N_7088,N_6981,N_6974);
nand U7089 (N_7089,N_6911,N_6951);
nand U7090 (N_7090,N_6985,N_6970);
and U7091 (N_7091,N_6978,N_6963);
nand U7092 (N_7092,N_6930,N_6936);
nor U7093 (N_7093,N_6941,N_6991);
and U7094 (N_7094,N_6910,N_6945);
and U7095 (N_7095,N_6911,N_6995);
nor U7096 (N_7096,N_6930,N_6967);
nand U7097 (N_7097,N_6968,N_6919);
and U7098 (N_7098,N_6912,N_6964);
nor U7099 (N_7099,N_6937,N_6982);
or U7100 (N_7100,N_7038,N_7012);
nor U7101 (N_7101,N_7092,N_7031);
and U7102 (N_7102,N_7097,N_7083);
and U7103 (N_7103,N_7042,N_7066);
nand U7104 (N_7104,N_7033,N_7007);
nand U7105 (N_7105,N_7063,N_7054);
and U7106 (N_7106,N_7029,N_7088);
and U7107 (N_7107,N_7094,N_7040);
or U7108 (N_7108,N_7014,N_7068);
nor U7109 (N_7109,N_7077,N_7000);
or U7110 (N_7110,N_7053,N_7087);
nand U7111 (N_7111,N_7041,N_7091);
or U7112 (N_7112,N_7004,N_7080);
nand U7113 (N_7113,N_7085,N_7065);
nor U7114 (N_7114,N_7084,N_7060);
nor U7115 (N_7115,N_7075,N_7081);
nand U7116 (N_7116,N_7003,N_7058);
and U7117 (N_7117,N_7072,N_7090);
and U7118 (N_7118,N_7017,N_7062);
nand U7119 (N_7119,N_7015,N_7079);
and U7120 (N_7120,N_7070,N_7026);
or U7121 (N_7121,N_7076,N_7055);
and U7122 (N_7122,N_7048,N_7098);
nor U7123 (N_7123,N_7046,N_7089);
and U7124 (N_7124,N_7074,N_7052);
or U7125 (N_7125,N_7005,N_7064);
nand U7126 (N_7126,N_7024,N_7011);
and U7127 (N_7127,N_7099,N_7082);
and U7128 (N_7128,N_7027,N_7071);
or U7129 (N_7129,N_7036,N_7009);
nor U7130 (N_7130,N_7013,N_7043);
nand U7131 (N_7131,N_7073,N_7086);
nor U7132 (N_7132,N_7006,N_7022);
and U7133 (N_7133,N_7049,N_7021);
nor U7134 (N_7134,N_7002,N_7023);
nor U7135 (N_7135,N_7044,N_7010);
or U7136 (N_7136,N_7008,N_7034);
and U7137 (N_7137,N_7078,N_7056);
or U7138 (N_7138,N_7032,N_7001);
nand U7139 (N_7139,N_7095,N_7018);
nand U7140 (N_7140,N_7019,N_7057);
and U7141 (N_7141,N_7067,N_7096);
and U7142 (N_7142,N_7016,N_7051);
or U7143 (N_7143,N_7039,N_7035);
nor U7144 (N_7144,N_7045,N_7037);
nor U7145 (N_7145,N_7047,N_7069);
nand U7146 (N_7146,N_7061,N_7020);
nand U7147 (N_7147,N_7093,N_7030);
nand U7148 (N_7148,N_7028,N_7050);
nand U7149 (N_7149,N_7059,N_7025);
and U7150 (N_7150,N_7039,N_7014);
or U7151 (N_7151,N_7046,N_7028);
and U7152 (N_7152,N_7067,N_7054);
and U7153 (N_7153,N_7072,N_7037);
nor U7154 (N_7154,N_7048,N_7070);
and U7155 (N_7155,N_7051,N_7006);
and U7156 (N_7156,N_7080,N_7050);
nand U7157 (N_7157,N_7061,N_7038);
nand U7158 (N_7158,N_7078,N_7051);
or U7159 (N_7159,N_7071,N_7028);
and U7160 (N_7160,N_7044,N_7095);
nand U7161 (N_7161,N_7041,N_7057);
nor U7162 (N_7162,N_7082,N_7080);
or U7163 (N_7163,N_7098,N_7074);
or U7164 (N_7164,N_7063,N_7029);
and U7165 (N_7165,N_7065,N_7082);
or U7166 (N_7166,N_7009,N_7053);
or U7167 (N_7167,N_7091,N_7013);
and U7168 (N_7168,N_7024,N_7062);
or U7169 (N_7169,N_7063,N_7084);
nor U7170 (N_7170,N_7017,N_7069);
nor U7171 (N_7171,N_7072,N_7007);
and U7172 (N_7172,N_7005,N_7062);
nand U7173 (N_7173,N_7092,N_7055);
and U7174 (N_7174,N_7004,N_7075);
and U7175 (N_7175,N_7020,N_7006);
nor U7176 (N_7176,N_7097,N_7081);
or U7177 (N_7177,N_7018,N_7086);
nand U7178 (N_7178,N_7038,N_7044);
or U7179 (N_7179,N_7070,N_7020);
nor U7180 (N_7180,N_7049,N_7098);
and U7181 (N_7181,N_7057,N_7085);
or U7182 (N_7182,N_7019,N_7079);
and U7183 (N_7183,N_7038,N_7047);
nand U7184 (N_7184,N_7057,N_7056);
nor U7185 (N_7185,N_7086,N_7013);
nor U7186 (N_7186,N_7087,N_7047);
nand U7187 (N_7187,N_7019,N_7045);
and U7188 (N_7188,N_7000,N_7022);
nor U7189 (N_7189,N_7041,N_7066);
nor U7190 (N_7190,N_7013,N_7011);
or U7191 (N_7191,N_7068,N_7050);
nand U7192 (N_7192,N_7004,N_7083);
nand U7193 (N_7193,N_7060,N_7053);
nor U7194 (N_7194,N_7029,N_7044);
and U7195 (N_7195,N_7078,N_7018);
or U7196 (N_7196,N_7025,N_7043);
or U7197 (N_7197,N_7034,N_7085);
nor U7198 (N_7198,N_7078,N_7091);
nand U7199 (N_7199,N_7045,N_7036);
xor U7200 (N_7200,N_7131,N_7157);
nand U7201 (N_7201,N_7132,N_7144);
or U7202 (N_7202,N_7137,N_7102);
or U7203 (N_7203,N_7178,N_7174);
nand U7204 (N_7204,N_7194,N_7155);
and U7205 (N_7205,N_7164,N_7182);
and U7206 (N_7206,N_7153,N_7159);
nor U7207 (N_7207,N_7126,N_7173);
or U7208 (N_7208,N_7172,N_7145);
or U7209 (N_7209,N_7192,N_7190);
nand U7210 (N_7210,N_7106,N_7107);
nor U7211 (N_7211,N_7130,N_7165);
nor U7212 (N_7212,N_7134,N_7195);
nor U7213 (N_7213,N_7152,N_7120);
nand U7214 (N_7214,N_7125,N_7127);
or U7215 (N_7215,N_7197,N_7109);
nor U7216 (N_7216,N_7167,N_7143);
and U7217 (N_7217,N_7147,N_7112);
nand U7218 (N_7218,N_7162,N_7111);
or U7219 (N_7219,N_7118,N_7140);
or U7220 (N_7220,N_7150,N_7141);
nor U7221 (N_7221,N_7105,N_7183);
xnor U7222 (N_7222,N_7198,N_7161);
or U7223 (N_7223,N_7199,N_7103);
nand U7224 (N_7224,N_7189,N_7191);
and U7225 (N_7225,N_7168,N_7196);
or U7226 (N_7226,N_7129,N_7186);
nor U7227 (N_7227,N_7166,N_7121);
or U7228 (N_7228,N_7160,N_7149);
and U7229 (N_7229,N_7181,N_7101);
or U7230 (N_7230,N_7177,N_7188);
nor U7231 (N_7231,N_7104,N_7110);
nor U7232 (N_7232,N_7139,N_7138);
nor U7233 (N_7233,N_7175,N_7193);
nor U7234 (N_7234,N_7142,N_7116);
xor U7235 (N_7235,N_7124,N_7122);
or U7236 (N_7236,N_7119,N_7135);
nand U7237 (N_7237,N_7115,N_7163);
nor U7238 (N_7238,N_7180,N_7146);
or U7239 (N_7239,N_7133,N_7123);
xnor U7240 (N_7240,N_7128,N_7187);
nor U7241 (N_7241,N_7184,N_7148);
nor U7242 (N_7242,N_7114,N_7136);
nand U7243 (N_7243,N_7156,N_7108);
nor U7244 (N_7244,N_7113,N_7170);
or U7245 (N_7245,N_7151,N_7117);
and U7246 (N_7246,N_7158,N_7100);
or U7247 (N_7247,N_7154,N_7185);
and U7248 (N_7248,N_7171,N_7176);
nand U7249 (N_7249,N_7169,N_7179);
nand U7250 (N_7250,N_7122,N_7118);
or U7251 (N_7251,N_7145,N_7132);
and U7252 (N_7252,N_7155,N_7185);
nor U7253 (N_7253,N_7142,N_7124);
and U7254 (N_7254,N_7174,N_7130);
nor U7255 (N_7255,N_7125,N_7107);
nand U7256 (N_7256,N_7178,N_7173);
and U7257 (N_7257,N_7147,N_7138);
nand U7258 (N_7258,N_7165,N_7150);
nand U7259 (N_7259,N_7137,N_7186);
nor U7260 (N_7260,N_7150,N_7149);
and U7261 (N_7261,N_7157,N_7172);
or U7262 (N_7262,N_7101,N_7159);
or U7263 (N_7263,N_7115,N_7109);
and U7264 (N_7264,N_7130,N_7158);
xor U7265 (N_7265,N_7198,N_7101);
and U7266 (N_7266,N_7173,N_7163);
nand U7267 (N_7267,N_7120,N_7116);
nor U7268 (N_7268,N_7191,N_7126);
nand U7269 (N_7269,N_7102,N_7173);
and U7270 (N_7270,N_7123,N_7160);
and U7271 (N_7271,N_7180,N_7187);
nand U7272 (N_7272,N_7149,N_7176);
and U7273 (N_7273,N_7104,N_7156);
and U7274 (N_7274,N_7152,N_7156);
nor U7275 (N_7275,N_7117,N_7129);
nand U7276 (N_7276,N_7199,N_7154);
and U7277 (N_7277,N_7162,N_7171);
nor U7278 (N_7278,N_7190,N_7111);
nand U7279 (N_7279,N_7181,N_7133);
and U7280 (N_7280,N_7110,N_7170);
nand U7281 (N_7281,N_7146,N_7183);
nand U7282 (N_7282,N_7175,N_7100);
and U7283 (N_7283,N_7139,N_7134);
and U7284 (N_7284,N_7173,N_7179);
nand U7285 (N_7285,N_7143,N_7140);
nand U7286 (N_7286,N_7199,N_7120);
and U7287 (N_7287,N_7153,N_7136);
nor U7288 (N_7288,N_7142,N_7140);
or U7289 (N_7289,N_7140,N_7174);
and U7290 (N_7290,N_7108,N_7131);
nand U7291 (N_7291,N_7179,N_7166);
nand U7292 (N_7292,N_7128,N_7176);
nand U7293 (N_7293,N_7172,N_7115);
nor U7294 (N_7294,N_7140,N_7163);
nand U7295 (N_7295,N_7123,N_7177);
nand U7296 (N_7296,N_7198,N_7152);
or U7297 (N_7297,N_7110,N_7105);
and U7298 (N_7298,N_7193,N_7146);
nand U7299 (N_7299,N_7140,N_7122);
and U7300 (N_7300,N_7200,N_7259);
or U7301 (N_7301,N_7230,N_7233);
nor U7302 (N_7302,N_7203,N_7224);
and U7303 (N_7303,N_7219,N_7216);
nor U7304 (N_7304,N_7244,N_7273);
nor U7305 (N_7305,N_7280,N_7238);
nor U7306 (N_7306,N_7227,N_7240);
nor U7307 (N_7307,N_7264,N_7232);
and U7308 (N_7308,N_7207,N_7250);
nand U7309 (N_7309,N_7297,N_7272);
or U7310 (N_7310,N_7206,N_7210);
or U7311 (N_7311,N_7288,N_7290);
nor U7312 (N_7312,N_7275,N_7293);
and U7313 (N_7313,N_7253,N_7249);
nand U7314 (N_7314,N_7204,N_7284);
or U7315 (N_7315,N_7211,N_7247);
and U7316 (N_7316,N_7292,N_7243);
nor U7317 (N_7317,N_7291,N_7298);
or U7318 (N_7318,N_7281,N_7271);
nor U7319 (N_7319,N_7262,N_7221);
nor U7320 (N_7320,N_7261,N_7248);
or U7321 (N_7321,N_7286,N_7283);
or U7322 (N_7322,N_7256,N_7220);
nand U7323 (N_7323,N_7289,N_7294);
nor U7324 (N_7324,N_7270,N_7217);
nand U7325 (N_7325,N_7285,N_7263);
nand U7326 (N_7326,N_7242,N_7214);
nor U7327 (N_7327,N_7299,N_7209);
and U7328 (N_7328,N_7208,N_7235);
nor U7329 (N_7329,N_7226,N_7237);
nand U7330 (N_7330,N_7222,N_7255);
or U7331 (N_7331,N_7260,N_7212);
nor U7332 (N_7332,N_7218,N_7228);
and U7333 (N_7333,N_7241,N_7251);
nor U7334 (N_7334,N_7201,N_7295);
nand U7335 (N_7335,N_7236,N_7229);
nor U7336 (N_7336,N_7268,N_7267);
nor U7337 (N_7337,N_7215,N_7282);
nor U7338 (N_7338,N_7279,N_7278);
or U7339 (N_7339,N_7274,N_7258);
or U7340 (N_7340,N_7239,N_7276);
or U7341 (N_7341,N_7245,N_7277);
or U7342 (N_7342,N_7266,N_7252);
or U7343 (N_7343,N_7213,N_7265);
or U7344 (N_7344,N_7296,N_7231);
nand U7345 (N_7345,N_7287,N_7254);
nand U7346 (N_7346,N_7257,N_7223);
nor U7347 (N_7347,N_7202,N_7234);
and U7348 (N_7348,N_7205,N_7269);
and U7349 (N_7349,N_7246,N_7225);
and U7350 (N_7350,N_7222,N_7260);
nand U7351 (N_7351,N_7238,N_7248);
nand U7352 (N_7352,N_7256,N_7210);
nor U7353 (N_7353,N_7294,N_7282);
and U7354 (N_7354,N_7253,N_7291);
nor U7355 (N_7355,N_7258,N_7289);
or U7356 (N_7356,N_7239,N_7252);
nand U7357 (N_7357,N_7202,N_7225);
nand U7358 (N_7358,N_7253,N_7296);
nand U7359 (N_7359,N_7200,N_7250);
or U7360 (N_7360,N_7210,N_7245);
xor U7361 (N_7361,N_7243,N_7200);
nand U7362 (N_7362,N_7213,N_7200);
nand U7363 (N_7363,N_7219,N_7257);
xor U7364 (N_7364,N_7267,N_7255);
and U7365 (N_7365,N_7239,N_7287);
nor U7366 (N_7366,N_7254,N_7276);
nand U7367 (N_7367,N_7200,N_7267);
nand U7368 (N_7368,N_7253,N_7257);
and U7369 (N_7369,N_7260,N_7214);
nor U7370 (N_7370,N_7259,N_7245);
and U7371 (N_7371,N_7233,N_7225);
or U7372 (N_7372,N_7266,N_7250);
nand U7373 (N_7373,N_7279,N_7219);
or U7374 (N_7374,N_7225,N_7265);
or U7375 (N_7375,N_7266,N_7251);
nor U7376 (N_7376,N_7270,N_7200);
nor U7377 (N_7377,N_7243,N_7229);
and U7378 (N_7378,N_7229,N_7266);
and U7379 (N_7379,N_7257,N_7241);
nand U7380 (N_7380,N_7209,N_7281);
or U7381 (N_7381,N_7202,N_7272);
or U7382 (N_7382,N_7280,N_7290);
nor U7383 (N_7383,N_7231,N_7226);
or U7384 (N_7384,N_7273,N_7238);
nor U7385 (N_7385,N_7281,N_7240);
nand U7386 (N_7386,N_7262,N_7290);
or U7387 (N_7387,N_7292,N_7254);
nor U7388 (N_7388,N_7249,N_7214);
or U7389 (N_7389,N_7200,N_7245);
or U7390 (N_7390,N_7289,N_7234);
nor U7391 (N_7391,N_7253,N_7274);
and U7392 (N_7392,N_7268,N_7287);
nand U7393 (N_7393,N_7268,N_7234);
or U7394 (N_7394,N_7241,N_7207);
or U7395 (N_7395,N_7288,N_7220);
nor U7396 (N_7396,N_7223,N_7270);
or U7397 (N_7397,N_7246,N_7257);
nor U7398 (N_7398,N_7297,N_7232);
nor U7399 (N_7399,N_7238,N_7253);
nand U7400 (N_7400,N_7358,N_7361);
and U7401 (N_7401,N_7334,N_7315);
and U7402 (N_7402,N_7303,N_7326);
and U7403 (N_7403,N_7341,N_7305);
and U7404 (N_7404,N_7316,N_7383);
nand U7405 (N_7405,N_7311,N_7364);
nand U7406 (N_7406,N_7332,N_7395);
nand U7407 (N_7407,N_7329,N_7393);
nand U7408 (N_7408,N_7338,N_7309);
or U7409 (N_7409,N_7318,N_7304);
and U7410 (N_7410,N_7378,N_7357);
nand U7411 (N_7411,N_7333,N_7386);
nand U7412 (N_7412,N_7392,N_7312);
nand U7413 (N_7413,N_7389,N_7300);
nand U7414 (N_7414,N_7371,N_7351);
or U7415 (N_7415,N_7323,N_7342);
nand U7416 (N_7416,N_7347,N_7313);
and U7417 (N_7417,N_7324,N_7336);
and U7418 (N_7418,N_7370,N_7346);
nand U7419 (N_7419,N_7397,N_7314);
nand U7420 (N_7420,N_7340,N_7385);
nand U7421 (N_7421,N_7330,N_7363);
and U7422 (N_7422,N_7327,N_7339);
nor U7423 (N_7423,N_7384,N_7373);
and U7424 (N_7424,N_7368,N_7319);
and U7425 (N_7425,N_7353,N_7382);
nor U7426 (N_7426,N_7356,N_7399);
nor U7427 (N_7427,N_7302,N_7317);
nor U7428 (N_7428,N_7354,N_7376);
nand U7429 (N_7429,N_7365,N_7377);
and U7430 (N_7430,N_7366,N_7398);
and U7431 (N_7431,N_7380,N_7306);
or U7432 (N_7432,N_7345,N_7308);
nand U7433 (N_7433,N_7322,N_7320);
nand U7434 (N_7434,N_7307,N_7352);
and U7435 (N_7435,N_7331,N_7372);
nand U7436 (N_7436,N_7396,N_7369);
nor U7437 (N_7437,N_7321,N_7355);
nor U7438 (N_7438,N_7359,N_7394);
and U7439 (N_7439,N_7343,N_7390);
or U7440 (N_7440,N_7387,N_7381);
or U7441 (N_7441,N_7379,N_7328);
or U7442 (N_7442,N_7325,N_7337);
and U7443 (N_7443,N_7335,N_7391);
or U7444 (N_7444,N_7350,N_7375);
nor U7445 (N_7445,N_7360,N_7374);
nand U7446 (N_7446,N_7388,N_7301);
nor U7447 (N_7447,N_7348,N_7344);
and U7448 (N_7448,N_7349,N_7310);
nor U7449 (N_7449,N_7367,N_7362);
and U7450 (N_7450,N_7386,N_7303);
nand U7451 (N_7451,N_7353,N_7312);
or U7452 (N_7452,N_7326,N_7376);
or U7453 (N_7453,N_7351,N_7341);
or U7454 (N_7454,N_7340,N_7368);
xnor U7455 (N_7455,N_7386,N_7392);
xnor U7456 (N_7456,N_7393,N_7359);
nor U7457 (N_7457,N_7333,N_7368);
nand U7458 (N_7458,N_7326,N_7396);
or U7459 (N_7459,N_7319,N_7347);
nand U7460 (N_7460,N_7356,N_7380);
nand U7461 (N_7461,N_7323,N_7367);
or U7462 (N_7462,N_7335,N_7385);
and U7463 (N_7463,N_7353,N_7303);
xnor U7464 (N_7464,N_7386,N_7338);
and U7465 (N_7465,N_7389,N_7369);
and U7466 (N_7466,N_7379,N_7393);
and U7467 (N_7467,N_7345,N_7318);
nor U7468 (N_7468,N_7335,N_7331);
and U7469 (N_7469,N_7314,N_7359);
or U7470 (N_7470,N_7357,N_7309);
or U7471 (N_7471,N_7383,N_7339);
or U7472 (N_7472,N_7396,N_7371);
xnor U7473 (N_7473,N_7315,N_7324);
and U7474 (N_7474,N_7331,N_7399);
nand U7475 (N_7475,N_7378,N_7398);
and U7476 (N_7476,N_7328,N_7397);
or U7477 (N_7477,N_7353,N_7352);
or U7478 (N_7478,N_7374,N_7385);
and U7479 (N_7479,N_7335,N_7377);
nand U7480 (N_7480,N_7309,N_7342);
nor U7481 (N_7481,N_7346,N_7362);
or U7482 (N_7482,N_7317,N_7301);
xnor U7483 (N_7483,N_7382,N_7371);
or U7484 (N_7484,N_7370,N_7344);
nand U7485 (N_7485,N_7361,N_7336);
nand U7486 (N_7486,N_7393,N_7328);
nor U7487 (N_7487,N_7340,N_7341);
nor U7488 (N_7488,N_7346,N_7371);
or U7489 (N_7489,N_7339,N_7346);
nor U7490 (N_7490,N_7301,N_7350);
and U7491 (N_7491,N_7340,N_7315);
nor U7492 (N_7492,N_7346,N_7388);
and U7493 (N_7493,N_7334,N_7345);
nand U7494 (N_7494,N_7381,N_7358);
nand U7495 (N_7495,N_7391,N_7386);
or U7496 (N_7496,N_7379,N_7381);
or U7497 (N_7497,N_7306,N_7382);
nor U7498 (N_7498,N_7323,N_7331);
nand U7499 (N_7499,N_7330,N_7327);
nor U7500 (N_7500,N_7467,N_7453);
nor U7501 (N_7501,N_7430,N_7428);
nand U7502 (N_7502,N_7436,N_7421);
and U7503 (N_7503,N_7424,N_7486);
nand U7504 (N_7504,N_7415,N_7441);
nand U7505 (N_7505,N_7426,N_7496);
nand U7506 (N_7506,N_7404,N_7490);
and U7507 (N_7507,N_7485,N_7495);
or U7508 (N_7508,N_7403,N_7482);
nor U7509 (N_7509,N_7413,N_7401);
nand U7510 (N_7510,N_7462,N_7484);
or U7511 (N_7511,N_7448,N_7452);
and U7512 (N_7512,N_7447,N_7481);
nand U7513 (N_7513,N_7498,N_7492);
nor U7514 (N_7514,N_7443,N_7473);
or U7515 (N_7515,N_7474,N_7497);
and U7516 (N_7516,N_7445,N_7414);
nand U7517 (N_7517,N_7418,N_7472);
or U7518 (N_7518,N_7480,N_7408);
and U7519 (N_7519,N_7499,N_7444);
nand U7520 (N_7520,N_7409,N_7478);
nand U7521 (N_7521,N_7451,N_7479);
nand U7522 (N_7522,N_7461,N_7411);
or U7523 (N_7523,N_7429,N_7469);
nand U7524 (N_7524,N_7442,N_7488);
nor U7525 (N_7525,N_7412,N_7458);
nor U7526 (N_7526,N_7417,N_7449);
nand U7527 (N_7527,N_7450,N_7420);
nor U7528 (N_7528,N_7494,N_7435);
or U7529 (N_7529,N_7468,N_7406);
and U7530 (N_7530,N_7434,N_7402);
nand U7531 (N_7531,N_7454,N_7455);
xnor U7532 (N_7532,N_7431,N_7437);
nor U7533 (N_7533,N_7459,N_7465);
and U7534 (N_7534,N_7416,N_7439);
nand U7535 (N_7535,N_7405,N_7475);
nor U7536 (N_7536,N_7423,N_7425);
or U7537 (N_7537,N_7470,N_7410);
nor U7538 (N_7538,N_7483,N_7456);
or U7539 (N_7539,N_7464,N_7407);
or U7540 (N_7540,N_7457,N_7438);
nor U7541 (N_7541,N_7432,N_7440);
or U7542 (N_7542,N_7477,N_7489);
or U7543 (N_7543,N_7446,N_7419);
and U7544 (N_7544,N_7422,N_7493);
or U7545 (N_7545,N_7471,N_7466);
nand U7546 (N_7546,N_7487,N_7400);
and U7547 (N_7547,N_7427,N_7463);
and U7548 (N_7548,N_7433,N_7476);
or U7549 (N_7549,N_7491,N_7460);
or U7550 (N_7550,N_7440,N_7406);
nand U7551 (N_7551,N_7497,N_7422);
nand U7552 (N_7552,N_7473,N_7458);
nor U7553 (N_7553,N_7474,N_7446);
and U7554 (N_7554,N_7445,N_7444);
nor U7555 (N_7555,N_7466,N_7439);
nand U7556 (N_7556,N_7470,N_7459);
and U7557 (N_7557,N_7439,N_7421);
nand U7558 (N_7558,N_7448,N_7443);
and U7559 (N_7559,N_7423,N_7490);
nand U7560 (N_7560,N_7435,N_7408);
nor U7561 (N_7561,N_7497,N_7431);
and U7562 (N_7562,N_7485,N_7470);
nor U7563 (N_7563,N_7453,N_7428);
nor U7564 (N_7564,N_7434,N_7493);
nor U7565 (N_7565,N_7498,N_7457);
or U7566 (N_7566,N_7483,N_7463);
nand U7567 (N_7567,N_7496,N_7433);
or U7568 (N_7568,N_7462,N_7465);
nand U7569 (N_7569,N_7440,N_7425);
and U7570 (N_7570,N_7464,N_7499);
xnor U7571 (N_7571,N_7453,N_7452);
nor U7572 (N_7572,N_7437,N_7452);
nor U7573 (N_7573,N_7419,N_7489);
nand U7574 (N_7574,N_7460,N_7421);
or U7575 (N_7575,N_7408,N_7405);
nand U7576 (N_7576,N_7426,N_7402);
or U7577 (N_7577,N_7492,N_7452);
nor U7578 (N_7578,N_7422,N_7490);
nor U7579 (N_7579,N_7424,N_7446);
or U7580 (N_7580,N_7402,N_7404);
nand U7581 (N_7581,N_7418,N_7431);
or U7582 (N_7582,N_7400,N_7426);
and U7583 (N_7583,N_7402,N_7491);
and U7584 (N_7584,N_7423,N_7451);
nor U7585 (N_7585,N_7436,N_7439);
or U7586 (N_7586,N_7420,N_7453);
and U7587 (N_7587,N_7487,N_7417);
and U7588 (N_7588,N_7425,N_7417);
or U7589 (N_7589,N_7472,N_7424);
nand U7590 (N_7590,N_7486,N_7439);
nor U7591 (N_7591,N_7420,N_7425);
nand U7592 (N_7592,N_7401,N_7415);
nor U7593 (N_7593,N_7489,N_7431);
nand U7594 (N_7594,N_7413,N_7431);
and U7595 (N_7595,N_7442,N_7447);
nand U7596 (N_7596,N_7407,N_7459);
and U7597 (N_7597,N_7405,N_7414);
xnor U7598 (N_7598,N_7445,N_7494);
and U7599 (N_7599,N_7477,N_7412);
nand U7600 (N_7600,N_7524,N_7558);
nor U7601 (N_7601,N_7574,N_7572);
and U7602 (N_7602,N_7521,N_7587);
nand U7603 (N_7603,N_7575,N_7545);
or U7604 (N_7604,N_7503,N_7567);
nand U7605 (N_7605,N_7551,N_7530);
nand U7606 (N_7606,N_7579,N_7509);
and U7607 (N_7607,N_7566,N_7578);
nand U7608 (N_7608,N_7510,N_7591);
or U7609 (N_7609,N_7541,N_7532);
nand U7610 (N_7610,N_7582,N_7556);
nand U7611 (N_7611,N_7581,N_7500);
nand U7612 (N_7612,N_7549,N_7515);
nand U7613 (N_7613,N_7569,N_7596);
or U7614 (N_7614,N_7522,N_7561);
xnor U7615 (N_7615,N_7546,N_7501);
and U7616 (N_7616,N_7590,N_7539);
nor U7617 (N_7617,N_7589,N_7517);
nor U7618 (N_7618,N_7542,N_7553);
xnor U7619 (N_7619,N_7504,N_7586);
nor U7620 (N_7620,N_7512,N_7525);
nand U7621 (N_7621,N_7554,N_7588);
nor U7622 (N_7622,N_7570,N_7597);
and U7623 (N_7623,N_7528,N_7508);
or U7624 (N_7624,N_7565,N_7571);
nor U7625 (N_7625,N_7533,N_7595);
nor U7626 (N_7626,N_7523,N_7514);
nand U7627 (N_7627,N_7583,N_7547);
nor U7628 (N_7628,N_7518,N_7516);
and U7629 (N_7629,N_7550,N_7552);
nor U7630 (N_7630,N_7598,N_7527);
or U7631 (N_7631,N_7543,N_7593);
nand U7632 (N_7632,N_7505,N_7519);
nand U7633 (N_7633,N_7564,N_7577);
and U7634 (N_7634,N_7513,N_7599);
or U7635 (N_7635,N_7548,N_7557);
nand U7636 (N_7636,N_7562,N_7573);
nand U7637 (N_7637,N_7560,N_7534);
or U7638 (N_7638,N_7555,N_7544);
nand U7639 (N_7639,N_7529,N_7511);
nor U7640 (N_7640,N_7592,N_7538);
or U7641 (N_7641,N_7507,N_7535);
or U7642 (N_7642,N_7594,N_7537);
and U7643 (N_7643,N_7559,N_7526);
or U7644 (N_7644,N_7584,N_7540);
nand U7645 (N_7645,N_7502,N_7563);
xnor U7646 (N_7646,N_7580,N_7585);
or U7647 (N_7647,N_7531,N_7520);
nor U7648 (N_7648,N_7568,N_7576);
or U7649 (N_7649,N_7536,N_7506);
and U7650 (N_7650,N_7510,N_7530);
or U7651 (N_7651,N_7527,N_7585);
nor U7652 (N_7652,N_7589,N_7547);
or U7653 (N_7653,N_7591,N_7564);
and U7654 (N_7654,N_7512,N_7511);
nand U7655 (N_7655,N_7533,N_7558);
nand U7656 (N_7656,N_7545,N_7501);
and U7657 (N_7657,N_7521,N_7512);
nor U7658 (N_7658,N_7515,N_7520);
nand U7659 (N_7659,N_7548,N_7531);
nand U7660 (N_7660,N_7519,N_7589);
xor U7661 (N_7661,N_7508,N_7521);
nand U7662 (N_7662,N_7572,N_7578);
nand U7663 (N_7663,N_7570,N_7544);
nand U7664 (N_7664,N_7511,N_7525);
or U7665 (N_7665,N_7561,N_7599);
or U7666 (N_7666,N_7561,N_7565);
and U7667 (N_7667,N_7569,N_7585);
and U7668 (N_7668,N_7589,N_7559);
nor U7669 (N_7669,N_7594,N_7540);
nand U7670 (N_7670,N_7552,N_7527);
or U7671 (N_7671,N_7550,N_7527);
nor U7672 (N_7672,N_7581,N_7598);
or U7673 (N_7673,N_7500,N_7574);
xor U7674 (N_7674,N_7560,N_7551);
nand U7675 (N_7675,N_7519,N_7585);
and U7676 (N_7676,N_7552,N_7559);
and U7677 (N_7677,N_7505,N_7529);
nor U7678 (N_7678,N_7504,N_7508);
and U7679 (N_7679,N_7502,N_7544);
nand U7680 (N_7680,N_7556,N_7580);
and U7681 (N_7681,N_7565,N_7580);
or U7682 (N_7682,N_7523,N_7526);
nand U7683 (N_7683,N_7569,N_7588);
nand U7684 (N_7684,N_7511,N_7577);
and U7685 (N_7685,N_7571,N_7518);
or U7686 (N_7686,N_7598,N_7501);
nor U7687 (N_7687,N_7588,N_7532);
and U7688 (N_7688,N_7542,N_7527);
nand U7689 (N_7689,N_7585,N_7599);
and U7690 (N_7690,N_7509,N_7505);
or U7691 (N_7691,N_7537,N_7513);
nand U7692 (N_7692,N_7565,N_7553);
nor U7693 (N_7693,N_7535,N_7542);
nor U7694 (N_7694,N_7512,N_7547);
and U7695 (N_7695,N_7526,N_7542);
nand U7696 (N_7696,N_7505,N_7553);
nand U7697 (N_7697,N_7592,N_7522);
nand U7698 (N_7698,N_7517,N_7515);
or U7699 (N_7699,N_7566,N_7537);
nand U7700 (N_7700,N_7615,N_7610);
and U7701 (N_7701,N_7639,N_7630);
and U7702 (N_7702,N_7649,N_7637);
nor U7703 (N_7703,N_7621,N_7697);
nand U7704 (N_7704,N_7674,N_7665);
nor U7705 (N_7705,N_7619,N_7641);
nor U7706 (N_7706,N_7670,N_7612);
nand U7707 (N_7707,N_7667,N_7695);
and U7708 (N_7708,N_7657,N_7689);
and U7709 (N_7709,N_7608,N_7618);
nand U7710 (N_7710,N_7614,N_7634);
or U7711 (N_7711,N_7661,N_7636);
and U7712 (N_7712,N_7633,N_7694);
nor U7713 (N_7713,N_7635,N_7622);
or U7714 (N_7714,N_7652,N_7651);
nor U7715 (N_7715,N_7690,N_7603);
nor U7716 (N_7716,N_7675,N_7600);
and U7717 (N_7717,N_7631,N_7607);
nand U7718 (N_7718,N_7602,N_7642);
nor U7719 (N_7719,N_7672,N_7678);
and U7720 (N_7720,N_7660,N_7623);
and U7721 (N_7721,N_7679,N_7653);
and U7722 (N_7722,N_7645,N_7605);
nor U7723 (N_7723,N_7659,N_7683);
and U7724 (N_7724,N_7668,N_7696);
or U7725 (N_7725,N_7648,N_7617);
nand U7726 (N_7726,N_7671,N_7682);
nand U7727 (N_7727,N_7688,N_7626);
nor U7728 (N_7728,N_7604,N_7620);
xor U7729 (N_7729,N_7681,N_7677);
nor U7730 (N_7730,N_7628,N_7647);
nor U7731 (N_7731,N_7673,N_7655);
xnor U7732 (N_7732,N_7664,N_7601);
nand U7733 (N_7733,N_7663,N_7656);
and U7734 (N_7734,N_7680,N_7625);
or U7735 (N_7735,N_7650,N_7646);
nand U7736 (N_7736,N_7616,N_7629);
nand U7737 (N_7737,N_7640,N_7684);
and U7738 (N_7738,N_7669,N_7698);
nand U7739 (N_7739,N_7654,N_7692);
or U7740 (N_7740,N_7691,N_7609);
and U7741 (N_7741,N_7632,N_7687);
nand U7742 (N_7742,N_7606,N_7685);
or U7743 (N_7743,N_7666,N_7676);
or U7744 (N_7744,N_7643,N_7699);
nand U7745 (N_7745,N_7611,N_7624);
nand U7746 (N_7746,N_7627,N_7662);
or U7747 (N_7747,N_7638,N_7658);
and U7748 (N_7748,N_7613,N_7693);
nand U7749 (N_7749,N_7686,N_7644);
nor U7750 (N_7750,N_7649,N_7625);
or U7751 (N_7751,N_7661,N_7603);
and U7752 (N_7752,N_7652,N_7640);
or U7753 (N_7753,N_7606,N_7617);
or U7754 (N_7754,N_7648,N_7666);
nand U7755 (N_7755,N_7642,N_7683);
and U7756 (N_7756,N_7614,N_7608);
nor U7757 (N_7757,N_7668,N_7643);
or U7758 (N_7758,N_7659,N_7648);
xor U7759 (N_7759,N_7626,N_7645);
nor U7760 (N_7760,N_7674,N_7669);
or U7761 (N_7761,N_7665,N_7669);
or U7762 (N_7762,N_7685,N_7621);
and U7763 (N_7763,N_7634,N_7610);
nand U7764 (N_7764,N_7654,N_7670);
and U7765 (N_7765,N_7692,N_7679);
nand U7766 (N_7766,N_7671,N_7623);
nor U7767 (N_7767,N_7647,N_7616);
and U7768 (N_7768,N_7639,N_7607);
nor U7769 (N_7769,N_7620,N_7659);
nand U7770 (N_7770,N_7668,N_7656);
xnor U7771 (N_7771,N_7682,N_7691);
or U7772 (N_7772,N_7698,N_7601);
nor U7773 (N_7773,N_7608,N_7672);
and U7774 (N_7774,N_7684,N_7679);
or U7775 (N_7775,N_7655,N_7650);
nor U7776 (N_7776,N_7625,N_7653);
or U7777 (N_7777,N_7647,N_7672);
and U7778 (N_7778,N_7641,N_7632);
nand U7779 (N_7779,N_7671,N_7658);
nor U7780 (N_7780,N_7609,N_7672);
or U7781 (N_7781,N_7694,N_7660);
nor U7782 (N_7782,N_7621,N_7678);
or U7783 (N_7783,N_7616,N_7613);
nand U7784 (N_7784,N_7688,N_7618);
nor U7785 (N_7785,N_7656,N_7657);
nand U7786 (N_7786,N_7602,N_7646);
nand U7787 (N_7787,N_7676,N_7640);
or U7788 (N_7788,N_7677,N_7603);
nor U7789 (N_7789,N_7692,N_7689);
nor U7790 (N_7790,N_7609,N_7688);
nand U7791 (N_7791,N_7685,N_7651);
and U7792 (N_7792,N_7681,N_7687);
nor U7793 (N_7793,N_7668,N_7679);
or U7794 (N_7794,N_7653,N_7665);
and U7795 (N_7795,N_7664,N_7657);
and U7796 (N_7796,N_7666,N_7652);
or U7797 (N_7797,N_7631,N_7699);
or U7798 (N_7798,N_7690,N_7697);
or U7799 (N_7799,N_7609,N_7664);
nand U7800 (N_7800,N_7743,N_7739);
nand U7801 (N_7801,N_7703,N_7781);
nand U7802 (N_7802,N_7791,N_7758);
nand U7803 (N_7803,N_7760,N_7799);
nor U7804 (N_7804,N_7735,N_7785);
or U7805 (N_7805,N_7746,N_7777);
and U7806 (N_7806,N_7779,N_7794);
nor U7807 (N_7807,N_7723,N_7786);
or U7808 (N_7808,N_7714,N_7789);
nor U7809 (N_7809,N_7783,N_7795);
nand U7810 (N_7810,N_7768,N_7774);
xor U7811 (N_7811,N_7793,N_7763);
nor U7812 (N_7812,N_7749,N_7790);
and U7813 (N_7813,N_7745,N_7796);
or U7814 (N_7814,N_7771,N_7737);
and U7815 (N_7815,N_7788,N_7766);
nand U7816 (N_7816,N_7761,N_7759);
xor U7817 (N_7817,N_7778,N_7754);
or U7818 (N_7818,N_7787,N_7712);
nand U7819 (N_7819,N_7770,N_7702);
nand U7820 (N_7820,N_7773,N_7717);
nor U7821 (N_7821,N_7757,N_7715);
nand U7822 (N_7822,N_7742,N_7730);
and U7823 (N_7823,N_7764,N_7744);
or U7824 (N_7824,N_7726,N_7767);
nand U7825 (N_7825,N_7747,N_7710);
nor U7826 (N_7826,N_7751,N_7748);
nand U7827 (N_7827,N_7755,N_7727);
nor U7828 (N_7828,N_7716,N_7784);
or U7829 (N_7829,N_7797,N_7750);
nor U7830 (N_7830,N_7708,N_7772);
or U7831 (N_7831,N_7792,N_7740);
and U7832 (N_7832,N_7706,N_7701);
or U7833 (N_7833,N_7752,N_7769);
or U7834 (N_7834,N_7725,N_7731);
and U7835 (N_7835,N_7728,N_7718);
xnor U7836 (N_7836,N_7782,N_7705);
nor U7837 (N_7837,N_7709,N_7734);
nor U7838 (N_7838,N_7721,N_7776);
nor U7839 (N_7839,N_7780,N_7765);
nand U7840 (N_7840,N_7775,N_7713);
or U7841 (N_7841,N_7719,N_7733);
nor U7842 (N_7842,N_7707,N_7729);
or U7843 (N_7843,N_7741,N_7753);
and U7844 (N_7844,N_7700,N_7724);
nor U7845 (N_7845,N_7762,N_7736);
nor U7846 (N_7846,N_7720,N_7732);
or U7847 (N_7847,N_7704,N_7798);
nand U7848 (N_7848,N_7756,N_7711);
or U7849 (N_7849,N_7722,N_7738);
nand U7850 (N_7850,N_7703,N_7723);
nor U7851 (N_7851,N_7796,N_7737);
and U7852 (N_7852,N_7777,N_7794);
or U7853 (N_7853,N_7703,N_7785);
nand U7854 (N_7854,N_7769,N_7722);
or U7855 (N_7855,N_7793,N_7798);
nor U7856 (N_7856,N_7739,N_7738);
and U7857 (N_7857,N_7753,N_7728);
and U7858 (N_7858,N_7784,N_7772);
and U7859 (N_7859,N_7706,N_7735);
and U7860 (N_7860,N_7761,N_7702);
nor U7861 (N_7861,N_7707,N_7702);
or U7862 (N_7862,N_7738,N_7716);
nor U7863 (N_7863,N_7794,N_7784);
nand U7864 (N_7864,N_7701,N_7747);
nor U7865 (N_7865,N_7767,N_7748);
or U7866 (N_7866,N_7741,N_7779);
nand U7867 (N_7867,N_7753,N_7720);
nor U7868 (N_7868,N_7759,N_7779);
or U7869 (N_7869,N_7788,N_7723);
nand U7870 (N_7870,N_7734,N_7723);
and U7871 (N_7871,N_7713,N_7784);
and U7872 (N_7872,N_7747,N_7729);
or U7873 (N_7873,N_7702,N_7717);
nor U7874 (N_7874,N_7755,N_7731);
nand U7875 (N_7875,N_7773,N_7785);
and U7876 (N_7876,N_7759,N_7758);
and U7877 (N_7877,N_7725,N_7718);
nor U7878 (N_7878,N_7744,N_7704);
or U7879 (N_7879,N_7765,N_7796);
nand U7880 (N_7880,N_7723,N_7727);
nor U7881 (N_7881,N_7744,N_7728);
nor U7882 (N_7882,N_7726,N_7717);
or U7883 (N_7883,N_7733,N_7747);
nand U7884 (N_7884,N_7744,N_7738);
and U7885 (N_7885,N_7727,N_7749);
and U7886 (N_7886,N_7704,N_7792);
or U7887 (N_7887,N_7703,N_7736);
xor U7888 (N_7888,N_7776,N_7750);
or U7889 (N_7889,N_7711,N_7738);
nor U7890 (N_7890,N_7751,N_7704);
and U7891 (N_7891,N_7700,N_7788);
nand U7892 (N_7892,N_7765,N_7737);
and U7893 (N_7893,N_7752,N_7777);
nand U7894 (N_7894,N_7737,N_7720);
and U7895 (N_7895,N_7701,N_7744);
and U7896 (N_7896,N_7709,N_7774);
nand U7897 (N_7897,N_7745,N_7731);
or U7898 (N_7898,N_7714,N_7740);
and U7899 (N_7899,N_7785,N_7725);
nor U7900 (N_7900,N_7819,N_7824);
nand U7901 (N_7901,N_7825,N_7837);
or U7902 (N_7902,N_7831,N_7810);
or U7903 (N_7903,N_7861,N_7807);
or U7904 (N_7904,N_7851,N_7879);
nor U7905 (N_7905,N_7880,N_7853);
or U7906 (N_7906,N_7863,N_7806);
or U7907 (N_7907,N_7892,N_7897);
or U7908 (N_7908,N_7842,N_7833);
or U7909 (N_7909,N_7894,N_7809);
nand U7910 (N_7910,N_7827,N_7848);
nor U7911 (N_7911,N_7822,N_7813);
and U7912 (N_7912,N_7801,N_7899);
nand U7913 (N_7913,N_7875,N_7828);
or U7914 (N_7914,N_7855,N_7852);
xnor U7915 (N_7915,N_7817,N_7808);
nor U7916 (N_7916,N_7839,N_7834);
or U7917 (N_7917,N_7846,N_7847);
and U7918 (N_7918,N_7886,N_7877);
nor U7919 (N_7919,N_7874,N_7845);
nor U7920 (N_7920,N_7812,N_7849);
nand U7921 (N_7921,N_7838,N_7805);
nor U7922 (N_7922,N_7882,N_7815);
nor U7923 (N_7923,N_7829,N_7864);
and U7924 (N_7924,N_7866,N_7878);
nor U7925 (N_7925,N_7865,N_7890);
and U7926 (N_7926,N_7803,N_7800);
nand U7927 (N_7927,N_7873,N_7844);
nor U7928 (N_7928,N_7891,N_7835);
nand U7929 (N_7929,N_7830,N_7859);
nand U7930 (N_7930,N_7883,N_7836);
and U7931 (N_7931,N_7881,N_7854);
nor U7932 (N_7932,N_7898,N_7816);
nor U7933 (N_7933,N_7887,N_7811);
xor U7934 (N_7934,N_7870,N_7889);
or U7935 (N_7935,N_7841,N_7820);
nand U7936 (N_7936,N_7862,N_7867);
nand U7937 (N_7937,N_7857,N_7868);
or U7938 (N_7938,N_7821,N_7823);
nand U7939 (N_7939,N_7826,N_7876);
or U7940 (N_7940,N_7832,N_7871);
nor U7941 (N_7941,N_7818,N_7884);
and U7942 (N_7942,N_7840,N_7856);
and U7943 (N_7943,N_7895,N_7802);
or U7944 (N_7944,N_7869,N_7896);
and U7945 (N_7945,N_7850,N_7843);
nor U7946 (N_7946,N_7804,N_7893);
nand U7947 (N_7947,N_7860,N_7814);
nand U7948 (N_7948,N_7888,N_7885);
or U7949 (N_7949,N_7872,N_7858);
and U7950 (N_7950,N_7865,N_7805);
nor U7951 (N_7951,N_7814,N_7882);
or U7952 (N_7952,N_7895,N_7804);
and U7953 (N_7953,N_7869,N_7858);
xor U7954 (N_7954,N_7877,N_7841);
nand U7955 (N_7955,N_7862,N_7850);
nor U7956 (N_7956,N_7803,N_7818);
and U7957 (N_7957,N_7857,N_7809);
nor U7958 (N_7958,N_7849,N_7828);
and U7959 (N_7959,N_7842,N_7804);
or U7960 (N_7960,N_7852,N_7810);
and U7961 (N_7961,N_7869,N_7890);
nand U7962 (N_7962,N_7820,N_7876);
or U7963 (N_7963,N_7828,N_7880);
nand U7964 (N_7964,N_7812,N_7889);
nor U7965 (N_7965,N_7824,N_7896);
or U7966 (N_7966,N_7884,N_7885);
nor U7967 (N_7967,N_7845,N_7856);
nand U7968 (N_7968,N_7855,N_7801);
nor U7969 (N_7969,N_7832,N_7869);
and U7970 (N_7970,N_7835,N_7873);
and U7971 (N_7971,N_7896,N_7860);
or U7972 (N_7972,N_7885,N_7873);
and U7973 (N_7973,N_7803,N_7896);
nor U7974 (N_7974,N_7831,N_7888);
or U7975 (N_7975,N_7886,N_7817);
nand U7976 (N_7976,N_7876,N_7812);
nor U7977 (N_7977,N_7800,N_7844);
nor U7978 (N_7978,N_7803,N_7801);
and U7979 (N_7979,N_7870,N_7863);
and U7980 (N_7980,N_7800,N_7883);
and U7981 (N_7981,N_7830,N_7833);
or U7982 (N_7982,N_7805,N_7826);
nand U7983 (N_7983,N_7866,N_7856);
nor U7984 (N_7984,N_7849,N_7866);
nor U7985 (N_7985,N_7826,N_7862);
or U7986 (N_7986,N_7897,N_7832);
nand U7987 (N_7987,N_7888,N_7816);
and U7988 (N_7988,N_7807,N_7806);
or U7989 (N_7989,N_7893,N_7884);
and U7990 (N_7990,N_7811,N_7851);
nor U7991 (N_7991,N_7859,N_7838);
nand U7992 (N_7992,N_7875,N_7894);
or U7993 (N_7993,N_7830,N_7823);
xnor U7994 (N_7994,N_7840,N_7804);
or U7995 (N_7995,N_7871,N_7883);
nand U7996 (N_7996,N_7803,N_7846);
or U7997 (N_7997,N_7825,N_7809);
nor U7998 (N_7998,N_7891,N_7865);
or U7999 (N_7999,N_7874,N_7889);
nor U8000 (N_8000,N_7927,N_7937);
nor U8001 (N_8001,N_7974,N_7998);
nor U8002 (N_8002,N_7906,N_7915);
nor U8003 (N_8003,N_7938,N_7908);
and U8004 (N_8004,N_7920,N_7980);
nor U8005 (N_8005,N_7971,N_7921);
or U8006 (N_8006,N_7918,N_7934);
nor U8007 (N_8007,N_7995,N_7994);
nor U8008 (N_8008,N_7904,N_7932);
or U8009 (N_8009,N_7956,N_7999);
nand U8010 (N_8010,N_7977,N_7954);
and U8011 (N_8011,N_7943,N_7953);
nand U8012 (N_8012,N_7973,N_7946);
or U8013 (N_8013,N_7901,N_7947);
nand U8014 (N_8014,N_7933,N_7982);
and U8015 (N_8015,N_7923,N_7996);
or U8016 (N_8016,N_7991,N_7959);
and U8017 (N_8017,N_7990,N_7986);
and U8018 (N_8018,N_7931,N_7910);
nor U8019 (N_8019,N_7936,N_7919);
nor U8020 (N_8020,N_7914,N_7961);
and U8021 (N_8021,N_7963,N_7922);
nor U8022 (N_8022,N_7968,N_7952);
or U8023 (N_8023,N_7907,N_7926);
nor U8024 (N_8024,N_7960,N_7972);
nor U8025 (N_8025,N_7979,N_7924);
nand U8026 (N_8026,N_7981,N_7966);
or U8027 (N_8027,N_7987,N_7942);
and U8028 (N_8028,N_7916,N_7917);
and U8029 (N_8029,N_7935,N_7902);
and U8030 (N_8030,N_7985,N_7984);
or U8031 (N_8031,N_7929,N_7993);
nand U8032 (N_8032,N_7989,N_7925);
nand U8033 (N_8033,N_7905,N_7939);
or U8034 (N_8034,N_7913,N_7957);
and U8035 (N_8035,N_7912,N_7951);
nand U8036 (N_8036,N_7909,N_7962);
or U8037 (N_8037,N_7941,N_7940);
nand U8038 (N_8038,N_7955,N_7976);
nand U8039 (N_8039,N_7948,N_7969);
nand U8040 (N_8040,N_7997,N_7970);
or U8041 (N_8041,N_7958,N_7964);
and U8042 (N_8042,N_7950,N_7944);
and U8043 (N_8043,N_7988,N_7911);
nor U8044 (N_8044,N_7967,N_7965);
and U8045 (N_8045,N_7992,N_7930);
nor U8046 (N_8046,N_7900,N_7945);
nand U8047 (N_8047,N_7975,N_7978);
nand U8048 (N_8048,N_7949,N_7983);
nand U8049 (N_8049,N_7928,N_7903);
nor U8050 (N_8050,N_7992,N_7978);
and U8051 (N_8051,N_7983,N_7921);
or U8052 (N_8052,N_7962,N_7960);
or U8053 (N_8053,N_7921,N_7907);
nor U8054 (N_8054,N_7988,N_7924);
nor U8055 (N_8055,N_7953,N_7983);
or U8056 (N_8056,N_7959,N_7967);
nand U8057 (N_8057,N_7940,N_7993);
and U8058 (N_8058,N_7902,N_7922);
nor U8059 (N_8059,N_7944,N_7943);
and U8060 (N_8060,N_7957,N_7958);
or U8061 (N_8061,N_7936,N_7948);
and U8062 (N_8062,N_7990,N_7931);
nor U8063 (N_8063,N_7956,N_7976);
and U8064 (N_8064,N_7973,N_7948);
or U8065 (N_8065,N_7946,N_7914);
nand U8066 (N_8066,N_7922,N_7961);
nor U8067 (N_8067,N_7958,N_7902);
or U8068 (N_8068,N_7918,N_7955);
nand U8069 (N_8069,N_7901,N_7937);
nand U8070 (N_8070,N_7995,N_7909);
nand U8071 (N_8071,N_7958,N_7904);
and U8072 (N_8072,N_7924,N_7937);
nand U8073 (N_8073,N_7935,N_7944);
nor U8074 (N_8074,N_7901,N_7955);
or U8075 (N_8075,N_7984,N_7995);
nor U8076 (N_8076,N_7979,N_7915);
or U8077 (N_8077,N_7994,N_7955);
nor U8078 (N_8078,N_7978,N_7901);
nand U8079 (N_8079,N_7906,N_7914);
nand U8080 (N_8080,N_7961,N_7978);
nor U8081 (N_8081,N_7935,N_7963);
and U8082 (N_8082,N_7925,N_7901);
nand U8083 (N_8083,N_7958,N_7975);
nor U8084 (N_8084,N_7915,N_7949);
and U8085 (N_8085,N_7973,N_7949);
nand U8086 (N_8086,N_7910,N_7960);
and U8087 (N_8087,N_7941,N_7976);
nor U8088 (N_8088,N_7984,N_7999);
nor U8089 (N_8089,N_7973,N_7951);
or U8090 (N_8090,N_7964,N_7994);
nand U8091 (N_8091,N_7941,N_7981);
and U8092 (N_8092,N_7957,N_7949);
nand U8093 (N_8093,N_7911,N_7973);
nand U8094 (N_8094,N_7902,N_7918);
nor U8095 (N_8095,N_7966,N_7994);
nand U8096 (N_8096,N_7964,N_7949);
nand U8097 (N_8097,N_7920,N_7931);
and U8098 (N_8098,N_7950,N_7977);
nand U8099 (N_8099,N_7936,N_7911);
or U8100 (N_8100,N_8053,N_8072);
or U8101 (N_8101,N_8063,N_8003);
nor U8102 (N_8102,N_8029,N_8020);
or U8103 (N_8103,N_8056,N_8070);
nand U8104 (N_8104,N_8077,N_8092);
nor U8105 (N_8105,N_8022,N_8016);
and U8106 (N_8106,N_8066,N_8019);
and U8107 (N_8107,N_8098,N_8034);
nand U8108 (N_8108,N_8046,N_8049);
or U8109 (N_8109,N_8050,N_8083);
or U8110 (N_8110,N_8051,N_8075);
nand U8111 (N_8111,N_8018,N_8027);
nor U8112 (N_8112,N_8073,N_8011);
nand U8113 (N_8113,N_8060,N_8064);
and U8114 (N_8114,N_8091,N_8086);
nor U8115 (N_8115,N_8094,N_8031);
nand U8116 (N_8116,N_8052,N_8026);
or U8117 (N_8117,N_8039,N_8041);
and U8118 (N_8118,N_8024,N_8081);
and U8119 (N_8119,N_8061,N_8028);
or U8120 (N_8120,N_8036,N_8042);
nor U8121 (N_8121,N_8000,N_8032);
and U8122 (N_8122,N_8005,N_8067);
and U8123 (N_8123,N_8084,N_8059);
nor U8124 (N_8124,N_8082,N_8078);
and U8125 (N_8125,N_8096,N_8030);
nand U8126 (N_8126,N_8047,N_8058);
nand U8127 (N_8127,N_8085,N_8001);
or U8128 (N_8128,N_8045,N_8089);
nor U8129 (N_8129,N_8044,N_8015);
nand U8130 (N_8130,N_8040,N_8037);
nor U8131 (N_8131,N_8057,N_8069);
xor U8132 (N_8132,N_8076,N_8055);
or U8133 (N_8133,N_8074,N_8048);
and U8134 (N_8134,N_8087,N_8002);
and U8135 (N_8135,N_8021,N_8080);
and U8136 (N_8136,N_8065,N_8035);
or U8137 (N_8137,N_8004,N_8099);
or U8138 (N_8138,N_8008,N_8013);
and U8139 (N_8139,N_8007,N_8068);
and U8140 (N_8140,N_8071,N_8088);
xor U8141 (N_8141,N_8014,N_8090);
and U8142 (N_8142,N_8017,N_8010);
nor U8143 (N_8143,N_8009,N_8038);
nand U8144 (N_8144,N_8054,N_8093);
nor U8145 (N_8145,N_8097,N_8062);
nor U8146 (N_8146,N_8012,N_8095);
xor U8147 (N_8147,N_8079,N_8043);
and U8148 (N_8148,N_8025,N_8006);
or U8149 (N_8149,N_8023,N_8033);
nor U8150 (N_8150,N_8070,N_8043);
nand U8151 (N_8151,N_8001,N_8051);
or U8152 (N_8152,N_8001,N_8043);
or U8153 (N_8153,N_8035,N_8072);
nor U8154 (N_8154,N_8052,N_8093);
and U8155 (N_8155,N_8011,N_8031);
and U8156 (N_8156,N_8046,N_8069);
and U8157 (N_8157,N_8058,N_8054);
nor U8158 (N_8158,N_8021,N_8083);
and U8159 (N_8159,N_8039,N_8006);
or U8160 (N_8160,N_8022,N_8021);
or U8161 (N_8161,N_8078,N_8075);
nand U8162 (N_8162,N_8019,N_8095);
or U8163 (N_8163,N_8036,N_8016);
nor U8164 (N_8164,N_8014,N_8018);
nor U8165 (N_8165,N_8045,N_8004);
nand U8166 (N_8166,N_8043,N_8055);
and U8167 (N_8167,N_8067,N_8064);
and U8168 (N_8168,N_8049,N_8033);
and U8169 (N_8169,N_8024,N_8048);
nor U8170 (N_8170,N_8046,N_8070);
and U8171 (N_8171,N_8098,N_8056);
and U8172 (N_8172,N_8087,N_8013);
and U8173 (N_8173,N_8052,N_8008);
nor U8174 (N_8174,N_8036,N_8021);
nand U8175 (N_8175,N_8005,N_8093);
nor U8176 (N_8176,N_8010,N_8028);
nand U8177 (N_8177,N_8063,N_8065);
or U8178 (N_8178,N_8078,N_8088);
nand U8179 (N_8179,N_8006,N_8071);
nor U8180 (N_8180,N_8020,N_8083);
and U8181 (N_8181,N_8090,N_8045);
xor U8182 (N_8182,N_8077,N_8097);
or U8183 (N_8183,N_8072,N_8038);
nor U8184 (N_8184,N_8071,N_8078);
and U8185 (N_8185,N_8057,N_8097);
and U8186 (N_8186,N_8036,N_8032);
nand U8187 (N_8187,N_8032,N_8092);
nand U8188 (N_8188,N_8034,N_8011);
or U8189 (N_8189,N_8014,N_8077);
and U8190 (N_8190,N_8078,N_8054);
nand U8191 (N_8191,N_8041,N_8035);
and U8192 (N_8192,N_8070,N_8080);
nand U8193 (N_8193,N_8059,N_8018);
and U8194 (N_8194,N_8035,N_8037);
nor U8195 (N_8195,N_8042,N_8053);
and U8196 (N_8196,N_8002,N_8003);
nand U8197 (N_8197,N_8026,N_8067);
nor U8198 (N_8198,N_8033,N_8008);
nand U8199 (N_8199,N_8024,N_8006);
or U8200 (N_8200,N_8136,N_8113);
or U8201 (N_8201,N_8166,N_8159);
nor U8202 (N_8202,N_8141,N_8198);
and U8203 (N_8203,N_8144,N_8178);
and U8204 (N_8204,N_8158,N_8139);
nand U8205 (N_8205,N_8101,N_8116);
or U8206 (N_8206,N_8138,N_8172);
nand U8207 (N_8207,N_8142,N_8102);
nand U8208 (N_8208,N_8130,N_8109);
and U8209 (N_8209,N_8192,N_8191);
and U8210 (N_8210,N_8104,N_8149);
nand U8211 (N_8211,N_8131,N_8157);
nand U8212 (N_8212,N_8134,N_8148);
nand U8213 (N_8213,N_8193,N_8133);
and U8214 (N_8214,N_8169,N_8185);
nor U8215 (N_8215,N_8161,N_8145);
nand U8216 (N_8216,N_8183,N_8160);
or U8217 (N_8217,N_8124,N_8187);
nand U8218 (N_8218,N_8117,N_8128);
or U8219 (N_8219,N_8107,N_8125);
nor U8220 (N_8220,N_8188,N_8171);
nor U8221 (N_8221,N_8112,N_8103);
xnor U8222 (N_8222,N_8162,N_8174);
nor U8223 (N_8223,N_8184,N_8170);
nand U8224 (N_8224,N_8180,N_8110);
nand U8225 (N_8225,N_8115,N_8190);
nand U8226 (N_8226,N_8147,N_8155);
nand U8227 (N_8227,N_8123,N_8122);
nand U8228 (N_8228,N_8175,N_8181);
and U8229 (N_8229,N_8150,N_8196);
and U8230 (N_8230,N_8120,N_8164);
and U8231 (N_8231,N_8167,N_8197);
nor U8232 (N_8232,N_8176,N_8189);
nand U8233 (N_8233,N_8151,N_8106);
xnor U8234 (N_8234,N_8119,N_8127);
or U8235 (N_8235,N_8177,N_8152);
nand U8236 (N_8236,N_8114,N_8195);
nor U8237 (N_8237,N_8168,N_8121);
nor U8238 (N_8238,N_8137,N_8126);
nor U8239 (N_8239,N_8146,N_8173);
and U8240 (N_8240,N_8111,N_8182);
or U8241 (N_8241,N_8154,N_8199);
nand U8242 (N_8242,N_8108,N_8186);
and U8243 (N_8243,N_8140,N_8179);
nor U8244 (N_8244,N_8156,N_8194);
nand U8245 (N_8245,N_8132,N_8163);
or U8246 (N_8246,N_8165,N_8129);
nor U8247 (N_8247,N_8105,N_8118);
or U8248 (N_8248,N_8143,N_8135);
nand U8249 (N_8249,N_8100,N_8153);
and U8250 (N_8250,N_8119,N_8139);
or U8251 (N_8251,N_8135,N_8196);
or U8252 (N_8252,N_8143,N_8194);
and U8253 (N_8253,N_8170,N_8122);
and U8254 (N_8254,N_8106,N_8160);
or U8255 (N_8255,N_8117,N_8138);
and U8256 (N_8256,N_8133,N_8113);
or U8257 (N_8257,N_8112,N_8116);
nand U8258 (N_8258,N_8196,N_8141);
and U8259 (N_8259,N_8157,N_8121);
nand U8260 (N_8260,N_8178,N_8117);
nand U8261 (N_8261,N_8194,N_8159);
or U8262 (N_8262,N_8164,N_8165);
and U8263 (N_8263,N_8155,N_8108);
nor U8264 (N_8264,N_8155,N_8189);
nor U8265 (N_8265,N_8124,N_8151);
and U8266 (N_8266,N_8105,N_8141);
and U8267 (N_8267,N_8146,N_8136);
nand U8268 (N_8268,N_8179,N_8194);
or U8269 (N_8269,N_8121,N_8138);
and U8270 (N_8270,N_8118,N_8102);
xnor U8271 (N_8271,N_8141,N_8108);
or U8272 (N_8272,N_8187,N_8132);
nor U8273 (N_8273,N_8116,N_8104);
and U8274 (N_8274,N_8122,N_8194);
nand U8275 (N_8275,N_8136,N_8186);
nand U8276 (N_8276,N_8146,N_8159);
nand U8277 (N_8277,N_8134,N_8185);
nand U8278 (N_8278,N_8193,N_8111);
and U8279 (N_8279,N_8141,N_8125);
and U8280 (N_8280,N_8145,N_8112);
and U8281 (N_8281,N_8150,N_8191);
and U8282 (N_8282,N_8104,N_8191);
nand U8283 (N_8283,N_8195,N_8158);
nand U8284 (N_8284,N_8120,N_8165);
or U8285 (N_8285,N_8128,N_8142);
nor U8286 (N_8286,N_8168,N_8188);
nand U8287 (N_8287,N_8112,N_8110);
and U8288 (N_8288,N_8122,N_8181);
nand U8289 (N_8289,N_8168,N_8119);
nand U8290 (N_8290,N_8100,N_8104);
and U8291 (N_8291,N_8152,N_8109);
and U8292 (N_8292,N_8142,N_8110);
nand U8293 (N_8293,N_8177,N_8121);
and U8294 (N_8294,N_8154,N_8130);
or U8295 (N_8295,N_8140,N_8129);
nand U8296 (N_8296,N_8162,N_8116);
nand U8297 (N_8297,N_8164,N_8176);
nand U8298 (N_8298,N_8138,N_8148);
and U8299 (N_8299,N_8121,N_8150);
or U8300 (N_8300,N_8295,N_8206);
and U8301 (N_8301,N_8246,N_8228);
and U8302 (N_8302,N_8248,N_8265);
and U8303 (N_8303,N_8261,N_8217);
or U8304 (N_8304,N_8288,N_8278);
or U8305 (N_8305,N_8290,N_8291);
or U8306 (N_8306,N_8255,N_8238);
or U8307 (N_8307,N_8233,N_8226);
nand U8308 (N_8308,N_8254,N_8281);
and U8309 (N_8309,N_8235,N_8214);
nor U8310 (N_8310,N_8285,N_8280);
or U8311 (N_8311,N_8251,N_8245);
nand U8312 (N_8312,N_8256,N_8283);
or U8313 (N_8313,N_8225,N_8216);
nor U8314 (N_8314,N_8211,N_8207);
or U8315 (N_8315,N_8298,N_8260);
nor U8316 (N_8316,N_8215,N_8271);
nor U8317 (N_8317,N_8275,N_8209);
nor U8318 (N_8318,N_8272,N_8223);
nand U8319 (N_8319,N_8230,N_8262);
or U8320 (N_8320,N_8244,N_8289);
xnor U8321 (N_8321,N_8284,N_8222);
nor U8322 (N_8322,N_8240,N_8210);
and U8323 (N_8323,N_8270,N_8220);
nor U8324 (N_8324,N_8286,N_8218);
nor U8325 (N_8325,N_8227,N_8257);
nand U8326 (N_8326,N_8294,N_8293);
and U8327 (N_8327,N_8297,N_8279);
and U8328 (N_8328,N_8202,N_8247);
nand U8329 (N_8329,N_8231,N_8243);
nand U8330 (N_8330,N_8269,N_8208);
nor U8331 (N_8331,N_8236,N_8258);
nand U8332 (N_8332,N_8229,N_8237);
nand U8333 (N_8333,N_8282,N_8259);
and U8334 (N_8334,N_8299,N_8212);
or U8335 (N_8335,N_8250,N_8204);
or U8336 (N_8336,N_8292,N_8200);
or U8337 (N_8337,N_8224,N_8249);
or U8338 (N_8338,N_8268,N_8273);
or U8339 (N_8339,N_8234,N_8276);
nor U8340 (N_8340,N_8203,N_8213);
and U8341 (N_8341,N_8267,N_8219);
or U8342 (N_8342,N_8242,N_8266);
nand U8343 (N_8343,N_8274,N_8253);
nand U8344 (N_8344,N_8287,N_8232);
or U8345 (N_8345,N_8201,N_8221);
or U8346 (N_8346,N_8252,N_8263);
nand U8347 (N_8347,N_8239,N_8205);
nand U8348 (N_8348,N_8277,N_8241);
and U8349 (N_8349,N_8264,N_8296);
nand U8350 (N_8350,N_8205,N_8222);
nand U8351 (N_8351,N_8255,N_8224);
and U8352 (N_8352,N_8258,N_8205);
or U8353 (N_8353,N_8262,N_8294);
nor U8354 (N_8354,N_8278,N_8226);
and U8355 (N_8355,N_8266,N_8298);
xnor U8356 (N_8356,N_8286,N_8235);
nor U8357 (N_8357,N_8266,N_8293);
and U8358 (N_8358,N_8231,N_8236);
and U8359 (N_8359,N_8251,N_8296);
and U8360 (N_8360,N_8222,N_8230);
nor U8361 (N_8361,N_8285,N_8251);
nand U8362 (N_8362,N_8245,N_8225);
and U8363 (N_8363,N_8287,N_8220);
or U8364 (N_8364,N_8239,N_8202);
nor U8365 (N_8365,N_8218,N_8261);
nand U8366 (N_8366,N_8209,N_8280);
and U8367 (N_8367,N_8275,N_8244);
xor U8368 (N_8368,N_8266,N_8213);
or U8369 (N_8369,N_8227,N_8261);
nor U8370 (N_8370,N_8281,N_8250);
and U8371 (N_8371,N_8287,N_8229);
and U8372 (N_8372,N_8292,N_8254);
nand U8373 (N_8373,N_8244,N_8220);
xor U8374 (N_8374,N_8204,N_8252);
nor U8375 (N_8375,N_8215,N_8238);
nor U8376 (N_8376,N_8224,N_8215);
and U8377 (N_8377,N_8244,N_8202);
nand U8378 (N_8378,N_8254,N_8213);
or U8379 (N_8379,N_8257,N_8259);
nand U8380 (N_8380,N_8288,N_8209);
nor U8381 (N_8381,N_8253,N_8217);
or U8382 (N_8382,N_8239,N_8229);
or U8383 (N_8383,N_8251,N_8207);
nand U8384 (N_8384,N_8232,N_8272);
nand U8385 (N_8385,N_8229,N_8231);
nand U8386 (N_8386,N_8281,N_8207);
nor U8387 (N_8387,N_8269,N_8264);
nor U8388 (N_8388,N_8220,N_8234);
or U8389 (N_8389,N_8200,N_8253);
nor U8390 (N_8390,N_8282,N_8204);
nor U8391 (N_8391,N_8269,N_8216);
and U8392 (N_8392,N_8297,N_8209);
nor U8393 (N_8393,N_8287,N_8293);
and U8394 (N_8394,N_8228,N_8208);
nand U8395 (N_8395,N_8206,N_8253);
nand U8396 (N_8396,N_8274,N_8232);
nor U8397 (N_8397,N_8246,N_8273);
nor U8398 (N_8398,N_8277,N_8256);
and U8399 (N_8399,N_8251,N_8284);
and U8400 (N_8400,N_8349,N_8386);
nor U8401 (N_8401,N_8359,N_8302);
nand U8402 (N_8402,N_8362,N_8305);
and U8403 (N_8403,N_8323,N_8365);
nand U8404 (N_8404,N_8354,N_8327);
and U8405 (N_8405,N_8363,N_8382);
nand U8406 (N_8406,N_8326,N_8311);
nor U8407 (N_8407,N_8330,N_8389);
nor U8408 (N_8408,N_8348,N_8338);
nor U8409 (N_8409,N_8336,N_8335);
xnor U8410 (N_8410,N_8345,N_8397);
xnor U8411 (N_8411,N_8391,N_8384);
nand U8412 (N_8412,N_8333,N_8399);
nor U8413 (N_8413,N_8317,N_8381);
nor U8414 (N_8414,N_8387,N_8321);
nand U8415 (N_8415,N_8377,N_8374);
nand U8416 (N_8416,N_8357,N_8315);
or U8417 (N_8417,N_8325,N_8319);
nor U8418 (N_8418,N_8383,N_8328);
and U8419 (N_8419,N_8300,N_8370);
and U8420 (N_8420,N_8392,N_8390);
nor U8421 (N_8421,N_8331,N_8395);
xor U8422 (N_8422,N_8343,N_8347);
and U8423 (N_8423,N_8356,N_8351);
nor U8424 (N_8424,N_8385,N_8316);
nor U8425 (N_8425,N_8307,N_8309);
nand U8426 (N_8426,N_8304,N_8310);
and U8427 (N_8427,N_8393,N_8380);
xnor U8428 (N_8428,N_8352,N_8366);
nand U8429 (N_8429,N_8346,N_8388);
or U8430 (N_8430,N_8313,N_8367);
and U8431 (N_8431,N_8364,N_8372);
nor U8432 (N_8432,N_8342,N_8337);
or U8433 (N_8433,N_8398,N_8340);
nand U8434 (N_8434,N_8332,N_8329);
and U8435 (N_8435,N_8312,N_8303);
or U8436 (N_8436,N_8318,N_8314);
nand U8437 (N_8437,N_8320,N_8324);
xnor U8438 (N_8438,N_8353,N_8339);
nand U8439 (N_8439,N_8396,N_8375);
or U8440 (N_8440,N_8369,N_8301);
nor U8441 (N_8441,N_8306,N_8379);
or U8442 (N_8442,N_8378,N_8376);
nor U8443 (N_8443,N_8334,N_8373);
nor U8444 (N_8444,N_8361,N_8360);
xnor U8445 (N_8445,N_8341,N_8344);
or U8446 (N_8446,N_8368,N_8394);
or U8447 (N_8447,N_8322,N_8350);
nand U8448 (N_8448,N_8308,N_8358);
and U8449 (N_8449,N_8371,N_8355);
and U8450 (N_8450,N_8390,N_8398);
nand U8451 (N_8451,N_8350,N_8348);
nand U8452 (N_8452,N_8357,N_8375);
or U8453 (N_8453,N_8327,N_8322);
nand U8454 (N_8454,N_8349,N_8324);
nor U8455 (N_8455,N_8307,N_8342);
xnor U8456 (N_8456,N_8333,N_8388);
and U8457 (N_8457,N_8370,N_8347);
nor U8458 (N_8458,N_8398,N_8311);
xor U8459 (N_8459,N_8343,N_8321);
and U8460 (N_8460,N_8342,N_8343);
or U8461 (N_8461,N_8329,N_8356);
or U8462 (N_8462,N_8334,N_8344);
or U8463 (N_8463,N_8347,N_8338);
nor U8464 (N_8464,N_8352,N_8320);
and U8465 (N_8465,N_8358,N_8304);
or U8466 (N_8466,N_8328,N_8342);
or U8467 (N_8467,N_8304,N_8342);
nor U8468 (N_8468,N_8359,N_8399);
nor U8469 (N_8469,N_8379,N_8351);
or U8470 (N_8470,N_8325,N_8336);
or U8471 (N_8471,N_8383,N_8358);
or U8472 (N_8472,N_8340,N_8359);
nand U8473 (N_8473,N_8374,N_8310);
and U8474 (N_8474,N_8383,N_8356);
nand U8475 (N_8475,N_8321,N_8397);
and U8476 (N_8476,N_8349,N_8325);
nand U8477 (N_8477,N_8317,N_8359);
nor U8478 (N_8478,N_8306,N_8392);
nand U8479 (N_8479,N_8326,N_8343);
nand U8480 (N_8480,N_8375,N_8376);
nand U8481 (N_8481,N_8365,N_8315);
nor U8482 (N_8482,N_8320,N_8361);
or U8483 (N_8483,N_8385,N_8338);
nor U8484 (N_8484,N_8393,N_8302);
nand U8485 (N_8485,N_8377,N_8365);
or U8486 (N_8486,N_8374,N_8330);
and U8487 (N_8487,N_8321,N_8339);
or U8488 (N_8488,N_8309,N_8340);
nand U8489 (N_8489,N_8385,N_8303);
nor U8490 (N_8490,N_8355,N_8352);
nor U8491 (N_8491,N_8308,N_8390);
and U8492 (N_8492,N_8318,N_8336);
nor U8493 (N_8493,N_8310,N_8340);
nor U8494 (N_8494,N_8339,N_8309);
or U8495 (N_8495,N_8374,N_8398);
nand U8496 (N_8496,N_8301,N_8353);
and U8497 (N_8497,N_8355,N_8347);
nor U8498 (N_8498,N_8385,N_8337);
nor U8499 (N_8499,N_8361,N_8376);
nand U8500 (N_8500,N_8491,N_8439);
and U8501 (N_8501,N_8463,N_8416);
nor U8502 (N_8502,N_8436,N_8482);
nor U8503 (N_8503,N_8479,N_8406);
nor U8504 (N_8504,N_8456,N_8475);
nor U8505 (N_8505,N_8454,N_8495);
or U8506 (N_8506,N_8401,N_8452);
nand U8507 (N_8507,N_8409,N_8499);
and U8508 (N_8508,N_8480,N_8498);
nor U8509 (N_8509,N_8451,N_8426);
or U8510 (N_8510,N_8432,N_8459);
nand U8511 (N_8511,N_8496,N_8472);
nand U8512 (N_8512,N_8407,N_8453);
nand U8513 (N_8513,N_8430,N_8490);
and U8514 (N_8514,N_8473,N_8469);
and U8515 (N_8515,N_8420,N_8467);
nand U8516 (N_8516,N_8444,N_8417);
or U8517 (N_8517,N_8429,N_8466);
or U8518 (N_8518,N_8489,N_8458);
or U8519 (N_8519,N_8457,N_8412);
nor U8520 (N_8520,N_8427,N_8421);
nand U8521 (N_8521,N_8435,N_8422);
nor U8522 (N_8522,N_8423,N_8419);
nand U8523 (N_8523,N_8424,N_8425);
and U8524 (N_8524,N_8470,N_8494);
nor U8525 (N_8525,N_8448,N_8474);
and U8526 (N_8526,N_8437,N_8487);
or U8527 (N_8527,N_8408,N_8450);
or U8528 (N_8528,N_8404,N_8477);
nand U8529 (N_8529,N_8400,N_8445);
nor U8530 (N_8530,N_8493,N_8485);
nor U8531 (N_8531,N_8414,N_8460);
and U8532 (N_8532,N_8433,N_8471);
nand U8533 (N_8533,N_8413,N_8465);
xor U8534 (N_8534,N_8405,N_8497);
and U8535 (N_8535,N_8481,N_8446);
nor U8536 (N_8536,N_8468,N_8441);
or U8537 (N_8537,N_8410,N_8440);
or U8538 (N_8538,N_8483,N_8449);
nand U8539 (N_8539,N_8431,N_8461);
or U8540 (N_8540,N_8488,N_8478);
nand U8541 (N_8541,N_8438,N_8486);
nand U8542 (N_8542,N_8403,N_8492);
nand U8543 (N_8543,N_8447,N_8434);
and U8544 (N_8544,N_8411,N_8442);
nand U8545 (N_8545,N_8415,N_8443);
nand U8546 (N_8546,N_8428,N_8402);
xnor U8547 (N_8547,N_8418,N_8464);
or U8548 (N_8548,N_8484,N_8455);
nor U8549 (N_8549,N_8476,N_8462);
nor U8550 (N_8550,N_8410,N_8454);
and U8551 (N_8551,N_8445,N_8448);
nand U8552 (N_8552,N_8442,N_8422);
nor U8553 (N_8553,N_8418,N_8487);
and U8554 (N_8554,N_8404,N_8463);
nor U8555 (N_8555,N_8402,N_8484);
and U8556 (N_8556,N_8489,N_8438);
xor U8557 (N_8557,N_8422,N_8430);
or U8558 (N_8558,N_8416,N_8400);
nand U8559 (N_8559,N_8465,N_8484);
nand U8560 (N_8560,N_8447,N_8402);
nor U8561 (N_8561,N_8474,N_8443);
and U8562 (N_8562,N_8430,N_8410);
nor U8563 (N_8563,N_8441,N_8407);
nor U8564 (N_8564,N_8466,N_8405);
nand U8565 (N_8565,N_8476,N_8465);
nand U8566 (N_8566,N_8447,N_8427);
and U8567 (N_8567,N_8406,N_8489);
nor U8568 (N_8568,N_8480,N_8406);
nor U8569 (N_8569,N_8469,N_8424);
and U8570 (N_8570,N_8435,N_8473);
nor U8571 (N_8571,N_8431,N_8465);
or U8572 (N_8572,N_8463,N_8441);
nand U8573 (N_8573,N_8495,N_8404);
nand U8574 (N_8574,N_8445,N_8411);
nor U8575 (N_8575,N_8428,N_8462);
or U8576 (N_8576,N_8446,N_8425);
nand U8577 (N_8577,N_8488,N_8410);
or U8578 (N_8578,N_8432,N_8426);
and U8579 (N_8579,N_8425,N_8481);
and U8580 (N_8580,N_8461,N_8406);
nor U8581 (N_8581,N_8408,N_8436);
nand U8582 (N_8582,N_8415,N_8499);
nand U8583 (N_8583,N_8400,N_8446);
or U8584 (N_8584,N_8412,N_8450);
and U8585 (N_8585,N_8445,N_8435);
nand U8586 (N_8586,N_8480,N_8487);
nand U8587 (N_8587,N_8410,N_8474);
and U8588 (N_8588,N_8479,N_8489);
nand U8589 (N_8589,N_8458,N_8496);
nand U8590 (N_8590,N_8452,N_8476);
nand U8591 (N_8591,N_8476,N_8454);
xnor U8592 (N_8592,N_8489,N_8421);
nor U8593 (N_8593,N_8477,N_8461);
or U8594 (N_8594,N_8410,N_8484);
nand U8595 (N_8595,N_8469,N_8453);
nand U8596 (N_8596,N_8480,N_8447);
nor U8597 (N_8597,N_8429,N_8481);
or U8598 (N_8598,N_8422,N_8494);
nor U8599 (N_8599,N_8491,N_8497);
nand U8600 (N_8600,N_8569,N_8590);
nand U8601 (N_8601,N_8517,N_8598);
and U8602 (N_8602,N_8538,N_8513);
nor U8603 (N_8603,N_8508,N_8545);
and U8604 (N_8604,N_8527,N_8580);
or U8605 (N_8605,N_8555,N_8522);
nor U8606 (N_8606,N_8574,N_8543);
nand U8607 (N_8607,N_8530,N_8525);
and U8608 (N_8608,N_8526,N_8529);
and U8609 (N_8609,N_8595,N_8503);
nand U8610 (N_8610,N_8592,N_8504);
or U8611 (N_8611,N_8509,N_8560);
or U8612 (N_8612,N_8581,N_8594);
nand U8613 (N_8613,N_8559,N_8553);
nand U8614 (N_8614,N_8516,N_8563);
nor U8615 (N_8615,N_8506,N_8505);
or U8616 (N_8616,N_8552,N_8501);
and U8617 (N_8617,N_8507,N_8584);
nand U8618 (N_8618,N_8524,N_8591);
nor U8619 (N_8619,N_8582,N_8568);
or U8620 (N_8620,N_8562,N_8533);
and U8621 (N_8621,N_8531,N_8572);
and U8622 (N_8622,N_8549,N_8589);
nand U8623 (N_8623,N_8587,N_8597);
nor U8624 (N_8624,N_8514,N_8532);
nor U8625 (N_8625,N_8518,N_8593);
nor U8626 (N_8626,N_8536,N_8539);
nor U8627 (N_8627,N_8565,N_8515);
and U8628 (N_8628,N_8547,N_8511);
or U8629 (N_8629,N_8567,N_8521);
nand U8630 (N_8630,N_8550,N_8558);
and U8631 (N_8631,N_8544,N_8556);
or U8632 (N_8632,N_8575,N_8523);
and U8633 (N_8633,N_8540,N_8546);
nor U8634 (N_8634,N_8519,N_8578);
or U8635 (N_8635,N_8510,N_8554);
nor U8636 (N_8636,N_8579,N_8500);
nand U8637 (N_8637,N_8588,N_8542);
nand U8638 (N_8638,N_8596,N_8561);
and U8639 (N_8639,N_8534,N_8586);
nand U8640 (N_8640,N_8576,N_8548);
or U8641 (N_8641,N_8541,N_8571);
nor U8642 (N_8642,N_8551,N_8564);
and U8643 (N_8643,N_8577,N_8502);
and U8644 (N_8644,N_8573,N_8566);
or U8645 (N_8645,N_8512,N_8599);
and U8646 (N_8646,N_8583,N_8570);
nor U8647 (N_8647,N_8520,N_8528);
nor U8648 (N_8648,N_8585,N_8537);
nor U8649 (N_8649,N_8557,N_8535);
nand U8650 (N_8650,N_8504,N_8549);
nand U8651 (N_8651,N_8523,N_8599);
or U8652 (N_8652,N_8580,N_8512);
or U8653 (N_8653,N_8543,N_8508);
nor U8654 (N_8654,N_8578,N_8570);
nor U8655 (N_8655,N_8522,N_8552);
and U8656 (N_8656,N_8503,N_8552);
and U8657 (N_8657,N_8583,N_8582);
or U8658 (N_8658,N_8556,N_8571);
nor U8659 (N_8659,N_8529,N_8542);
and U8660 (N_8660,N_8599,N_8538);
and U8661 (N_8661,N_8522,N_8537);
nor U8662 (N_8662,N_8594,N_8536);
or U8663 (N_8663,N_8566,N_8594);
or U8664 (N_8664,N_8558,N_8560);
nand U8665 (N_8665,N_8551,N_8508);
and U8666 (N_8666,N_8547,N_8516);
or U8667 (N_8667,N_8520,N_8512);
nor U8668 (N_8668,N_8569,N_8511);
nor U8669 (N_8669,N_8535,N_8504);
xnor U8670 (N_8670,N_8587,N_8586);
nand U8671 (N_8671,N_8545,N_8575);
nand U8672 (N_8672,N_8594,N_8578);
or U8673 (N_8673,N_8553,N_8520);
nand U8674 (N_8674,N_8549,N_8571);
and U8675 (N_8675,N_8596,N_8503);
nand U8676 (N_8676,N_8576,N_8588);
or U8677 (N_8677,N_8506,N_8580);
xnor U8678 (N_8678,N_8505,N_8504);
nand U8679 (N_8679,N_8532,N_8589);
and U8680 (N_8680,N_8537,N_8514);
or U8681 (N_8681,N_8571,N_8501);
or U8682 (N_8682,N_8525,N_8522);
nand U8683 (N_8683,N_8551,N_8568);
nor U8684 (N_8684,N_8539,N_8510);
nor U8685 (N_8685,N_8558,N_8583);
nand U8686 (N_8686,N_8520,N_8544);
or U8687 (N_8687,N_8544,N_8590);
nand U8688 (N_8688,N_8514,N_8574);
nor U8689 (N_8689,N_8538,N_8554);
and U8690 (N_8690,N_8542,N_8599);
or U8691 (N_8691,N_8521,N_8561);
xnor U8692 (N_8692,N_8591,N_8532);
or U8693 (N_8693,N_8578,N_8581);
nor U8694 (N_8694,N_8542,N_8512);
nand U8695 (N_8695,N_8504,N_8537);
or U8696 (N_8696,N_8589,N_8554);
and U8697 (N_8697,N_8537,N_8560);
or U8698 (N_8698,N_8528,N_8554);
nand U8699 (N_8699,N_8516,N_8566);
and U8700 (N_8700,N_8681,N_8641);
nand U8701 (N_8701,N_8691,N_8649);
or U8702 (N_8702,N_8615,N_8647);
or U8703 (N_8703,N_8621,N_8659);
nand U8704 (N_8704,N_8631,N_8673);
nand U8705 (N_8705,N_8657,N_8636);
nand U8706 (N_8706,N_8695,N_8697);
and U8707 (N_8707,N_8624,N_8613);
and U8708 (N_8708,N_8643,N_8686);
nand U8709 (N_8709,N_8611,N_8626);
nand U8710 (N_8710,N_8690,N_8646);
nor U8711 (N_8711,N_8692,N_8604);
and U8712 (N_8712,N_8635,N_8616);
nand U8713 (N_8713,N_8656,N_8637);
nand U8714 (N_8714,N_8655,N_8694);
or U8715 (N_8715,N_8628,N_8618);
nand U8716 (N_8716,N_8632,N_8672);
nand U8717 (N_8717,N_8670,N_8689);
nand U8718 (N_8718,N_8609,N_8660);
or U8719 (N_8719,N_8627,N_8696);
or U8720 (N_8720,N_8601,N_8612);
xnor U8721 (N_8721,N_8650,N_8625);
nor U8722 (N_8722,N_8607,N_8653);
nand U8723 (N_8723,N_8661,N_8684);
or U8724 (N_8724,N_8638,N_8619);
nor U8725 (N_8725,N_8663,N_8639);
and U8726 (N_8726,N_8668,N_8654);
and U8727 (N_8727,N_8633,N_8606);
or U8728 (N_8728,N_8687,N_8662);
or U8729 (N_8729,N_8630,N_8640);
or U8730 (N_8730,N_8685,N_8602);
nand U8731 (N_8731,N_8644,N_8680);
nand U8732 (N_8732,N_8671,N_8667);
nor U8733 (N_8733,N_8608,N_8675);
and U8734 (N_8734,N_8600,N_8665);
or U8735 (N_8735,N_8674,N_8629);
nand U8736 (N_8736,N_8610,N_8605);
and U8737 (N_8737,N_8683,N_8669);
nor U8738 (N_8738,N_8676,N_8658);
or U8739 (N_8739,N_8603,N_8693);
or U8740 (N_8740,N_8678,N_8622);
nand U8741 (N_8741,N_8645,N_8620);
nor U8742 (N_8742,N_8623,N_8617);
nor U8743 (N_8743,N_8688,N_8679);
or U8744 (N_8744,N_8648,N_8642);
nand U8745 (N_8745,N_8682,N_8652);
nor U8746 (N_8746,N_8677,N_8699);
nand U8747 (N_8747,N_8614,N_8664);
and U8748 (N_8748,N_8698,N_8634);
nand U8749 (N_8749,N_8651,N_8666);
or U8750 (N_8750,N_8640,N_8641);
or U8751 (N_8751,N_8694,N_8682);
or U8752 (N_8752,N_8632,N_8634);
or U8753 (N_8753,N_8670,N_8654);
or U8754 (N_8754,N_8623,N_8632);
and U8755 (N_8755,N_8641,N_8611);
and U8756 (N_8756,N_8617,N_8619);
nor U8757 (N_8757,N_8665,N_8605);
and U8758 (N_8758,N_8696,N_8604);
or U8759 (N_8759,N_8680,N_8620);
or U8760 (N_8760,N_8699,N_8660);
nand U8761 (N_8761,N_8627,N_8684);
or U8762 (N_8762,N_8648,N_8661);
and U8763 (N_8763,N_8649,N_8656);
xnor U8764 (N_8764,N_8644,N_8664);
or U8765 (N_8765,N_8612,N_8638);
nand U8766 (N_8766,N_8667,N_8619);
and U8767 (N_8767,N_8640,N_8623);
nor U8768 (N_8768,N_8648,N_8691);
and U8769 (N_8769,N_8657,N_8653);
xor U8770 (N_8770,N_8679,N_8640);
nand U8771 (N_8771,N_8600,N_8608);
and U8772 (N_8772,N_8629,N_8616);
nand U8773 (N_8773,N_8602,N_8613);
or U8774 (N_8774,N_8670,N_8646);
or U8775 (N_8775,N_8693,N_8671);
nand U8776 (N_8776,N_8654,N_8651);
or U8777 (N_8777,N_8638,N_8679);
and U8778 (N_8778,N_8627,N_8674);
or U8779 (N_8779,N_8691,N_8678);
nand U8780 (N_8780,N_8626,N_8643);
and U8781 (N_8781,N_8633,N_8637);
nand U8782 (N_8782,N_8623,N_8600);
nand U8783 (N_8783,N_8608,N_8646);
nand U8784 (N_8784,N_8622,N_8667);
and U8785 (N_8785,N_8629,N_8683);
nand U8786 (N_8786,N_8677,N_8607);
and U8787 (N_8787,N_8667,N_8627);
or U8788 (N_8788,N_8668,N_8640);
or U8789 (N_8789,N_8629,N_8630);
or U8790 (N_8790,N_8689,N_8634);
nor U8791 (N_8791,N_8636,N_8622);
or U8792 (N_8792,N_8664,N_8609);
nand U8793 (N_8793,N_8645,N_8676);
and U8794 (N_8794,N_8686,N_8631);
and U8795 (N_8795,N_8632,N_8622);
nand U8796 (N_8796,N_8623,N_8692);
nor U8797 (N_8797,N_8666,N_8661);
nor U8798 (N_8798,N_8699,N_8671);
nand U8799 (N_8799,N_8655,N_8668);
and U8800 (N_8800,N_8725,N_8721);
and U8801 (N_8801,N_8757,N_8788);
nor U8802 (N_8802,N_8752,N_8731);
or U8803 (N_8803,N_8732,N_8700);
xnor U8804 (N_8804,N_8715,N_8764);
and U8805 (N_8805,N_8741,N_8782);
and U8806 (N_8806,N_8756,N_8747);
or U8807 (N_8807,N_8720,N_8706);
nor U8808 (N_8808,N_8761,N_8762);
nand U8809 (N_8809,N_8745,N_8763);
xor U8810 (N_8810,N_8701,N_8717);
nor U8811 (N_8811,N_8794,N_8733);
or U8812 (N_8812,N_8718,N_8736);
nand U8813 (N_8813,N_8716,N_8726);
nor U8814 (N_8814,N_8777,N_8743);
nor U8815 (N_8815,N_8769,N_8751);
nor U8816 (N_8816,N_8771,N_8798);
and U8817 (N_8817,N_8750,N_8765);
nor U8818 (N_8818,N_8702,N_8713);
and U8819 (N_8819,N_8760,N_8709);
nand U8820 (N_8820,N_8767,N_8746);
or U8821 (N_8821,N_8719,N_8722);
and U8822 (N_8822,N_8799,N_8710);
or U8823 (N_8823,N_8783,N_8758);
and U8824 (N_8824,N_8795,N_8707);
nor U8825 (N_8825,N_8753,N_8779);
or U8826 (N_8826,N_8778,N_8748);
or U8827 (N_8827,N_8704,N_8712);
nor U8828 (N_8828,N_8791,N_8755);
nand U8829 (N_8829,N_8776,N_8770);
or U8830 (N_8830,N_8728,N_8773);
or U8831 (N_8831,N_8737,N_8724);
xnor U8832 (N_8832,N_8723,N_8797);
and U8833 (N_8833,N_8790,N_8708);
nor U8834 (N_8834,N_8734,N_8789);
nor U8835 (N_8835,N_8739,N_8729);
nand U8836 (N_8836,N_8766,N_8727);
or U8837 (N_8837,N_8703,N_8768);
and U8838 (N_8838,N_8774,N_8775);
and U8839 (N_8839,N_8744,N_8792);
and U8840 (N_8840,N_8786,N_8735);
nor U8841 (N_8841,N_8772,N_8780);
or U8842 (N_8842,N_8793,N_8740);
nor U8843 (N_8843,N_8730,N_8749);
nor U8844 (N_8844,N_8781,N_8714);
nand U8845 (N_8845,N_8742,N_8796);
and U8846 (N_8846,N_8759,N_8785);
nand U8847 (N_8847,N_8705,N_8711);
and U8848 (N_8848,N_8738,N_8784);
nor U8849 (N_8849,N_8787,N_8754);
nor U8850 (N_8850,N_8773,N_8742);
and U8851 (N_8851,N_8722,N_8736);
nand U8852 (N_8852,N_8760,N_8798);
nand U8853 (N_8853,N_8782,N_8703);
nor U8854 (N_8854,N_8726,N_8798);
or U8855 (N_8855,N_8738,N_8770);
nand U8856 (N_8856,N_8731,N_8711);
or U8857 (N_8857,N_8777,N_8762);
nor U8858 (N_8858,N_8717,N_8709);
nor U8859 (N_8859,N_8755,N_8771);
and U8860 (N_8860,N_8764,N_8782);
nor U8861 (N_8861,N_8745,N_8708);
nor U8862 (N_8862,N_8720,N_8745);
or U8863 (N_8863,N_8785,N_8724);
nor U8864 (N_8864,N_8704,N_8793);
or U8865 (N_8865,N_8740,N_8777);
nor U8866 (N_8866,N_8709,N_8732);
and U8867 (N_8867,N_8713,N_8721);
or U8868 (N_8868,N_8731,N_8786);
nor U8869 (N_8869,N_8715,N_8723);
and U8870 (N_8870,N_8735,N_8757);
nor U8871 (N_8871,N_8769,N_8774);
nand U8872 (N_8872,N_8783,N_8706);
nor U8873 (N_8873,N_8793,N_8748);
nor U8874 (N_8874,N_8775,N_8756);
and U8875 (N_8875,N_8701,N_8755);
nor U8876 (N_8876,N_8712,N_8787);
and U8877 (N_8877,N_8710,N_8702);
or U8878 (N_8878,N_8793,N_8749);
nand U8879 (N_8879,N_8754,N_8746);
nand U8880 (N_8880,N_8786,N_8734);
and U8881 (N_8881,N_8761,N_8727);
and U8882 (N_8882,N_8743,N_8778);
nor U8883 (N_8883,N_8720,N_8725);
nand U8884 (N_8884,N_8709,N_8747);
and U8885 (N_8885,N_8723,N_8784);
or U8886 (N_8886,N_8735,N_8795);
nand U8887 (N_8887,N_8709,N_8773);
nand U8888 (N_8888,N_8727,N_8749);
or U8889 (N_8889,N_8754,N_8793);
and U8890 (N_8890,N_8791,N_8787);
nor U8891 (N_8891,N_8789,N_8776);
nor U8892 (N_8892,N_8796,N_8753);
xor U8893 (N_8893,N_8792,N_8709);
nor U8894 (N_8894,N_8723,N_8777);
nor U8895 (N_8895,N_8799,N_8762);
nand U8896 (N_8896,N_8781,N_8799);
or U8897 (N_8897,N_8728,N_8729);
nor U8898 (N_8898,N_8714,N_8749);
and U8899 (N_8899,N_8721,N_8771);
or U8900 (N_8900,N_8845,N_8836);
or U8901 (N_8901,N_8841,N_8858);
nand U8902 (N_8902,N_8869,N_8815);
nor U8903 (N_8903,N_8814,N_8811);
and U8904 (N_8904,N_8847,N_8853);
and U8905 (N_8905,N_8817,N_8849);
and U8906 (N_8906,N_8832,N_8877);
nand U8907 (N_8907,N_8868,N_8804);
or U8908 (N_8908,N_8862,N_8843);
or U8909 (N_8909,N_8865,N_8840);
nand U8910 (N_8910,N_8897,N_8889);
or U8911 (N_8911,N_8895,N_8827);
and U8912 (N_8912,N_8833,N_8828);
nor U8913 (N_8913,N_8805,N_8850);
nand U8914 (N_8914,N_8857,N_8881);
or U8915 (N_8915,N_8892,N_8854);
and U8916 (N_8916,N_8874,N_8873);
nand U8917 (N_8917,N_8826,N_8848);
and U8918 (N_8918,N_8878,N_8834);
or U8919 (N_8919,N_8801,N_8896);
and U8920 (N_8920,N_8837,N_8838);
nand U8921 (N_8921,N_8818,N_8898);
and U8922 (N_8922,N_8880,N_8863);
and U8923 (N_8923,N_8856,N_8890);
nor U8924 (N_8924,N_8846,N_8887);
xor U8925 (N_8925,N_8871,N_8866);
or U8926 (N_8926,N_8852,N_8851);
and U8927 (N_8927,N_8807,N_8816);
or U8928 (N_8928,N_8830,N_8806);
nand U8929 (N_8929,N_8813,N_8809);
nor U8930 (N_8930,N_8844,N_8886);
or U8931 (N_8931,N_8860,N_8859);
nor U8932 (N_8932,N_8870,N_8891);
nand U8933 (N_8933,N_8822,N_8831);
nor U8934 (N_8934,N_8894,N_8835);
or U8935 (N_8935,N_8893,N_8810);
nor U8936 (N_8936,N_8879,N_8800);
nor U8937 (N_8937,N_8861,N_8820);
and U8938 (N_8938,N_8803,N_8864);
and U8939 (N_8939,N_8855,N_8885);
and U8940 (N_8940,N_8884,N_8825);
nor U8941 (N_8941,N_8883,N_8808);
or U8942 (N_8942,N_8899,N_8839);
and U8943 (N_8943,N_8888,N_8829);
nand U8944 (N_8944,N_8824,N_8876);
or U8945 (N_8945,N_8802,N_8875);
or U8946 (N_8946,N_8872,N_8821);
and U8947 (N_8947,N_8867,N_8819);
nor U8948 (N_8948,N_8812,N_8823);
or U8949 (N_8949,N_8882,N_8842);
nand U8950 (N_8950,N_8891,N_8864);
and U8951 (N_8951,N_8876,N_8853);
and U8952 (N_8952,N_8836,N_8806);
or U8953 (N_8953,N_8834,N_8818);
xnor U8954 (N_8954,N_8810,N_8872);
nand U8955 (N_8955,N_8826,N_8849);
or U8956 (N_8956,N_8843,N_8811);
nand U8957 (N_8957,N_8853,N_8863);
nor U8958 (N_8958,N_8868,N_8859);
nand U8959 (N_8959,N_8871,N_8875);
nand U8960 (N_8960,N_8817,N_8883);
nor U8961 (N_8961,N_8893,N_8812);
and U8962 (N_8962,N_8818,N_8864);
nor U8963 (N_8963,N_8814,N_8813);
xor U8964 (N_8964,N_8801,N_8841);
nand U8965 (N_8965,N_8815,N_8814);
nor U8966 (N_8966,N_8877,N_8860);
or U8967 (N_8967,N_8879,N_8893);
nor U8968 (N_8968,N_8888,N_8800);
and U8969 (N_8969,N_8812,N_8869);
nand U8970 (N_8970,N_8843,N_8858);
and U8971 (N_8971,N_8832,N_8801);
nand U8972 (N_8972,N_8806,N_8832);
and U8973 (N_8973,N_8895,N_8875);
nor U8974 (N_8974,N_8808,N_8875);
nand U8975 (N_8975,N_8813,N_8810);
nand U8976 (N_8976,N_8841,N_8873);
and U8977 (N_8977,N_8893,N_8863);
or U8978 (N_8978,N_8855,N_8801);
nor U8979 (N_8979,N_8828,N_8868);
or U8980 (N_8980,N_8824,N_8804);
or U8981 (N_8981,N_8884,N_8805);
and U8982 (N_8982,N_8820,N_8842);
nor U8983 (N_8983,N_8857,N_8809);
nor U8984 (N_8984,N_8848,N_8803);
nor U8985 (N_8985,N_8897,N_8822);
nand U8986 (N_8986,N_8857,N_8824);
nor U8987 (N_8987,N_8845,N_8886);
nor U8988 (N_8988,N_8828,N_8832);
nor U8989 (N_8989,N_8839,N_8820);
nor U8990 (N_8990,N_8889,N_8887);
and U8991 (N_8991,N_8858,N_8864);
nor U8992 (N_8992,N_8859,N_8828);
nand U8993 (N_8993,N_8845,N_8864);
nor U8994 (N_8994,N_8807,N_8810);
and U8995 (N_8995,N_8814,N_8894);
and U8996 (N_8996,N_8801,N_8851);
nor U8997 (N_8997,N_8885,N_8816);
nor U8998 (N_8998,N_8895,N_8828);
and U8999 (N_8999,N_8851,N_8885);
and U9000 (N_9000,N_8954,N_8987);
or U9001 (N_9001,N_8956,N_8969);
nor U9002 (N_9002,N_8916,N_8927);
nor U9003 (N_9003,N_8926,N_8925);
nor U9004 (N_9004,N_8904,N_8915);
and U9005 (N_9005,N_8951,N_8995);
nor U9006 (N_9006,N_8962,N_8974);
or U9007 (N_9007,N_8931,N_8923);
nor U9008 (N_9008,N_8944,N_8943);
nor U9009 (N_9009,N_8936,N_8976);
nor U9010 (N_9010,N_8938,N_8972);
nand U9011 (N_9011,N_8953,N_8913);
xor U9012 (N_9012,N_8947,N_8975);
nor U9013 (N_9013,N_8961,N_8966);
nor U9014 (N_9014,N_8930,N_8901);
or U9015 (N_9015,N_8914,N_8919);
nor U9016 (N_9016,N_8998,N_8932);
nor U9017 (N_9017,N_8984,N_8909);
and U9018 (N_9018,N_8902,N_8989);
or U9019 (N_9019,N_8973,N_8999);
and U9020 (N_9020,N_8977,N_8964);
nor U9021 (N_9021,N_8991,N_8979);
xor U9022 (N_9022,N_8946,N_8935);
and U9023 (N_9023,N_8957,N_8942);
nand U9024 (N_9024,N_8934,N_8908);
and U9025 (N_9025,N_8970,N_8996);
and U9026 (N_9026,N_8903,N_8980);
nand U9027 (N_9027,N_8960,N_8929);
nor U9028 (N_9028,N_8985,N_8922);
nor U9029 (N_9029,N_8941,N_8990);
or U9030 (N_9030,N_8949,N_8986);
or U9031 (N_9031,N_8965,N_8993);
and U9032 (N_9032,N_8907,N_8918);
or U9033 (N_9033,N_8940,N_8968);
nand U9034 (N_9034,N_8933,N_8982);
or U9035 (N_9035,N_8945,N_8988);
nand U9036 (N_9036,N_8920,N_8924);
and U9037 (N_9037,N_8971,N_8910);
or U9038 (N_9038,N_8921,N_8967);
nor U9039 (N_9039,N_8981,N_8994);
nor U9040 (N_9040,N_8912,N_8900);
nor U9041 (N_9041,N_8997,N_8978);
nor U9042 (N_9042,N_8905,N_8959);
nand U9043 (N_9043,N_8992,N_8937);
nor U9044 (N_9044,N_8983,N_8952);
nor U9045 (N_9045,N_8955,N_8948);
and U9046 (N_9046,N_8939,N_8950);
nor U9047 (N_9047,N_8911,N_8958);
or U9048 (N_9048,N_8928,N_8906);
and U9049 (N_9049,N_8917,N_8963);
nor U9050 (N_9050,N_8969,N_8971);
and U9051 (N_9051,N_8901,N_8969);
xor U9052 (N_9052,N_8918,N_8983);
and U9053 (N_9053,N_8915,N_8989);
nor U9054 (N_9054,N_8922,N_8997);
nor U9055 (N_9055,N_8926,N_8995);
or U9056 (N_9056,N_8957,N_8941);
nand U9057 (N_9057,N_8913,N_8916);
or U9058 (N_9058,N_8937,N_8990);
nand U9059 (N_9059,N_8989,N_8986);
or U9060 (N_9060,N_8958,N_8900);
and U9061 (N_9061,N_8918,N_8966);
nand U9062 (N_9062,N_8900,N_8915);
or U9063 (N_9063,N_8959,N_8902);
and U9064 (N_9064,N_8959,N_8966);
nand U9065 (N_9065,N_8982,N_8946);
nor U9066 (N_9066,N_8908,N_8957);
nor U9067 (N_9067,N_8907,N_8917);
and U9068 (N_9068,N_8903,N_8905);
nand U9069 (N_9069,N_8999,N_8994);
nand U9070 (N_9070,N_8920,N_8949);
nor U9071 (N_9071,N_8993,N_8928);
or U9072 (N_9072,N_8994,N_8931);
xnor U9073 (N_9073,N_8982,N_8948);
nor U9074 (N_9074,N_8966,N_8919);
and U9075 (N_9075,N_8921,N_8961);
and U9076 (N_9076,N_8924,N_8983);
nor U9077 (N_9077,N_8967,N_8907);
and U9078 (N_9078,N_8944,N_8961);
nand U9079 (N_9079,N_8902,N_8956);
xnor U9080 (N_9080,N_8956,N_8927);
or U9081 (N_9081,N_8924,N_8917);
or U9082 (N_9082,N_8951,N_8963);
and U9083 (N_9083,N_8985,N_8977);
and U9084 (N_9084,N_8948,N_8990);
nor U9085 (N_9085,N_8977,N_8981);
xnor U9086 (N_9086,N_8913,N_8904);
nand U9087 (N_9087,N_8975,N_8974);
xnor U9088 (N_9088,N_8907,N_8985);
nand U9089 (N_9089,N_8948,N_8932);
nor U9090 (N_9090,N_8995,N_8990);
and U9091 (N_9091,N_8936,N_8918);
nor U9092 (N_9092,N_8900,N_8916);
nand U9093 (N_9093,N_8913,N_8943);
nand U9094 (N_9094,N_8989,N_8984);
nor U9095 (N_9095,N_8950,N_8981);
nor U9096 (N_9096,N_8997,N_8991);
nand U9097 (N_9097,N_8936,N_8999);
or U9098 (N_9098,N_8989,N_8947);
and U9099 (N_9099,N_8934,N_8952);
and U9100 (N_9100,N_9046,N_9043);
or U9101 (N_9101,N_9094,N_9027);
nand U9102 (N_9102,N_9018,N_9047);
nand U9103 (N_9103,N_9070,N_9089);
nor U9104 (N_9104,N_9034,N_9056);
nor U9105 (N_9105,N_9055,N_9085);
or U9106 (N_9106,N_9037,N_9024);
nand U9107 (N_9107,N_9010,N_9050);
xor U9108 (N_9108,N_9068,N_9090);
or U9109 (N_9109,N_9038,N_9076);
nor U9110 (N_9110,N_9006,N_9019);
nor U9111 (N_9111,N_9045,N_9028);
and U9112 (N_9112,N_9051,N_9000);
nand U9113 (N_9113,N_9007,N_9087);
nand U9114 (N_9114,N_9078,N_9030);
and U9115 (N_9115,N_9016,N_9048);
nand U9116 (N_9116,N_9063,N_9025);
and U9117 (N_9117,N_9069,N_9044);
nand U9118 (N_9118,N_9035,N_9029);
nor U9119 (N_9119,N_9088,N_9036);
nand U9120 (N_9120,N_9005,N_9004);
nor U9121 (N_9121,N_9023,N_9093);
and U9122 (N_9122,N_9021,N_9058);
and U9123 (N_9123,N_9092,N_9059);
or U9124 (N_9124,N_9091,N_9008);
nand U9125 (N_9125,N_9039,N_9084);
nand U9126 (N_9126,N_9049,N_9026);
nor U9127 (N_9127,N_9097,N_9098);
or U9128 (N_9128,N_9017,N_9062);
and U9129 (N_9129,N_9003,N_9080);
and U9130 (N_9130,N_9081,N_9052);
and U9131 (N_9131,N_9057,N_9061);
or U9132 (N_9132,N_9053,N_9060);
or U9133 (N_9133,N_9072,N_9014);
nor U9134 (N_9134,N_9067,N_9032);
nand U9135 (N_9135,N_9064,N_9015);
or U9136 (N_9136,N_9075,N_9083);
nand U9137 (N_9137,N_9011,N_9042);
nor U9138 (N_9138,N_9001,N_9033);
or U9139 (N_9139,N_9071,N_9077);
xnor U9140 (N_9140,N_9054,N_9066);
or U9141 (N_9141,N_9041,N_9096);
nand U9142 (N_9142,N_9073,N_9020);
and U9143 (N_9143,N_9002,N_9082);
nand U9144 (N_9144,N_9086,N_9074);
or U9145 (N_9145,N_9095,N_9040);
xnor U9146 (N_9146,N_9065,N_9022);
or U9147 (N_9147,N_9013,N_9099);
nor U9148 (N_9148,N_9009,N_9012);
or U9149 (N_9149,N_9079,N_9031);
nand U9150 (N_9150,N_9066,N_9002);
xnor U9151 (N_9151,N_9056,N_9072);
and U9152 (N_9152,N_9044,N_9026);
nand U9153 (N_9153,N_9043,N_9034);
xor U9154 (N_9154,N_9038,N_9029);
and U9155 (N_9155,N_9046,N_9021);
nand U9156 (N_9156,N_9074,N_9002);
nand U9157 (N_9157,N_9034,N_9090);
nor U9158 (N_9158,N_9032,N_9078);
and U9159 (N_9159,N_9061,N_9078);
xnor U9160 (N_9160,N_9042,N_9003);
and U9161 (N_9161,N_9058,N_9071);
nor U9162 (N_9162,N_9041,N_9006);
and U9163 (N_9163,N_9080,N_9001);
nor U9164 (N_9164,N_9011,N_9060);
and U9165 (N_9165,N_9051,N_9020);
nor U9166 (N_9166,N_9062,N_9086);
nand U9167 (N_9167,N_9081,N_9040);
nor U9168 (N_9168,N_9074,N_9016);
and U9169 (N_9169,N_9090,N_9063);
nor U9170 (N_9170,N_9084,N_9020);
or U9171 (N_9171,N_9011,N_9028);
nor U9172 (N_9172,N_9009,N_9085);
nor U9173 (N_9173,N_9065,N_9062);
nand U9174 (N_9174,N_9078,N_9039);
nor U9175 (N_9175,N_9099,N_9034);
or U9176 (N_9176,N_9027,N_9081);
nand U9177 (N_9177,N_9008,N_9055);
and U9178 (N_9178,N_9051,N_9072);
and U9179 (N_9179,N_9030,N_9059);
and U9180 (N_9180,N_9052,N_9050);
or U9181 (N_9181,N_9062,N_9011);
nand U9182 (N_9182,N_9091,N_9061);
or U9183 (N_9183,N_9099,N_9014);
nor U9184 (N_9184,N_9001,N_9084);
nor U9185 (N_9185,N_9097,N_9012);
and U9186 (N_9186,N_9019,N_9096);
or U9187 (N_9187,N_9024,N_9027);
nor U9188 (N_9188,N_9083,N_9071);
nand U9189 (N_9189,N_9046,N_9098);
nor U9190 (N_9190,N_9070,N_9056);
or U9191 (N_9191,N_9048,N_9054);
and U9192 (N_9192,N_9018,N_9028);
nand U9193 (N_9193,N_9006,N_9089);
or U9194 (N_9194,N_9008,N_9084);
and U9195 (N_9195,N_9027,N_9042);
nor U9196 (N_9196,N_9041,N_9043);
nor U9197 (N_9197,N_9028,N_9049);
nor U9198 (N_9198,N_9071,N_9098);
nor U9199 (N_9199,N_9029,N_9007);
or U9200 (N_9200,N_9159,N_9107);
nor U9201 (N_9201,N_9186,N_9194);
and U9202 (N_9202,N_9195,N_9133);
and U9203 (N_9203,N_9135,N_9119);
and U9204 (N_9204,N_9189,N_9157);
nor U9205 (N_9205,N_9126,N_9134);
nor U9206 (N_9206,N_9150,N_9192);
nor U9207 (N_9207,N_9122,N_9104);
and U9208 (N_9208,N_9130,N_9121);
nor U9209 (N_9209,N_9116,N_9144);
nor U9210 (N_9210,N_9124,N_9110);
and U9211 (N_9211,N_9147,N_9118);
nor U9212 (N_9212,N_9129,N_9160);
or U9213 (N_9213,N_9145,N_9162);
nand U9214 (N_9214,N_9113,N_9103);
and U9215 (N_9215,N_9188,N_9137);
and U9216 (N_9216,N_9117,N_9155);
nor U9217 (N_9217,N_9173,N_9132);
or U9218 (N_9218,N_9182,N_9164);
nand U9219 (N_9219,N_9158,N_9105);
nor U9220 (N_9220,N_9136,N_9112);
nand U9221 (N_9221,N_9161,N_9100);
nor U9222 (N_9222,N_9167,N_9153);
or U9223 (N_9223,N_9177,N_9111);
and U9224 (N_9224,N_9138,N_9183);
or U9225 (N_9225,N_9175,N_9190);
and U9226 (N_9226,N_9152,N_9156);
or U9227 (N_9227,N_9115,N_9184);
nand U9228 (N_9228,N_9109,N_9151);
and U9229 (N_9229,N_9140,N_9148);
and U9230 (N_9230,N_9106,N_9128);
and U9231 (N_9231,N_9187,N_9197);
and U9232 (N_9232,N_9139,N_9142);
nand U9233 (N_9233,N_9170,N_9141);
nand U9234 (N_9234,N_9120,N_9176);
and U9235 (N_9235,N_9169,N_9178);
nand U9236 (N_9236,N_9191,N_9108);
and U9237 (N_9237,N_9193,N_9180);
and U9238 (N_9238,N_9131,N_9102);
or U9239 (N_9239,N_9163,N_9165);
and U9240 (N_9240,N_9146,N_9171);
or U9241 (N_9241,N_9123,N_9196);
or U9242 (N_9242,N_9127,N_9179);
nor U9243 (N_9243,N_9199,N_9166);
or U9244 (N_9244,N_9198,N_9154);
nand U9245 (N_9245,N_9114,N_9143);
nand U9246 (N_9246,N_9185,N_9125);
xnor U9247 (N_9247,N_9101,N_9168);
or U9248 (N_9248,N_9149,N_9181);
and U9249 (N_9249,N_9172,N_9174);
or U9250 (N_9250,N_9181,N_9109);
nor U9251 (N_9251,N_9151,N_9104);
and U9252 (N_9252,N_9159,N_9142);
and U9253 (N_9253,N_9192,N_9169);
nand U9254 (N_9254,N_9160,N_9153);
nor U9255 (N_9255,N_9187,N_9122);
nor U9256 (N_9256,N_9128,N_9133);
nand U9257 (N_9257,N_9162,N_9177);
nand U9258 (N_9258,N_9196,N_9199);
and U9259 (N_9259,N_9183,N_9168);
or U9260 (N_9260,N_9137,N_9106);
and U9261 (N_9261,N_9126,N_9164);
nand U9262 (N_9262,N_9143,N_9182);
nand U9263 (N_9263,N_9115,N_9157);
or U9264 (N_9264,N_9134,N_9186);
or U9265 (N_9265,N_9182,N_9107);
nand U9266 (N_9266,N_9193,N_9126);
nand U9267 (N_9267,N_9117,N_9108);
or U9268 (N_9268,N_9170,N_9150);
nor U9269 (N_9269,N_9147,N_9173);
nand U9270 (N_9270,N_9178,N_9125);
xor U9271 (N_9271,N_9122,N_9158);
nor U9272 (N_9272,N_9109,N_9184);
nor U9273 (N_9273,N_9161,N_9132);
and U9274 (N_9274,N_9163,N_9191);
or U9275 (N_9275,N_9144,N_9130);
nand U9276 (N_9276,N_9110,N_9181);
nor U9277 (N_9277,N_9184,N_9153);
nand U9278 (N_9278,N_9164,N_9125);
nor U9279 (N_9279,N_9128,N_9127);
or U9280 (N_9280,N_9178,N_9185);
nand U9281 (N_9281,N_9162,N_9128);
or U9282 (N_9282,N_9187,N_9168);
or U9283 (N_9283,N_9193,N_9112);
nand U9284 (N_9284,N_9198,N_9111);
or U9285 (N_9285,N_9159,N_9155);
or U9286 (N_9286,N_9198,N_9129);
nand U9287 (N_9287,N_9125,N_9194);
nand U9288 (N_9288,N_9128,N_9191);
nor U9289 (N_9289,N_9132,N_9163);
nand U9290 (N_9290,N_9171,N_9142);
and U9291 (N_9291,N_9119,N_9105);
or U9292 (N_9292,N_9118,N_9111);
or U9293 (N_9293,N_9171,N_9183);
and U9294 (N_9294,N_9160,N_9131);
or U9295 (N_9295,N_9196,N_9143);
and U9296 (N_9296,N_9188,N_9164);
or U9297 (N_9297,N_9185,N_9161);
nor U9298 (N_9298,N_9114,N_9135);
nand U9299 (N_9299,N_9109,N_9169);
and U9300 (N_9300,N_9233,N_9297);
and U9301 (N_9301,N_9273,N_9287);
nor U9302 (N_9302,N_9296,N_9200);
and U9303 (N_9303,N_9222,N_9229);
nor U9304 (N_9304,N_9276,N_9241);
nand U9305 (N_9305,N_9268,N_9207);
nor U9306 (N_9306,N_9205,N_9245);
or U9307 (N_9307,N_9293,N_9292);
and U9308 (N_9308,N_9239,N_9262);
nand U9309 (N_9309,N_9203,N_9257);
and U9310 (N_9310,N_9211,N_9219);
or U9311 (N_9311,N_9288,N_9232);
or U9312 (N_9312,N_9235,N_9277);
nand U9313 (N_9313,N_9281,N_9243);
nor U9314 (N_9314,N_9242,N_9230);
or U9315 (N_9315,N_9261,N_9254);
and U9316 (N_9316,N_9249,N_9206);
nand U9317 (N_9317,N_9215,N_9265);
or U9318 (N_9318,N_9269,N_9255);
or U9319 (N_9319,N_9266,N_9208);
or U9320 (N_9320,N_9283,N_9285);
or U9321 (N_9321,N_9271,N_9278);
nor U9322 (N_9322,N_9221,N_9260);
nand U9323 (N_9323,N_9202,N_9214);
nand U9324 (N_9324,N_9246,N_9256);
nor U9325 (N_9325,N_9290,N_9201);
or U9326 (N_9326,N_9251,N_9279);
nand U9327 (N_9327,N_9234,N_9218);
nand U9328 (N_9328,N_9212,N_9280);
nand U9329 (N_9329,N_9217,N_9289);
or U9330 (N_9330,N_9253,N_9225);
nor U9331 (N_9331,N_9226,N_9220);
or U9332 (N_9332,N_9240,N_9236);
nand U9333 (N_9333,N_9282,N_9291);
nor U9334 (N_9334,N_9223,N_9227);
nor U9335 (N_9335,N_9210,N_9259);
nor U9336 (N_9336,N_9267,N_9216);
or U9337 (N_9337,N_9247,N_9213);
or U9338 (N_9338,N_9275,N_9272);
xor U9339 (N_9339,N_9299,N_9274);
xor U9340 (N_9340,N_9286,N_9228);
nand U9341 (N_9341,N_9298,N_9224);
nor U9342 (N_9342,N_9258,N_9250);
nor U9343 (N_9343,N_9264,N_9244);
and U9344 (N_9344,N_9263,N_9294);
or U9345 (N_9345,N_9252,N_9248);
nand U9346 (N_9346,N_9238,N_9270);
or U9347 (N_9347,N_9295,N_9204);
nor U9348 (N_9348,N_9237,N_9209);
nor U9349 (N_9349,N_9231,N_9284);
and U9350 (N_9350,N_9252,N_9291);
or U9351 (N_9351,N_9225,N_9242);
nor U9352 (N_9352,N_9269,N_9243);
xnor U9353 (N_9353,N_9216,N_9256);
nand U9354 (N_9354,N_9251,N_9250);
and U9355 (N_9355,N_9264,N_9269);
nor U9356 (N_9356,N_9204,N_9282);
nand U9357 (N_9357,N_9294,N_9258);
or U9358 (N_9358,N_9251,N_9215);
nand U9359 (N_9359,N_9224,N_9243);
and U9360 (N_9360,N_9289,N_9283);
nor U9361 (N_9361,N_9261,N_9265);
or U9362 (N_9362,N_9280,N_9239);
nand U9363 (N_9363,N_9274,N_9272);
nor U9364 (N_9364,N_9219,N_9213);
nor U9365 (N_9365,N_9212,N_9241);
and U9366 (N_9366,N_9293,N_9265);
or U9367 (N_9367,N_9255,N_9236);
and U9368 (N_9368,N_9256,N_9244);
and U9369 (N_9369,N_9216,N_9210);
and U9370 (N_9370,N_9204,N_9268);
or U9371 (N_9371,N_9236,N_9203);
nor U9372 (N_9372,N_9265,N_9223);
nand U9373 (N_9373,N_9255,N_9266);
nor U9374 (N_9374,N_9297,N_9255);
nor U9375 (N_9375,N_9288,N_9213);
nand U9376 (N_9376,N_9297,N_9205);
and U9377 (N_9377,N_9297,N_9235);
nor U9378 (N_9378,N_9204,N_9252);
nor U9379 (N_9379,N_9257,N_9267);
nor U9380 (N_9380,N_9222,N_9237);
nand U9381 (N_9381,N_9252,N_9295);
and U9382 (N_9382,N_9256,N_9206);
nand U9383 (N_9383,N_9271,N_9206);
or U9384 (N_9384,N_9240,N_9256);
nor U9385 (N_9385,N_9247,N_9273);
and U9386 (N_9386,N_9222,N_9278);
nor U9387 (N_9387,N_9236,N_9272);
or U9388 (N_9388,N_9289,N_9215);
and U9389 (N_9389,N_9238,N_9204);
nand U9390 (N_9390,N_9263,N_9295);
and U9391 (N_9391,N_9299,N_9220);
nor U9392 (N_9392,N_9290,N_9216);
and U9393 (N_9393,N_9266,N_9272);
and U9394 (N_9394,N_9242,N_9202);
or U9395 (N_9395,N_9283,N_9280);
nand U9396 (N_9396,N_9275,N_9243);
nor U9397 (N_9397,N_9261,N_9206);
or U9398 (N_9398,N_9232,N_9200);
nand U9399 (N_9399,N_9238,N_9201);
or U9400 (N_9400,N_9337,N_9347);
and U9401 (N_9401,N_9379,N_9380);
xor U9402 (N_9402,N_9353,N_9384);
nor U9403 (N_9403,N_9340,N_9316);
and U9404 (N_9404,N_9378,N_9303);
or U9405 (N_9405,N_9365,N_9394);
nand U9406 (N_9406,N_9359,N_9322);
nor U9407 (N_9407,N_9317,N_9306);
or U9408 (N_9408,N_9351,N_9357);
and U9409 (N_9409,N_9315,N_9331);
nand U9410 (N_9410,N_9301,N_9355);
nand U9411 (N_9411,N_9362,N_9393);
nand U9412 (N_9412,N_9390,N_9319);
nand U9413 (N_9413,N_9300,N_9326);
nor U9414 (N_9414,N_9302,N_9318);
and U9415 (N_9415,N_9314,N_9352);
or U9416 (N_9416,N_9367,N_9361);
nand U9417 (N_9417,N_9313,N_9376);
nand U9418 (N_9418,N_9396,N_9369);
nand U9419 (N_9419,N_9385,N_9372);
and U9420 (N_9420,N_9375,N_9323);
xnor U9421 (N_9421,N_9341,N_9387);
nor U9422 (N_9422,N_9320,N_9345);
or U9423 (N_9423,N_9307,N_9343);
nor U9424 (N_9424,N_9321,N_9324);
and U9425 (N_9425,N_9346,N_9338);
nor U9426 (N_9426,N_9356,N_9309);
or U9427 (N_9427,N_9391,N_9368);
nand U9428 (N_9428,N_9381,N_9364);
nand U9429 (N_9429,N_9334,N_9363);
and U9430 (N_9430,N_9344,N_9370);
nor U9431 (N_9431,N_9354,N_9311);
and U9432 (N_9432,N_9310,N_9366);
or U9433 (N_9433,N_9328,N_9327);
nand U9434 (N_9434,N_9388,N_9360);
nand U9435 (N_9435,N_9389,N_9308);
or U9436 (N_9436,N_9399,N_9305);
nor U9437 (N_9437,N_9312,N_9377);
nand U9438 (N_9438,N_9358,N_9392);
and U9439 (N_9439,N_9395,N_9371);
nor U9440 (N_9440,N_9329,N_9304);
nor U9441 (N_9441,N_9373,N_9325);
or U9442 (N_9442,N_9398,N_9382);
nor U9443 (N_9443,N_9335,N_9342);
or U9444 (N_9444,N_9333,N_9336);
nand U9445 (N_9445,N_9330,N_9386);
or U9446 (N_9446,N_9383,N_9349);
nor U9447 (N_9447,N_9348,N_9350);
and U9448 (N_9448,N_9339,N_9397);
or U9449 (N_9449,N_9374,N_9332);
or U9450 (N_9450,N_9326,N_9308);
and U9451 (N_9451,N_9370,N_9363);
nand U9452 (N_9452,N_9382,N_9338);
or U9453 (N_9453,N_9340,N_9378);
nand U9454 (N_9454,N_9300,N_9316);
and U9455 (N_9455,N_9344,N_9324);
nor U9456 (N_9456,N_9392,N_9330);
or U9457 (N_9457,N_9391,N_9359);
and U9458 (N_9458,N_9312,N_9384);
or U9459 (N_9459,N_9359,N_9317);
or U9460 (N_9460,N_9321,N_9378);
nand U9461 (N_9461,N_9317,N_9388);
or U9462 (N_9462,N_9357,N_9367);
nor U9463 (N_9463,N_9354,N_9378);
or U9464 (N_9464,N_9342,N_9373);
xnor U9465 (N_9465,N_9301,N_9395);
nor U9466 (N_9466,N_9394,N_9366);
and U9467 (N_9467,N_9306,N_9352);
nand U9468 (N_9468,N_9310,N_9362);
and U9469 (N_9469,N_9399,N_9343);
nand U9470 (N_9470,N_9383,N_9309);
and U9471 (N_9471,N_9366,N_9315);
nand U9472 (N_9472,N_9399,N_9393);
nor U9473 (N_9473,N_9315,N_9398);
and U9474 (N_9474,N_9355,N_9388);
or U9475 (N_9475,N_9320,N_9343);
nor U9476 (N_9476,N_9338,N_9356);
or U9477 (N_9477,N_9332,N_9361);
nor U9478 (N_9478,N_9322,N_9351);
nand U9479 (N_9479,N_9336,N_9364);
and U9480 (N_9480,N_9384,N_9362);
and U9481 (N_9481,N_9326,N_9374);
or U9482 (N_9482,N_9392,N_9391);
and U9483 (N_9483,N_9397,N_9393);
nand U9484 (N_9484,N_9327,N_9382);
nand U9485 (N_9485,N_9369,N_9381);
and U9486 (N_9486,N_9301,N_9344);
nand U9487 (N_9487,N_9337,N_9308);
nor U9488 (N_9488,N_9322,N_9371);
nor U9489 (N_9489,N_9326,N_9396);
nand U9490 (N_9490,N_9384,N_9350);
nor U9491 (N_9491,N_9364,N_9387);
and U9492 (N_9492,N_9369,N_9345);
nor U9493 (N_9493,N_9328,N_9345);
nor U9494 (N_9494,N_9311,N_9368);
and U9495 (N_9495,N_9392,N_9367);
nand U9496 (N_9496,N_9337,N_9309);
nand U9497 (N_9497,N_9357,N_9383);
nor U9498 (N_9498,N_9324,N_9372);
or U9499 (N_9499,N_9315,N_9388);
nor U9500 (N_9500,N_9447,N_9406);
nor U9501 (N_9501,N_9450,N_9471);
or U9502 (N_9502,N_9454,N_9445);
nor U9503 (N_9503,N_9446,N_9459);
nand U9504 (N_9504,N_9462,N_9418);
or U9505 (N_9505,N_9494,N_9496);
nor U9506 (N_9506,N_9405,N_9475);
and U9507 (N_9507,N_9497,N_9419);
and U9508 (N_9508,N_9473,N_9490);
nor U9509 (N_9509,N_9439,N_9424);
and U9510 (N_9510,N_9434,N_9493);
and U9511 (N_9511,N_9408,N_9440);
nand U9512 (N_9512,N_9432,N_9448);
and U9513 (N_9513,N_9441,N_9469);
and U9514 (N_9514,N_9489,N_9423);
or U9515 (N_9515,N_9400,N_9435);
nor U9516 (N_9516,N_9427,N_9498);
nor U9517 (N_9517,N_9437,N_9422);
xor U9518 (N_9518,N_9492,N_9455);
nor U9519 (N_9519,N_9453,N_9478);
and U9520 (N_9520,N_9463,N_9438);
nand U9521 (N_9521,N_9425,N_9409);
and U9522 (N_9522,N_9480,N_9429);
nand U9523 (N_9523,N_9468,N_9414);
and U9524 (N_9524,N_9402,N_9464);
nand U9525 (N_9525,N_9484,N_9458);
and U9526 (N_9526,N_9495,N_9499);
nor U9527 (N_9527,N_9460,N_9465);
or U9528 (N_9528,N_9482,N_9428);
nor U9529 (N_9529,N_9443,N_9470);
nand U9530 (N_9530,N_9485,N_9413);
and U9531 (N_9531,N_9410,N_9404);
or U9532 (N_9532,N_9436,N_9415);
nand U9533 (N_9533,N_9444,N_9472);
or U9534 (N_9534,N_9401,N_9451);
nand U9535 (N_9535,N_9461,N_9466);
nand U9536 (N_9536,N_9476,N_9426);
nor U9537 (N_9537,N_9431,N_9483);
nor U9538 (N_9538,N_9491,N_9412);
nand U9539 (N_9539,N_9474,N_9477);
nand U9540 (N_9540,N_9486,N_9481);
and U9541 (N_9541,N_9442,N_9417);
nand U9542 (N_9542,N_9467,N_9449);
nand U9543 (N_9543,N_9487,N_9420);
and U9544 (N_9544,N_9479,N_9456);
nor U9545 (N_9545,N_9488,N_9411);
or U9546 (N_9546,N_9403,N_9421);
nand U9547 (N_9547,N_9416,N_9433);
nand U9548 (N_9548,N_9407,N_9457);
nor U9549 (N_9549,N_9430,N_9452);
or U9550 (N_9550,N_9447,N_9410);
or U9551 (N_9551,N_9477,N_9409);
nor U9552 (N_9552,N_9489,N_9477);
nand U9553 (N_9553,N_9404,N_9488);
and U9554 (N_9554,N_9449,N_9471);
and U9555 (N_9555,N_9474,N_9439);
and U9556 (N_9556,N_9415,N_9485);
nand U9557 (N_9557,N_9418,N_9466);
and U9558 (N_9558,N_9410,N_9475);
xnor U9559 (N_9559,N_9451,N_9478);
nor U9560 (N_9560,N_9466,N_9499);
nor U9561 (N_9561,N_9416,N_9408);
nor U9562 (N_9562,N_9458,N_9482);
nand U9563 (N_9563,N_9403,N_9409);
or U9564 (N_9564,N_9423,N_9407);
or U9565 (N_9565,N_9442,N_9489);
or U9566 (N_9566,N_9426,N_9492);
nand U9567 (N_9567,N_9484,N_9415);
and U9568 (N_9568,N_9437,N_9410);
and U9569 (N_9569,N_9495,N_9489);
xnor U9570 (N_9570,N_9477,N_9415);
nand U9571 (N_9571,N_9427,N_9424);
or U9572 (N_9572,N_9445,N_9481);
or U9573 (N_9573,N_9446,N_9473);
nand U9574 (N_9574,N_9491,N_9477);
nor U9575 (N_9575,N_9410,N_9467);
nor U9576 (N_9576,N_9457,N_9414);
nor U9577 (N_9577,N_9489,N_9451);
nand U9578 (N_9578,N_9402,N_9479);
or U9579 (N_9579,N_9443,N_9486);
and U9580 (N_9580,N_9495,N_9411);
and U9581 (N_9581,N_9425,N_9458);
and U9582 (N_9582,N_9455,N_9460);
nand U9583 (N_9583,N_9411,N_9462);
or U9584 (N_9584,N_9421,N_9463);
or U9585 (N_9585,N_9409,N_9435);
and U9586 (N_9586,N_9463,N_9465);
and U9587 (N_9587,N_9419,N_9484);
nand U9588 (N_9588,N_9444,N_9496);
or U9589 (N_9589,N_9457,N_9441);
nand U9590 (N_9590,N_9487,N_9401);
nand U9591 (N_9591,N_9491,N_9471);
or U9592 (N_9592,N_9433,N_9471);
nor U9593 (N_9593,N_9409,N_9474);
nor U9594 (N_9594,N_9453,N_9468);
nor U9595 (N_9595,N_9431,N_9442);
and U9596 (N_9596,N_9499,N_9412);
nor U9597 (N_9597,N_9405,N_9449);
nand U9598 (N_9598,N_9467,N_9486);
and U9599 (N_9599,N_9443,N_9412);
and U9600 (N_9600,N_9596,N_9563);
or U9601 (N_9601,N_9578,N_9534);
and U9602 (N_9602,N_9546,N_9583);
and U9603 (N_9603,N_9577,N_9528);
or U9604 (N_9604,N_9530,N_9586);
nand U9605 (N_9605,N_9574,N_9514);
and U9606 (N_9606,N_9590,N_9544);
and U9607 (N_9607,N_9597,N_9543);
nor U9608 (N_9608,N_9562,N_9553);
or U9609 (N_9609,N_9592,N_9554);
nand U9610 (N_9610,N_9556,N_9510);
and U9611 (N_9611,N_9505,N_9567);
nand U9612 (N_9612,N_9513,N_9575);
xnor U9613 (N_9613,N_9519,N_9584);
nor U9614 (N_9614,N_9509,N_9570);
and U9615 (N_9615,N_9542,N_9595);
nand U9616 (N_9616,N_9520,N_9581);
or U9617 (N_9617,N_9555,N_9517);
nor U9618 (N_9618,N_9536,N_9593);
nand U9619 (N_9619,N_9591,N_9532);
nor U9620 (N_9620,N_9540,N_9525);
and U9621 (N_9621,N_9535,N_9568);
nand U9622 (N_9622,N_9569,N_9518);
nand U9623 (N_9623,N_9582,N_9557);
or U9624 (N_9624,N_9522,N_9539);
xor U9625 (N_9625,N_9526,N_9560);
nor U9626 (N_9626,N_9571,N_9566);
and U9627 (N_9627,N_9580,N_9527);
nand U9628 (N_9628,N_9588,N_9523);
or U9629 (N_9629,N_9524,N_9552);
and U9630 (N_9630,N_9558,N_9594);
and U9631 (N_9631,N_9598,N_9599);
nor U9632 (N_9632,N_9529,N_9585);
and U9633 (N_9633,N_9589,N_9500);
nor U9634 (N_9634,N_9515,N_9506);
and U9635 (N_9635,N_9502,N_9508);
or U9636 (N_9636,N_9561,N_9576);
nand U9637 (N_9637,N_9573,N_9511);
or U9638 (N_9638,N_9507,N_9533);
or U9639 (N_9639,N_9572,N_9521);
and U9640 (N_9640,N_9512,N_9564);
nand U9641 (N_9641,N_9541,N_9503);
and U9642 (N_9642,N_9545,N_9516);
nand U9643 (N_9643,N_9587,N_9579);
and U9644 (N_9644,N_9538,N_9504);
nor U9645 (N_9645,N_9537,N_9565);
nand U9646 (N_9646,N_9501,N_9549);
or U9647 (N_9647,N_9559,N_9547);
nand U9648 (N_9648,N_9550,N_9551);
nor U9649 (N_9649,N_9548,N_9531);
nand U9650 (N_9650,N_9578,N_9553);
nor U9651 (N_9651,N_9576,N_9523);
or U9652 (N_9652,N_9579,N_9576);
nor U9653 (N_9653,N_9526,N_9513);
nor U9654 (N_9654,N_9572,N_9516);
nand U9655 (N_9655,N_9538,N_9536);
nor U9656 (N_9656,N_9544,N_9525);
or U9657 (N_9657,N_9527,N_9598);
xnor U9658 (N_9658,N_9529,N_9507);
nor U9659 (N_9659,N_9517,N_9536);
nor U9660 (N_9660,N_9580,N_9514);
nor U9661 (N_9661,N_9587,N_9569);
nor U9662 (N_9662,N_9512,N_9591);
nand U9663 (N_9663,N_9540,N_9596);
nor U9664 (N_9664,N_9523,N_9579);
nand U9665 (N_9665,N_9573,N_9546);
or U9666 (N_9666,N_9525,N_9557);
xor U9667 (N_9667,N_9532,N_9542);
and U9668 (N_9668,N_9570,N_9510);
nand U9669 (N_9669,N_9593,N_9528);
nor U9670 (N_9670,N_9568,N_9592);
nor U9671 (N_9671,N_9591,N_9520);
nand U9672 (N_9672,N_9584,N_9520);
nor U9673 (N_9673,N_9523,N_9567);
and U9674 (N_9674,N_9543,N_9548);
or U9675 (N_9675,N_9515,N_9559);
nand U9676 (N_9676,N_9553,N_9534);
and U9677 (N_9677,N_9572,N_9507);
or U9678 (N_9678,N_9578,N_9567);
nor U9679 (N_9679,N_9530,N_9538);
or U9680 (N_9680,N_9515,N_9522);
nand U9681 (N_9681,N_9593,N_9567);
or U9682 (N_9682,N_9559,N_9516);
or U9683 (N_9683,N_9586,N_9578);
or U9684 (N_9684,N_9587,N_9556);
nand U9685 (N_9685,N_9555,N_9542);
nand U9686 (N_9686,N_9560,N_9545);
or U9687 (N_9687,N_9593,N_9543);
xor U9688 (N_9688,N_9594,N_9504);
nand U9689 (N_9689,N_9524,N_9537);
or U9690 (N_9690,N_9567,N_9551);
and U9691 (N_9691,N_9514,N_9598);
nor U9692 (N_9692,N_9599,N_9511);
xor U9693 (N_9693,N_9529,N_9570);
nor U9694 (N_9694,N_9575,N_9538);
nand U9695 (N_9695,N_9574,N_9569);
or U9696 (N_9696,N_9561,N_9572);
or U9697 (N_9697,N_9522,N_9599);
nor U9698 (N_9698,N_9588,N_9551);
nand U9699 (N_9699,N_9510,N_9504);
nor U9700 (N_9700,N_9673,N_9698);
nor U9701 (N_9701,N_9635,N_9610);
or U9702 (N_9702,N_9615,N_9674);
and U9703 (N_9703,N_9617,N_9622);
nand U9704 (N_9704,N_9600,N_9616);
nand U9705 (N_9705,N_9631,N_9644);
and U9706 (N_9706,N_9697,N_9661);
nand U9707 (N_9707,N_9602,N_9647);
nand U9708 (N_9708,N_9672,N_9684);
nand U9709 (N_9709,N_9607,N_9683);
or U9710 (N_9710,N_9660,N_9687);
nand U9711 (N_9711,N_9652,N_9629);
nand U9712 (N_9712,N_9667,N_9628);
nor U9713 (N_9713,N_9664,N_9696);
nor U9714 (N_9714,N_9653,N_9680);
nand U9715 (N_9715,N_9638,N_9608);
nor U9716 (N_9716,N_9605,N_9636);
and U9717 (N_9717,N_9686,N_9682);
or U9718 (N_9718,N_9675,N_9627);
or U9719 (N_9719,N_9601,N_9625);
xnor U9720 (N_9720,N_9630,N_9655);
nand U9721 (N_9721,N_9671,N_9603);
nor U9722 (N_9722,N_9695,N_9663);
nor U9723 (N_9723,N_9621,N_9678);
nand U9724 (N_9724,N_9699,N_9623);
nand U9725 (N_9725,N_9609,N_9619);
nor U9726 (N_9726,N_9659,N_9688);
and U9727 (N_9727,N_9606,N_9618);
or U9728 (N_9728,N_9692,N_9677);
or U9729 (N_9729,N_9694,N_9668);
xnor U9730 (N_9730,N_9611,N_9657);
or U9731 (N_9731,N_9689,N_9658);
and U9732 (N_9732,N_9633,N_9650);
nand U9733 (N_9733,N_9639,N_9666);
nor U9734 (N_9734,N_9651,N_9679);
and U9735 (N_9735,N_9656,N_9648);
and U9736 (N_9736,N_9640,N_9690);
or U9737 (N_9737,N_9614,N_9670);
nand U9738 (N_9738,N_9685,N_9612);
and U9739 (N_9739,N_9676,N_9646);
and U9740 (N_9740,N_9654,N_9634);
and U9741 (N_9741,N_9669,N_9649);
nand U9742 (N_9742,N_9613,N_9665);
and U9743 (N_9743,N_9645,N_9641);
and U9744 (N_9744,N_9620,N_9624);
and U9745 (N_9745,N_9662,N_9643);
and U9746 (N_9746,N_9637,N_9604);
nor U9747 (N_9747,N_9693,N_9626);
nor U9748 (N_9748,N_9642,N_9681);
and U9749 (N_9749,N_9632,N_9691);
nand U9750 (N_9750,N_9655,N_9644);
or U9751 (N_9751,N_9616,N_9601);
nor U9752 (N_9752,N_9652,N_9637);
nor U9753 (N_9753,N_9686,N_9681);
or U9754 (N_9754,N_9603,N_9670);
nand U9755 (N_9755,N_9604,N_9648);
and U9756 (N_9756,N_9649,N_9661);
or U9757 (N_9757,N_9698,N_9643);
nor U9758 (N_9758,N_9686,N_9658);
and U9759 (N_9759,N_9651,N_9615);
nor U9760 (N_9760,N_9618,N_9634);
nand U9761 (N_9761,N_9678,N_9647);
or U9762 (N_9762,N_9636,N_9611);
or U9763 (N_9763,N_9664,N_9612);
nand U9764 (N_9764,N_9646,N_9615);
and U9765 (N_9765,N_9605,N_9607);
nor U9766 (N_9766,N_9653,N_9691);
nand U9767 (N_9767,N_9604,N_9619);
or U9768 (N_9768,N_9602,N_9648);
or U9769 (N_9769,N_9623,N_9686);
xnor U9770 (N_9770,N_9673,N_9605);
or U9771 (N_9771,N_9676,N_9628);
or U9772 (N_9772,N_9623,N_9679);
or U9773 (N_9773,N_9637,N_9649);
or U9774 (N_9774,N_9631,N_9614);
nor U9775 (N_9775,N_9628,N_9695);
and U9776 (N_9776,N_9644,N_9621);
nand U9777 (N_9777,N_9671,N_9655);
nor U9778 (N_9778,N_9692,N_9603);
nor U9779 (N_9779,N_9643,N_9644);
nor U9780 (N_9780,N_9648,N_9654);
or U9781 (N_9781,N_9632,N_9642);
or U9782 (N_9782,N_9689,N_9650);
or U9783 (N_9783,N_9637,N_9618);
nor U9784 (N_9784,N_9652,N_9610);
nand U9785 (N_9785,N_9638,N_9676);
nor U9786 (N_9786,N_9662,N_9698);
nor U9787 (N_9787,N_9697,N_9635);
nor U9788 (N_9788,N_9682,N_9664);
nand U9789 (N_9789,N_9678,N_9639);
nand U9790 (N_9790,N_9616,N_9644);
and U9791 (N_9791,N_9671,N_9696);
and U9792 (N_9792,N_9639,N_9654);
nand U9793 (N_9793,N_9659,N_9668);
and U9794 (N_9794,N_9615,N_9675);
or U9795 (N_9795,N_9630,N_9658);
and U9796 (N_9796,N_9657,N_9689);
nor U9797 (N_9797,N_9633,N_9667);
nor U9798 (N_9798,N_9693,N_9621);
and U9799 (N_9799,N_9661,N_9692);
and U9800 (N_9800,N_9746,N_9726);
and U9801 (N_9801,N_9790,N_9753);
nor U9802 (N_9802,N_9757,N_9798);
nor U9803 (N_9803,N_9719,N_9724);
and U9804 (N_9804,N_9727,N_9720);
nand U9805 (N_9805,N_9789,N_9766);
nand U9806 (N_9806,N_9763,N_9751);
or U9807 (N_9807,N_9742,N_9799);
nor U9808 (N_9808,N_9722,N_9732);
nor U9809 (N_9809,N_9749,N_9796);
and U9810 (N_9810,N_9738,N_9750);
or U9811 (N_9811,N_9736,N_9785);
or U9812 (N_9812,N_9780,N_9723);
or U9813 (N_9813,N_9755,N_9758);
or U9814 (N_9814,N_9787,N_9747);
nand U9815 (N_9815,N_9729,N_9756);
nor U9816 (N_9816,N_9769,N_9706);
or U9817 (N_9817,N_9725,N_9788);
nand U9818 (N_9818,N_9733,N_9784);
or U9819 (N_9819,N_9771,N_9794);
or U9820 (N_9820,N_9739,N_9793);
or U9821 (N_9821,N_9744,N_9707);
or U9822 (N_9822,N_9735,N_9705);
nor U9823 (N_9823,N_9792,N_9737);
or U9824 (N_9824,N_9700,N_9712);
or U9825 (N_9825,N_9731,N_9743);
nand U9826 (N_9826,N_9754,N_9734);
nand U9827 (N_9827,N_9721,N_9762);
nand U9828 (N_9828,N_9709,N_9718);
nand U9829 (N_9829,N_9759,N_9777);
nand U9830 (N_9830,N_9761,N_9702);
and U9831 (N_9831,N_9740,N_9748);
nor U9832 (N_9832,N_9713,N_9770);
nor U9833 (N_9833,N_9710,N_9781);
and U9834 (N_9834,N_9714,N_9768);
and U9835 (N_9835,N_9717,N_9773);
nor U9836 (N_9836,N_9730,N_9765);
or U9837 (N_9837,N_9752,N_9779);
nand U9838 (N_9838,N_9711,N_9786);
or U9839 (N_9839,N_9745,N_9795);
and U9840 (N_9840,N_9791,N_9704);
nor U9841 (N_9841,N_9716,N_9775);
nand U9842 (N_9842,N_9772,N_9767);
or U9843 (N_9843,N_9741,N_9797);
nand U9844 (N_9844,N_9776,N_9728);
nand U9845 (N_9845,N_9778,N_9708);
nor U9846 (N_9846,N_9701,N_9760);
or U9847 (N_9847,N_9715,N_9783);
nand U9848 (N_9848,N_9764,N_9774);
nor U9849 (N_9849,N_9703,N_9782);
nand U9850 (N_9850,N_9733,N_9799);
or U9851 (N_9851,N_9767,N_9795);
and U9852 (N_9852,N_9783,N_9794);
and U9853 (N_9853,N_9724,N_9705);
nand U9854 (N_9854,N_9722,N_9753);
nor U9855 (N_9855,N_9717,N_9780);
or U9856 (N_9856,N_9738,N_9705);
nand U9857 (N_9857,N_9793,N_9794);
and U9858 (N_9858,N_9780,N_9788);
nand U9859 (N_9859,N_9792,N_9755);
or U9860 (N_9860,N_9782,N_9763);
and U9861 (N_9861,N_9720,N_9733);
or U9862 (N_9862,N_9707,N_9713);
nor U9863 (N_9863,N_9796,N_9759);
and U9864 (N_9864,N_9727,N_9738);
or U9865 (N_9865,N_9714,N_9730);
nand U9866 (N_9866,N_9774,N_9737);
nor U9867 (N_9867,N_9761,N_9778);
and U9868 (N_9868,N_9794,N_9738);
nor U9869 (N_9869,N_9761,N_9730);
or U9870 (N_9870,N_9731,N_9720);
nand U9871 (N_9871,N_9711,N_9701);
nor U9872 (N_9872,N_9704,N_9773);
or U9873 (N_9873,N_9795,N_9751);
nor U9874 (N_9874,N_9719,N_9785);
or U9875 (N_9875,N_9784,N_9751);
or U9876 (N_9876,N_9765,N_9798);
nor U9877 (N_9877,N_9718,N_9793);
nor U9878 (N_9878,N_9780,N_9790);
nand U9879 (N_9879,N_9772,N_9779);
xnor U9880 (N_9880,N_9784,N_9745);
nor U9881 (N_9881,N_9724,N_9756);
xnor U9882 (N_9882,N_9785,N_9765);
or U9883 (N_9883,N_9786,N_9731);
nor U9884 (N_9884,N_9753,N_9760);
and U9885 (N_9885,N_9765,N_9745);
nor U9886 (N_9886,N_9765,N_9799);
or U9887 (N_9887,N_9782,N_9759);
nand U9888 (N_9888,N_9770,N_9731);
and U9889 (N_9889,N_9730,N_9721);
or U9890 (N_9890,N_9706,N_9732);
nor U9891 (N_9891,N_9789,N_9742);
nor U9892 (N_9892,N_9765,N_9750);
or U9893 (N_9893,N_9734,N_9767);
nor U9894 (N_9894,N_9702,N_9756);
and U9895 (N_9895,N_9797,N_9788);
or U9896 (N_9896,N_9720,N_9791);
nand U9897 (N_9897,N_9760,N_9710);
and U9898 (N_9898,N_9740,N_9757);
nand U9899 (N_9899,N_9720,N_9708);
and U9900 (N_9900,N_9815,N_9810);
or U9901 (N_9901,N_9807,N_9863);
or U9902 (N_9902,N_9864,N_9893);
nor U9903 (N_9903,N_9817,N_9845);
and U9904 (N_9904,N_9891,N_9876);
or U9905 (N_9905,N_9899,N_9895);
nor U9906 (N_9906,N_9882,N_9883);
nand U9907 (N_9907,N_9805,N_9831);
or U9908 (N_9908,N_9875,N_9846);
nand U9909 (N_9909,N_9861,N_9833);
and U9910 (N_9910,N_9854,N_9821);
nand U9911 (N_9911,N_9851,N_9850);
nor U9912 (N_9912,N_9824,N_9849);
nor U9913 (N_9913,N_9859,N_9887);
or U9914 (N_9914,N_9865,N_9852);
nor U9915 (N_9915,N_9812,N_9803);
and U9916 (N_9916,N_9808,N_9804);
nand U9917 (N_9917,N_9890,N_9809);
and U9918 (N_9918,N_9870,N_9838);
nand U9919 (N_9919,N_9836,N_9889);
and U9920 (N_9920,N_9878,N_9813);
nor U9921 (N_9921,N_9818,N_9869);
or U9922 (N_9922,N_9877,N_9829);
nand U9923 (N_9923,N_9819,N_9844);
or U9924 (N_9924,N_9847,N_9832);
or U9925 (N_9925,N_9814,N_9885);
nor U9926 (N_9926,N_9834,N_9879);
or U9927 (N_9927,N_9894,N_9839);
and U9928 (N_9928,N_9873,N_9841);
nand U9929 (N_9929,N_9886,N_9897);
and U9930 (N_9930,N_9880,N_9896);
or U9931 (N_9931,N_9881,N_9872);
and U9932 (N_9932,N_9858,N_9806);
and U9933 (N_9933,N_9842,N_9898);
nor U9934 (N_9934,N_9825,N_9840);
nand U9935 (N_9935,N_9828,N_9826);
nand U9936 (N_9936,N_9827,N_9800);
or U9937 (N_9937,N_9862,N_9892);
nor U9938 (N_9938,N_9822,N_9811);
nor U9939 (N_9939,N_9866,N_9837);
nor U9940 (N_9940,N_9867,N_9856);
nand U9941 (N_9941,N_9843,N_9874);
nand U9942 (N_9942,N_9830,N_9820);
nand U9943 (N_9943,N_9888,N_9801);
nand U9944 (N_9944,N_9855,N_9860);
and U9945 (N_9945,N_9853,N_9835);
or U9946 (N_9946,N_9868,N_9848);
nor U9947 (N_9947,N_9823,N_9871);
or U9948 (N_9948,N_9884,N_9802);
nand U9949 (N_9949,N_9816,N_9857);
nor U9950 (N_9950,N_9859,N_9806);
or U9951 (N_9951,N_9881,N_9873);
nor U9952 (N_9952,N_9803,N_9842);
and U9953 (N_9953,N_9837,N_9819);
xor U9954 (N_9954,N_9889,N_9839);
and U9955 (N_9955,N_9885,N_9812);
and U9956 (N_9956,N_9871,N_9869);
xnor U9957 (N_9957,N_9871,N_9809);
nor U9958 (N_9958,N_9815,N_9892);
or U9959 (N_9959,N_9890,N_9862);
nor U9960 (N_9960,N_9866,N_9863);
or U9961 (N_9961,N_9809,N_9826);
or U9962 (N_9962,N_9827,N_9851);
or U9963 (N_9963,N_9803,N_9872);
xnor U9964 (N_9964,N_9851,N_9848);
and U9965 (N_9965,N_9855,N_9834);
nand U9966 (N_9966,N_9840,N_9873);
nand U9967 (N_9967,N_9804,N_9815);
or U9968 (N_9968,N_9834,N_9870);
and U9969 (N_9969,N_9807,N_9820);
and U9970 (N_9970,N_9831,N_9881);
and U9971 (N_9971,N_9829,N_9845);
nor U9972 (N_9972,N_9840,N_9866);
nand U9973 (N_9973,N_9899,N_9853);
and U9974 (N_9974,N_9812,N_9865);
nor U9975 (N_9975,N_9803,N_9809);
nand U9976 (N_9976,N_9800,N_9896);
and U9977 (N_9977,N_9878,N_9852);
and U9978 (N_9978,N_9881,N_9854);
or U9979 (N_9979,N_9850,N_9806);
xnor U9980 (N_9980,N_9845,N_9897);
or U9981 (N_9981,N_9817,N_9814);
or U9982 (N_9982,N_9857,N_9820);
nand U9983 (N_9983,N_9883,N_9862);
nor U9984 (N_9984,N_9848,N_9864);
nand U9985 (N_9985,N_9893,N_9851);
or U9986 (N_9986,N_9814,N_9858);
nor U9987 (N_9987,N_9802,N_9821);
and U9988 (N_9988,N_9868,N_9880);
xnor U9989 (N_9989,N_9895,N_9873);
nor U9990 (N_9990,N_9879,N_9893);
and U9991 (N_9991,N_9854,N_9893);
nand U9992 (N_9992,N_9849,N_9800);
and U9993 (N_9993,N_9859,N_9889);
nand U9994 (N_9994,N_9883,N_9821);
and U9995 (N_9995,N_9830,N_9823);
and U9996 (N_9996,N_9835,N_9802);
nor U9997 (N_9997,N_9821,N_9839);
xnor U9998 (N_9998,N_9846,N_9816);
nor U9999 (N_9999,N_9898,N_9888);
nor UO_0 (O_0,N_9938,N_9918);
nor UO_1 (O_1,N_9994,N_9991);
and UO_2 (O_2,N_9959,N_9951);
and UO_3 (O_3,N_9921,N_9913);
or UO_4 (O_4,N_9929,N_9956);
or UO_5 (O_5,N_9923,N_9903);
nand UO_6 (O_6,N_9963,N_9926);
nor UO_7 (O_7,N_9946,N_9932);
xor UO_8 (O_8,N_9949,N_9933);
nor UO_9 (O_9,N_9955,N_9945);
and UO_10 (O_10,N_9998,N_9999);
nand UO_11 (O_11,N_9941,N_9964);
and UO_12 (O_12,N_9937,N_9967);
and UO_13 (O_13,N_9952,N_9920);
nand UO_14 (O_14,N_9906,N_9900);
or UO_15 (O_15,N_9960,N_9910);
and UO_16 (O_16,N_9993,N_9931);
and UO_17 (O_17,N_9977,N_9995);
and UO_18 (O_18,N_9904,N_9980);
nor UO_19 (O_19,N_9939,N_9979);
or UO_20 (O_20,N_9901,N_9916);
or UO_21 (O_21,N_9909,N_9930);
or UO_22 (O_22,N_9953,N_9992);
or UO_23 (O_23,N_9975,N_9950);
nand UO_24 (O_24,N_9917,N_9924);
nor UO_25 (O_25,N_9987,N_9912);
or UO_26 (O_26,N_9982,N_9974);
nand UO_27 (O_27,N_9997,N_9905);
nand UO_28 (O_28,N_9973,N_9957);
and UO_29 (O_29,N_9915,N_9971);
nor UO_30 (O_30,N_9948,N_9947);
nand UO_31 (O_31,N_9970,N_9976);
or UO_32 (O_32,N_9928,N_9943);
or UO_33 (O_33,N_9968,N_9940);
nor UO_34 (O_34,N_9966,N_9908);
or UO_35 (O_35,N_9914,N_9907);
nor UO_36 (O_36,N_9983,N_9935);
and UO_37 (O_37,N_9936,N_9965);
nor UO_38 (O_38,N_9988,N_9981);
nor UO_39 (O_39,N_9927,N_9962);
or UO_40 (O_40,N_9984,N_9911);
or UO_41 (O_41,N_9919,N_9961);
or UO_42 (O_42,N_9958,N_9972);
or UO_43 (O_43,N_9902,N_9978);
nand UO_44 (O_44,N_9942,N_9954);
nor UO_45 (O_45,N_9934,N_9969);
or UO_46 (O_46,N_9985,N_9925);
and UO_47 (O_47,N_9989,N_9986);
nor UO_48 (O_48,N_9944,N_9990);
and UO_49 (O_49,N_9996,N_9922);
or UO_50 (O_50,N_9932,N_9985);
nand UO_51 (O_51,N_9994,N_9941);
nand UO_52 (O_52,N_9943,N_9965);
nor UO_53 (O_53,N_9951,N_9969);
or UO_54 (O_54,N_9954,N_9952);
nand UO_55 (O_55,N_9966,N_9991);
and UO_56 (O_56,N_9923,N_9988);
or UO_57 (O_57,N_9966,N_9996);
and UO_58 (O_58,N_9942,N_9982);
nand UO_59 (O_59,N_9973,N_9974);
nand UO_60 (O_60,N_9954,N_9939);
or UO_61 (O_61,N_9936,N_9969);
or UO_62 (O_62,N_9952,N_9991);
and UO_63 (O_63,N_9944,N_9953);
nand UO_64 (O_64,N_9976,N_9919);
and UO_65 (O_65,N_9962,N_9973);
xor UO_66 (O_66,N_9965,N_9935);
and UO_67 (O_67,N_9971,N_9950);
nand UO_68 (O_68,N_9912,N_9996);
and UO_69 (O_69,N_9944,N_9972);
nand UO_70 (O_70,N_9900,N_9927);
or UO_71 (O_71,N_9975,N_9920);
or UO_72 (O_72,N_9992,N_9970);
and UO_73 (O_73,N_9982,N_9997);
nand UO_74 (O_74,N_9910,N_9920);
nor UO_75 (O_75,N_9993,N_9988);
nand UO_76 (O_76,N_9990,N_9954);
nand UO_77 (O_77,N_9967,N_9906);
nand UO_78 (O_78,N_9951,N_9949);
and UO_79 (O_79,N_9963,N_9990);
nand UO_80 (O_80,N_9968,N_9900);
or UO_81 (O_81,N_9938,N_9961);
nor UO_82 (O_82,N_9996,N_9987);
nor UO_83 (O_83,N_9975,N_9932);
nand UO_84 (O_84,N_9921,N_9949);
or UO_85 (O_85,N_9946,N_9949);
and UO_86 (O_86,N_9908,N_9955);
nor UO_87 (O_87,N_9962,N_9996);
nor UO_88 (O_88,N_9969,N_9948);
nand UO_89 (O_89,N_9990,N_9927);
and UO_90 (O_90,N_9946,N_9927);
nand UO_91 (O_91,N_9960,N_9956);
and UO_92 (O_92,N_9904,N_9901);
xnor UO_93 (O_93,N_9913,N_9984);
nand UO_94 (O_94,N_9907,N_9936);
and UO_95 (O_95,N_9945,N_9916);
or UO_96 (O_96,N_9943,N_9974);
and UO_97 (O_97,N_9912,N_9960);
and UO_98 (O_98,N_9938,N_9928);
or UO_99 (O_99,N_9979,N_9905);
or UO_100 (O_100,N_9971,N_9933);
nor UO_101 (O_101,N_9903,N_9937);
and UO_102 (O_102,N_9969,N_9984);
nand UO_103 (O_103,N_9952,N_9906);
or UO_104 (O_104,N_9962,N_9904);
and UO_105 (O_105,N_9947,N_9999);
and UO_106 (O_106,N_9999,N_9955);
and UO_107 (O_107,N_9933,N_9929);
or UO_108 (O_108,N_9909,N_9911);
xor UO_109 (O_109,N_9977,N_9955);
and UO_110 (O_110,N_9914,N_9947);
or UO_111 (O_111,N_9997,N_9957);
or UO_112 (O_112,N_9945,N_9914);
nand UO_113 (O_113,N_9991,N_9919);
nand UO_114 (O_114,N_9951,N_9942);
nand UO_115 (O_115,N_9900,N_9985);
and UO_116 (O_116,N_9909,N_9971);
nand UO_117 (O_117,N_9949,N_9945);
nand UO_118 (O_118,N_9946,N_9992);
nor UO_119 (O_119,N_9903,N_9913);
nor UO_120 (O_120,N_9952,N_9932);
nor UO_121 (O_121,N_9915,N_9980);
nand UO_122 (O_122,N_9946,N_9987);
nor UO_123 (O_123,N_9976,N_9903);
or UO_124 (O_124,N_9977,N_9926);
and UO_125 (O_125,N_9998,N_9946);
or UO_126 (O_126,N_9964,N_9987);
and UO_127 (O_127,N_9956,N_9948);
nor UO_128 (O_128,N_9996,N_9951);
or UO_129 (O_129,N_9944,N_9986);
nor UO_130 (O_130,N_9946,N_9938);
or UO_131 (O_131,N_9932,N_9990);
xnor UO_132 (O_132,N_9964,N_9914);
and UO_133 (O_133,N_9940,N_9912);
or UO_134 (O_134,N_9967,N_9924);
or UO_135 (O_135,N_9963,N_9985);
and UO_136 (O_136,N_9962,N_9966);
nand UO_137 (O_137,N_9937,N_9981);
nand UO_138 (O_138,N_9935,N_9905);
or UO_139 (O_139,N_9952,N_9992);
or UO_140 (O_140,N_9987,N_9989);
and UO_141 (O_141,N_9942,N_9925);
or UO_142 (O_142,N_9905,N_9901);
or UO_143 (O_143,N_9995,N_9991);
xor UO_144 (O_144,N_9978,N_9956);
and UO_145 (O_145,N_9961,N_9977);
nand UO_146 (O_146,N_9947,N_9966);
nand UO_147 (O_147,N_9947,N_9949);
or UO_148 (O_148,N_9950,N_9946);
nor UO_149 (O_149,N_9918,N_9920);
nor UO_150 (O_150,N_9921,N_9972);
nor UO_151 (O_151,N_9917,N_9999);
and UO_152 (O_152,N_9990,N_9900);
nand UO_153 (O_153,N_9939,N_9984);
xnor UO_154 (O_154,N_9900,N_9989);
and UO_155 (O_155,N_9960,N_9911);
nand UO_156 (O_156,N_9911,N_9964);
nand UO_157 (O_157,N_9957,N_9940);
nor UO_158 (O_158,N_9958,N_9994);
nor UO_159 (O_159,N_9940,N_9948);
nor UO_160 (O_160,N_9983,N_9945);
nor UO_161 (O_161,N_9910,N_9955);
or UO_162 (O_162,N_9981,N_9942);
nor UO_163 (O_163,N_9912,N_9958);
or UO_164 (O_164,N_9954,N_9959);
or UO_165 (O_165,N_9992,N_9965);
nand UO_166 (O_166,N_9944,N_9985);
and UO_167 (O_167,N_9946,N_9901);
nand UO_168 (O_168,N_9930,N_9926);
nor UO_169 (O_169,N_9976,N_9942);
nor UO_170 (O_170,N_9968,N_9999);
nor UO_171 (O_171,N_9907,N_9960);
nand UO_172 (O_172,N_9956,N_9925);
nand UO_173 (O_173,N_9971,N_9910);
and UO_174 (O_174,N_9979,N_9901);
and UO_175 (O_175,N_9988,N_9990);
nor UO_176 (O_176,N_9988,N_9955);
and UO_177 (O_177,N_9943,N_9927);
nor UO_178 (O_178,N_9985,N_9913);
nand UO_179 (O_179,N_9989,N_9907);
and UO_180 (O_180,N_9967,N_9909);
xnor UO_181 (O_181,N_9970,N_9969);
and UO_182 (O_182,N_9981,N_9966);
nor UO_183 (O_183,N_9979,N_9953);
nand UO_184 (O_184,N_9902,N_9982);
nor UO_185 (O_185,N_9983,N_9950);
nand UO_186 (O_186,N_9909,N_9910);
xor UO_187 (O_187,N_9933,N_9934);
or UO_188 (O_188,N_9951,N_9945);
nand UO_189 (O_189,N_9962,N_9992);
nor UO_190 (O_190,N_9902,N_9912);
nand UO_191 (O_191,N_9981,N_9918);
nand UO_192 (O_192,N_9975,N_9936);
or UO_193 (O_193,N_9993,N_9920);
or UO_194 (O_194,N_9958,N_9936);
and UO_195 (O_195,N_9910,N_9956);
and UO_196 (O_196,N_9964,N_9948);
nor UO_197 (O_197,N_9910,N_9970);
and UO_198 (O_198,N_9983,N_9967);
nand UO_199 (O_199,N_9949,N_9944);
nand UO_200 (O_200,N_9919,N_9964);
nor UO_201 (O_201,N_9967,N_9996);
nand UO_202 (O_202,N_9905,N_9987);
nand UO_203 (O_203,N_9959,N_9934);
nor UO_204 (O_204,N_9973,N_9950);
or UO_205 (O_205,N_9941,N_9912);
nor UO_206 (O_206,N_9923,N_9909);
nor UO_207 (O_207,N_9949,N_9909);
or UO_208 (O_208,N_9988,N_9926);
nor UO_209 (O_209,N_9966,N_9976);
nand UO_210 (O_210,N_9997,N_9932);
nand UO_211 (O_211,N_9986,N_9930);
or UO_212 (O_212,N_9965,N_9914);
nand UO_213 (O_213,N_9937,N_9949);
nand UO_214 (O_214,N_9936,N_9922);
or UO_215 (O_215,N_9969,N_9965);
and UO_216 (O_216,N_9939,N_9911);
and UO_217 (O_217,N_9923,N_9920);
or UO_218 (O_218,N_9975,N_9927);
and UO_219 (O_219,N_9985,N_9951);
and UO_220 (O_220,N_9977,N_9917);
nor UO_221 (O_221,N_9904,N_9995);
or UO_222 (O_222,N_9982,N_9985);
nor UO_223 (O_223,N_9943,N_9935);
nand UO_224 (O_224,N_9989,N_9939);
nor UO_225 (O_225,N_9939,N_9921);
nor UO_226 (O_226,N_9989,N_9990);
or UO_227 (O_227,N_9998,N_9902);
or UO_228 (O_228,N_9984,N_9926);
nand UO_229 (O_229,N_9908,N_9954);
or UO_230 (O_230,N_9925,N_9971);
or UO_231 (O_231,N_9941,N_9989);
or UO_232 (O_232,N_9925,N_9910);
nor UO_233 (O_233,N_9994,N_9943);
nand UO_234 (O_234,N_9974,N_9933);
or UO_235 (O_235,N_9975,N_9956);
and UO_236 (O_236,N_9963,N_9922);
nor UO_237 (O_237,N_9939,N_9918);
and UO_238 (O_238,N_9964,N_9900);
nor UO_239 (O_239,N_9998,N_9961);
nor UO_240 (O_240,N_9948,N_9972);
or UO_241 (O_241,N_9966,N_9935);
nand UO_242 (O_242,N_9975,N_9968);
nor UO_243 (O_243,N_9967,N_9970);
nor UO_244 (O_244,N_9916,N_9992);
or UO_245 (O_245,N_9901,N_9920);
nor UO_246 (O_246,N_9973,N_9903);
and UO_247 (O_247,N_9905,N_9967);
xnor UO_248 (O_248,N_9911,N_9973);
and UO_249 (O_249,N_9991,N_9906);
nor UO_250 (O_250,N_9964,N_9983);
nand UO_251 (O_251,N_9901,N_9902);
nor UO_252 (O_252,N_9988,N_9978);
and UO_253 (O_253,N_9999,N_9990);
nor UO_254 (O_254,N_9942,N_9966);
nand UO_255 (O_255,N_9980,N_9956);
nor UO_256 (O_256,N_9956,N_9981);
nand UO_257 (O_257,N_9937,N_9902);
nand UO_258 (O_258,N_9984,N_9973);
and UO_259 (O_259,N_9954,N_9927);
nor UO_260 (O_260,N_9976,N_9953);
nor UO_261 (O_261,N_9919,N_9939);
nand UO_262 (O_262,N_9924,N_9952);
nand UO_263 (O_263,N_9989,N_9954);
or UO_264 (O_264,N_9934,N_9925);
and UO_265 (O_265,N_9904,N_9931);
and UO_266 (O_266,N_9915,N_9963);
nand UO_267 (O_267,N_9986,N_9903);
nand UO_268 (O_268,N_9957,N_9955);
nor UO_269 (O_269,N_9967,N_9961);
nor UO_270 (O_270,N_9984,N_9946);
and UO_271 (O_271,N_9912,N_9980);
and UO_272 (O_272,N_9904,N_9985);
nand UO_273 (O_273,N_9927,N_9921);
and UO_274 (O_274,N_9967,N_9974);
or UO_275 (O_275,N_9993,N_9999);
and UO_276 (O_276,N_9969,N_9980);
nor UO_277 (O_277,N_9907,N_9963);
nand UO_278 (O_278,N_9989,N_9977);
xor UO_279 (O_279,N_9925,N_9991);
xor UO_280 (O_280,N_9918,N_9928);
or UO_281 (O_281,N_9979,N_9971);
or UO_282 (O_282,N_9922,N_9984);
nor UO_283 (O_283,N_9997,N_9966);
nor UO_284 (O_284,N_9925,N_9974);
or UO_285 (O_285,N_9925,N_9906);
nor UO_286 (O_286,N_9927,N_9903);
nor UO_287 (O_287,N_9923,N_9928);
and UO_288 (O_288,N_9904,N_9920);
nor UO_289 (O_289,N_9904,N_9954);
nand UO_290 (O_290,N_9962,N_9906);
and UO_291 (O_291,N_9969,N_9944);
and UO_292 (O_292,N_9965,N_9930);
nand UO_293 (O_293,N_9983,N_9966);
nor UO_294 (O_294,N_9914,N_9998);
or UO_295 (O_295,N_9928,N_9984);
or UO_296 (O_296,N_9912,N_9975);
or UO_297 (O_297,N_9908,N_9998);
and UO_298 (O_298,N_9936,N_9914);
or UO_299 (O_299,N_9931,N_9974);
nand UO_300 (O_300,N_9953,N_9915);
nand UO_301 (O_301,N_9918,N_9976);
nor UO_302 (O_302,N_9938,N_9966);
and UO_303 (O_303,N_9916,N_9928);
and UO_304 (O_304,N_9992,N_9907);
and UO_305 (O_305,N_9941,N_9932);
nor UO_306 (O_306,N_9939,N_9978);
nand UO_307 (O_307,N_9929,N_9905);
nor UO_308 (O_308,N_9937,N_9987);
and UO_309 (O_309,N_9973,N_9901);
nor UO_310 (O_310,N_9966,N_9931);
nand UO_311 (O_311,N_9982,N_9988);
or UO_312 (O_312,N_9962,N_9965);
nor UO_313 (O_313,N_9958,N_9930);
nand UO_314 (O_314,N_9923,N_9930);
xnor UO_315 (O_315,N_9913,N_9941);
nand UO_316 (O_316,N_9900,N_9991);
or UO_317 (O_317,N_9959,N_9946);
nand UO_318 (O_318,N_9956,N_9924);
nor UO_319 (O_319,N_9923,N_9996);
or UO_320 (O_320,N_9962,N_9993);
xor UO_321 (O_321,N_9985,N_9942);
nor UO_322 (O_322,N_9999,N_9988);
or UO_323 (O_323,N_9930,N_9917);
or UO_324 (O_324,N_9965,N_9929);
nand UO_325 (O_325,N_9915,N_9997);
and UO_326 (O_326,N_9900,N_9914);
or UO_327 (O_327,N_9956,N_9977);
nand UO_328 (O_328,N_9942,N_9973);
and UO_329 (O_329,N_9998,N_9971);
nor UO_330 (O_330,N_9939,N_9953);
or UO_331 (O_331,N_9933,N_9904);
or UO_332 (O_332,N_9965,N_9975);
and UO_333 (O_333,N_9976,N_9996);
and UO_334 (O_334,N_9912,N_9948);
nand UO_335 (O_335,N_9938,N_9925);
nor UO_336 (O_336,N_9908,N_9946);
nand UO_337 (O_337,N_9963,N_9961);
and UO_338 (O_338,N_9986,N_9908);
nand UO_339 (O_339,N_9906,N_9956);
nand UO_340 (O_340,N_9960,N_9928);
nand UO_341 (O_341,N_9909,N_9960);
nor UO_342 (O_342,N_9976,N_9928);
and UO_343 (O_343,N_9999,N_9979);
nor UO_344 (O_344,N_9993,N_9958);
and UO_345 (O_345,N_9961,N_9904);
or UO_346 (O_346,N_9946,N_9931);
or UO_347 (O_347,N_9906,N_9963);
xnor UO_348 (O_348,N_9974,N_9991);
and UO_349 (O_349,N_9958,N_9999);
or UO_350 (O_350,N_9929,N_9921);
nand UO_351 (O_351,N_9984,N_9991);
and UO_352 (O_352,N_9951,N_9917);
nor UO_353 (O_353,N_9977,N_9959);
nand UO_354 (O_354,N_9973,N_9923);
and UO_355 (O_355,N_9990,N_9986);
and UO_356 (O_356,N_9900,N_9980);
nor UO_357 (O_357,N_9936,N_9972);
nand UO_358 (O_358,N_9982,N_9945);
and UO_359 (O_359,N_9968,N_9949);
or UO_360 (O_360,N_9988,N_9966);
or UO_361 (O_361,N_9956,N_9938);
or UO_362 (O_362,N_9913,N_9990);
and UO_363 (O_363,N_9935,N_9913);
xor UO_364 (O_364,N_9983,N_9986);
nor UO_365 (O_365,N_9920,N_9971);
or UO_366 (O_366,N_9953,N_9912);
or UO_367 (O_367,N_9949,N_9964);
nand UO_368 (O_368,N_9911,N_9913);
and UO_369 (O_369,N_9953,N_9921);
nand UO_370 (O_370,N_9968,N_9943);
nand UO_371 (O_371,N_9919,N_9981);
nand UO_372 (O_372,N_9992,N_9932);
nor UO_373 (O_373,N_9969,N_9915);
nor UO_374 (O_374,N_9970,N_9909);
and UO_375 (O_375,N_9916,N_9943);
or UO_376 (O_376,N_9957,N_9989);
nor UO_377 (O_377,N_9964,N_9917);
nand UO_378 (O_378,N_9962,N_9980);
nand UO_379 (O_379,N_9993,N_9916);
xnor UO_380 (O_380,N_9940,N_9927);
and UO_381 (O_381,N_9907,N_9929);
nor UO_382 (O_382,N_9903,N_9987);
and UO_383 (O_383,N_9960,N_9992);
and UO_384 (O_384,N_9923,N_9967);
and UO_385 (O_385,N_9968,N_9954);
nor UO_386 (O_386,N_9993,N_9976);
or UO_387 (O_387,N_9991,N_9997);
and UO_388 (O_388,N_9964,N_9906);
or UO_389 (O_389,N_9968,N_9948);
or UO_390 (O_390,N_9931,N_9963);
nor UO_391 (O_391,N_9988,N_9987);
or UO_392 (O_392,N_9944,N_9924);
or UO_393 (O_393,N_9957,N_9920);
or UO_394 (O_394,N_9911,N_9920);
nand UO_395 (O_395,N_9952,N_9943);
or UO_396 (O_396,N_9970,N_9957);
nor UO_397 (O_397,N_9924,N_9906);
and UO_398 (O_398,N_9946,N_9990);
and UO_399 (O_399,N_9958,N_9965);
nor UO_400 (O_400,N_9930,N_9918);
or UO_401 (O_401,N_9965,N_9967);
or UO_402 (O_402,N_9981,N_9913);
and UO_403 (O_403,N_9929,N_9993);
nor UO_404 (O_404,N_9965,N_9957);
and UO_405 (O_405,N_9969,N_9979);
and UO_406 (O_406,N_9998,N_9972);
and UO_407 (O_407,N_9935,N_9992);
nand UO_408 (O_408,N_9999,N_9977);
or UO_409 (O_409,N_9942,N_9927);
or UO_410 (O_410,N_9918,N_9963);
or UO_411 (O_411,N_9975,N_9914);
and UO_412 (O_412,N_9985,N_9979);
and UO_413 (O_413,N_9946,N_9920);
and UO_414 (O_414,N_9950,N_9947);
and UO_415 (O_415,N_9996,N_9964);
or UO_416 (O_416,N_9947,N_9906);
or UO_417 (O_417,N_9990,N_9929);
or UO_418 (O_418,N_9916,N_9973);
nand UO_419 (O_419,N_9960,N_9923);
nor UO_420 (O_420,N_9922,N_9928);
nand UO_421 (O_421,N_9928,N_9989);
or UO_422 (O_422,N_9988,N_9917);
and UO_423 (O_423,N_9917,N_9981);
nand UO_424 (O_424,N_9973,N_9932);
or UO_425 (O_425,N_9942,N_9943);
nor UO_426 (O_426,N_9902,N_9940);
nand UO_427 (O_427,N_9903,N_9934);
nor UO_428 (O_428,N_9990,N_9977);
nand UO_429 (O_429,N_9944,N_9966);
and UO_430 (O_430,N_9975,N_9905);
nand UO_431 (O_431,N_9921,N_9901);
and UO_432 (O_432,N_9903,N_9935);
or UO_433 (O_433,N_9927,N_9978);
and UO_434 (O_434,N_9919,N_9910);
and UO_435 (O_435,N_9920,N_9961);
and UO_436 (O_436,N_9933,N_9930);
nand UO_437 (O_437,N_9935,N_9936);
nand UO_438 (O_438,N_9930,N_9978);
nor UO_439 (O_439,N_9964,N_9972);
nor UO_440 (O_440,N_9976,N_9989);
and UO_441 (O_441,N_9924,N_9908);
and UO_442 (O_442,N_9922,N_9949);
nand UO_443 (O_443,N_9924,N_9922);
and UO_444 (O_444,N_9937,N_9955);
or UO_445 (O_445,N_9924,N_9936);
and UO_446 (O_446,N_9941,N_9945);
and UO_447 (O_447,N_9965,N_9973);
xnor UO_448 (O_448,N_9901,N_9909);
or UO_449 (O_449,N_9977,N_9927);
or UO_450 (O_450,N_9984,N_9931);
and UO_451 (O_451,N_9971,N_9912);
xor UO_452 (O_452,N_9955,N_9992);
and UO_453 (O_453,N_9907,N_9930);
nor UO_454 (O_454,N_9950,N_9918);
nand UO_455 (O_455,N_9950,N_9925);
and UO_456 (O_456,N_9987,N_9916);
nor UO_457 (O_457,N_9963,N_9998);
nand UO_458 (O_458,N_9975,N_9976);
nor UO_459 (O_459,N_9902,N_9931);
nor UO_460 (O_460,N_9961,N_9935);
and UO_461 (O_461,N_9955,N_9995);
and UO_462 (O_462,N_9927,N_9957);
nand UO_463 (O_463,N_9981,N_9997);
and UO_464 (O_464,N_9910,N_9952);
xor UO_465 (O_465,N_9975,N_9996);
or UO_466 (O_466,N_9960,N_9990);
nand UO_467 (O_467,N_9974,N_9922);
nand UO_468 (O_468,N_9985,N_9983);
nor UO_469 (O_469,N_9943,N_9939);
nor UO_470 (O_470,N_9917,N_9971);
and UO_471 (O_471,N_9946,N_9981);
xor UO_472 (O_472,N_9913,N_9923);
or UO_473 (O_473,N_9955,N_9926);
nand UO_474 (O_474,N_9981,N_9962);
nand UO_475 (O_475,N_9974,N_9947);
nor UO_476 (O_476,N_9922,N_9935);
nand UO_477 (O_477,N_9968,N_9956);
and UO_478 (O_478,N_9968,N_9911);
nor UO_479 (O_479,N_9975,N_9915);
nor UO_480 (O_480,N_9935,N_9946);
nand UO_481 (O_481,N_9997,N_9944);
and UO_482 (O_482,N_9906,N_9985);
or UO_483 (O_483,N_9904,N_9964);
and UO_484 (O_484,N_9978,N_9904);
xor UO_485 (O_485,N_9935,N_9970);
nand UO_486 (O_486,N_9914,N_9989);
nor UO_487 (O_487,N_9963,N_9934);
nor UO_488 (O_488,N_9938,N_9902);
nand UO_489 (O_489,N_9986,N_9911);
nor UO_490 (O_490,N_9989,N_9961);
nand UO_491 (O_491,N_9941,N_9948);
or UO_492 (O_492,N_9907,N_9993);
nand UO_493 (O_493,N_9930,N_9911);
xor UO_494 (O_494,N_9937,N_9905);
nand UO_495 (O_495,N_9926,N_9909);
or UO_496 (O_496,N_9985,N_9960);
and UO_497 (O_497,N_9942,N_9958);
nor UO_498 (O_498,N_9958,N_9995);
and UO_499 (O_499,N_9985,N_9991);
nand UO_500 (O_500,N_9950,N_9984);
or UO_501 (O_501,N_9961,N_9982);
nand UO_502 (O_502,N_9929,N_9959);
nor UO_503 (O_503,N_9904,N_9965);
or UO_504 (O_504,N_9984,N_9930);
nor UO_505 (O_505,N_9991,N_9921);
and UO_506 (O_506,N_9911,N_9948);
and UO_507 (O_507,N_9942,N_9993);
nand UO_508 (O_508,N_9962,N_9907);
or UO_509 (O_509,N_9947,N_9988);
nor UO_510 (O_510,N_9920,N_9968);
and UO_511 (O_511,N_9973,N_9983);
or UO_512 (O_512,N_9946,N_9912);
nand UO_513 (O_513,N_9904,N_9928);
and UO_514 (O_514,N_9959,N_9906);
nand UO_515 (O_515,N_9992,N_9929);
nor UO_516 (O_516,N_9927,N_9968);
xor UO_517 (O_517,N_9942,N_9957);
nor UO_518 (O_518,N_9936,N_9948);
and UO_519 (O_519,N_9948,N_9955);
nand UO_520 (O_520,N_9961,N_9986);
or UO_521 (O_521,N_9970,N_9925);
nor UO_522 (O_522,N_9921,N_9968);
or UO_523 (O_523,N_9905,N_9966);
or UO_524 (O_524,N_9957,N_9933);
or UO_525 (O_525,N_9924,N_9905);
nor UO_526 (O_526,N_9938,N_9924);
nor UO_527 (O_527,N_9951,N_9908);
nor UO_528 (O_528,N_9901,N_9922);
nand UO_529 (O_529,N_9988,N_9952);
nor UO_530 (O_530,N_9910,N_9958);
nand UO_531 (O_531,N_9993,N_9989);
or UO_532 (O_532,N_9951,N_9925);
or UO_533 (O_533,N_9982,N_9929);
nand UO_534 (O_534,N_9954,N_9950);
nor UO_535 (O_535,N_9901,N_9944);
or UO_536 (O_536,N_9967,N_9982);
or UO_537 (O_537,N_9965,N_9964);
nor UO_538 (O_538,N_9920,N_9958);
nor UO_539 (O_539,N_9942,N_9974);
or UO_540 (O_540,N_9988,N_9912);
or UO_541 (O_541,N_9917,N_9944);
nor UO_542 (O_542,N_9999,N_9937);
nor UO_543 (O_543,N_9910,N_9926);
nand UO_544 (O_544,N_9950,N_9934);
or UO_545 (O_545,N_9980,N_9958);
and UO_546 (O_546,N_9918,N_9985);
nand UO_547 (O_547,N_9966,N_9922);
and UO_548 (O_548,N_9952,N_9958);
nand UO_549 (O_549,N_9910,N_9967);
and UO_550 (O_550,N_9906,N_9926);
and UO_551 (O_551,N_9926,N_9920);
or UO_552 (O_552,N_9952,N_9990);
nor UO_553 (O_553,N_9909,N_9936);
xnor UO_554 (O_554,N_9935,N_9950);
nand UO_555 (O_555,N_9901,N_9967);
or UO_556 (O_556,N_9903,N_9910);
nand UO_557 (O_557,N_9981,N_9938);
and UO_558 (O_558,N_9967,N_9913);
nor UO_559 (O_559,N_9910,N_9906);
nand UO_560 (O_560,N_9948,N_9927);
nand UO_561 (O_561,N_9911,N_9914);
nor UO_562 (O_562,N_9900,N_9938);
or UO_563 (O_563,N_9959,N_9968);
nor UO_564 (O_564,N_9924,N_9969);
nand UO_565 (O_565,N_9946,N_9915);
or UO_566 (O_566,N_9974,N_9906);
or UO_567 (O_567,N_9962,N_9908);
and UO_568 (O_568,N_9906,N_9960);
and UO_569 (O_569,N_9987,N_9948);
nor UO_570 (O_570,N_9945,N_9959);
nand UO_571 (O_571,N_9919,N_9987);
and UO_572 (O_572,N_9977,N_9963);
nor UO_573 (O_573,N_9978,N_9925);
nand UO_574 (O_574,N_9931,N_9900);
nor UO_575 (O_575,N_9974,N_9910);
nand UO_576 (O_576,N_9943,N_9980);
nand UO_577 (O_577,N_9923,N_9945);
nor UO_578 (O_578,N_9944,N_9970);
or UO_579 (O_579,N_9981,N_9995);
nor UO_580 (O_580,N_9944,N_9999);
or UO_581 (O_581,N_9949,N_9990);
or UO_582 (O_582,N_9911,N_9977);
nand UO_583 (O_583,N_9974,N_9953);
nor UO_584 (O_584,N_9934,N_9952);
nand UO_585 (O_585,N_9960,N_9980);
nor UO_586 (O_586,N_9935,N_9981);
nor UO_587 (O_587,N_9958,N_9901);
nor UO_588 (O_588,N_9980,N_9984);
and UO_589 (O_589,N_9967,N_9992);
and UO_590 (O_590,N_9991,N_9973);
and UO_591 (O_591,N_9960,N_9943);
nand UO_592 (O_592,N_9940,N_9933);
or UO_593 (O_593,N_9977,N_9973);
and UO_594 (O_594,N_9955,N_9969);
nor UO_595 (O_595,N_9901,N_9976);
nor UO_596 (O_596,N_9917,N_9985);
or UO_597 (O_597,N_9922,N_9946);
nor UO_598 (O_598,N_9975,N_9921);
or UO_599 (O_599,N_9978,N_9973);
and UO_600 (O_600,N_9914,N_9995);
nor UO_601 (O_601,N_9983,N_9902);
or UO_602 (O_602,N_9975,N_9985);
nor UO_603 (O_603,N_9927,N_9947);
and UO_604 (O_604,N_9938,N_9958);
or UO_605 (O_605,N_9994,N_9938);
and UO_606 (O_606,N_9915,N_9927);
or UO_607 (O_607,N_9936,N_9979);
xnor UO_608 (O_608,N_9997,N_9959);
and UO_609 (O_609,N_9992,N_9983);
or UO_610 (O_610,N_9997,N_9939);
or UO_611 (O_611,N_9930,N_9941);
nor UO_612 (O_612,N_9901,N_9940);
nand UO_613 (O_613,N_9940,N_9947);
or UO_614 (O_614,N_9943,N_9918);
nor UO_615 (O_615,N_9913,N_9956);
or UO_616 (O_616,N_9949,N_9941);
nor UO_617 (O_617,N_9986,N_9985);
nand UO_618 (O_618,N_9916,N_9982);
nor UO_619 (O_619,N_9958,N_9905);
nand UO_620 (O_620,N_9982,N_9941);
nor UO_621 (O_621,N_9961,N_9962);
and UO_622 (O_622,N_9988,N_9967);
and UO_623 (O_623,N_9939,N_9974);
or UO_624 (O_624,N_9944,N_9938);
and UO_625 (O_625,N_9983,N_9922);
nand UO_626 (O_626,N_9938,N_9951);
and UO_627 (O_627,N_9971,N_9906);
nand UO_628 (O_628,N_9918,N_9970);
and UO_629 (O_629,N_9996,N_9921);
and UO_630 (O_630,N_9990,N_9903);
nor UO_631 (O_631,N_9922,N_9951);
nand UO_632 (O_632,N_9933,N_9944);
or UO_633 (O_633,N_9906,N_9945);
or UO_634 (O_634,N_9959,N_9983);
nand UO_635 (O_635,N_9908,N_9964);
or UO_636 (O_636,N_9918,N_9988);
nor UO_637 (O_637,N_9946,N_9960);
and UO_638 (O_638,N_9948,N_9946);
and UO_639 (O_639,N_9983,N_9900);
and UO_640 (O_640,N_9919,N_9901);
nand UO_641 (O_641,N_9990,N_9998);
and UO_642 (O_642,N_9971,N_9968);
or UO_643 (O_643,N_9950,N_9915);
and UO_644 (O_644,N_9923,N_9949);
nand UO_645 (O_645,N_9962,N_9982);
nor UO_646 (O_646,N_9922,N_9925);
or UO_647 (O_647,N_9935,N_9949);
or UO_648 (O_648,N_9981,N_9989);
and UO_649 (O_649,N_9908,N_9911);
nand UO_650 (O_650,N_9931,N_9986);
and UO_651 (O_651,N_9966,N_9967);
or UO_652 (O_652,N_9970,N_9946);
or UO_653 (O_653,N_9991,N_9908);
nand UO_654 (O_654,N_9935,N_9940);
and UO_655 (O_655,N_9990,N_9901);
and UO_656 (O_656,N_9984,N_9974);
nor UO_657 (O_657,N_9981,N_9963);
or UO_658 (O_658,N_9930,N_9931);
and UO_659 (O_659,N_9929,N_9957);
or UO_660 (O_660,N_9910,N_9992);
or UO_661 (O_661,N_9935,N_9904);
nand UO_662 (O_662,N_9960,N_9904);
xnor UO_663 (O_663,N_9982,N_9923);
or UO_664 (O_664,N_9930,N_9989);
nand UO_665 (O_665,N_9924,N_9966);
nor UO_666 (O_666,N_9907,N_9945);
nand UO_667 (O_667,N_9922,N_9937);
nor UO_668 (O_668,N_9938,N_9922);
or UO_669 (O_669,N_9987,N_9917);
and UO_670 (O_670,N_9920,N_9973);
nand UO_671 (O_671,N_9984,N_9953);
nand UO_672 (O_672,N_9907,N_9938);
nand UO_673 (O_673,N_9929,N_9925);
and UO_674 (O_674,N_9908,N_9989);
nand UO_675 (O_675,N_9997,N_9928);
nand UO_676 (O_676,N_9987,N_9971);
nand UO_677 (O_677,N_9963,N_9914);
nor UO_678 (O_678,N_9970,N_9902);
nand UO_679 (O_679,N_9968,N_9992);
and UO_680 (O_680,N_9962,N_9928);
nand UO_681 (O_681,N_9981,N_9931);
nand UO_682 (O_682,N_9949,N_9930);
nor UO_683 (O_683,N_9998,N_9918);
nand UO_684 (O_684,N_9920,N_9943);
and UO_685 (O_685,N_9900,N_9976);
or UO_686 (O_686,N_9970,N_9923);
or UO_687 (O_687,N_9915,N_9985);
or UO_688 (O_688,N_9905,N_9989);
and UO_689 (O_689,N_9944,N_9959);
nor UO_690 (O_690,N_9971,N_9900);
nor UO_691 (O_691,N_9998,N_9939);
nand UO_692 (O_692,N_9984,N_9903);
and UO_693 (O_693,N_9901,N_9964);
and UO_694 (O_694,N_9919,N_9941);
and UO_695 (O_695,N_9989,N_9913);
nor UO_696 (O_696,N_9905,N_9981);
or UO_697 (O_697,N_9918,N_9942);
and UO_698 (O_698,N_9991,N_9968);
nand UO_699 (O_699,N_9911,N_9966);
nand UO_700 (O_700,N_9933,N_9996);
nand UO_701 (O_701,N_9953,N_9987);
and UO_702 (O_702,N_9931,N_9953);
or UO_703 (O_703,N_9914,N_9955);
nand UO_704 (O_704,N_9957,N_9906);
and UO_705 (O_705,N_9942,N_9903);
or UO_706 (O_706,N_9969,N_9985);
nand UO_707 (O_707,N_9930,N_9946);
or UO_708 (O_708,N_9941,N_9937);
and UO_709 (O_709,N_9962,N_9952);
and UO_710 (O_710,N_9935,N_9939);
and UO_711 (O_711,N_9994,N_9917);
nand UO_712 (O_712,N_9990,N_9982);
and UO_713 (O_713,N_9948,N_9944);
nor UO_714 (O_714,N_9925,N_9981);
or UO_715 (O_715,N_9935,N_9930);
nor UO_716 (O_716,N_9960,N_9999);
and UO_717 (O_717,N_9964,N_9947);
nand UO_718 (O_718,N_9949,N_9914);
nor UO_719 (O_719,N_9903,N_9944);
nor UO_720 (O_720,N_9990,N_9934);
and UO_721 (O_721,N_9927,N_9986);
and UO_722 (O_722,N_9957,N_9926);
and UO_723 (O_723,N_9954,N_9910);
xnor UO_724 (O_724,N_9987,N_9967);
nor UO_725 (O_725,N_9984,N_9952);
or UO_726 (O_726,N_9920,N_9959);
nor UO_727 (O_727,N_9918,N_9944);
nor UO_728 (O_728,N_9955,N_9978);
nand UO_729 (O_729,N_9955,N_9904);
xor UO_730 (O_730,N_9982,N_9905);
nand UO_731 (O_731,N_9914,N_9967);
nand UO_732 (O_732,N_9999,N_9938);
nor UO_733 (O_733,N_9992,N_9905);
and UO_734 (O_734,N_9953,N_9901);
nor UO_735 (O_735,N_9959,N_9907);
xnor UO_736 (O_736,N_9981,N_9973);
nand UO_737 (O_737,N_9976,N_9971);
and UO_738 (O_738,N_9975,N_9907);
nand UO_739 (O_739,N_9956,N_9918);
nor UO_740 (O_740,N_9929,N_9953);
nand UO_741 (O_741,N_9920,N_9915);
nor UO_742 (O_742,N_9925,N_9933);
nor UO_743 (O_743,N_9927,N_9988);
nor UO_744 (O_744,N_9939,N_9962);
or UO_745 (O_745,N_9956,N_9999);
or UO_746 (O_746,N_9995,N_9903);
nor UO_747 (O_747,N_9968,N_9947);
nand UO_748 (O_748,N_9917,N_9995);
nand UO_749 (O_749,N_9980,N_9991);
or UO_750 (O_750,N_9938,N_9903);
or UO_751 (O_751,N_9987,N_9940);
nand UO_752 (O_752,N_9921,N_9993);
nor UO_753 (O_753,N_9905,N_9908);
nor UO_754 (O_754,N_9903,N_9969);
and UO_755 (O_755,N_9991,N_9911);
or UO_756 (O_756,N_9942,N_9914);
nor UO_757 (O_757,N_9929,N_9967);
or UO_758 (O_758,N_9991,N_9955);
or UO_759 (O_759,N_9987,N_9915);
nor UO_760 (O_760,N_9975,N_9977);
and UO_761 (O_761,N_9942,N_9930);
nand UO_762 (O_762,N_9906,N_9992);
or UO_763 (O_763,N_9971,N_9980);
and UO_764 (O_764,N_9913,N_9982);
xnor UO_765 (O_765,N_9950,N_9909);
or UO_766 (O_766,N_9955,N_9919);
or UO_767 (O_767,N_9982,N_9930);
or UO_768 (O_768,N_9939,N_9917);
or UO_769 (O_769,N_9988,N_9997);
nor UO_770 (O_770,N_9972,N_9941);
nand UO_771 (O_771,N_9900,N_9992);
and UO_772 (O_772,N_9907,N_9946);
nor UO_773 (O_773,N_9948,N_9978);
and UO_774 (O_774,N_9976,N_9973);
and UO_775 (O_775,N_9998,N_9974);
nand UO_776 (O_776,N_9918,N_9929);
nor UO_777 (O_777,N_9950,N_9981);
nand UO_778 (O_778,N_9925,N_9963);
nor UO_779 (O_779,N_9930,N_9905);
nor UO_780 (O_780,N_9978,N_9938);
nand UO_781 (O_781,N_9956,N_9907);
nand UO_782 (O_782,N_9939,N_9975);
nor UO_783 (O_783,N_9935,N_9911);
nor UO_784 (O_784,N_9918,N_9975);
or UO_785 (O_785,N_9930,N_9950);
xnor UO_786 (O_786,N_9955,N_9917);
nand UO_787 (O_787,N_9903,N_9982);
nand UO_788 (O_788,N_9915,N_9966);
or UO_789 (O_789,N_9948,N_9967);
or UO_790 (O_790,N_9911,N_9970);
nand UO_791 (O_791,N_9912,N_9928);
nor UO_792 (O_792,N_9930,N_9985);
nand UO_793 (O_793,N_9972,N_9938);
xor UO_794 (O_794,N_9953,N_9913);
nor UO_795 (O_795,N_9970,N_9975);
and UO_796 (O_796,N_9977,N_9939);
nor UO_797 (O_797,N_9967,N_9928);
or UO_798 (O_798,N_9954,N_9928);
nor UO_799 (O_799,N_9930,N_9919);
and UO_800 (O_800,N_9964,N_9910);
nor UO_801 (O_801,N_9980,N_9927);
nor UO_802 (O_802,N_9994,N_9933);
or UO_803 (O_803,N_9986,N_9915);
nor UO_804 (O_804,N_9944,N_9996);
nor UO_805 (O_805,N_9923,N_9972);
and UO_806 (O_806,N_9911,N_9951);
and UO_807 (O_807,N_9986,N_9926);
nor UO_808 (O_808,N_9949,N_9966);
nand UO_809 (O_809,N_9983,N_9941);
nand UO_810 (O_810,N_9967,N_9934);
and UO_811 (O_811,N_9911,N_9958);
and UO_812 (O_812,N_9989,N_9942);
and UO_813 (O_813,N_9962,N_9978);
nand UO_814 (O_814,N_9939,N_9936);
and UO_815 (O_815,N_9914,N_9957);
nand UO_816 (O_816,N_9973,N_9913);
or UO_817 (O_817,N_9930,N_9953);
nand UO_818 (O_818,N_9948,N_9921);
nand UO_819 (O_819,N_9994,N_9929);
and UO_820 (O_820,N_9964,N_9971);
or UO_821 (O_821,N_9995,N_9905);
nor UO_822 (O_822,N_9960,N_9915);
nand UO_823 (O_823,N_9991,N_9993);
nor UO_824 (O_824,N_9972,N_9903);
nor UO_825 (O_825,N_9993,N_9982);
nand UO_826 (O_826,N_9907,N_9905);
nor UO_827 (O_827,N_9956,N_9915);
and UO_828 (O_828,N_9963,N_9968);
nor UO_829 (O_829,N_9960,N_9994);
and UO_830 (O_830,N_9904,N_9941);
nor UO_831 (O_831,N_9930,N_9910);
or UO_832 (O_832,N_9952,N_9904);
nand UO_833 (O_833,N_9917,N_9954);
nor UO_834 (O_834,N_9930,N_9999);
or UO_835 (O_835,N_9903,N_9922);
or UO_836 (O_836,N_9991,N_9946);
nor UO_837 (O_837,N_9950,N_9941);
nor UO_838 (O_838,N_9916,N_9939);
or UO_839 (O_839,N_9957,N_9960);
nor UO_840 (O_840,N_9978,N_9935);
or UO_841 (O_841,N_9900,N_9925);
nand UO_842 (O_842,N_9992,N_9947);
nand UO_843 (O_843,N_9973,N_9971);
nor UO_844 (O_844,N_9985,N_9901);
nor UO_845 (O_845,N_9932,N_9983);
nand UO_846 (O_846,N_9916,N_9932);
or UO_847 (O_847,N_9994,N_9916);
nand UO_848 (O_848,N_9909,N_9987);
nand UO_849 (O_849,N_9994,N_9992);
nor UO_850 (O_850,N_9961,N_9960);
nor UO_851 (O_851,N_9926,N_9939);
nand UO_852 (O_852,N_9929,N_9998);
or UO_853 (O_853,N_9959,N_9953);
nor UO_854 (O_854,N_9913,N_9934);
nor UO_855 (O_855,N_9964,N_9942);
and UO_856 (O_856,N_9905,N_9985);
and UO_857 (O_857,N_9933,N_9920);
nor UO_858 (O_858,N_9979,N_9954);
nand UO_859 (O_859,N_9993,N_9979);
nor UO_860 (O_860,N_9916,N_9927);
nand UO_861 (O_861,N_9949,N_9943);
nand UO_862 (O_862,N_9969,N_9939);
nor UO_863 (O_863,N_9942,N_9917);
or UO_864 (O_864,N_9972,N_9993);
and UO_865 (O_865,N_9965,N_9968);
nand UO_866 (O_866,N_9960,N_9984);
or UO_867 (O_867,N_9986,N_9957);
nor UO_868 (O_868,N_9965,N_9976);
nand UO_869 (O_869,N_9944,N_9998);
and UO_870 (O_870,N_9933,N_9900);
xnor UO_871 (O_871,N_9923,N_9943);
and UO_872 (O_872,N_9988,N_9913);
or UO_873 (O_873,N_9923,N_9989);
xor UO_874 (O_874,N_9937,N_9962);
xor UO_875 (O_875,N_9922,N_9967);
or UO_876 (O_876,N_9957,N_9909);
nand UO_877 (O_877,N_9924,N_9977);
and UO_878 (O_878,N_9943,N_9925);
nor UO_879 (O_879,N_9945,N_9976);
nand UO_880 (O_880,N_9967,N_9945);
xnor UO_881 (O_881,N_9945,N_9968);
and UO_882 (O_882,N_9941,N_9947);
xnor UO_883 (O_883,N_9927,N_9944);
or UO_884 (O_884,N_9993,N_9978);
xnor UO_885 (O_885,N_9953,N_9910);
nor UO_886 (O_886,N_9915,N_9983);
nor UO_887 (O_887,N_9943,N_9903);
and UO_888 (O_888,N_9959,N_9996);
nor UO_889 (O_889,N_9959,N_9909);
and UO_890 (O_890,N_9984,N_9978);
xnor UO_891 (O_891,N_9904,N_9900);
and UO_892 (O_892,N_9970,N_9922);
and UO_893 (O_893,N_9929,N_9987);
nand UO_894 (O_894,N_9926,N_9994);
nor UO_895 (O_895,N_9929,N_9986);
or UO_896 (O_896,N_9946,N_9951);
nor UO_897 (O_897,N_9955,N_9920);
nand UO_898 (O_898,N_9936,N_9908);
nor UO_899 (O_899,N_9913,N_9974);
nand UO_900 (O_900,N_9959,N_9910);
or UO_901 (O_901,N_9924,N_9988);
nor UO_902 (O_902,N_9901,N_9984);
or UO_903 (O_903,N_9980,N_9917);
nand UO_904 (O_904,N_9972,N_9953);
nor UO_905 (O_905,N_9966,N_9933);
nand UO_906 (O_906,N_9902,N_9908);
and UO_907 (O_907,N_9978,N_9944);
or UO_908 (O_908,N_9924,N_9996);
nand UO_909 (O_909,N_9969,N_9900);
or UO_910 (O_910,N_9903,N_9925);
nand UO_911 (O_911,N_9990,N_9993);
and UO_912 (O_912,N_9923,N_9944);
nor UO_913 (O_913,N_9918,N_9906);
nor UO_914 (O_914,N_9909,N_9994);
nand UO_915 (O_915,N_9933,N_9995);
nor UO_916 (O_916,N_9901,N_9926);
or UO_917 (O_917,N_9927,N_9933);
and UO_918 (O_918,N_9961,N_9987);
or UO_919 (O_919,N_9994,N_9959);
nand UO_920 (O_920,N_9925,N_9959);
and UO_921 (O_921,N_9917,N_9956);
or UO_922 (O_922,N_9914,N_9992);
or UO_923 (O_923,N_9919,N_9915);
nand UO_924 (O_924,N_9997,N_9938);
nand UO_925 (O_925,N_9934,N_9996);
xor UO_926 (O_926,N_9977,N_9932);
or UO_927 (O_927,N_9989,N_9971);
and UO_928 (O_928,N_9917,N_9983);
or UO_929 (O_929,N_9977,N_9997);
xor UO_930 (O_930,N_9933,N_9916);
xnor UO_931 (O_931,N_9992,N_9903);
nand UO_932 (O_932,N_9931,N_9956);
nand UO_933 (O_933,N_9930,N_9967);
nor UO_934 (O_934,N_9929,N_9964);
or UO_935 (O_935,N_9900,N_9986);
nor UO_936 (O_936,N_9928,N_9946);
nand UO_937 (O_937,N_9915,N_9961);
or UO_938 (O_938,N_9926,N_9922);
or UO_939 (O_939,N_9992,N_9918);
and UO_940 (O_940,N_9996,N_9947);
nor UO_941 (O_941,N_9914,N_9941);
nor UO_942 (O_942,N_9990,N_9967);
nor UO_943 (O_943,N_9959,N_9957);
nor UO_944 (O_944,N_9973,N_9924);
nand UO_945 (O_945,N_9989,N_9943);
nand UO_946 (O_946,N_9950,N_9993);
nand UO_947 (O_947,N_9960,N_9959);
nand UO_948 (O_948,N_9908,N_9906);
nor UO_949 (O_949,N_9914,N_9987);
nor UO_950 (O_950,N_9924,N_9954);
nand UO_951 (O_951,N_9948,N_9991);
nor UO_952 (O_952,N_9904,N_9976);
or UO_953 (O_953,N_9993,N_9945);
or UO_954 (O_954,N_9919,N_9907);
nand UO_955 (O_955,N_9977,N_9943);
or UO_956 (O_956,N_9965,N_9932);
or UO_957 (O_957,N_9996,N_9907);
and UO_958 (O_958,N_9912,N_9909);
nor UO_959 (O_959,N_9997,N_9924);
nand UO_960 (O_960,N_9931,N_9962);
and UO_961 (O_961,N_9965,N_9988);
nor UO_962 (O_962,N_9912,N_9991);
and UO_963 (O_963,N_9920,N_9969);
or UO_964 (O_964,N_9990,N_9973);
nand UO_965 (O_965,N_9983,N_9947);
or UO_966 (O_966,N_9942,N_9936);
nand UO_967 (O_967,N_9954,N_9948);
or UO_968 (O_968,N_9967,N_9964);
and UO_969 (O_969,N_9998,N_9931);
nand UO_970 (O_970,N_9966,N_9904);
and UO_971 (O_971,N_9923,N_9927);
nand UO_972 (O_972,N_9916,N_9948);
and UO_973 (O_973,N_9972,N_9910);
and UO_974 (O_974,N_9963,N_9983);
and UO_975 (O_975,N_9936,N_9912);
or UO_976 (O_976,N_9962,N_9945);
and UO_977 (O_977,N_9931,N_9967);
and UO_978 (O_978,N_9907,N_9947);
or UO_979 (O_979,N_9947,N_9917);
xnor UO_980 (O_980,N_9962,N_9951);
or UO_981 (O_981,N_9941,N_9980);
nor UO_982 (O_982,N_9972,N_9949);
nand UO_983 (O_983,N_9909,N_9921);
or UO_984 (O_984,N_9929,N_9961);
nand UO_985 (O_985,N_9982,N_9971);
nand UO_986 (O_986,N_9976,N_9990);
and UO_987 (O_987,N_9999,N_9964);
nor UO_988 (O_988,N_9918,N_9912);
and UO_989 (O_989,N_9996,N_9950);
nand UO_990 (O_990,N_9939,N_9966);
and UO_991 (O_991,N_9995,N_9920);
nand UO_992 (O_992,N_9933,N_9991);
nand UO_993 (O_993,N_9939,N_9938);
nor UO_994 (O_994,N_9927,N_9941);
or UO_995 (O_995,N_9928,N_9941);
and UO_996 (O_996,N_9944,N_9920);
and UO_997 (O_997,N_9934,N_9954);
and UO_998 (O_998,N_9935,N_9910);
and UO_999 (O_999,N_9957,N_9937);
or UO_1000 (O_1000,N_9927,N_9981);
and UO_1001 (O_1001,N_9970,N_9948);
and UO_1002 (O_1002,N_9986,N_9966);
or UO_1003 (O_1003,N_9908,N_9942);
nor UO_1004 (O_1004,N_9921,N_9976);
nand UO_1005 (O_1005,N_9945,N_9913);
or UO_1006 (O_1006,N_9924,N_9940);
or UO_1007 (O_1007,N_9988,N_9963);
nand UO_1008 (O_1008,N_9972,N_9901);
nand UO_1009 (O_1009,N_9963,N_9982);
nand UO_1010 (O_1010,N_9941,N_9996);
nor UO_1011 (O_1011,N_9909,N_9974);
nor UO_1012 (O_1012,N_9945,N_9944);
xor UO_1013 (O_1013,N_9974,N_9965);
or UO_1014 (O_1014,N_9909,N_9958);
and UO_1015 (O_1015,N_9916,N_9952);
or UO_1016 (O_1016,N_9938,N_9980);
and UO_1017 (O_1017,N_9968,N_9942);
nand UO_1018 (O_1018,N_9924,N_9976);
xnor UO_1019 (O_1019,N_9949,N_9938);
nor UO_1020 (O_1020,N_9948,N_9996);
and UO_1021 (O_1021,N_9975,N_9909);
or UO_1022 (O_1022,N_9915,N_9999);
nor UO_1023 (O_1023,N_9979,N_9942);
and UO_1024 (O_1024,N_9991,N_9944);
or UO_1025 (O_1025,N_9937,N_9926);
or UO_1026 (O_1026,N_9983,N_9974);
nand UO_1027 (O_1027,N_9912,N_9973);
nand UO_1028 (O_1028,N_9965,N_9984);
and UO_1029 (O_1029,N_9937,N_9978);
nor UO_1030 (O_1030,N_9904,N_9944);
or UO_1031 (O_1031,N_9907,N_9982);
and UO_1032 (O_1032,N_9956,N_9942);
nor UO_1033 (O_1033,N_9977,N_9978);
nand UO_1034 (O_1034,N_9905,N_9912);
or UO_1035 (O_1035,N_9934,N_9965);
nand UO_1036 (O_1036,N_9953,N_9935);
and UO_1037 (O_1037,N_9993,N_9910);
nand UO_1038 (O_1038,N_9922,N_9980);
nand UO_1039 (O_1039,N_9944,N_9914);
nand UO_1040 (O_1040,N_9973,N_9922);
nor UO_1041 (O_1041,N_9958,N_9921);
and UO_1042 (O_1042,N_9900,N_9901);
or UO_1043 (O_1043,N_9978,N_9981);
xor UO_1044 (O_1044,N_9982,N_9943);
and UO_1045 (O_1045,N_9972,N_9971);
or UO_1046 (O_1046,N_9937,N_9909);
and UO_1047 (O_1047,N_9966,N_9955);
and UO_1048 (O_1048,N_9921,N_9955);
or UO_1049 (O_1049,N_9926,N_9943);
or UO_1050 (O_1050,N_9908,N_9961);
or UO_1051 (O_1051,N_9969,N_9921);
nor UO_1052 (O_1052,N_9990,N_9910);
and UO_1053 (O_1053,N_9913,N_9907);
nor UO_1054 (O_1054,N_9959,N_9981);
or UO_1055 (O_1055,N_9975,N_9986);
nand UO_1056 (O_1056,N_9986,N_9951);
nand UO_1057 (O_1057,N_9925,N_9948);
or UO_1058 (O_1058,N_9913,N_9902);
nand UO_1059 (O_1059,N_9964,N_9905);
nand UO_1060 (O_1060,N_9980,N_9959);
nor UO_1061 (O_1061,N_9940,N_9943);
and UO_1062 (O_1062,N_9928,N_9917);
or UO_1063 (O_1063,N_9970,N_9956);
nor UO_1064 (O_1064,N_9940,N_9907);
or UO_1065 (O_1065,N_9922,N_9921);
or UO_1066 (O_1066,N_9972,N_9934);
and UO_1067 (O_1067,N_9983,N_9994);
nor UO_1068 (O_1068,N_9945,N_9957);
nor UO_1069 (O_1069,N_9959,N_9982);
nand UO_1070 (O_1070,N_9911,N_9955);
and UO_1071 (O_1071,N_9953,N_9936);
or UO_1072 (O_1072,N_9998,N_9979);
nor UO_1073 (O_1073,N_9993,N_9961);
nor UO_1074 (O_1074,N_9941,N_9967);
nor UO_1075 (O_1075,N_9970,N_9907);
or UO_1076 (O_1076,N_9958,N_9947);
nand UO_1077 (O_1077,N_9948,N_9922);
nor UO_1078 (O_1078,N_9929,N_9976);
nor UO_1079 (O_1079,N_9949,N_9985);
nor UO_1080 (O_1080,N_9920,N_9924);
nand UO_1081 (O_1081,N_9960,N_9926);
and UO_1082 (O_1082,N_9992,N_9957);
nor UO_1083 (O_1083,N_9989,N_9918);
nand UO_1084 (O_1084,N_9917,N_9925);
nor UO_1085 (O_1085,N_9929,N_9913);
xnor UO_1086 (O_1086,N_9936,N_9973);
xor UO_1087 (O_1087,N_9942,N_9904);
nor UO_1088 (O_1088,N_9979,N_9981);
or UO_1089 (O_1089,N_9917,N_9918);
and UO_1090 (O_1090,N_9975,N_9908);
nor UO_1091 (O_1091,N_9965,N_9942);
nand UO_1092 (O_1092,N_9929,N_9916);
nor UO_1093 (O_1093,N_9931,N_9906);
or UO_1094 (O_1094,N_9959,N_9974);
and UO_1095 (O_1095,N_9974,N_9945);
nor UO_1096 (O_1096,N_9922,N_9923);
and UO_1097 (O_1097,N_9958,N_9913);
nand UO_1098 (O_1098,N_9988,N_9991);
and UO_1099 (O_1099,N_9947,N_9931);
nand UO_1100 (O_1100,N_9942,N_9986);
or UO_1101 (O_1101,N_9974,N_9995);
nand UO_1102 (O_1102,N_9968,N_9918);
nand UO_1103 (O_1103,N_9976,N_9994);
or UO_1104 (O_1104,N_9948,N_9965);
nand UO_1105 (O_1105,N_9952,N_9901);
or UO_1106 (O_1106,N_9970,N_9958);
or UO_1107 (O_1107,N_9929,N_9927);
or UO_1108 (O_1108,N_9992,N_9934);
nand UO_1109 (O_1109,N_9963,N_9948);
nor UO_1110 (O_1110,N_9976,N_9986);
nor UO_1111 (O_1111,N_9943,N_9919);
xor UO_1112 (O_1112,N_9970,N_9926);
nand UO_1113 (O_1113,N_9975,N_9946);
and UO_1114 (O_1114,N_9925,N_9958);
nand UO_1115 (O_1115,N_9966,N_9913);
xnor UO_1116 (O_1116,N_9900,N_9997);
nand UO_1117 (O_1117,N_9989,N_9924);
nor UO_1118 (O_1118,N_9926,N_9972);
and UO_1119 (O_1119,N_9983,N_9958);
nand UO_1120 (O_1120,N_9934,N_9953);
and UO_1121 (O_1121,N_9965,N_9902);
nor UO_1122 (O_1122,N_9963,N_9917);
and UO_1123 (O_1123,N_9932,N_9905);
or UO_1124 (O_1124,N_9968,N_9905);
nand UO_1125 (O_1125,N_9976,N_9915);
and UO_1126 (O_1126,N_9996,N_9970);
or UO_1127 (O_1127,N_9901,N_9933);
or UO_1128 (O_1128,N_9967,N_9977);
nand UO_1129 (O_1129,N_9915,N_9907);
or UO_1130 (O_1130,N_9909,N_9992);
nor UO_1131 (O_1131,N_9990,N_9974);
or UO_1132 (O_1132,N_9971,N_9903);
xor UO_1133 (O_1133,N_9975,N_9925);
nor UO_1134 (O_1134,N_9966,N_9973);
or UO_1135 (O_1135,N_9989,N_9935);
nand UO_1136 (O_1136,N_9968,N_9912);
nor UO_1137 (O_1137,N_9952,N_9918);
or UO_1138 (O_1138,N_9933,N_9902);
and UO_1139 (O_1139,N_9966,N_9925);
nor UO_1140 (O_1140,N_9940,N_9959);
nor UO_1141 (O_1141,N_9921,N_9944);
nand UO_1142 (O_1142,N_9954,N_9935);
or UO_1143 (O_1143,N_9999,N_9989);
nor UO_1144 (O_1144,N_9909,N_9953);
xnor UO_1145 (O_1145,N_9985,N_9973);
nor UO_1146 (O_1146,N_9922,N_9982);
nor UO_1147 (O_1147,N_9971,N_9938);
nand UO_1148 (O_1148,N_9959,N_9922);
nor UO_1149 (O_1149,N_9991,N_9918);
nand UO_1150 (O_1150,N_9980,N_9955);
or UO_1151 (O_1151,N_9931,N_9928);
nor UO_1152 (O_1152,N_9961,N_9947);
nand UO_1153 (O_1153,N_9928,N_9935);
nor UO_1154 (O_1154,N_9997,N_9986);
and UO_1155 (O_1155,N_9905,N_9998);
and UO_1156 (O_1156,N_9968,N_9982);
nand UO_1157 (O_1157,N_9909,N_9952);
nor UO_1158 (O_1158,N_9977,N_9972);
nand UO_1159 (O_1159,N_9945,N_9988);
nand UO_1160 (O_1160,N_9977,N_9953);
or UO_1161 (O_1161,N_9909,N_9982);
nand UO_1162 (O_1162,N_9929,N_9904);
nor UO_1163 (O_1163,N_9964,N_9940);
nand UO_1164 (O_1164,N_9979,N_9949);
nand UO_1165 (O_1165,N_9998,N_9921);
or UO_1166 (O_1166,N_9938,N_9917);
or UO_1167 (O_1167,N_9941,N_9973);
nor UO_1168 (O_1168,N_9914,N_9982);
nor UO_1169 (O_1169,N_9980,N_9932);
or UO_1170 (O_1170,N_9943,N_9963);
or UO_1171 (O_1171,N_9966,N_9923);
and UO_1172 (O_1172,N_9947,N_9994);
nor UO_1173 (O_1173,N_9935,N_9979);
nor UO_1174 (O_1174,N_9911,N_9905);
or UO_1175 (O_1175,N_9995,N_9921);
and UO_1176 (O_1176,N_9970,N_9940);
or UO_1177 (O_1177,N_9915,N_9934);
nand UO_1178 (O_1178,N_9999,N_9994);
and UO_1179 (O_1179,N_9985,N_9978);
nor UO_1180 (O_1180,N_9942,N_9924);
nor UO_1181 (O_1181,N_9986,N_9996);
nor UO_1182 (O_1182,N_9995,N_9928);
or UO_1183 (O_1183,N_9932,N_9939);
nor UO_1184 (O_1184,N_9901,N_9969);
nand UO_1185 (O_1185,N_9944,N_9900);
nand UO_1186 (O_1186,N_9933,N_9976);
nand UO_1187 (O_1187,N_9975,N_9902);
or UO_1188 (O_1188,N_9949,N_9950);
nand UO_1189 (O_1189,N_9945,N_9910);
nand UO_1190 (O_1190,N_9928,N_9993);
nor UO_1191 (O_1191,N_9916,N_9974);
nand UO_1192 (O_1192,N_9938,N_9930);
and UO_1193 (O_1193,N_9988,N_9911);
and UO_1194 (O_1194,N_9952,N_9912);
nand UO_1195 (O_1195,N_9937,N_9946);
nor UO_1196 (O_1196,N_9932,N_9959);
nor UO_1197 (O_1197,N_9962,N_9948);
and UO_1198 (O_1198,N_9953,N_9949);
or UO_1199 (O_1199,N_9948,N_9976);
or UO_1200 (O_1200,N_9922,N_9913);
nand UO_1201 (O_1201,N_9960,N_9934);
and UO_1202 (O_1202,N_9928,N_9909);
and UO_1203 (O_1203,N_9910,N_9968);
or UO_1204 (O_1204,N_9909,N_9935);
or UO_1205 (O_1205,N_9994,N_9972);
and UO_1206 (O_1206,N_9956,N_9905);
xnor UO_1207 (O_1207,N_9971,N_9921);
nor UO_1208 (O_1208,N_9925,N_9928);
and UO_1209 (O_1209,N_9919,N_9973);
nand UO_1210 (O_1210,N_9954,N_9906);
or UO_1211 (O_1211,N_9939,N_9903);
and UO_1212 (O_1212,N_9911,N_9921);
nand UO_1213 (O_1213,N_9985,N_9945);
or UO_1214 (O_1214,N_9998,N_9941);
nand UO_1215 (O_1215,N_9974,N_9920);
and UO_1216 (O_1216,N_9968,N_9946);
or UO_1217 (O_1217,N_9909,N_9944);
or UO_1218 (O_1218,N_9923,N_9916);
nand UO_1219 (O_1219,N_9973,N_9918);
and UO_1220 (O_1220,N_9906,N_9977);
nand UO_1221 (O_1221,N_9944,N_9992);
nor UO_1222 (O_1222,N_9985,N_9909);
nor UO_1223 (O_1223,N_9970,N_9983);
nor UO_1224 (O_1224,N_9990,N_9958);
nor UO_1225 (O_1225,N_9969,N_9949);
xor UO_1226 (O_1226,N_9987,N_9934);
nor UO_1227 (O_1227,N_9943,N_9912);
xor UO_1228 (O_1228,N_9988,N_9972);
nand UO_1229 (O_1229,N_9940,N_9950);
or UO_1230 (O_1230,N_9952,N_9975);
or UO_1231 (O_1231,N_9901,N_9943);
or UO_1232 (O_1232,N_9995,N_9969);
nor UO_1233 (O_1233,N_9953,N_9916);
and UO_1234 (O_1234,N_9906,N_9998);
nor UO_1235 (O_1235,N_9925,N_9980);
and UO_1236 (O_1236,N_9953,N_9904);
and UO_1237 (O_1237,N_9965,N_9993);
nor UO_1238 (O_1238,N_9984,N_9963);
nor UO_1239 (O_1239,N_9941,N_9963);
or UO_1240 (O_1240,N_9956,N_9955);
nor UO_1241 (O_1241,N_9967,N_9999);
or UO_1242 (O_1242,N_9950,N_9967);
nor UO_1243 (O_1243,N_9986,N_9956);
nand UO_1244 (O_1244,N_9950,N_9974);
nor UO_1245 (O_1245,N_9957,N_9985);
nor UO_1246 (O_1246,N_9948,N_9932);
and UO_1247 (O_1247,N_9977,N_9947);
or UO_1248 (O_1248,N_9932,N_9954);
and UO_1249 (O_1249,N_9919,N_9954);
or UO_1250 (O_1250,N_9947,N_9936);
and UO_1251 (O_1251,N_9945,N_9981);
nor UO_1252 (O_1252,N_9905,N_9960);
nand UO_1253 (O_1253,N_9900,N_9978);
or UO_1254 (O_1254,N_9927,N_9936);
or UO_1255 (O_1255,N_9983,N_9905);
nand UO_1256 (O_1256,N_9999,N_9929);
or UO_1257 (O_1257,N_9911,N_9996);
or UO_1258 (O_1258,N_9931,N_9911);
and UO_1259 (O_1259,N_9987,N_9920);
or UO_1260 (O_1260,N_9902,N_9995);
and UO_1261 (O_1261,N_9966,N_9902);
or UO_1262 (O_1262,N_9986,N_9965);
nand UO_1263 (O_1263,N_9972,N_9979);
nand UO_1264 (O_1264,N_9945,N_9975);
nand UO_1265 (O_1265,N_9934,N_9997);
or UO_1266 (O_1266,N_9950,N_9990);
nand UO_1267 (O_1267,N_9984,N_9967);
nand UO_1268 (O_1268,N_9955,N_9964);
nor UO_1269 (O_1269,N_9959,N_9948);
nor UO_1270 (O_1270,N_9981,N_9965);
or UO_1271 (O_1271,N_9990,N_9904);
or UO_1272 (O_1272,N_9916,N_9942);
nor UO_1273 (O_1273,N_9973,N_9987);
nor UO_1274 (O_1274,N_9915,N_9990);
or UO_1275 (O_1275,N_9946,N_9954);
and UO_1276 (O_1276,N_9976,N_9906);
nor UO_1277 (O_1277,N_9931,N_9944);
nand UO_1278 (O_1278,N_9975,N_9990);
nor UO_1279 (O_1279,N_9991,N_9922);
nand UO_1280 (O_1280,N_9983,N_9909);
nor UO_1281 (O_1281,N_9918,N_9937);
and UO_1282 (O_1282,N_9960,N_9970);
nor UO_1283 (O_1283,N_9958,N_9931);
nor UO_1284 (O_1284,N_9992,N_9928);
or UO_1285 (O_1285,N_9908,N_9996);
xor UO_1286 (O_1286,N_9976,N_9912);
nor UO_1287 (O_1287,N_9950,N_9906);
nor UO_1288 (O_1288,N_9964,N_9994);
nand UO_1289 (O_1289,N_9922,N_9964);
nand UO_1290 (O_1290,N_9955,N_9913);
and UO_1291 (O_1291,N_9901,N_9995);
xnor UO_1292 (O_1292,N_9923,N_9915);
or UO_1293 (O_1293,N_9908,N_9918);
nand UO_1294 (O_1294,N_9972,N_9924);
nand UO_1295 (O_1295,N_9963,N_9932);
or UO_1296 (O_1296,N_9991,N_9979);
and UO_1297 (O_1297,N_9926,N_9905);
nor UO_1298 (O_1298,N_9957,N_9977);
or UO_1299 (O_1299,N_9932,N_9930);
nor UO_1300 (O_1300,N_9945,N_9965);
and UO_1301 (O_1301,N_9900,N_9926);
nor UO_1302 (O_1302,N_9918,N_9972);
nand UO_1303 (O_1303,N_9958,N_9950);
nand UO_1304 (O_1304,N_9943,N_9936);
nor UO_1305 (O_1305,N_9985,N_9933);
and UO_1306 (O_1306,N_9957,N_9983);
nor UO_1307 (O_1307,N_9986,N_9991);
nand UO_1308 (O_1308,N_9983,N_9937);
nor UO_1309 (O_1309,N_9912,N_9932);
or UO_1310 (O_1310,N_9987,N_9906);
nand UO_1311 (O_1311,N_9923,N_9942);
nor UO_1312 (O_1312,N_9995,N_9931);
or UO_1313 (O_1313,N_9994,N_9942);
and UO_1314 (O_1314,N_9943,N_9993);
or UO_1315 (O_1315,N_9948,N_9935);
or UO_1316 (O_1316,N_9936,N_9918);
xnor UO_1317 (O_1317,N_9978,N_9936);
nand UO_1318 (O_1318,N_9967,N_9968);
or UO_1319 (O_1319,N_9911,N_9953);
or UO_1320 (O_1320,N_9961,N_9959);
xor UO_1321 (O_1321,N_9987,N_9960);
and UO_1322 (O_1322,N_9962,N_9921);
or UO_1323 (O_1323,N_9941,N_9992);
nand UO_1324 (O_1324,N_9914,N_9976);
nor UO_1325 (O_1325,N_9924,N_9939);
or UO_1326 (O_1326,N_9956,N_9912);
or UO_1327 (O_1327,N_9969,N_9922);
nand UO_1328 (O_1328,N_9986,N_9932);
or UO_1329 (O_1329,N_9923,N_9906);
or UO_1330 (O_1330,N_9988,N_9962);
nand UO_1331 (O_1331,N_9992,N_9943);
nor UO_1332 (O_1332,N_9971,N_9936);
and UO_1333 (O_1333,N_9937,N_9950);
and UO_1334 (O_1334,N_9915,N_9937);
or UO_1335 (O_1335,N_9904,N_9974);
nor UO_1336 (O_1336,N_9992,N_9993);
nand UO_1337 (O_1337,N_9972,N_9957);
or UO_1338 (O_1338,N_9973,N_9925);
nand UO_1339 (O_1339,N_9993,N_9975);
or UO_1340 (O_1340,N_9940,N_9920);
nand UO_1341 (O_1341,N_9917,N_9973);
or UO_1342 (O_1342,N_9917,N_9989);
and UO_1343 (O_1343,N_9973,N_9928);
or UO_1344 (O_1344,N_9962,N_9995);
nand UO_1345 (O_1345,N_9982,N_9983);
or UO_1346 (O_1346,N_9971,N_9908);
nand UO_1347 (O_1347,N_9960,N_9901);
nand UO_1348 (O_1348,N_9928,N_9974);
nand UO_1349 (O_1349,N_9977,N_9915);
or UO_1350 (O_1350,N_9971,N_9948);
nor UO_1351 (O_1351,N_9904,N_9909);
xor UO_1352 (O_1352,N_9980,N_9987);
nor UO_1353 (O_1353,N_9965,N_9913);
and UO_1354 (O_1354,N_9922,N_9918);
and UO_1355 (O_1355,N_9958,N_9963);
or UO_1356 (O_1356,N_9918,N_9933);
or UO_1357 (O_1357,N_9982,N_9904);
or UO_1358 (O_1358,N_9972,N_9997);
or UO_1359 (O_1359,N_9917,N_9950);
and UO_1360 (O_1360,N_9984,N_9968);
nor UO_1361 (O_1361,N_9976,N_9940);
or UO_1362 (O_1362,N_9919,N_9984);
nor UO_1363 (O_1363,N_9910,N_9976);
and UO_1364 (O_1364,N_9958,N_9969);
and UO_1365 (O_1365,N_9985,N_9996);
nand UO_1366 (O_1366,N_9976,N_9920);
nand UO_1367 (O_1367,N_9982,N_9946);
and UO_1368 (O_1368,N_9926,N_9946);
and UO_1369 (O_1369,N_9911,N_9900);
and UO_1370 (O_1370,N_9919,N_9935);
xnor UO_1371 (O_1371,N_9925,N_9916);
and UO_1372 (O_1372,N_9935,N_9908);
nor UO_1373 (O_1373,N_9967,N_9939);
xor UO_1374 (O_1374,N_9914,N_9983);
nand UO_1375 (O_1375,N_9958,N_9940);
or UO_1376 (O_1376,N_9925,N_9939);
and UO_1377 (O_1377,N_9921,N_9923);
nor UO_1378 (O_1378,N_9987,N_9954);
or UO_1379 (O_1379,N_9981,N_9947);
or UO_1380 (O_1380,N_9924,N_9941);
and UO_1381 (O_1381,N_9975,N_9966);
and UO_1382 (O_1382,N_9970,N_9919);
xor UO_1383 (O_1383,N_9929,N_9942);
nand UO_1384 (O_1384,N_9912,N_9911);
nor UO_1385 (O_1385,N_9973,N_9938);
nor UO_1386 (O_1386,N_9926,N_9933);
nand UO_1387 (O_1387,N_9997,N_9904);
xor UO_1388 (O_1388,N_9922,N_9956);
nor UO_1389 (O_1389,N_9926,N_9962);
or UO_1390 (O_1390,N_9961,N_9909);
and UO_1391 (O_1391,N_9973,N_9954);
and UO_1392 (O_1392,N_9988,N_9951);
nand UO_1393 (O_1393,N_9970,N_9932);
or UO_1394 (O_1394,N_9987,N_9982);
nor UO_1395 (O_1395,N_9941,N_9921);
nor UO_1396 (O_1396,N_9937,N_9976);
or UO_1397 (O_1397,N_9993,N_9904);
nor UO_1398 (O_1398,N_9988,N_9949);
nor UO_1399 (O_1399,N_9922,N_9941);
or UO_1400 (O_1400,N_9984,N_9906);
nand UO_1401 (O_1401,N_9961,N_9956);
or UO_1402 (O_1402,N_9928,N_9950);
and UO_1403 (O_1403,N_9911,N_9949);
nand UO_1404 (O_1404,N_9931,N_9971);
and UO_1405 (O_1405,N_9960,N_9962);
and UO_1406 (O_1406,N_9981,N_9975);
nor UO_1407 (O_1407,N_9911,N_9956);
nor UO_1408 (O_1408,N_9960,N_9968);
or UO_1409 (O_1409,N_9922,N_9972);
or UO_1410 (O_1410,N_9902,N_9906);
nor UO_1411 (O_1411,N_9926,N_9908);
or UO_1412 (O_1412,N_9989,N_9916);
nor UO_1413 (O_1413,N_9940,N_9936);
nand UO_1414 (O_1414,N_9962,N_9943);
nand UO_1415 (O_1415,N_9949,N_9920);
and UO_1416 (O_1416,N_9918,N_9959);
nand UO_1417 (O_1417,N_9967,N_9907);
nand UO_1418 (O_1418,N_9990,N_9956);
and UO_1419 (O_1419,N_9921,N_9904);
nand UO_1420 (O_1420,N_9978,N_9976);
nand UO_1421 (O_1421,N_9906,N_9958);
nand UO_1422 (O_1422,N_9902,N_9930);
nand UO_1423 (O_1423,N_9925,N_9952);
or UO_1424 (O_1424,N_9949,N_9936);
nand UO_1425 (O_1425,N_9949,N_9997);
or UO_1426 (O_1426,N_9979,N_9916);
nor UO_1427 (O_1427,N_9941,N_9910);
nor UO_1428 (O_1428,N_9976,N_9917);
and UO_1429 (O_1429,N_9969,N_9977);
and UO_1430 (O_1430,N_9966,N_9968);
and UO_1431 (O_1431,N_9998,N_9975);
nand UO_1432 (O_1432,N_9934,N_9904);
and UO_1433 (O_1433,N_9904,N_9924);
nor UO_1434 (O_1434,N_9985,N_9907);
nand UO_1435 (O_1435,N_9900,N_9942);
or UO_1436 (O_1436,N_9970,N_9995);
nand UO_1437 (O_1437,N_9920,N_9913);
nand UO_1438 (O_1438,N_9943,N_9972);
and UO_1439 (O_1439,N_9976,N_9908);
or UO_1440 (O_1440,N_9966,N_9980);
nand UO_1441 (O_1441,N_9994,N_9902);
nor UO_1442 (O_1442,N_9994,N_9975);
nand UO_1443 (O_1443,N_9916,N_9903);
and UO_1444 (O_1444,N_9945,N_9921);
and UO_1445 (O_1445,N_9981,N_9906);
nor UO_1446 (O_1446,N_9976,N_9959);
nor UO_1447 (O_1447,N_9968,N_9979);
nand UO_1448 (O_1448,N_9908,N_9919);
nand UO_1449 (O_1449,N_9976,N_9950);
nand UO_1450 (O_1450,N_9905,N_9919);
nor UO_1451 (O_1451,N_9962,N_9979);
nand UO_1452 (O_1452,N_9992,N_9980);
nor UO_1453 (O_1453,N_9960,N_9988);
or UO_1454 (O_1454,N_9959,N_9989);
and UO_1455 (O_1455,N_9998,N_9957);
nor UO_1456 (O_1456,N_9944,N_9934);
or UO_1457 (O_1457,N_9941,N_9936);
nand UO_1458 (O_1458,N_9914,N_9915);
nor UO_1459 (O_1459,N_9914,N_9968);
nand UO_1460 (O_1460,N_9960,N_9922);
or UO_1461 (O_1461,N_9960,N_9981);
or UO_1462 (O_1462,N_9902,N_9929);
or UO_1463 (O_1463,N_9972,N_9959);
nor UO_1464 (O_1464,N_9914,N_9952);
or UO_1465 (O_1465,N_9964,N_9913);
or UO_1466 (O_1466,N_9994,N_9919);
or UO_1467 (O_1467,N_9968,N_9922);
or UO_1468 (O_1468,N_9902,N_9963);
nor UO_1469 (O_1469,N_9974,N_9970);
or UO_1470 (O_1470,N_9973,N_9945);
nor UO_1471 (O_1471,N_9916,N_9911);
nor UO_1472 (O_1472,N_9920,N_9925);
nor UO_1473 (O_1473,N_9974,N_9956);
nor UO_1474 (O_1474,N_9953,N_9961);
nand UO_1475 (O_1475,N_9934,N_9998);
nand UO_1476 (O_1476,N_9971,N_9985);
nand UO_1477 (O_1477,N_9917,N_9996);
nor UO_1478 (O_1478,N_9919,N_9978);
nand UO_1479 (O_1479,N_9933,N_9987);
and UO_1480 (O_1480,N_9948,N_9974);
or UO_1481 (O_1481,N_9927,N_9914);
nor UO_1482 (O_1482,N_9927,N_9935);
nand UO_1483 (O_1483,N_9957,N_9941);
nor UO_1484 (O_1484,N_9904,N_9914);
nor UO_1485 (O_1485,N_9911,N_9995);
and UO_1486 (O_1486,N_9948,N_9960);
or UO_1487 (O_1487,N_9910,N_9948);
or UO_1488 (O_1488,N_9945,N_9977);
nor UO_1489 (O_1489,N_9957,N_9954);
and UO_1490 (O_1490,N_9950,N_9945);
or UO_1491 (O_1491,N_9982,N_9966);
nor UO_1492 (O_1492,N_9959,N_9904);
nor UO_1493 (O_1493,N_9945,N_9972);
nor UO_1494 (O_1494,N_9931,N_9912);
or UO_1495 (O_1495,N_9948,N_9951);
nand UO_1496 (O_1496,N_9910,N_9933);
or UO_1497 (O_1497,N_9921,N_9937);
and UO_1498 (O_1498,N_9930,N_9981);
and UO_1499 (O_1499,N_9985,N_9922);
endmodule