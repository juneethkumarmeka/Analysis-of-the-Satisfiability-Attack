module basic_2000_20000_2500_4_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1972,In_368);
xnor U1 (N_1,In_1290,In_1547);
nor U2 (N_2,In_242,In_361);
and U3 (N_3,In_1429,In_232);
nor U4 (N_4,In_739,In_550);
xor U5 (N_5,In_1339,In_1563);
nor U6 (N_6,In_1103,In_829);
xor U7 (N_7,In_1546,In_1461);
nor U8 (N_8,In_209,In_1861);
nand U9 (N_9,In_1557,In_236);
xnor U10 (N_10,In_1196,In_1410);
nor U11 (N_11,In_435,In_1492);
xnor U12 (N_12,In_668,In_987);
xnor U13 (N_13,In_1783,In_1488);
and U14 (N_14,In_589,In_1685);
xnor U15 (N_15,In_455,In_643);
and U16 (N_16,In_1954,In_59);
nor U17 (N_17,In_304,In_385);
nand U18 (N_18,In_1905,In_146);
xor U19 (N_19,In_960,In_1633);
xor U20 (N_20,In_1042,In_1171);
nand U21 (N_21,In_1707,In_579);
xor U22 (N_22,In_655,In_1239);
nor U23 (N_23,In_339,In_1072);
xnor U24 (N_24,In_111,In_1654);
or U25 (N_25,In_805,In_1074);
or U26 (N_26,In_724,In_605);
or U27 (N_27,In_645,In_1335);
nand U28 (N_28,In_1832,In_1266);
nor U29 (N_29,In_491,In_119);
nand U30 (N_30,In_1645,In_1516);
nor U31 (N_31,In_810,In_623);
nand U32 (N_32,In_1804,In_892);
nor U33 (N_33,In_1921,In_649);
nand U34 (N_34,In_174,In_15);
and U35 (N_35,In_1694,In_944);
nand U36 (N_36,In_858,In_1132);
or U37 (N_37,In_1404,In_969);
and U38 (N_38,In_726,In_1887);
nand U39 (N_39,In_716,In_1891);
nand U40 (N_40,In_1270,In_101);
nand U41 (N_41,In_1330,In_1774);
and U42 (N_42,In_761,In_907);
nand U43 (N_43,In_364,In_603);
or U44 (N_44,In_950,In_1641);
or U45 (N_45,In_1926,In_1279);
and U46 (N_46,In_1894,In_590);
or U47 (N_47,In_483,In_432);
and U48 (N_48,In_1400,In_1054);
nand U49 (N_49,In_79,In_722);
xnor U50 (N_50,In_168,In_1088);
nand U51 (N_51,In_87,In_863);
nor U52 (N_52,In_777,In_67);
nor U53 (N_53,In_417,In_395);
nor U54 (N_54,In_654,In_1969);
nor U55 (N_55,In_1112,In_154);
xor U56 (N_56,In_81,In_1948);
nand U57 (N_57,In_1441,In_1847);
nand U58 (N_58,In_1843,In_634);
xor U59 (N_59,In_865,In_1952);
nand U60 (N_60,In_1159,In_1003);
and U61 (N_61,In_1373,In_1147);
nand U62 (N_62,In_854,In_1082);
nand U63 (N_63,In_6,In_343);
xnor U64 (N_64,In_995,In_1477);
xor U65 (N_65,In_1995,In_1919);
nor U66 (N_66,In_1220,In_1028);
nor U67 (N_67,In_538,In_1090);
and U68 (N_68,In_1217,In_1188);
nand U69 (N_69,In_319,In_793);
nor U70 (N_70,In_307,In_516);
xor U71 (N_71,In_1369,In_115);
or U72 (N_72,In_1793,In_1652);
and U73 (N_73,In_529,In_1614);
and U74 (N_74,In_171,In_1539);
nand U75 (N_75,In_949,In_819);
nor U76 (N_76,In_690,In_331);
nand U77 (N_77,In_1284,In_184);
and U78 (N_78,In_796,In_1045);
or U79 (N_79,In_1880,In_162);
nand U80 (N_80,In_1796,In_815);
xor U81 (N_81,In_1838,In_992);
nor U82 (N_82,In_1318,In_797);
nand U83 (N_83,In_1288,In_1935);
or U84 (N_84,In_720,In_947);
nor U85 (N_85,In_1970,In_1473);
xor U86 (N_86,In_51,In_939);
and U87 (N_87,In_412,In_1937);
or U88 (N_88,In_1742,In_117);
nor U89 (N_89,In_475,In_1570);
or U90 (N_90,In_1665,In_135);
nor U91 (N_91,In_549,In_24);
nand U92 (N_92,In_1020,In_129);
nand U93 (N_93,In_1133,In_1272);
xnor U94 (N_94,In_779,In_98);
and U95 (N_95,In_677,In_1192);
and U96 (N_96,In_57,In_1658);
or U97 (N_97,In_1567,In_1609);
or U98 (N_98,In_1190,In_575);
nor U99 (N_99,In_465,In_457);
and U100 (N_100,In_803,In_1008);
and U101 (N_101,In_225,In_635);
or U102 (N_102,In_1485,In_1022);
nor U103 (N_103,In_1223,In_1786);
and U104 (N_104,In_1913,In_835);
and U105 (N_105,In_956,In_888);
nor U106 (N_106,In_1390,In_1210);
and U107 (N_107,In_1924,In_1545);
or U108 (N_108,In_1690,In_340);
nand U109 (N_109,In_1490,In_91);
nor U110 (N_110,In_394,In_1755);
xnor U111 (N_111,In_1237,In_261);
nor U112 (N_112,In_1585,In_825);
and U113 (N_113,In_1635,In_1012);
and U114 (N_114,In_229,In_1494);
or U115 (N_115,In_164,In_186);
nand U116 (N_116,In_1602,In_1256);
nand U117 (N_117,In_1254,In_822);
and U118 (N_118,In_638,In_1476);
xnor U119 (N_119,In_1606,In_99);
nand U120 (N_120,In_1401,In_192);
and U121 (N_121,In_1138,In_561);
or U122 (N_122,In_29,In_856);
and U123 (N_123,In_790,In_109);
or U124 (N_124,In_1696,In_287);
and U125 (N_125,In_1487,In_1077);
or U126 (N_126,In_673,In_305);
or U127 (N_127,In_1912,In_1358);
xnor U128 (N_128,In_1992,In_1039);
nor U129 (N_129,In_734,In_1918);
and U130 (N_130,In_1505,In_1999);
xor U131 (N_131,In_134,In_130);
xnor U132 (N_132,In_1174,In_1693);
nand U133 (N_133,In_272,In_723);
and U134 (N_134,In_1803,In_985);
nand U135 (N_135,In_1666,In_826);
or U136 (N_136,In_861,In_1826);
nor U137 (N_137,In_131,In_539);
or U138 (N_138,In_1058,In_180);
nor U139 (N_139,In_1961,In_1509);
and U140 (N_140,In_1865,In_970);
or U141 (N_141,In_884,In_660);
and U142 (N_142,In_317,In_398);
xor U143 (N_143,In_872,In_1319);
and U144 (N_144,In_1885,In_1517);
nand U145 (N_145,In_1756,In_1303);
nand U146 (N_146,In_1914,In_1428);
xnor U147 (N_147,In_1399,In_1361);
and U148 (N_148,In_836,In_844);
nand U149 (N_149,In_1483,In_243);
nand U150 (N_150,In_85,In_1357);
nand U151 (N_151,In_1629,In_363);
xnor U152 (N_152,In_1260,In_818);
or U153 (N_153,In_619,In_1382);
xnor U154 (N_154,In_569,In_1586);
xnor U155 (N_155,In_837,In_166);
and U156 (N_156,In_1548,In_1197);
xnor U157 (N_157,In_568,In_1491);
and U158 (N_158,In_543,In_778);
nand U159 (N_159,In_1562,In_606);
nor U160 (N_160,In_1148,In_1381);
xor U161 (N_161,In_631,In_1640);
or U162 (N_162,In_1285,In_1314);
nand U163 (N_163,In_239,In_9);
and U164 (N_164,In_766,In_1734);
nand U165 (N_165,In_1458,In_1018);
or U166 (N_166,In_915,In_507);
nand U167 (N_167,In_1255,In_775);
nor U168 (N_168,In_625,In_306);
or U169 (N_169,In_1544,In_1376);
nor U170 (N_170,In_592,In_1471);
nor U171 (N_171,In_1438,In_883);
nor U172 (N_172,In_185,In_757);
or U173 (N_173,In_452,In_1317);
xnor U174 (N_174,In_1202,In_383);
nor U175 (N_175,In_1825,In_1713);
or U176 (N_176,In_1501,In_867);
and U177 (N_177,In_403,In_782);
nor U178 (N_178,In_1868,In_687);
nor U179 (N_179,In_324,In_1819);
nand U180 (N_180,In_1712,In_714);
or U181 (N_181,In_1437,In_429);
or U182 (N_182,In_629,In_509);
nor U183 (N_183,In_1958,In_431);
nor U184 (N_184,In_372,In_1730);
and U185 (N_185,In_293,In_1026);
and U186 (N_186,In_842,In_1176);
and U187 (N_187,In_83,In_1522);
nand U188 (N_188,In_1396,In_441);
or U189 (N_189,In_551,In_1642);
nor U190 (N_190,In_212,In_1809);
or U191 (N_191,In_1289,In_160);
or U192 (N_192,In_1834,In_418);
and U193 (N_193,In_375,In_607);
and U194 (N_194,In_273,In_1007);
or U195 (N_195,In_1717,In_968);
and U196 (N_196,In_1205,In_128);
nor U197 (N_197,In_963,In_313);
and U198 (N_198,In_1247,In_1909);
nand U199 (N_199,In_444,In_315);
and U200 (N_200,In_1395,In_546);
or U201 (N_201,In_1189,In_1157);
and U202 (N_202,In_989,In_641);
or U203 (N_203,In_898,In_20);
nand U204 (N_204,In_1449,In_637);
nor U205 (N_205,In_27,In_1346);
nand U206 (N_206,In_1542,In_1497);
or U207 (N_207,In_528,In_682);
xor U208 (N_208,In_1768,In_1788);
and U209 (N_209,In_505,In_70);
xor U210 (N_210,In_1735,In_337);
or U211 (N_211,In_750,In_536);
or U212 (N_212,In_1676,In_1044);
xnor U213 (N_213,In_1597,In_1725);
and U214 (N_214,In_1340,In_1244);
xnor U215 (N_215,In_1662,In_857);
or U216 (N_216,In_1064,In_489);
nand U217 (N_217,In_1114,In_1309);
nor U218 (N_218,In_1455,In_280);
or U219 (N_219,In_1448,In_1822);
xor U220 (N_220,In_1594,In_769);
and U221 (N_221,In_86,In_1257);
nand U222 (N_222,In_903,In_610);
and U223 (N_223,In_1384,In_1840);
nor U224 (N_224,In_500,In_233);
nand U225 (N_225,In_1776,In_584);
nor U226 (N_226,In_646,In_650);
nand U227 (N_227,In_1737,In_1094);
nand U228 (N_228,In_1038,In_1718);
nand U229 (N_229,In_367,In_787);
or U230 (N_230,In_1475,In_833);
nand U231 (N_231,In_583,In_34);
nor U232 (N_232,In_1261,In_602);
or U233 (N_233,In_1632,In_1910);
nand U234 (N_234,In_295,In_1356);
nand U235 (N_235,In_1278,In_449);
nor U236 (N_236,In_1808,In_917);
or U237 (N_237,In_1086,In_627);
nor U238 (N_238,In_308,In_406);
nor U239 (N_239,In_399,In_674);
or U240 (N_240,In_920,In_1502);
or U241 (N_241,In_862,In_1705);
and U242 (N_242,In_1785,In_227);
and U243 (N_243,In_824,In_215);
nand U244 (N_244,In_1343,In_1017);
or U245 (N_245,In_934,In_1554);
nand U246 (N_246,In_1025,In_1328);
xnor U247 (N_247,In_1418,In_163);
nand U248 (N_248,In_1583,In_26);
xor U249 (N_249,In_1050,In_1081);
and U250 (N_250,In_453,In_585);
xor U251 (N_251,In_1160,In_1375);
nor U252 (N_252,In_1150,In_1234);
and U253 (N_253,In_1230,In_43);
nand U254 (N_254,In_1224,In_1552);
xor U255 (N_255,In_515,In_176);
nand U256 (N_256,In_159,In_699);
or U257 (N_257,In_1214,In_999);
nor U258 (N_258,In_1744,In_1681);
and U259 (N_259,In_1656,In_1127);
nor U260 (N_260,In_1538,In_1610);
xnor U261 (N_261,In_143,In_1365);
nor U262 (N_262,In_1582,In_876);
and U263 (N_263,In_990,In_541);
and U264 (N_264,In_1442,In_1432);
or U265 (N_265,In_942,In_1839);
nand U266 (N_266,In_1794,In_523);
nor U267 (N_267,In_1049,In_289);
and U268 (N_268,In_95,In_1252);
nand U269 (N_269,In_878,In_1967);
nor U270 (N_270,In_19,In_731);
nand U271 (N_271,In_1661,In_746);
and U272 (N_272,In_1630,In_1218);
nor U273 (N_273,In_1648,In_1782);
xnor U274 (N_274,In_1499,In_203);
nor U275 (N_275,In_423,In_710);
and U276 (N_276,In_460,In_1878);
or U277 (N_277,In_852,In_1055);
nand U278 (N_278,In_1144,In_1638);
xor U279 (N_279,In_997,In_1037);
and U280 (N_280,In_1164,In_977);
nor U281 (N_281,In_61,In_44);
and U282 (N_282,In_1061,In_198);
or U283 (N_283,In_576,In_381);
and U284 (N_284,In_1312,In_1805);
and U285 (N_285,In_821,In_1882);
nand U286 (N_286,In_1033,In_150);
nor U287 (N_287,In_1659,In_1149);
and U288 (N_288,In_378,In_598);
nor U289 (N_289,In_1864,In_1075);
nor U290 (N_290,In_1298,In_1875);
and U291 (N_291,In_329,In_595);
nand U292 (N_292,In_1116,In_632);
nand U293 (N_293,In_50,In_1079);
and U294 (N_294,In_369,In_1683);
and U295 (N_295,In_902,In_848);
or U296 (N_296,In_18,In_374);
and U297 (N_297,In_1564,In_1519);
xnor U298 (N_298,In_330,In_1844);
nand U299 (N_299,In_284,In_873);
nand U300 (N_300,In_38,In_1431);
or U301 (N_301,In_1985,In_952);
and U302 (N_302,In_401,In_1355);
nand U303 (N_303,In_1593,In_1953);
nand U304 (N_304,In_662,In_1308);
nor U305 (N_305,In_653,In_1946);
or U306 (N_306,In_1753,In_113);
nand U307 (N_307,In_1615,In_341);
xor U308 (N_308,In_809,In_554);
nor U309 (N_309,In_1858,In_1812);
nand U310 (N_310,In_1463,In_820);
nand U311 (N_311,In_1626,In_633);
or U312 (N_312,In_925,In_1345);
or U313 (N_313,In_735,In_1076);
or U314 (N_314,In_1336,In_588);
or U315 (N_315,In_1657,In_1708);
nor U316 (N_316,In_889,In_1169);
xnor U317 (N_317,In_1349,In_1293);
or U318 (N_318,In_1670,In_1010);
nand U319 (N_319,In_88,In_139);
and U320 (N_320,In_1226,In_1925);
and U321 (N_321,In_1679,In_748);
and U322 (N_322,In_376,In_182);
or U323 (N_323,In_651,In_1903);
and U324 (N_324,In_1684,In_1265);
or U325 (N_325,In_832,In_379);
and U326 (N_326,In_1286,In_122);
and U327 (N_327,In_234,In_350);
and U328 (N_328,In_336,In_979);
nor U329 (N_329,In_183,In_303);
nand U330 (N_330,In_228,In_428);
nor U331 (N_331,In_194,In_1013);
and U332 (N_332,In_1801,In_1974);
or U333 (N_333,In_998,In_351);
nand U334 (N_334,In_165,In_1815);
nor U335 (N_335,In_933,In_1886);
or U336 (N_336,In_278,In_1555);
and U337 (N_337,In_1019,In_1850);
nand U338 (N_338,In_1321,In_1829);
and U339 (N_339,In_1740,In_1398);
and U340 (N_340,In_108,In_1813);
or U341 (N_341,In_1917,In_1470);
nor U342 (N_342,In_614,In_244);
or U343 (N_343,In_807,In_846);
nor U344 (N_344,In_1631,In_1978);
nand U345 (N_345,In_1599,In_1514);
nor U346 (N_346,In_1619,In_1622);
nand U347 (N_347,In_1863,In_657);
nand U348 (N_348,In_1818,In_1739);
and U349 (N_349,In_359,In_1367);
and U350 (N_350,In_1040,In_78);
nor U351 (N_351,In_525,In_1559);
xor U352 (N_352,In_1093,In_1062);
and U353 (N_353,In_25,In_1498);
and U354 (N_354,In_436,In_235);
or U355 (N_355,In_488,In_1787);
xnor U356 (N_356,In_1763,In_1089);
nor U357 (N_357,In_864,In_1837);
or U358 (N_358,In_1922,In_768);
nor U359 (N_359,In_1806,In_1830);
xnor U360 (N_360,In_1268,In_537);
or U361 (N_361,In_397,In_1853);
nand U362 (N_362,In_1080,In_1927);
nand U363 (N_363,In_1173,In_972);
or U364 (N_364,In_895,In_695);
and U365 (N_365,In_301,In_1817);
or U366 (N_366,In_971,In_388);
and U367 (N_367,In_811,In_532);
and U368 (N_368,In_258,In_1030);
xnor U369 (N_369,In_1551,In_1047);
and U370 (N_370,In_260,In_1469);
or U371 (N_371,In_249,In_1294);
and U372 (N_372,In_953,In_1024);
nor U373 (N_373,In_238,In_1348);
or U374 (N_374,In_207,In_1493);
nor U375 (N_375,In_446,In_574);
and U376 (N_376,In_210,In_22);
nand U377 (N_377,In_1736,In_983);
or U378 (N_378,In_23,In_1206);
or U379 (N_379,In_202,In_1137);
nor U380 (N_380,In_1411,In_149);
and U381 (N_381,In_1747,In_1452);
nand U382 (N_382,In_591,In_580);
nor U383 (N_383,In_1757,In_1553);
or U384 (N_384,In_1561,In_494);
nor U385 (N_385,In_1084,In_36);
xnor U386 (N_386,In_615,In_103);
nand U387 (N_387,In_1253,In_840);
xnor U388 (N_388,In_1417,In_599);
nand U389 (N_389,In_1118,In_1750);
or U390 (N_390,In_497,In_503);
or U391 (N_391,In_1211,In_1415);
or U392 (N_392,In_937,In_1179);
nand U393 (N_393,In_1503,In_1621);
nor U394 (N_394,In_1569,In_175);
or U395 (N_395,In_611,In_573);
and U396 (N_396,In_1724,In_1456);
nor U397 (N_397,In_1238,In_422);
nand U398 (N_398,In_1034,In_326);
nand U399 (N_399,In_335,In_1233);
nor U400 (N_400,In_1109,In_439);
nor U401 (N_401,In_1784,In_1091);
nor U402 (N_402,In_252,In_1986);
nand U403 (N_403,In_1264,In_1678);
and U404 (N_404,In_984,In_754);
or U405 (N_405,In_530,In_365);
nand U406 (N_406,In_1393,In_1126);
or U407 (N_407,In_64,In_269);
nand U408 (N_408,In_430,In_373);
nor U409 (N_409,In_1354,In_725);
nor U410 (N_410,In_962,In_996);
nand U411 (N_411,In_1532,In_948);
or U412 (N_412,In_1352,In_743);
nor U413 (N_413,In_2,In_706);
or U414 (N_414,In_679,In_1957);
xnor U415 (N_415,In_594,In_1916);
nand U416 (N_416,In_112,In_981);
xor U417 (N_417,In_749,In_348);
nor U418 (N_418,In_1388,In_262);
nor U419 (N_419,In_389,In_1588);
nand U420 (N_420,In_954,In_945);
or U421 (N_421,In_425,In_1027);
nor U422 (N_422,In_1960,In_358);
or U423 (N_423,In_1966,In_717);
nor U424 (N_424,In_562,In_1980);
or U425 (N_425,In_104,In_776);
and U426 (N_426,In_416,In_991);
xnor U427 (N_427,In_1625,In_63);
or U428 (N_428,In_461,In_1835);
nor U429 (N_429,In_1623,In_1883);
or U430 (N_430,In_66,In_675);
nand U431 (N_431,In_738,In_410);
nor U432 (N_432,In_1472,In_181);
and U433 (N_433,In_1928,In_1484);
or U434 (N_434,In_1125,In_1406);
and U435 (N_435,In_493,In_1950);
xor U436 (N_436,In_97,In_292);
or U437 (N_437,In_1011,In_1711);
nand U438 (N_438,In_581,In_1496);
nor U439 (N_439,In_46,In_297);
and U440 (N_440,In_1274,In_451);
nor U441 (N_441,In_666,In_285);
nor U442 (N_442,In_1892,In_386);
or U443 (N_443,In_147,In_1325);
xor U444 (N_444,In_1113,In_1479);
nand U445 (N_445,In_762,In_1489);
nand U446 (N_446,In_1549,In_1823);
and U447 (N_447,In_886,In_900);
nand U448 (N_448,In_1647,In_563);
or U449 (N_449,In_1703,In_1246);
or U450 (N_450,In_676,In_770);
nand U451 (N_451,In_1001,In_800);
nor U452 (N_452,In_978,In_1162);
or U453 (N_453,In_1453,In_1624);
nor U454 (N_454,In_1715,In_1200);
nor U455 (N_455,In_1754,In_681);
nor U456 (N_456,In_231,In_535);
and U457 (N_457,In_1212,In_1964);
nand U458 (N_458,In_1752,In_1041);
or U459 (N_459,In_1374,In_760);
and U460 (N_460,In_1122,In_1984);
nand U461 (N_461,In_327,In_1566);
nor U462 (N_462,In_193,In_780);
and U463 (N_463,In_890,In_736);
or U464 (N_464,In_555,In_1771);
nor U465 (N_465,In_189,In_1152);
xor U466 (N_466,In_459,In_72);
and U467 (N_467,In_314,In_853);
nor U468 (N_468,In_464,In_1899);
and U469 (N_469,In_290,In_642);
xnor U470 (N_470,In_1603,In_524);
or U471 (N_471,In_1136,In_1414);
or U472 (N_472,In_578,In_1379);
and U473 (N_473,In_1889,In_908);
and U474 (N_474,In_941,In_1722);
or U475 (N_475,In_121,In_1762);
nand U476 (N_476,In_1009,In_909);
xor U477 (N_477,In_1616,In_1350);
or U478 (N_478,In_434,In_1102);
or U479 (N_479,In_1764,In_709);
and U480 (N_480,In_1720,In_893);
nand U481 (N_481,In_1031,In_37);
and U482 (N_482,In_448,In_1550);
nor U483 (N_483,In_1675,In_1191);
or U484 (N_484,In_1856,In_1135);
or U485 (N_485,In_1478,In_1228);
and U486 (N_486,In_1251,In_1976);
xor U487 (N_487,In_1920,In_1153);
or U488 (N_488,In_47,In_201);
or U489 (N_489,In_1576,In_366);
or U490 (N_490,In_966,In_798);
nor U491 (N_491,In_1209,In_703);
and U492 (N_492,In_698,In_744);
nand U493 (N_493,In_1636,In_1151);
nor U494 (N_494,In_1460,In_1650);
xnor U495 (N_495,In_700,In_799);
and U496 (N_496,In_1526,In_1177);
and U497 (N_497,In_1474,In_849);
nor U498 (N_498,In_254,In_1291);
or U499 (N_499,In_1423,In_1944);
nor U500 (N_500,In_1016,In_1262);
or U501 (N_501,In_1110,In_1165);
and U502 (N_502,In_82,In_414);
or U503 (N_503,In_622,In_1271);
nand U504 (N_504,In_318,In_302);
or U505 (N_505,In_1095,In_1997);
or U506 (N_506,In_1377,In_683);
nor U507 (N_507,In_1653,In_1777);
nor U508 (N_508,In_1486,In_1901);
nand U509 (N_509,In_1575,In_114);
nand U510 (N_510,In_1359,In_1433);
and U511 (N_511,In_964,In_499);
and U512 (N_512,In_71,In_1107);
or U513 (N_513,In_609,In_1389);
nand U514 (N_514,In_1897,In_344);
and U515 (N_515,In_1236,In_771);
and U516 (N_516,In_1962,In_473);
and U517 (N_517,In_1723,In_1518);
nand U518 (N_518,In_1341,In_899);
and U519 (N_519,In_1930,In_1536);
or U520 (N_520,In_1700,In_880);
nor U521 (N_521,In_355,In_1193);
nor U522 (N_522,In_1326,In_1971);
or U523 (N_523,In_1344,In_172);
xor U524 (N_524,In_1385,In_237);
nor U525 (N_525,In_1605,In_747);
nand U526 (N_526,In_1166,In_16);
or U527 (N_527,In_1911,In_1070);
nor U528 (N_528,In_173,In_1836);
and U529 (N_529,In_35,In_1316);
and U530 (N_530,In_851,In_1408);
and U531 (N_531,In_1945,In_794);
or U532 (N_532,In_567,In_1896);
and U533 (N_533,In_1380,In_5);
or U534 (N_534,In_1120,In_792);
and U535 (N_535,In_1881,In_409);
xor U536 (N_536,In_1347,In_100);
and U537 (N_537,In_76,In_456);
or U538 (N_538,In_1668,In_808);
nor U539 (N_539,In_152,In_1180);
nand U540 (N_540,In_1426,In_1989);
nand U541 (N_541,In_1577,In_496);
xnor U542 (N_542,In_1871,In_138);
nor U543 (N_543,In_795,In_906);
and U544 (N_544,In_10,In_1994);
nor U545 (N_545,In_1904,In_268);
nand U546 (N_546,In_1391,In_1006);
or U547 (N_547,In_1851,In_1759);
or U548 (N_548,In_1761,In_1129);
or U549 (N_549,In_1436,In_391);
nand U550 (N_550,In_1184,In_380);
or U551 (N_551,In_1821,In_1592);
or U552 (N_552,In_1424,In_582);
or U553 (N_553,In_600,In_1387);
nor U554 (N_554,In_407,In_993);
or U555 (N_555,In_466,In_1158);
or U556 (N_556,In_1056,In_1186);
or U557 (N_557,In_1249,In_156);
nand U558 (N_558,In_1140,In_501);
nand U559 (N_559,In_1620,In_360);
nor U560 (N_560,In_1363,In_1907);
and U561 (N_561,In_1760,In_74);
and U562 (N_562,In_1955,In_1595);
and U563 (N_563,In_267,In_1541);
nand U564 (N_564,In_1331,In_1182);
and U565 (N_565,In_1779,In_932);
and U566 (N_566,In_1168,In_765);
xor U567 (N_567,In_1568,In_1324);
or U568 (N_568,In_891,In_1301);
nor U569 (N_569,In_691,In_1259);
and U570 (N_570,In_357,In_1227);
and U571 (N_571,In_1726,In_1686);
nand U572 (N_572,In_1500,In_1195);
or U573 (N_573,In_1134,In_255);
nor U574 (N_574,In_640,In_479);
xor U575 (N_575,In_190,In_1530);
nor U576 (N_576,In_1248,In_120);
xor U577 (N_577,In_1746,In_1307);
and U578 (N_578,In_1420,In_316);
and U579 (N_579,In_45,In_197);
xor U580 (N_580,In_294,In_1059);
or U581 (N_581,In_125,In_859);
and U582 (N_582,In_1982,In_1695);
nand U583 (N_583,In_450,In_1691);
and U584 (N_584,In_392,In_1680);
nand U585 (N_585,In_1183,In_241);
nand U586 (N_586,In_1213,In_1895);
nand U587 (N_587,In_1280,In_1612);
or U588 (N_588,In_1032,In_843);
or U589 (N_589,In_1991,In_1397);
and U590 (N_590,In_253,In_106);
nand U591 (N_591,In_879,In_1807);
and U592 (N_592,In_245,In_427);
nand U593 (N_593,In_1462,In_1527);
nor U594 (N_594,In_1877,In_1512);
or U595 (N_595,In_1101,In_1596);
or U596 (N_596,In_542,In_141);
nand U597 (N_597,In_916,In_105);
and U598 (N_598,In_1827,In_1071);
or U599 (N_599,In_564,In_1731);
nor U600 (N_600,In_1281,In_1313);
nand U601 (N_601,In_1673,In_613);
nand U602 (N_602,In_12,In_264);
and U603 (N_603,In_930,In_404);
nand U604 (N_604,In_1204,In_58);
or U605 (N_605,In_547,In_1445);
and U606 (N_606,In_155,In_1579);
nor U607 (N_607,In_1578,In_1781);
nand U608 (N_608,In_759,In_785);
nand U609 (N_609,In_957,In_1879);
nor U610 (N_610,In_1353,In_1600);
nand U611 (N_611,In_1772,In_847);
nor U612 (N_612,In_1310,In_1123);
xor U613 (N_613,In_1304,In_1671);
nand U614 (N_614,In_1323,In_1608);
and U615 (N_615,In_1506,In_1692);
or U616 (N_616,In_151,In_1275);
and U617 (N_617,In_680,In_1156);
and U618 (N_618,In_1300,In_1508);
nand U619 (N_619,In_1015,In_636);
and U620 (N_620,In_310,In_1085);
nor U621 (N_621,In_1060,In_1743);
xnor U622 (N_622,In_887,In_323);
and U623 (N_623,In_299,In_1874);
and U624 (N_624,In_1951,In_974);
and U625 (N_625,In_756,In_572);
and U626 (N_626,In_158,In_1117);
and U627 (N_627,In_733,In_1528);
nand U628 (N_628,In_177,In_1959);
nor U629 (N_629,In_338,In_552);
or U630 (N_630,In_1852,In_8);
nor U631 (N_631,In_1601,In_387);
nand U632 (N_632,In_1131,In_1245);
nor U633 (N_633,In_1128,In_30);
or U634 (N_634,In_1667,In_1322);
or U635 (N_635,In_1721,In_1689);
and U636 (N_636,In_871,In_896);
or U637 (N_637,In_630,In_1701);
nor U638 (N_638,In_1185,In_1524);
or U639 (N_639,In_1523,In_1175);
and U640 (N_640,In_571,In_89);
nand U641 (N_641,In_1208,In_692);
or U642 (N_642,In_1362,In_1146);
and U643 (N_643,In_1219,In_1464);
nand U644 (N_644,In_943,In_1933);
nor U645 (N_645,In_1956,In_1811);
or U646 (N_646,In_1097,In_1360);
nand U647 (N_647,In_148,In_1590);
and U648 (N_648,In_1078,In_1338);
nor U649 (N_649,In_828,In_877);
and U650 (N_650,In_1607,In_1987);
or U651 (N_651,In_712,In_553);
or U652 (N_652,In_188,In_411);
nand U653 (N_653,In_226,In_926);
nor U654 (N_654,In_923,In_144);
nor U655 (N_655,In_1993,In_1366);
nand U656 (N_656,In_170,In_628);
or U657 (N_657,In_1857,In_624);
nand U658 (N_658,In_965,In_1687);
nand U659 (N_659,In_1697,In_1073);
or U660 (N_660,In_1108,In_931);
or U661 (N_661,In_1949,In_526);
nor U662 (N_662,In_1181,In_1198);
nand U663 (N_663,In_413,In_1005);
nand U664 (N_664,In_1828,In_975);
xor U665 (N_665,In_1651,In_65);
nand U666 (N_666,In_1618,In_498);
or U667 (N_667,In_755,In_586);
nand U668 (N_668,In_684,In_283);
and U669 (N_669,In_1143,In_1450);
and U670 (N_670,In_322,In_77);
and U671 (N_671,In_1565,In_958);
and U672 (N_672,In_1728,In_764);
nor U673 (N_673,In_1051,In_1466);
nand U674 (N_674,In_727,In_558);
nand U675 (N_675,In_474,In_1351);
nor U676 (N_676,In_1422,In_1067);
nand U677 (N_677,In_1515,In_309);
nand U678 (N_678,In_1407,In_1646);
nand U679 (N_679,In_1704,In_1589);
or U680 (N_680,In_13,In_685);
xor U681 (N_681,In_342,In_534);
or U682 (N_682,In_885,In_982);
xnor U683 (N_683,In_905,In_1121);
or U684 (N_684,In_1446,In_772);
nor U685 (N_685,In_270,In_1792);
or U686 (N_686,In_266,In_1163);
nand U687 (N_687,In_626,In_1482);
or U688 (N_688,In_663,In_1447);
xor U689 (N_689,In_1888,In_352);
or U690 (N_690,In_1273,In_1370);
nand U691 (N_691,In_482,In_904);
nand U692 (N_692,In_263,In_545);
or U693 (N_693,In_1002,In_223);
and U694 (N_694,In_393,In_328);
nor U695 (N_695,In_90,In_1800);
or U696 (N_696,In_195,In_1591);
and U697 (N_697,In_565,In_277);
nor U698 (N_698,In_39,In_831);
and U699 (N_699,In_659,In_702);
and U700 (N_700,In_897,In_1587);
and U701 (N_701,In_1664,In_1021);
nor U702 (N_702,In_1241,In_1315);
nor U703 (N_703,In_502,In_478);
xnor U704 (N_704,In_929,In_214);
nand U705 (N_705,In_251,In_1797);
nor U706 (N_706,In_31,In_69);
nor U707 (N_707,In_531,In_1604);
xnor U708 (N_708,In_1915,In_1543);
nor U709 (N_709,In_1104,In_813);
nor U710 (N_710,In_1378,In_1581);
nor U711 (N_711,In_1029,In_80);
or U712 (N_712,In_806,In_689);
xnor U713 (N_713,In_1766,In_577);
nand U714 (N_714,In_1444,In_1520);
or U715 (N_715,In_1232,In_1048);
and U716 (N_716,In_462,In_356);
and U717 (N_717,In_737,In_1337);
nand U718 (N_718,In_1816,In_1057);
nor U719 (N_719,In_1403,In_935);
and U720 (N_720,In_719,In_205);
and U721 (N_721,In_1611,In_652);
or U722 (N_722,In_53,In_1710);
xor U723 (N_723,In_1627,In_219);
or U724 (N_724,In_415,In_1714);
nand U725 (N_725,In_1155,In_1833);
and U726 (N_726,In_84,In_1867);
nand U727 (N_727,In_21,In_298);
xnor U728 (N_728,In_40,In_276);
and U729 (N_729,In_447,In_1440);
and U730 (N_730,In_882,In_1068);
xnor U731 (N_731,In_1296,In_1225);
or U732 (N_732,In_1859,In_14);
nor U733 (N_733,In_566,In_639);
and U734 (N_734,In_1412,In_914);
and U735 (N_735,In_783,In_1709);
nand U736 (N_736,In_533,In_1299);
nor U737 (N_737,In_1820,In_1170);
nand U738 (N_738,In_729,In_1855);
nand U739 (N_739,In_1556,In_490);
nor U740 (N_740,In_1814,In_596);
or U741 (N_741,In_587,In_132);
nand U742 (N_742,In_1977,In_522);
or U743 (N_743,In_850,In_52);
nor U744 (N_744,In_901,In_325);
nor U745 (N_745,In_157,In_213);
or U746 (N_746,In_1222,In_938);
and U747 (N_747,In_495,In_257);
and U748 (N_748,In_838,In_894);
nor U749 (N_749,In_1035,In_1457);
or U750 (N_750,In_1053,In_1111);
and U751 (N_751,In_463,In_1902);
nor U752 (N_752,In_1405,In_1332);
nor U753 (N_753,In_1965,In_230);
nand U754 (N_754,In_767,In_711);
or U755 (N_755,In_1574,In_1751);
and U756 (N_756,In_1119,In_196);
or U757 (N_757,In_1719,In_616);
or U758 (N_758,In_845,In_1099);
xor U759 (N_759,In_1311,In_480);
nand U760 (N_760,In_922,In_1884);
and U761 (N_761,In_140,In_275);
or U762 (N_762,In_1167,In_1791);
xnor U763 (N_763,In_199,In_1936);
and U764 (N_764,In_1115,In_694);
or U765 (N_765,In_951,In_918);
and U766 (N_766,In_752,In_520);
nor U767 (N_767,In_1923,In_116);
nand U768 (N_768,In_707,In_1229);
nor U769 (N_769,In_454,In_1846);
nand U770 (N_770,In_3,In_1706);
or U771 (N_771,In_443,In_1802);
or U772 (N_772,In_1467,In_1748);
or U773 (N_773,In_7,In_708);
nand U774 (N_774,In_1947,In_1529);
or U775 (N_775,In_644,In_704);
nor U776 (N_776,In_1287,In_870);
nor U777 (N_777,In_1451,In_320);
xor U778 (N_778,In_1320,In_1283);
nand U779 (N_779,In_127,In_1409);
or U780 (N_780,In_426,In_1908);
nor U781 (N_781,In_468,In_1824);
nand U782 (N_782,In_286,In_910);
nand U783 (N_783,In_1534,In_955);
nand U784 (N_784,In_1014,In_1617);
or U785 (N_785,In_1780,In_521);
nand U786 (N_786,In_142,In_1990);
and U787 (N_787,In_559,In_1799);
or U788 (N_788,In_1682,In_486);
and U789 (N_789,In_1106,In_1773);
nor U790 (N_790,In_370,In_1573);
and U791 (N_791,In_1327,In_153);
and U792 (N_792,In_1770,In_48);
and U793 (N_793,In_476,In_178);
or U794 (N_794,In_1968,In_208);
and U795 (N_795,In_1201,In_1672);
nor U796 (N_796,In_382,In_93);
nor U797 (N_797,In_1943,In_492);
and U798 (N_798,In_1277,In_1);
and U799 (N_799,In_994,In_656);
and U800 (N_800,In_1386,In_216);
nand U801 (N_801,In_669,In_1963);
nor U802 (N_802,In_869,In_1372);
nand U803 (N_803,In_1677,In_1975);
or U804 (N_804,In_1216,In_1465);
and U805 (N_805,In_1983,In_73);
nand U806 (N_806,In_224,In_556);
nor U807 (N_807,In_1235,In_1434);
nand U808 (N_808,In_333,In_671);
nor U809 (N_809,In_1000,In_672);
and U810 (N_810,In_874,In_1934);
nand U811 (N_811,In_54,In_321);
and U812 (N_812,In_265,In_1540);
nor U813 (N_813,In_1297,In_256);
and U814 (N_814,In_508,In_1087);
or U815 (N_815,In_485,In_1854);
xnor U816 (N_816,In_697,In_1130);
or U817 (N_817,In_220,In_927);
and U818 (N_818,In_940,In_1810);
xnor U819 (N_819,In_1942,In_300);
xnor U820 (N_820,In_1481,In_353);
nor U821 (N_821,In_1269,In_211);
nor U822 (N_822,In_1525,In_1243);
nand U823 (N_823,In_118,In_1402);
and U824 (N_824,In_1172,In_728);
nand U825 (N_825,In_1276,In_973);
or U826 (N_826,In_1267,In_1727);
nand U827 (N_827,In_647,In_601);
or U828 (N_828,In_161,In_1221);
or U829 (N_829,In_1758,In_980);
nand U830 (N_830,In_620,In_248);
and U831 (N_831,In_511,In_126);
nand U832 (N_832,In_467,In_812);
or U833 (N_833,In_1906,In_390);
and U834 (N_834,In_1207,In_1383);
nand U835 (N_835,In_1639,In_1124);
and U836 (N_836,In_1394,In_259);
xor U837 (N_837,In_1749,In_597);
nand U838 (N_838,In_1778,In_402);
or U839 (N_839,In_1900,In_788);
nand U840 (N_840,In_32,In_1870);
nor U841 (N_841,In_1872,In_621);
nand U842 (N_842,In_1741,In_1511);
or U843 (N_843,In_274,In_107);
or U844 (N_844,In_1250,In_1427);
nand U845 (N_845,In_312,In_701);
and U846 (N_846,In_124,In_1775);
and U847 (N_847,In_961,In_472);
and U848 (N_848,In_1425,In_247);
or U849 (N_849,In_911,In_1092);
xor U850 (N_850,In_802,In_1535);
and U851 (N_851,In_804,In_763);
xor U852 (N_852,In_1178,In_354);
xor U853 (N_853,In_1215,In_217);
nand U854 (N_854,In_741,In_1435);
nand U855 (N_855,In_967,In_1860);
and U856 (N_856,In_1795,In_271);
nor U857 (N_857,In_688,In_713);
and U858 (N_858,In_1558,In_433);
nand U859 (N_859,In_200,In_1765);
nand U860 (N_860,In_41,In_222);
nand U861 (N_861,In_123,In_834);
nand U862 (N_862,In_1613,In_1932);
and U863 (N_863,In_740,In_512);
and U864 (N_864,In_1981,In_1674);
and U865 (N_865,In_1069,In_868);
xor U866 (N_866,In_718,In_1100);
and U867 (N_867,In_1584,In_1258);
and U868 (N_868,In_1729,In_1716);
nor U869 (N_869,In_408,In_218);
xor U870 (N_870,In_470,In_1702);
xnor U871 (N_871,In_191,In_1798);
and U872 (N_872,In_618,In_1142);
or U873 (N_873,In_514,In_540);
or U874 (N_874,In_693,In_875);
nor U875 (N_875,In_686,In_936);
nor U876 (N_876,In_946,In_1628);
and U877 (N_877,In_221,In_347);
xor U878 (N_878,In_55,In_0);
nand U879 (N_879,In_1413,In_570);
and U880 (N_880,In_445,In_830);
or U881 (N_881,In_1890,In_1295);
xnor U882 (N_882,In_919,In_419);
nand U883 (N_883,In_506,In_1733);
or U884 (N_884,In_1510,In_1831);
nand U885 (N_885,In_1979,In_1507);
or U886 (N_886,In_477,In_786);
nand U887 (N_887,In_167,In_240);
and U888 (N_888,In_481,In_1789);
and U889 (N_889,In_371,In_421);
and U890 (N_890,In_1660,In_742);
and U891 (N_891,In_1096,In_1052);
or U892 (N_892,In_1521,In_593);
or U893 (N_893,In_732,In_1698);
nor U894 (N_894,In_400,In_924);
nor U895 (N_895,In_1841,In_1199);
and U896 (N_896,In_544,In_1845);
or U897 (N_897,In_1419,In_1580);
nand U898 (N_898,In_246,In_437);
or U899 (N_899,In_1898,In_1893);
and U900 (N_900,In_1043,In_548);
nand U901 (N_901,In_696,In_137);
nand U902 (N_902,In_1572,In_291);
and U903 (N_903,In_1392,In_49);
and U904 (N_904,In_1848,In_1537);
or U905 (N_905,In_1066,In_1939);
xnor U906 (N_906,In_866,In_1098);
nor U907 (N_907,In_661,In_1988);
nand U908 (N_908,In_557,In_396);
and U909 (N_909,In_1154,In_334);
or U910 (N_910,In_204,In_384);
xnor U911 (N_911,In_1329,In_1421);
nand U912 (N_912,In_206,In_362);
or U913 (N_913,In_1141,In_1416);
nor U914 (N_914,In_1459,In_841);
and U915 (N_915,In_179,In_1842);
and U916 (N_916,In_773,In_658);
and U917 (N_917,In_1036,In_721);
or U918 (N_918,In_484,In_1065);
and U919 (N_919,In_1263,In_1866);
or U920 (N_920,In_518,In_133);
and U921 (N_921,In_513,In_110);
nor U922 (N_922,In_1699,In_487);
nand U923 (N_923,In_1430,In_1306);
nor U924 (N_924,In_1480,In_816);
nor U925 (N_925,In_560,In_791);
nand U926 (N_926,In_1849,In_855);
xor U927 (N_927,In_33,In_730);
and U928 (N_928,In_420,In_1745);
nand U929 (N_929,In_1873,In_928);
and U930 (N_930,In_442,In_1139);
and U931 (N_931,In_1371,In_1333);
nand U932 (N_932,In_774,In_881);
nand U933 (N_933,In_617,In_1083);
nor U934 (N_934,In_1292,In_1203);
or U935 (N_935,In_753,In_281);
or U936 (N_936,In_751,In_1996);
and U937 (N_937,In_976,In_1941);
nor U938 (N_938,In_28,In_1938);
xor U939 (N_939,In_1663,In_187);
or U940 (N_940,In_801,In_1998);
nand U941 (N_941,In_527,In_664);
or U942 (N_942,In_279,In_1187);
nor U943 (N_943,In_405,In_1732);
nand U944 (N_944,In_517,In_823);
nor U945 (N_945,In_648,In_504);
or U946 (N_946,In_1302,In_510);
and U947 (N_947,In_781,In_1240);
or U948 (N_948,In_1454,In_670);
nand U949 (N_949,In_288,In_1004);
nor U950 (N_950,In_68,In_912);
nand U951 (N_951,In_250,In_469);
xnor U952 (N_952,In_311,In_1334);
xor U953 (N_953,In_11,In_1533);
nand U954 (N_954,In_665,In_705);
nor U955 (N_955,In_60,In_1443);
or U956 (N_956,In_440,In_438);
nand U957 (N_957,In_1504,In_745);
nand U958 (N_958,In_986,In_1046);
or U959 (N_959,In_345,In_1973);
or U960 (N_960,In_169,In_62);
nand U961 (N_961,In_1637,In_519);
and U962 (N_962,In_1862,In_377);
or U963 (N_963,In_1242,In_1869);
xnor U964 (N_964,In_282,In_92);
or U965 (N_965,In_817,In_1876);
or U966 (N_966,In_1023,In_1105);
and U967 (N_967,In_604,In_1644);
or U968 (N_968,In_1364,In_17);
xnor U969 (N_969,In_1634,In_608);
xor U970 (N_970,In_827,In_678);
or U971 (N_971,In_458,In_471);
nand U972 (N_972,In_94,In_1931);
nor U973 (N_973,In_1769,In_1194);
or U974 (N_974,In_346,In_96);
or U975 (N_975,In_1342,In_1649);
nor U976 (N_976,In_4,In_1439);
xor U977 (N_977,In_42,In_1282);
nor U978 (N_978,In_1598,In_758);
and U979 (N_979,In_56,In_1643);
and U980 (N_980,In_1305,In_75);
nand U981 (N_981,In_1231,In_1688);
and U982 (N_982,In_296,In_1513);
nand U983 (N_983,In_1571,In_1767);
or U984 (N_984,In_1790,In_860);
and U985 (N_985,In_102,In_1669);
nand U986 (N_986,In_913,In_1161);
and U987 (N_987,In_1940,In_814);
nor U988 (N_988,In_1145,In_1468);
or U989 (N_989,In_1738,In_332);
xor U990 (N_990,In_136,In_145);
and U991 (N_991,In_1655,In_667);
and U992 (N_992,In_424,In_715);
nand U993 (N_993,In_789,In_1063);
or U994 (N_994,In_1368,In_1929);
and U995 (N_995,In_839,In_988);
nor U996 (N_996,In_1531,In_784);
nor U997 (N_997,In_349,In_612);
nor U998 (N_998,In_921,In_1560);
or U999 (N_999,In_1495,In_959);
nand U1000 (N_1000,In_479,In_1343);
nand U1001 (N_1001,In_1284,In_770);
nor U1002 (N_1002,In_1864,In_1928);
and U1003 (N_1003,In_377,In_933);
or U1004 (N_1004,In_1939,In_1573);
nor U1005 (N_1005,In_1614,In_1179);
nor U1006 (N_1006,In_422,In_400);
and U1007 (N_1007,In_158,In_907);
or U1008 (N_1008,In_1712,In_166);
and U1009 (N_1009,In_1971,In_1452);
or U1010 (N_1010,In_847,In_604);
nand U1011 (N_1011,In_633,In_916);
nor U1012 (N_1012,In_262,In_138);
and U1013 (N_1013,In_1389,In_917);
nand U1014 (N_1014,In_605,In_1383);
nand U1015 (N_1015,In_1381,In_1617);
nor U1016 (N_1016,In_420,In_309);
xor U1017 (N_1017,In_837,In_1935);
nand U1018 (N_1018,In_561,In_153);
or U1019 (N_1019,In_1656,In_292);
nor U1020 (N_1020,In_1044,In_969);
or U1021 (N_1021,In_409,In_1674);
nor U1022 (N_1022,In_317,In_1253);
or U1023 (N_1023,In_462,In_1133);
nand U1024 (N_1024,In_683,In_911);
nor U1025 (N_1025,In_1548,In_1488);
nor U1026 (N_1026,In_1706,In_1472);
or U1027 (N_1027,In_1935,In_189);
nand U1028 (N_1028,In_1400,In_1639);
nand U1029 (N_1029,In_1940,In_1197);
and U1030 (N_1030,In_375,In_609);
nand U1031 (N_1031,In_962,In_127);
and U1032 (N_1032,In_1745,In_1200);
nand U1033 (N_1033,In_337,In_23);
or U1034 (N_1034,In_545,In_876);
nor U1035 (N_1035,In_591,In_1136);
nand U1036 (N_1036,In_499,In_513);
nand U1037 (N_1037,In_1403,In_1479);
and U1038 (N_1038,In_1450,In_1025);
and U1039 (N_1039,In_949,In_377);
xnor U1040 (N_1040,In_1958,In_472);
and U1041 (N_1041,In_65,In_620);
nand U1042 (N_1042,In_759,In_256);
or U1043 (N_1043,In_383,In_879);
xor U1044 (N_1044,In_937,In_14);
and U1045 (N_1045,In_1079,In_41);
and U1046 (N_1046,In_700,In_419);
nor U1047 (N_1047,In_1453,In_737);
nor U1048 (N_1048,In_456,In_892);
or U1049 (N_1049,In_505,In_1558);
nor U1050 (N_1050,In_1107,In_416);
and U1051 (N_1051,In_748,In_240);
or U1052 (N_1052,In_731,In_1118);
or U1053 (N_1053,In_1648,In_543);
or U1054 (N_1054,In_736,In_349);
or U1055 (N_1055,In_738,In_1554);
nand U1056 (N_1056,In_1133,In_9);
or U1057 (N_1057,In_692,In_194);
nand U1058 (N_1058,In_845,In_1158);
nand U1059 (N_1059,In_1872,In_1664);
nor U1060 (N_1060,In_1475,In_265);
or U1061 (N_1061,In_9,In_1548);
and U1062 (N_1062,In_56,In_6);
xor U1063 (N_1063,In_394,In_1763);
or U1064 (N_1064,In_33,In_1713);
nor U1065 (N_1065,In_847,In_1962);
or U1066 (N_1066,In_1031,In_79);
or U1067 (N_1067,In_1001,In_1036);
and U1068 (N_1068,In_1789,In_114);
or U1069 (N_1069,In_3,In_1501);
nand U1070 (N_1070,In_1746,In_920);
nor U1071 (N_1071,In_191,In_1277);
nand U1072 (N_1072,In_1208,In_1122);
and U1073 (N_1073,In_424,In_895);
or U1074 (N_1074,In_53,In_1554);
and U1075 (N_1075,In_813,In_804);
nand U1076 (N_1076,In_1039,In_822);
nor U1077 (N_1077,In_1586,In_1225);
nand U1078 (N_1078,In_1055,In_1409);
and U1079 (N_1079,In_1174,In_1835);
nor U1080 (N_1080,In_366,In_1491);
and U1081 (N_1081,In_1353,In_1378);
xnor U1082 (N_1082,In_437,In_245);
nor U1083 (N_1083,In_1702,In_649);
xnor U1084 (N_1084,In_558,In_816);
or U1085 (N_1085,In_307,In_800);
and U1086 (N_1086,In_1481,In_392);
nand U1087 (N_1087,In_1186,In_1117);
or U1088 (N_1088,In_672,In_1249);
or U1089 (N_1089,In_1521,In_1639);
and U1090 (N_1090,In_804,In_235);
nor U1091 (N_1091,In_108,In_963);
nand U1092 (N_1092,In_768,In_1817);
and U1093 (N_1093,In_1103,In_555);
or U1094 (N_1094,In_532,In_459);
or U1095 (N_1095,In_771,In_1002);
and U1096 (N_1096,In_1570,In_1554);
nor U1097 (N_1097,In_167,In_1776);
nor U1098 (N_1098,In_1575,In_369);
nand U1099 (N_1099,In_754,In_1592);
or U1100 (N_1100,In_1229,In_5);
and U1101 (N_1101,In_528,In_214);
nor U1102 (N_1102,In_1525,In_424);
and U1103 (N_1103,In_1004,In_1196);
or U1104 (N_1104,In_454,In_722);
nor U1105 (N_1105,In_766,In_1253);
and U1106 (N_1106,In_1174,In_203);
nor U1107 (N_1107,In_649,In_826);
and U1108 (N_1108,In_489,In_77);
nand U1109 (N_1109,In_619,In_1835);
nand U1110 (N_1110,In_218,In_791);
nor U1111 (N_1111,In_1075,In_1093);
nand U1112 (N_1112,In_1777,In_1200);
nor U1113 (N_1113,In_687,In_1560);
nand U1114 (N_1114,In_1773,In_485);
xnor U1115 (N_1115,In_100,In_436);
and U1116 (N_1116,In_1240,In_1349);
and U1117 (N_1117,In_582,In_1742);
xnor U1118 (N_1118,In_1425,In_1257);
and U1119 (N_1119,In_1744,In_632);
nor U1120 (N_1120,In_1447,In_960);
and U1121 (N_1121,In_440,In_1095);
or U1122 (N_1122,In_50,In_891);
xnor U1123 (N_1123,In_1046,In_1329);
nor U1124 (N_1124,In_585,In_1867);
and U1125 (N_1125,In_94,In_406);
or U1126 (N_1126,In_1317,In_82);
and U1127 (N_1127,In_913,In_1847);
nor U1128 (N_1128,In_936,In_517);
nor U1129 (N_1129,In_480,In_1146);
nor U1130 (N_1130,In_1,In_433);
or U1131 (N_1131,In_219,In_612);
and U1132 (N_1132,In_29,In_1052);
nor U1133 (N_1133,In_1530,In_1145);
and U1134 (N_1134,In_1133,In_1711);
nor U1135 (N_1135,In_161,In_1690);
nand U1136 (N_1136,In_176,In_13);
nor U1137 (N_1137,In_1957,In_457);
nor U1138 (N_1138,In_1698,In_533);
nor U1139 (N_1139,In_1170,In_33);
xor U1140 (N_1140,In_1744,In_1344);
or U1141 (N_1141,In_266,In_1853);
and U1142 (N_1142,In_1750,In_797);
nor U1143 (N_1143,In_978,In_1396);
and U1144 (N_1144,In_1142,In_229);
or U1145 (N_1145,In_813,In_1102);
nor U1146 (N_1146,In_635,In_358);
and U1147 (N_1147,In_872,In_864);
nand U1148 (N_1148,In_1924,In_1950);
or U1149 (N_1149,In_1776,In_34);
nor U1150 (N_1150,In_548,In_364);
nand U1151 (N_1151,In_1437,In_1412);
and U1152 (N_1152,In_580,In_482);
nor U1153 (N_1153,In_1952,In_75);
nor U1154 (N_1154,In_109,In_466);
or U1155 (N_1155,In_1972,In_1721);
or U1156 (N_1156,In_372,In_1431);
nor U1157 (N_1157,In_222,In_962);
nand U1158 (N_1158,In_1870,In_640);
nand U1159 (N_1159,In_37,In_715);
nor U1160 (N_1160,In_1752,In_1619);
and U1161 (N_1161,In_642,In_367);
and U1162 (N_1162,In_1559,In_274);
or U1163 (N_1163,In_1669,In_1602);
nand U1164 (N_1164,In_270,In_1615);
nor U1165 (N_1165,In_1869,In_574);
xor U1166 (N_1166,In_1400,In_1153);
nor U1167 (N_1167,In_1841,In_1594);
or U1168 (N_1168,In_1878,In_906);
nand U1169 (N_1169,In_324,In_601);
nor U1170 (N_1170,In_11,In_1987);
nand U1171 (N_1171,In_1246,In_1871);
nor U1172 (N_1172,In_20,In_371);
or U1173 (N_1173,In_299,In_1513);
nor U1174 (N_1174,In_1491,In_743);
nand U1175 (N_1175,In_1066,In_1919);
or U1176 (N_1176,In_1475,In_327);
or U1177 (N_1177,In_1748,In_620);
nor U1178 (N_1178,In_1025,In_1760);
and U1179 (N_1179,In_955,In_139);
or U1180 (N_1180,In_1740,In_123);
nand U1181 (N_1181,In_42,In_44);
and U1182 (N_1182,In_180,In_1777);
and U1183 (N_1183,In_220,In_1984);
nor U1184 (N_1184,In_714,In_1144);
nor U1185 (N_1185,In_1490,In_656);
nand U1186 (N_1186,In_1627,In_1500);
nand U1187 (N_1187,In_1877,In_1198);
nand U1188 (N_1188,In_67,In_1541);
or U1189 (N_1189,In_598,In_1905);
nand U1190 (N_1190,In_538,In_1415);
or U1191 (N_1191,In_1360,In_1041);
or U1192 (N_1192,In_150,In_1408);
or U1193 (N_1193,In_60,In_1049);
nand U1194 (N_1194,In_1163,In_913);
and U1195 (N_1195,In_1103,In_14);
and U1196 (N_1196,In_406,In_1277);
or U1197 (N_1197,In_954,In_547);
nor U1198 (N_1198,In_1419,In_1945);
nand U1199 (N_1199,In_654,In_1560);
xnor U1200 (N_1200,In_1378,In_634);
or U1201 (N_1201,In_776,In_1557);
nand U1202 (N_1202,In_891,In_1865);
nand U1203 (N_1203,In_1990,In_1980);
nor U1204 (N_1204,In_1746,In_1827);
nor U1205 (N_1205,In_710,In_1410);
nor U1206 (N_1206,In_1638,In_552);
or U1207 (N_1207,In_980,In_525);
nor U1208 (N_1208,In_1279,In_1723);
and U1209 (N_1209,In_1603,In_179);
or U1210 (N_1210,In_1413,In_1428);
nand U1211 (N_1211,In_1136,In_431);
or U1212 (N_1212,In_1829,In_202);
and U1213 (N_1213,In_537,In_181);
or U1214 (N_1214,In_532,In_292);
nand U1215 (N_1215,In_374,In_579);
nor U1216 (N_1216,In_549,In_1316);
xnor U1217 (N_1217,In_1314,In_1927);
nand U1218 (N_1218,In_706,In_911);
nand U1219 (N_1219,In_1488,In_1799);
or U1220 (N_1220,In_1178,In_1550);
nor U1221 (N_1221,In_1487,In_842);
nor U1222 (N_1222,In_61,In_631);
xnor U1223 (N_1223,In_1134,In_284);
nand U1224 (N_1224,In_1686,In_940);
and U1225 (N_1225,In_1793,In_1851);
or U1226 (N_1226,In_600,In_748);
nand U1227 (N_1227,In_378,In_375);
nor U1228 (N_1228,In_248,In_709);
and U1229 (N_1229,In_387,In_339);
and U1230 (N_1230,In_1119,In_341);
nand U1231 (N_1231,In_42,In_1425);
nor U1232 (N_1232,In_1026,In_1157);
nor U1233 (N_1233,In_465,In_1934);
nand U1234 (N_1234,In_462,In_354);
and U1235 (N_1235,In_757,In_1193);
and U1236 (N_1236,In_517,In_333);
and U1237 (N_1237,In_686,In_1950);
or U1238 (N_1238,In_267,In_1076);
and U1239 (N_1239,In_858,In_394);
and U1240 (N_1240,In_1613,In_109);
xor U1241 (N_1241,In_1178,In_266);
or U1242 (N_1242,In_841,In_606);
or U1243 (N_1243,In_1535,In_54);
or U1244 (N_1244,In_361,In_313);
nor U1245 (N_1245,In_936,In_691);
nor U1246 (N_1246,In_571,In_1790);
or U1247 (N_1247,In_1563,In_1809);
nor U1248 (N_1248,In_451,In_338);
nand U1249 (N_1249,In_382,In_1792);
and U1250 (N_1250,In_665,In_1157);
xnor U1251 (N_1251,In_1171,In_1269);
or U1252 (N_1252,In_863,In_1072);
and U1253 (N_1253,In_1197,In_1550);
or U1254 (N_1254,In_1139,In_1302);
and U1255 (N_1255,In_1628,In_1911);
and U1256 (N_1256,In_899,In_1775);
and U1257 (N_1257,In_1749,In_1222);
nand U1258 (N_1258,In_1993,In_109);
nand U1259 (N_1259,In_1417,In_1319);
and U1260 (N_1260,In_1830,In_611);
nand U1261 (N_1261,In_1263,In_149);
nand U1262 (N_1262,In_1201,In_1086);
or U1263 (N_1263,In_1349,In_387);
nand U1264 (N_1264,In_1698,In_996);
xor U1265 (N_1265,In_344,In_139);
and U1266 (N_1266,In_1477,In_1603);
or U1267 (N_1267,In_1222,In_288);
nand U1268 (N_1268,In_298,In_1221);
nor U1269 (N_1269,In_1455,In_1682);
or U1270 (N_1270,In_1211,In_220);
and U1271 (N_1271,In_1070,In_473);
nor U1272 (N_1272,In_1478,In_106);
nor U1273 (N_1273,In_221,In_1309);
nor U1274 (N_1274,In_430,In_1214);
or U1275 (N_1275,In_833,In_678);
nand U1276 (N_1276,In_889,In_1811);
nand U1277 (N_1277,In_965,In_1898);
nand U1278 (N_1278,In_1564,In_1821);
or U1279 (N_1279,In_399,In_1650);
and U1280 (N_1280,In_427,In_1948);
xor U1281 (N_1281,In_941,In_424);
or U1282 (N_1282,In_493,In_1853);
or U1283 (N_1283,In_1269,In_1307);
xnor U1284 (N_1284,In_500,In_1856);
or U1285 (N_1285,In_1584,In_1618);
or U1286 (N_1286,In_1736,In_1831);
nand U1287 (N_1287,In_810,In_1703);
nand U1288 (N_1288,In_1448,In_1547);
nor U1289 (N_1289,In_243,In_488);
and U1290 (N_1290,In_928,In_1861);
or U1291 (N_1291,In_380,In_1487);
or U1292 (N_1292,In_928,In_1213);
and U1293 (N_1293,In_1746,In_240);
nor U1294 (N_1294,In_439,In_1130);
and U1295 (N_1295,In_1182,In_608);
nand U1296 (N_1296,In_1386,In_219);
nor U1297 (N_1297,In_428,In_1196);
nor U1298 (N_1298,In_684,In_386);
or U1299 (N_1299,In_298,In_433);
or U1300 (N_1300,In_1699,In_1787);
nor U1301 (N_1301,In_1189,In_1322);
xnor U1302 (N_1302,In_451,In_1742);
nor U1303 (N_1303,In_1894,In_1954);
nand U1304 (N_1304,In_900,In_540);
xor U1305 (N_1305,In_1921,In_1862);
or U1306 (N_1306,In_26,In_1387);
nor U1307 (N_1307,In_1441,In_322);
nand U1308 (N_1308,In_775,In_541);
xor U1309 (N_1309,In_1851,In_1488);
or U1310 (N_1310,In_1979,In_1011);
and U1311 (N_1311,In_864,In_1799);
or U1312 (N_1312,In_718,In_1468);
xor U1313 (N_1313,In_223,In_1052);
and U1314 (N_1314,In_1265,In_147);
nor U1315 (N_1315,In_1650,In_1153);
nor U1316 (N_1316,In_1950,In_1525);
and U1317 (N_1317,In_1783,In_1953);
nor U1318 (N_1318,In_1307,In_1052);
and U1319 (N_1319,In_1159,In_1278);
and U1320 (N_1320,In_958,In_374);
xnor U1321 (N_1321,In_47,In_364);
or U1322 (N_1322,In_1121,In_1525);
nor U1323 (N_1323,In_382,In_547);
nand U1324 (N_1324,In_1351,In_382);
xor U1325 (N_1325,In_352,In_396);
nand U1326 (N_1326,In_1514,In_1338);
or U1327 (N_1327,In_1903,In_378);
nor U1328 (N_1328,In_827,In_475);
and U1329 (N_1329,In_920,In_1220);
or U1330 (N_1330,In_677,In_1172);
xnor U1331 (N_1331,In_866,In_1561);
and U1332 (N_1332,In_1300,In_682);
xnor U1333 (N_1333,In_1661,In_819);
nor U1334 (N_1334,In_1612,In_1583);
and U1335 (N_1335,In_819,In_1881);
and U1336 (N_1336,In_272,In_65);
and U1337 (N_1337,In_1408,In_768);
or U1338 (N_1338,In_366,In_1620);
nor U1339 (N_1339,In_613,In_1762);
and U1340 (N_1340,In_1436,In_675);
nand U1341 (N_1341,In_773,In_1639);
or U1342 (N_1342,In_1984,In_1653);
or U1343 (N_1343,In_1318,In_1790);
nor U1344 (N_1344,In_169,In_647);
xor U1345 (N_1345,In_1029,In_872);
xnor U1346 (N_1346,In_1866,In_674);
nand U1347 (N_1347,In_474,In_1525);
nand U1348 (N_1348,In_879,In_858);
and U1349 (N_1349,In_1486,In_1450);
and U1350 (N_1350,In_752,In_1803);
nor U1351 (N_1351,In_1089,In_1124);
nand U1352 (N_1352,In_1836,In_1113);
or U1353 (N_1353,In_1844,In_745);
nand U1354 (N_1354,In_1413,In_1940);
nor U1355 (N_1355,In_447,In_1081);
xnor U1356 (N_1356,In_1037,In_65);
xnor U1357 (N_1357,In_533,In_908);
and U1358 (N_1358,In_131,In_1928);
and U1359 (N_1359,In_510,In_339);
and U1360 (N_1360,In_227,In_22);
or U1361 (N_1361,In_1288,In_755);
nor U1362 (N_1362,In_1363,In_699);
and U1363 (N_1363,In_338,In_557);
and U1364 (N_1364,In_1929,In_1775);
nand U1365 (N_1365,In_1028,In_634);
nand U1366 (N_1366,In_1136,In_192);
nor U1367 (N_1367,In_1109,In_678);
and U1368 (N_1368,In_1272,In_1625);
or U1369 (N_1369,In_281,In_101);
and U1370 (N_1370,In_491,In_228);
xor U1371 (N_1371,In_1409,In_886);
and U1372 (N_1372,In_1306,In_385);
or U1373 (N_1373,In_1966,In_210);
or U1374 (N_1374,In_76,In_1798);
nand U1375 (N_1375,In_217,In_115);
nor U1376 (N_1376,In_1689,In_1124);
and U1377 (N_1377,In_1605,In_482);
and U1378 (N_1378,In_154,In_1407);
and U1379 (N_1379,In_1258,In_1373);
and U1380 (N_1380,In_1289,In_622);
and U1381 (N_1381,In_1222,In_1864);
nand U1382 (N_1382,In_998,In_1980);
nor U1383 (N_1383,In_453,In_597);
and U1384 (N_1384,In_13,In_127);
nand U1385 (N_1385,In_1460,In_1811);
or U1386 (N_1386,In_1892,In_959);
or U1387 (N_1387,In_481,In_1069);
xor U1388 (N_1388,In_295,In_243);
and U1389 (N_1389,In_973,In_1345);
nor U1390 (N_1390,In_178,In_586);
and U1391 (N_1391,In_1923,In_1703);
and U1392 (N_1392,In_374,In_1810);
nor U1393 (N_1393,In_720,In_1204);
nor U1394 (N_1394,In_1283,In_1977);
and U1395 (N_1395,In_1835,In_1456);
or U1396 (N_1396,In_1884,In_1107);
or U1397 (N_1397,In_915,In_1257);
nand U1398 (N_1398,In_262,In_1856);
nor U1399 (N_1399,In_683,In_1965);
nand U1400 (N_1400,In_1354,In_1455);
xor U1401 (N_1401,In_1990,In_281);
and U1402 (N_1402,In_1149,In_200);
nor U1403 (N_1403,In_373,In_968);
nand U1404 (N_1404,In_740,In_1045);
and U1405 (N_1405,In_1253,In_1478);
or U1406 (N_1406,In_864,In_1509);
nor U1407 (N_1407,In_1339,In_1453);
or U1408 (N_1408,In_1149,In_186);
nor U1409 (N_1409,In_1024,In_1122);
nor U1410 (N_1410,In_165,In_863);
nand U1411 (N_1411,In_664,In_863);
or U1412 (N_1412,In_1920,In_633);
or U1413 (N_1413,In_850,In_1327);
or U1414 (N_1414,In_929,In_1001);
xnor U1415 (N_1415,In_117,In_1124);
and U1416 (N_1416,In_226,In_402);
nor U1417 (N_1417,In_1095,In_424);
and U1418 (N_1418,In_705,In_282);
and U1419 (N_1419,In_484,In_979);
nand U1420 (N_1420,In_1767,In_183);
xnor U1421 (N_1421,In_133,In_864);
nor U1422 (N_1422,In_896,In_121);
nand U1423 (N_1423,In_959,In_645);
or U1424 (N_1424,In_499,In_1739);
nor U1425 (N_1425,In_1422,In_1715);
xor U1426 (N_1426,In_113,In_610);
xor U1427 (N_1427,In_584,In_1451);
nand U1428 (N_1428,In_1495,In_1887);
nand U1429 (N_1429,In_371,In_451);
nand U1430 (N_1430,In_1032,In_1179);
and U1431 (N_1431,In_1017,In_137);
xnor U1432 (N_1432,In_1282,In_311);
and U1433 (N_1433,In_1245,In_1225);
nand U1434 (N_1434,In_1821,In_830);
or U1435 (N_1435,In_1745,In_881);
or U1436 (N_1436,In_1056,In_140);
nor U1437 (N_1437,In_1036,In_875);
or U1438 (N_1438,In_1639,In_1347);
and U1439 (N_1439,In_1376,In_425);
nor U1440 (N_1440,In_1699,In_673);
and U1441 (N_1441,In_1861,In_356);
or U1442 (N_1442,In_904,In_492);
or U1443 (N_1443,In_336,In_1492);
nand U1444 (N_1444,In_924,In_1935);
nand U1445 (N_1445,In_1798,In_1908);
xor U1446 (N_1446,In_1384,In_1281);
or U1447 (N_1447,In_38,In_1780);
nand U1448 (N_1448,In_866,In_1748);
nand U1449 (N_1449,In_256,In_508);
nand U1450 (N_1450,In_974,In_884);
nand U1451 (N_1451,In_829,In_1312);
nor U1452 (N_1452,In_1230,In_627);
xor U1453 (N_1453,In_177,In_155);
or U1454 (N_1454,In_1997,In_289);
or U1455 (N_1455,In_376,In_1571);
nand U1456 (N_1456,In_520,In_64);
nor U1457 (N_1457,In_1673,In_1179);
or U1458 (N_1458,In_296,In_1499);
or U1459 (N_1459,In_1986,In_1014);
or U1460 (N_1460,In_673,In_685);
or U1461 (N_1461,In_591,In_788);
xnor U1462 (N_1462,In_1758,In_1888);
nor U1463 (N_1463,In_149,In_1743);
or U1464 (N_1464,In_1870,In_75);
or U1465 (N_1465,In_415,In_1277);
xor U1466 (N_1466,In_1916,In_830);
nand U1467 (N_1467,In_118,In_1636);
nor U1468 (N_1468,In_451,In_1806);
or U1469 (N_1469,In_470,In_1930);
and U1470 (N_1470,In_718,In_761);
and U1471 (N_1471,In_1445,In_1106);
or U1472 (N_1472,In_1963,In_1252);
xor U1473 (N_1473,In_1075,In_1361);
nor U1474 (N_1474,In_142,In_1668);
and U1475 (N_1475,In_1412,In_641);
xnor U1476 (N_1476,In_1625,In_1173);
nand U1477 (N_1477,In_1568,In_803);
and U1478 (N_1478,In_1768,In_60);
or U1479 (N_1479,In_609,In_1856);
nor U1480 (N_1480,In_1123,In_453);
or U1481 (N_1481,In_527,In_1234);
and U1482 (N_1482,In_1231,In_1643);
or U1483 (N_1483,In_753,In_1346);
or U1484 (N_1484,In_630,In_985);
or U1485 (N_1485,In_1523,In_253);
nor U1486 (N_1486,In_1359,In_1408);
nand U1487 (N_1487,In_1660,In_296);
and U1488 (N_1488,In_30,In_1448);
nand U1489 (N_1489,In_538,In_1177);
or U1490 (N_1490,In_404,In_313);
and U1491 (N_1491,In_1372,In_1039);
nor U1492 (N_1492,In_587,In_1413);
and U1493 (N_1493,In_693,In_1087);
and U1494 (N_1494,In_1081,In_1631);
nand U1495 (N_1495,In_1040,In_1981);
nand U1496 (N_1496,In_1329,In_61);
or U1497 (N_1497,In_1028,In_24);
or U1498 (N_1498,In_162,In_1522);
or U1499 (N_1499,In_1416,In_1147);
or U1500 (N_1500,In_1513,In_444);
nor U1501 (N_1501,In_1073,In_781);
nand U1502 (N_1502,In_1232,In_851);
nand U1503 (N_1503,In_641,In_1805);
and U1504 (N_1504,In_1571,In_1990);
nand U1505 (N_1505,In_140,In_1513);
nor U1506 (N_1506,In_553,In_893);
and U1507 (N_1507,In_822,In_740);
xor U1508 (N_1508,In_1594,In_342);
nand U1509 (N_1509,In_469,In_174);
or U1510 (N_1510,In_739,In_1655);
nand U1511 (N_1511,In_1098,In_564);
nor U1512 (N_1512,In_1937,In_964);
nor U1513 (N_1513,In_591,In_1909);
or U1514 (N_1514,In_1404,In_812);
and U1515 (N_1515,In_743,In_580);
or U1516 (N_1516,In_1634,In_1194);
nor U1517 (N_1517,In_1151,In_1332);
or U1518 (N_1518,In_1487,In_246);
or U1519 (N_1519,In_1022,In_468);
and U1520 (N_1520,In_683,In_655);
or U1521 (N_1521,In_1371,In_1270);
xor U1522 (N_1522,In_1334,In_120);
nor U1523 (N_1523,In_668,In_1373);
or U1524 (N_1524,In_19,In_1731);
nand U1525 (N_1525,In_497,In_881);
nand U1526 (N_1526,In_1022,In_491);
or U1527 (N_1527,In_42,In_653);
nor U1528 (N_1528,In_1720,In_1695);
or U1529 (N_1529,In_1811,In_922);
nor U1530 (N_1530,In_281,In_1921);
or U1531 (N_1531,In_1905,In_542);
nor U1532 (N_1532,In_1159,In_832);
nand U1533 (N_1533,In_328,In_854);
nand U1534 (N_1534,In_780,In_410);
and U1535 (N_1535,In_5,In_1838);
nor U1536 (N_1536,In_542,In_1832);
nand U1537 (N_1537,In_1538,In_1375);
xnor U1538 (N_1538,In_1225,In_1113);
or U1539 (N_1539,In_1125,In_1893);
nor U1540 (N_1540,In_1110,In_130);
nand U1541 (N_1541,In_545,In_550);
or U1542 (N_1542,In_1527,In_314);
nand U1543 (N_1543,In_854,In_550);
and U1544 (N_1544,In_606,In_1447);
xnor U1545 (N_1545,In_980,In_703);
nor U1546 (N_1546,In_1224,In_766);
nand U1547 (N_1547,In_790,In_1426);
and U1548 (N_1548,In_377,In_563);
or U1549 (N_1549,In_398,In_1562);
or U1550 (N_1550,In_1711,In_1577);
or U1551 (N_1551,In_417,In_1771);
or U1552 (N_1552,In_1787,In_663);
or U1553 (N_1553,In_1802,In_1057);
or U1554 (N_1554,In_518,In_752);
nor U1555 (N_1555,In_371,In_546);
or U1556 (N_1556,In_1246,In_1560);
and U1557 (N_1557,In_906,In_1334);
or U1558 (N_1558,In_1014,In_579);
and U1559 (N_1559,In_730,In_1171);
and U1560 (N_1560,In_46,In_870);
nand U1561 (N_1561,In_883,In_1819);
and U1562 (N_1562,In_531,In_837);
and U1563 (N_1563,In_476,In_969);
or U1564 (N_1564,In_1609,In_375);
nor U1565 (N_1565,In_1492,In_300);
nand U1566 (N_1566,In_1504,In_1943);
nor U1567 (N_1567,In_1701,In_1739);
or U1568 (N_1568,In_227,In_684);
and U1569 (N_1569,In_529,In_377);
nand U1570 (N_1570,In_929,In_1939);
or U1571 (N_1571,In_1051,In_1770);
nor U1572 (N_1572,In_1580,In_339);
nor U1573 (N_1573,In_493,In_778);
nand U1574 (N_1574,In_880,In_869);
or U1575 (N_1575,In_1784,In_16);
or U1576 (N_1576,In_138,In_504);
nand U1577 (N_1577,In_465,In_812);
nand U1578 (N_1578,In_864,In_1109);
nand U1579 (N_1579,In_1654,In_1663);
and U1580 (N_1580,In_1635,In_26);
and U1581 (N_1581,In_1993,In_381);
xnor U1582 (N_1582,In_737,In_1327);
nor U1583 (N_1583,In_324,In_487);
nor U1584 (N_1584,In_897,In_433);
nand U1585 (N_1585,In_1726,In_246);
nor U1586 (N_1586,In_1900,In_874);
nand U1587 (N_1587,In_247,In_1607);
xor U1588 (N_1588,In_1981,In_1003);
nor U1589 (N_1589,In_47,In_1009);
nand U1590 (N_1590,In_1990,In_212);
nor U1591 (N_1591,In_729,In_355);
xnor U1592 (N_1592,In_1741,In_586);
nor U1593 (N_1593,In_1470,In_658);
xor U1594 (N_1594,In_218,In_739);
nand U1595 (N_1595,In_1346,In_431);
and U1596 (N_1596,In_57,In_79);
and U1597 (N_1597,In_1498,In_259);
nand U1598 (N_1598,In_37,In_1966);
and U1599 (N_1599,In_1062,In_679);
xnor U1600 (N_1600,In_1302,In_1378);
nand U1601 (N_1601,In_612,In_635);
and U1602 (N_1602,In_90,In_1641);
nor U1603 (N_1603,In_1081,In_690);
xnor U1604 (N_1604,In_1223,In_856);
xor U1605 (N_1605,In_612,In_1905);
and U1606 (N_1606,In_350,In_541);
nor U1607 (N_1607,In_1830,In_483);
or U1608 (N_1608,In_472,In_1641);
and U1609 (N_1609,In_1662,In_1999);
nor U1610 (N_1610,In_876,In_1115);
nand U1611 (N_1611,In_403,In_1367);
and U1612 (N_1612,In_624,In_1176);
and U1613 (N_1613,In_1018,In_80);
or U1614 (N_1614,In_1994,In_876);
nand U1615 (N_1615,In_264,In_1424);
and U1616 (N_1616,In_695,In_492);
nor U1617 (N_1617,In_923,In_687);
nand U1618 (N_1618,In_1916,In_112);
and U1619 (N_1619,In_154,In_227);
nor U1620 (N_1620,In_919,In_189);
or U1621 (N_1621,In_1923,In_989);
nor U1622 (N_1622,In_95,In_1574);
and U1623 (N_1623,In_346,In_1803);
xnor U1624 (N_1624,In_369,In_814);
nor U1625 (N_1625,In_1693,In_1444);
nor U1626 (N_1626,In_1302,In_1264);
xor U1627 (N_1627,In_1819,In_70);
and U1628 (N_1628,In_544,In_424);
nand U1629 (N_1629,In_329,In_849);
nor U1630 (N_1630,In_1881,In_221);
nand U1631 (N_1631,In_1550,In_698);
nor U1632 (N_1632,In_27,In_1491);
and U1633 (N_1633,In_49,In_399);
nor U1634 (N_1634,In_692,In_1103);
nor U1635 (N_1635,In_300,In_197);
nand U1636 (N_1636,In_166,In_497);
nand U1637 (N_1637,In_9,In_354);
and U1638 (N_1638,In_123,In_565);
nand U1639 (N_1639,In_468,In_204);
nand U1640 (N_1640,In_474,In_911);
xnor U1641 (N_1641,In_855,In_0);
nand U1642 (N_1642,In_1946,In_1607);
and U1643 (N_1643,In_1377,In_1272);
nor U1644 (N_1644,In_1078,In_1755);
or U1645 (N_1645,In_1375,In_498);
nor U1646 (N_1646,In_1471,In_736);
nor U1647 (N_1647,In_1378,In_1960);
nand U1648 (N_1648,In_83,In_795);
xor U1649 (N_1649,In_1287,In_675);
and U1650 (N_1650,In_209,In_902);
and U1651 (N_1651,In_597,In_1021);
nor U1652 (N_1652,In_1930,In_1470);
nand U1653 (N_1653,In_1062,In_1848);
and U1654 (N_1654,In_262,In_1117);
or U1655 (N_1655,In_885,In_750);
and U1656 (N_1656,In_1330,In_766);
or U1657 (N_1657,In_1759,In_1972);
and U1658 (N_1658,In_1584,In_1170);
or U1659 (N_1659,In_210,In_10);
and U1660 (N_1660,In_852,In_552);
nand U1661 (N_1661,In_1516,In_1344);
and U1662 (N_1662,In_1527,In_757);
nor U1663 (N_1663,In_1360,In_1506);
nor U1664 (N_1664,In_466,In_557);
xor U1665 (N_1665,In_809,In_530);
or U1666 (N_1666,In_1245,In_1841);
and U1667 (N_1667,In_1231,In_1433);
nor U1668 (N_1668,In_1825,In_555);
nand U1669 (N_1669,In_889,In_336);
or U1670 (N_1670,In_1784,In_1785);
and U1671 (N_1671,In_743,In_1227);
or U1672 (N_1672,In_85,In_1747);
and U1673 (N_1673,In_1823,In_1909);
nand U1674 (N_1674,In_649,In_599);
and U1675 (N_1675,In_1253,In_36);
and U1676 (N_1676,In_554,In_687);
or U1677 (N_1677,In_320,In_1250);
nor U1678 (N_1678,In_1855,In_1968);
nor U1679 (N_1679,In_1466,In_186);
or U1680 (N_1680,In_635,In_305);
and U1681 (N_1681,In_870,In_576);
nand U1682 (N_1682,In_905,In_68);
and U1683 (N_1683,In_1965,In_1874);
xnor U1684 (N_1684,In_1108,In_720);
nand U1685 (N_1685,In_1605,In_1364);
nor U1686 (N_1686,In_244,In_683);
and U1687 (N_1687,In_667,In_1169);
or U1688 (N_1688,In_507,In_170);
or U1689 (N_1689,In_359,In_1477);
nand U1690 (N_1690,In_1144,In_761);
and U1691 (N_1691,In_1564,In_592);
and U1692 (N_1692,In_1944,In_683);
or U1693 (N_1693,In_834,In_268);
or U1694 (N_1694,In_1271,In_619);
and U1695 (N_1695,In_1125,In_1425);
xor U1696 (N_1696,In_1430,In_1234);
or U1697 (N_1697,In_1179,In_623);
or U1698 (N_1698,In_928,In_184);
nand U1699 (N_1699,In_833,In_913);
or U1700 (N_1700,In_685,In_1972);
nor U1701 (N_1701,In_1863,In_469);
nand U1702 (N_1702,In_1997,In_1585);
and U1703 (N_1703,In_198,In_970);
or U1704 (N_1704,In_50,In_1259);
nand U1705 (N_1705,In_57,In_1746);
nand U1706 (N_1706,In_173,In_191);
nand U1707 (N_1707,In_1735,In_427);
or U1708 (N_1708,In_416,In_1821);
nor U1709 (N_1709,In_458,In_1998);
nor U1710 (N_1710,In_1999,In_1470);
or U1711 (N_1711,In_1969,In_1163);
and U1712 (N_1712,In_1830,In_215);
and U1713 (N_1713,In_446,In_1957);
nor U1714 (N_1714,In_665,In_462);
or U1715 (N_1715,In_1661,In_1493);
or U1716 (N_1716,In_721,In_1835);
nor U1717 (N_1717,In_622,In_1465);
or U1718 (N_1718,In_1728,In_1044);
xnor U1719 (N_1719,In_241,In_811);
nor U1720 (N_1720,In_181,In_1068);
and U1721 (N_1721,In_81,In_10);
xnor U1722 (N_1722,In_1165,In_1843);
nor U1723 (N_1723,In_1201,In_519);
xor U1724 (N_1724,In_55,In_35);
or U1725 (N_1725,In_1875,In_498);
nand U1726 (N_1726,In_1041,In_1906);
nand U1727 (N_1727,In_1055,In_1906);
xnor U1728 (N_1728,In_1602,In_1592);
nand U1729 (N_1729,In_286,In_1357);
or U1730 (N_1730,In_1571,In_688);
nand U1731 (N_1731,In_1918,In_1985);
xnor U1732 (N_1732,In_1654,In_471);
nor U1733 (N_1733,In_418,In_1583);
xor U1734 (N_1734,In_1341,In_1864);
and U1735 (N_1735,In_648,In_8);
xnor U1736 (N_1736,In_530,In_1221);
xor U1737 (N_1737,In_1487,In_254);
and U1738 (N_1738,In_748,In_959);
or U1739 (N_1739,In_133,In_1766);
or U1740 (N_1740,In_1147,In_1374);
or U1741 (N_1741,In_452,In_263);
and U1742 (N_1742,In_258,In_1333);
and U1743 (N_1743,In_476,In_1651);
nand U1744 (N_1744,In_396,In_817);
or U1745 (N_1745,In_671,In_655);
nand U1746 (N_1746,In_1694,In_1202);
nand U1747 (N_1747,In_709,In_63);
or U1748 (N_1748,In_674,In_977);
or U1749 (N_1749,In_209,In_1169);
or U1750 (N_1750,In_1755,In_1593);
nand U1751 (N_1751,In_1195,In_1774);
or U1752 (N_1752,In_223,In_484);
nor U1753 (N_1753,In_364,In_1577);
nand U1754 (N_1754,In_531,In_749);
or U1755 (N_1755,In_443,In_667);
nand U1756 (N_1756,In_575,In_249);
xnor U1757 (N_1757,In_571,In_143);
and U1758 (N_1758,In_826,In_728);
nor U1759 (N_1759,In_1154,In_177);
nand U1760 (N_1760,In_1617,In_150);
or U1761 (N_1761,In_170,In_1825);
and U1762 (N_1762,In_981,In_842);
or U1763 (N_1763,In_841,In_324);
and U1764 (N_1764,In_281,In_144);
nor U1765 (N_1765,In_792,In_1391);
and U1766 (N_1766,In_1681,In_1364);
and U1767 (N_1767,In_182,In_364);
or U1768 (N_1768,In_183,In_529);
and U1769 (N_1769,In_1689,In_1005);
nand U1770 (N_1770,In_1180,In_510);
nand U1771 (N_1771,In_1124,In_464);
nand U1772 (N_1772,In_1255,In_1736);
nor U1773 (N_1773,In_412,In_640);
and U1774 (N_1774,In_1892,In_289);
nand U1775 (N_1775,In_1957,In_263);
or U1776 (N_1776,In_1883,In_1784);
nor U1777 (N_1777,In_80,In_646);
or U1778 (N_1778,In_1966,In_1952);
and U1779 (N_1779,In_288,In_1693);
or U1780 (N_1780,In_1214,In_1170);
or U1781 (N_1781,In_1761,In_462);
and U1782 (N_1782,In_27,In_291);
and U1783 (N_1783,In_714,In_830);
and U1784 (N_1784,In_1916,In_753);
xnor U1785 (N_1785,In_1479,In_1070);
nand U1786 (N_1786,In_1223,In_1141);
or U1787 (N_1787,In_878,In_594);
nor U1788 (N_1788,In_1097,In_1034);
nor U1789 (N_1789,In_1103,In_1092);
nor U1790 (N_1790,In_1748,In_905);
or U1791 (N_1791,In_985,In_599);
nand U1792 (N_1792,In_1942,In_880);
or U1793 (N_1793,In_256,In_650);
and U1794 (N_1794,In_1133,In_1136);
nand U1795 (N_1795,In_936,In_1868);
nor U1796 (N_1796,In_1186,In_717);
or U1797 (N_1797,In_895,In_1069);
xor U1798 (N_1798,In_333,In_1603);
nand U1799 (N_1799,In_801,In_262);
nor U1800 (N_1800,In_142,In_925);
or U1801 (N_1801,In_86,In_1318);
or U1802 (N_1802,In_1251,In_241);
and U1803 (N_1803,In_1500,In_436);
and U1804 (N_1804,In_240,In_585);
or U1805 (N_1805,In_1874,In_1854);
or U1806 (N_1806,In_1021,In_1924);
nor U1807 (N_1807,In_227,In_297);
nand U1808 (N_1808,In_1104,In_786);
nand U1809 (N_1809,In_573,In_467);
and U1810 (N_1810,In_1212,In_283);
nor U1811 (N_1811,In_376,In_135);
and U1812 (N_1812,In_550,In_483);
xnor U1813 (N_1813,In_71,In_58);
nand U1814 (N_1814,In_121,In_1862);
nand U1815 (N_1815,In_107,In_1459);
xnor U1816 (N_1816,In_1529,In_254);
and U1817 (N_1817,In_1077,In_1319);
nor U1818 (N_1818,In_517,In_589);
nor U1819 (N_1819,In_834,In_156);
nand U1820 (N_1820,In_820,In_550);
nor U1821 (N_1821,In_1406,In_586);
or U1822 (N_1822,In_1801,In_309);
or U1823 (N_1823,In_1503,In_326);
nand U1824 (N_1824,In_1093,In_1873);
nand U1825 (N_1825,In_191,In_1524);
nor U1826 (N_1826,In_1623,In_1298);
and U1827 (N_1827,In_1537,In_626);
and U1828 (N_1828,In_928,In_900);
nand U1829 (N_1829,In_965,In_1616);
and U1830 (N_1830,In_736,In_594);
and U1831 (N_1831,In_864,In_1751);
nor U1832 (N_1832,In_1472,In_391);
and U1833 (N_1833,In_1602,In_1505);
nand U1834 (N_1834,In_825,In_522);
nand U1835 (N_1835,In_722,In_1402);
or U1836 (N_1836,In_1236,In_1876);
and U1837 (N_1837,In_413,In_189);
or U1838 (N_1838,In_1936,In_453);
nand U1839 (N_1839,In_869,In_1436);
nand U1840 (N_1840,In_104,In_114);
and U1841 (N_1841,In_1983,In_216);
and U1842 (N_1842,In_292,In_1212);
or U1843 (N_1843,In_1181,In_598);
nand U1844 (N_1844,In_1363,In_994);
or U1845 (N_1845,In_542,In_906);
nor U1846 (N_1846,In_1274,In_1389);
nor U1847 (N_1847,In_883,In_1279);
nor U1848 (N_1848,In_1792,In_1685);
or U1849 (N_1849,In_143,In_1097);
nand U1850 (N_1850,In_1991,In_385);
nand U1851 (N_1851,In_1095,In_1320);
nand U1852 (N_1852,In_1337,In_1884);
nand U1853 (N_1853,In_1146,In_1241);
or U1854 (N_1854,In_697,In_378);
and U1855 (N_1855,In_1768,In_1925);
or U1856 (N_1856,In_926,In_288);
nor U1857 (N_1857,In_1206,In_1729);
xnor U1858 (N_1858,In_183,In_15);
or U1859 (N_1859,In_971,In_130);
nand U1860 (N_1860,In_826,In_352);
nand U1861 (N_1861,In_1008,In_1415);
xnor U1862 (N_1862,In_1833,In_1266);
nor U1863 (N_1863,In_1719,In_41);
nand U1864 (N_1864,In_922,In_942);
and U1865 (N_1865,In_1914,In_440);
or U1866 (N_1866,In_1332,In_1834);
nand U1867 (N_1867,In_799,In_729);
or U1868 (N_1868,In_1833,In_1352);
nand U1869 (N_1869,In_887,In_191);
nor U1870 (N_1870,In_721,In_831);
nand U1871 (N_1871,In_134,In_1401);
or U1872 (N_1872,In_789,In_890);
nand U1873 (N_1873,In_1494,In_1416);
nand U1874 (N_1874,In_1555,In_1630);
and U1875 (N_1875,In_77,In_1095);
and U1876 (N_1876,In_214,In_849);
or U1877 (N_1877,In_1263,In_329);
nor U1878 (N_1878,In_824,In_1622);
and U1879 (N_1879,In_202,In_1589);
xnor U1880 (N_1880,In_791,In_1965);
nand U1881 (N_1881,In_1657,In_1223);
and U1882 (N_1882,In_1902,In_351);
or U1883 (N_1883,In_601,In_906);
nor U1884 (N_1884,In_1726,In_1228);
nand U1885 (N_1885,In_1414,In_821);
or U1886 (N_1886,In_758,In_13);
nand U1887 (N_1887,In_460,In_1223);
nor U1888 (N_1888,In_305,In_1622);
xor U1889 (N_1889,In_1277,In_1035);
xnor U1890 (N_1890,In_164,In_510);
nand U1891 (N_1891,In_748,In_1388);
or U1892 (N_1892,In_1513,In_1805);
or U1893 (N_1893,In_238,In_1802);
and U1894 (N_1894,In_11,In_106);
or U1895 (N_1895,In_832,In_21);
or U1896 (N_1896,In_1498,In_738);
xor U1897 (N_1897,In_444,In_957);
nand U1898 (N_1898,In_1150,In_447);
nor U1899 (N_1899,In_1464,In_337);
xor U1900 (N_1900,In_94,In_522);
nor U1901 (N_1901,In_1758,In_1468);
and U1902 (N_1902,In_1155,In_212);
nor U1903 (N_1903,In_1253,In_619);
nand U1904 (N_1904,In_572,In_735);
or U1905 (N_1905,In_1522,In_904);
nand U1906 (N_1906,In_863,In_952);
and U1907 (N_1907,In_1296,In_1852);
nand U1908 (N_1908,In_1434,In_1539);
and U1909 (N_1909,In_525,In_158);
and U1910 (N_1910,In_1451,In_1839);
and U1911 (N_1911,In_916,In_96);
nand U1912 (N_1912,In_1778,In_1301);
nand U1913 (N_1913,In_1461,In_793);
nand U1914 (N_1914,In_1974,In_1323);
or U1915 (N_1915,In_142,In_1615);
and U1916 (N_1916,In_998,In_968);
nand U1917 (N_1917,In_685,In_1955);
nand U1918 (N_1918,In_356,In_1027);
nor U1919 (N_1919,In_1394,In_417);
or U1920 (N_1920,In_526,In_1095);
or U1921 (N_1921,In_323,In_1224);
or U1922 (N_1922,In_1600,In_1311);
and U1923 (N_1923,In_1835,In_1563);
or U1924 (N_1924,In_556,In_1230);
and U1925 (N_1925,In_320,In_919);
and U1926 (N_1926,In_1738,In_921);
or U1927 (N_1927,In_1297,In_1758);
nand U1928 (N_1928,In_788,In_157);
or U1929 (N_1929,In_707,In_690);
nand U1930 (N_1930,In_613,In_929);
nand U1931 (N_1931,In_1303,In_146);
nor U1932 (N_1932,In_429,In_774);
nor U1933 (N_1933,In_156,In_669);
nor U1934 (N_1934,In_584,In_1267);
or U1935 (N_1935,In_296,In_1036);
and U1936 (N_1936,In_1295,In_1706);
nor U1937 (N_1937,In_23,In_199);
nor U1938 (N_1938,In_64,In_258);
xor U1939 (N_1939,In_565,In_1750);
and U1940 (N_1940,In_1972,In_1697);
nor U1941 (N_1941,In_1806,In_84);
and U1942 (N_1942,In_355,In_1846);
and U1943 (N_1943,In_1543,In_785);
xor U1944 (N_1944,In_82,In_179);
nor U1945 (N_1945,In_351,In_1139);
nor U1946 (N_1946,In_353,In_1379);
and U1947 (N_1947,In_1485,In_189);
or U1948 (N_1948,In_1298,In_1612);
or U1949 (N_1949,In_1558,In_1902);
or U1950 (N_1950,In_1306,In_1950);
nor U1951 (N_1951,In_390,In_1480);
nand U1952 (N_1952,In_1682,In_1170);
nor U1953 (N_1953,In_452,In_1739);
nor U1954 (N_1954,In_760,In_699);
nand U1955 (N_1955,In_953,In_1105);
nand U1956 (N_1956,In_1536,In_1725);
xor U1957 (N_1957,In_1115,In_1084);
nand U1958 (N_1958,In_1471,In_75);
xnor U1959 (N_1959,In_831,In_1395);
nand U1960 (N_1960,In_1490,In_1493);
nor U1961 (N_1961,In_1936,In_1246);
and U1962 (N_1962,In_1040,In_1809);
or U1963 (N_1963,In_1334,In_1665);
nor U1964 (N_1964,In_222,In_249);
and U1965 (N_1965,In_1427,In_1681);
nand U1966 (N_1966,In_498,In_232);
nor U1967 (N_1967,In_566,In_1391);
nand U1968 (N_1968,In_45,In_16);
nand U1969 (N_1969,In_1629,In_1112);
xor U1970 (N_1970,In_607,In_1638);
nor U1971 (N_1971,In_960,In_1867);
or U1972 (N_1972,In_1852,In_825);
or U1973 (N_1973,In_1488,In_405);
or U1974 (N_1974,In_1781,In_1783);
nor U1975 (N_1975,In_1425,In_767);
or U1976 (N_1976,In_1591,In_280);
nor U1977 (N_1977,In_1978,In_1361);
nand U1978 (N_1978,In_1436,In_1069);
xnor U1979 (N_1979,In_743,In_1961);
or U1980 (N_1980,In_1285,In_1700);
nand U1981 (N_1981,In_858,In_1821);
nor U1982 (N_1982,In_600,In_1957);
or U1983 (N_1983,In_940,In_852);
and U1984 (N_1984,In_1315,In_1358);
nand U1985 (N_1985,In_993,In_222);
nand U1986 (N_1986,In_502,In_1094);
and U1987 (N_1987,In_835,In_1693);
and U1988 (N_1988,In_419,In_495);
nor U1989 (N_1989,In_464,In_79);
or U1990 (N_1990,In_1807,In_169);
nor U1991 (N_1991,In_1554,In_1114);
and U1992 (N_1992,In_1913,In_189);
and U1993 (N_1993,In_301,In_442);
and U1994 (N_1994,In_1360,In_685);
nand U1995 (N_1995,In_913,In_1676);
or U1996 (N_1996,In_306,In_1748);
nor U1997 (N_1997,In_950,In_1630);
or U1998 (N_1998,In_1327,In_64);
or U1999 (N_1999,In_1824,In_1149);
xor U2000 (N_2000,In_423,In_780);
xor U2001 (N_2001,In_1296,In_653);
nand U2002 (N_2002,In_1185,In_816);
and U2003 (N_2003,In_784,In_1429);
nand U2004 (N_2004,In_295,In_1048);
nand U2005 (N_2005,In_185,In_1276);
nand U2006 (N_2006,In_1775,In_1642);
nand U2007 (N_2007,In_1031,In_235);
or U2008 (N_2008,In_907,In_1673);
nand U2009 (N_2009,In_844,In_1128);
nand U2010 (N_2010,In_935,In_652);
and U2011 (N_2011,In_1301,In_316);
and U2012 (N_2012,In_1863,In_1505);
or U2013 (N_2013,In_801,In_1884);
and U2014 (N_2014,In_943,In_492);
and U2015 (N_2015,In_1332,In_1523);
or U2016 (N_2016,In_1524,In_902);
nand U2017 (N_2017,In_1825,In_1793);
nor U2018 (N_2018,In_1283,In_1941);
nor U2019 (N_2019,In_423,In_315);
nor U2020 (N_2020,In_381,In_670);
or U2021 (N_2021,In_1918,In_1813);
nor U2022 (N_2022,In_1768,In_172);
nand U2023 (N_2023,In_1780,In_855);
nand U2024 (N_2024,In_1822,In_159);
nor U2025 (N_2025,In_1690,In_1774);
nor U2026 (N_2026,In_1593,In_564);
or U2027 (N_2027,In_333,In_1229);
or U2028 (N_2028,In_1065,In_1809);
nand U2029 (N_2029,In_538,In_147);
or U2030 (N_2030,In_1148,In_373);
and U2031 (N_2031,In_572,In_1602);
nand U2032 (N_2032,In_1152,In_900);
and U2033 (N_2033,In_1878,In_943);
xor U2034 (N_2034,In_139,In_516);
and U2035 (N_2035,In_759,In_649);
nor U2036 (N_2036,In_834,In_1366);
or U2037 (N_2037,In_302,In_104);
nor U2038 (N_2038,In_120,In_711);
or U2039 (N_2039,In_980,In_1346);
nand U2040 (N_2040,In_678,In_1064);
and U2041 (N_2041,In_1566,In_1945);
and U2042 (N_2042,In_1007,In_95);
nor U2043 (N_2043,In_52,In_887);
xor U2044 (N_2044,In_824,In_747);
and U2045 (N_2045,In_592,In_303);
nor U2046 (N_2046,In_655,In_1065);
xnor U2047 (N_2047,In_909,In_482);
and U2048 (N_2048,In_756,In_1723);
or U2049 (N_2049,In_1435,In_1625);
or U2050 (N_2050,In_74,In_209);
and U2051 (N_2051,In_1726,In_190);
nand U2052 (N_2052,In_544,In_922);
and U2053 (N_2053,In_824,In_18);
nand U2054 (N_2054,In_588,In_1697);
and U2055 (N_2055,In_419,In_1918);
xor U2056 (N_2056,In_360,In_1369);
and U2057 (N_2057,In_1631,In_1189);
nand U2058 (N_2058,In_1946,In_129);
nand U2059 (N_2059,In_1127,In_1795);
nand U2060 (N_2060,In_810,In_267);
nand U2061 (N_2061,In_1877,In_1606);
and U2062 (N_2062,In_72,In_1455);
xnor U2063 (N_2063,In_581,In_430);
nor U2064 (N_2064,In_114,In_503);
nor U2065 (N_2065,In_975,In_849);
nor U2066 (N_2066,In_1652,In_805);
and U2067 (N_2067,In_1163,In_1177);
xnor U2068 (N_2068,In_1945,In_1334);
or U2069 (N_2069,In_1831,In_1355);
and U2070 (N_2070,In_745,In_572);
xnor U2071 (N_2071,In_1631,In_305);
and U2072 (N_2072,In_1513,In_1691);
or U2073 (N_2073,In_1752,In_276);
nor U2074 (N_2074,In_1921,In_895);
or U2075 (N_2075,In_838,In_175);
and U2076 (N_2076,In_702,In_1915);
or U2077 (N_2077,In_63,In_1299);
nand U2078 (N_2078,In_1210,In_945);
or U2079 (N_2079,In_1078,In_575);
or U2080 (N_2080,In_1256,In_1275);
and U2081 (N_2081,In_1343,In_981);
and U2082 (N_2082,In_453,In_10);
nor U2083 (N_2083,In_10,In_1795);
or U2084 (N_2084,In_1389,In_313);
or U2085 (N_2085,In_1210,In_1671);
nand U2086 (N_2086,In_1981,In_1405);
and U2087 (N_2087,In_1428,In_1760);
nor U2088 (N_2088,In_1287,In_520);
and U2089 (N_2089,In_790,In_1163);
and U2090 (N_2090,In_513,In_278);
nor U2091 (N_2091,In_299,In_1297);
nor U2092 (N_2092,In_1110,In_845);
nor U2093 (N_2093,In_939,In_577);
and U2094 (N_2094,In_1371,In_452);
and U2095 (N_2095,In_617,In_244);
and U2096 (N_2096,In_1414,In_978);
or U2097 (N_2097,In_1972,In_937);
or U2098 (N_2098,In_1746,In_1333);
and U2099 (N_2099,In_803,In_333);
nand U2100 (N_2100,In_1464,In_1739);
or U2101 (N_2101,In_1067,In_48);
nor U2102 (N_2102,In_1510,In_483);
xnor U2103 (N_2103,In_472,In_1997);
nor U2104 (N_2104,In_1232,In_1503);
nand U2105 (N_2105,In_616,In_1199);
xor U2106 (N_2106,In_243,In_1986);
or U2107 (N_2107,In_1237,In_1453);
or U2108 (N_2108,In_1172,In_837);
or U2109 (N_2109,In_843,In_51);
xor U2110 (N_2110,In_1990,In_1202);
nand U2111 (N_2111,In_861,In_562);
nand U2112 (N_2112,In_954,In_809);
nor U2113 (N_2113,In_860,In_1123);
and U2114 (N_2114,In_1373,In_38);
and U2115 (N_2115,In_364,In_925);
or U2116 (N_2116,In_299,In_1811);
and U2117 (N_2117,In_1236,In_241);
and U2118 (N_2118,In_1242,In_1709);
and U2119 (N_2119,In_874,In_1374);
and U2120 (N_2120,In_758,In_1520);
or U2121 (N_2121,In_1641,In_1329);
and U2122 (N_2122,In_1102,In_732);
and U2123 (N_2123,In_1855,In_228);
nor U2124 (N_2124,In_346,In_625);
and U2125 (N_2125,In_285,In_1688);
xor U2126 (N_2126,In_1603,In_674);
and U2127 (N_2127,In_1620,In_97);
or U2128 (N_2128,In_1184,In_660);
or U2129 (N_2129,In_1694,In_1710);
or U2130 (N_2130,In_1913,In_738);
xnor U2131 (N_2131,In_69,In_324);
nand U2132 (N_2132,In_1770,In_346);
or U2133 (N_2133,In_1614,In_1495);
and U2134 (N_2134,In_606,In_1835);
nor U2135 (N_2135,In_1932,In_1957);
or U2136 (N_2136,In_99,In_411);
nand U2137 (N_2137,In_1003,In_772);
nand U2138 (N_2138,In_1186,In_801);
nor U2139 (N_2139,In_344,In_1829);
and U2140 (N_2140,In_551,In_1986);
nand U2141 (N_2141,In_139,In_1594);
and U2142 (N_2142,In_1852,In_989);
nor U2143 (N_2143,In_507,In_636);
nor U2144 (N_2144,In_1898,In_1119);
xor U2145 (N_2145,In_1659,In_932);
or U2146 (N_2146,In_322,In_1225);
nand U2147 (N_2147,In_836,In_1208);
or U2148 (N_2148,In_1021,In_1604);
nor U2149 (N_2149,In_1490,In_258);
and U2150 (N_2150,In_1440,In_759);
and U2151 (N_2151,In_851,In_1360);
nand U2152 (N_2152,In_617,In_1579);
nor U2153 (N_2153,In_1099,In_959);
or U2154 (N_2154,In_1615,In_276);
or U2155 (N_2155,In_375,In_836);
nor U2156 (N_2156,In_1130,In_801);
or U2157 (N_2157,In_1690,In_130);
or U2158 (N_2158,In_94,In_26);
nand U2159 (N_2159,In_571,In_519);
and U2160 (N_2160,In_1702,In_1287);
nor U2161 (N_2161,In_751,In_1388);
xnor U2162 (N_2162,In_286,In_801);
nor U2163 (N_2163,In_871,In_1547);
nor U2164 (N_2164,In_555,In_1184);
and U2165 (N_2165,In_662,In_599);
nor U2166 (N_2166,In_389,In_1950);
or U2167 (N_2167,In_684,In_397);
or U2168 (N_2168,In_773,In_1253);
nand U2169 (N_2169,In_1475,In_1778);
and U2170 (N_2170,In_1909,In_813);
and U2171 (N_2171,In_1930,In_5);
nand U2172 (N_2172,In_804,In_1200);
or U2173 (N_2173,In_1327,In_1448);
nor U2174 (N_2174,In_303,In_1788);
and U2175 (N_2175,In_1765,In_1807);
nand U2176 (N_2176,In_1304,In_1693);
nor U2177 (N_2177,In_364,In_1105);
nor U2178 (N_2178,In_262,In_1860);
xnor U2179 (N_2179,In_406,In_844);
xor U2180 (N_2180,In_1372,In_1358);
nand U2181 (N_2181,In_1473,In_32);
nor U2182 (N_2182,In_1992,In_817);
nand U2183 (N_2183,In_1914,In_991);
nor U2184 (N_2184,In_721,In_740);
nand U2185 (N_2185,In_1510,In_1995);
and U2186 (N_2186,In_836,In_1353);
or U2187 (N_2187,In_409,In_1174);
or U2188 (N_2188,In_1936,In_433);
nand U2189 (N_2189,In_733,In_249);
or U2190 (N_2190,In_1707,In_652);
and U2191 (N_2191,In_180,In_439);
xnor U2192 (N_2192,In_1012,In_420);
and U2193 (N_2193,In_372,In_1813);
and U2194 (N_2194,In_1026,In_1924);
nor U2195 (N_2195,In_1950,In_1237);
and U2196 (N_2196,In_1090,In_772);
xnor U2197 (N_2197,In_1615,In_1010);
or U2198 (N_2198,In_1263,In_891);
and U2199 (N_2199,In_694,In_1178);
and U2200 (N_2200,In_288,In_811);
nor U2201 (N_2201,In_1559,In_1460);
nand U2202 (N_2202,In_1208,In_1359);
or U2203 (N_2203,In_1262,In_1851);
and U2204 (N_2204,In_926,In_1814);
and U2205 (N_2205,In_1228,In_1982);
and U2206 (N_2206,In_971,In_1760);
and U2207 (N_2207,In_323,In_1492);
and U2208 (N_2208,In_71,In_1008);
nand U2209 (N_2209,In_142,In_39);
nor U2210 (N_2210,In_1649,In_1292);
xnor U2211 (N_2211,In_663,In_908);
nand U2212 (N_2212,In_1608,In_1803);
nand U2213 (N_2213,In_1324,In_932);
and U2214 (N_2214,In_652,In_1373);
and U2215 (N_2215,In_1784,In_1155);
or U2216 (N_2216,In_1973,In_146);
and U2217 (N_2217,In_1134,In_1770);
nor U2218 (N_2218,In_1980,In_1348);
and U2219 (N_2219,In_734,In_1034);
and U2220 (N_2220,In_1485,In_1352);
nand U2221 (N_2221,In_646,In_327);
nand U2222 (N_2222,In_1325,In_33);
nor U2223 (N_2223,In_421,In_18);
nand U2224 (N_2224,In_818,In_1826);
nand U2225 (N_2225,In_1303,In_1625);
or U2226 (N_2226,In_973,In_1837);
or U2227 (N_2227,In_1741,In_1179);
or U2228 (N_2228,In_960,In_800);
or U2229 (N_2229,In_1122,In_237);
and U2230 (N_2230,In_1265,In_568);
nor U2231 (N_2231,In_1902,In_1145);
and U2232 (N_2232,In_1984,In_401);
or U2233 (N_2233,In_906,In_1832);
or U2234 (N_2234,In_474,In_316);
nand U2235 (N_2235,In_1530,In_633);
nor U2236 (N_2236,In_268,In_0);
or U2237 (N_2237,In_917,In_561);
nor U2238 (N_2238,In_1358,In_1319);
nand U2239 (N_2239,In_382,In_832);
xnor U2240 (N_2240,In_1161,In_834);
xnor U2241 (N_2241,In_11,In_1583);
nand U2242 (N_2242,In_310,In_1266);
or U2243 (N_2243,In_504,In_913);
nand U2244 (N_2244,In_341,In_1865);
nor U2245 (N_2245,In_1836,In_610);
nor U2246 (N_2246,In_425,In_745);
nand U2247 (N_2247,In_1355,In_1821);
nor U2248 (N_2248,In_360,In_1747);
and U2249 (N_2249,In_1623,In_851);
nor U2250 (N_2250,In_1064,In_1437);
nand U2251 (N_2251,In_1878,In_1744);
nand U2252 (N_2252,In_1727,In_1005);
or U2253 (N_2253,In_1458,In_465);
or U2254 (N_2254,In_257,In_603);
xnor U2255 (N_2255,In_1812,In_168);
nor U2256 (N_2256,In_27,In_83);
nor U2257 (N_2257,In_1718,In_833);
or U2258 (N_2258,In_14,In_247);
xor U2259 (N_2259,In_480,In_664);
or U2260 (N_2260,In_819,In_751);
or U2261 (N_2261,In_639,In_1352);
nand U2262 (N_2262,In_86,In_821);
or U2263 (N_2263,In_1953,In_536);
and U2264 (N_2264,In_905,In_1951);
nand U2265 (N_2265,In_428,In_1422);
nor U2266 (N_2266,In_1500,In_1594);
or U2267 (N_2267,In_167,In_1085);
nor U2268 (N_2268,In_1299,In_528);
or U2269 (N_2269,In_1475,In_1502);
xor U2270 (N_2270,In_917,In_110);
nor U2271 (N_2271,In_666,In_1131);
nand U2272 (N_2272,In_1614,In_893);
nand U2273 (N_2273,In_1751,In_981);
or U2274 (N_2274,In_1841,In_798);
nand U2275 (N_2275,In_1039,In_1287);
nor U2276 (N_2276,In_130,In_295);
or U2277 (N_2277,In_567,In_1957);
and U2278 (N_2278,In_499,In_1248);
xnor U2279 (N_2279,In_971,In_179);
or U2280 (N_2280,In_5,In_268);
or U2281 (N_2281,In_1891,In_1776);
or U2282 (N_2282,In_708,In_847);
nor U2283 (N_2283,In_363,In_711);
and U2284 (N_2284,In_830,In_136);
nand U2285 (N_2285,In_1542,In_1552);
nor U2286 (N_2286,In_1889,In_422);
nor U2287 (N_2287,In_44,In_748);
and U2288 (N_2288,In_35,In_1484);
xor U2289 (N_2289,In_1368,In_1818);
xor U2290 (N_2290,In_1080,In_476);
and U2291 (N_2291,In_1417,In_900);
nand U2292 (N_2292,In_1259,In_122);
or U2293 (N_2293,In_1449,In_1363);
or U2294 (N_2294,In_595,In_1051);
or U2295 (N_2295,In_1575,In_435);
nand U2296 (N_2296,In_1817,In_1248);
nor U2297 (N_2297,In_261,In_1505);
xor U2298 (N_2298,In_664,In_225);
or U2299 (N_2299,In_1740,In_1627);
nand U2300 (N_2300,In_389,In_1282);
nor U2301 (N_2301,In_1790,In_1337);
and U2302 (N_2302,In_958,In_483);
nand U2303 (N_2303,In_519,In_1379);
and U2304 (N_2304,In_1881,In_521);
nand U2305 (N_2305,In_1809,In_505);
nand U2306 (N_2306,In_507,In_141);
nor U2307 (N_2307,In_1074,In_709);
xor U2308 (N_2308,In_207,In_452);
and U2309 (N_2309,In_1568,In_521);
nand U2310 (N_2310,In_1866,In_169);
or U2311 (N_2311,In_1199,In_327);
or U2312 (N_2312,In_1053,In_981);
and U2313 (N_2313,In_1184,In_1922);
and U2314 (N_2314,In_1312,In_22);
xnor U2315 (N_2315,In_1060,In_1588);
or U2316 (N_2316,In_629,In_1021);
or U2317 (N_2317,In_246,In_344);
and U2318 (N_2318,In_1924,In_260);
and U2319 (N_2319,In_955,In_1642);
or U2320 (N_2320,In_1109,In_1620);
nand U2321 (N_2321,In_123,In_1827);
or U2322 (N_2322,In_761,In_596);
or U2323 (N_2323,In_1129,In_1463);
xnor U2324 (N_2324,In_1609,In_299);
nor U2325 (N_2325,In_1042,In_1169);
xnor U2326 (N_2326,In_1188,In_613);
and U2327 (N_2327,In_1005,In_695);
xnor U2328 (N_2328,In_1714,In_1176);
nand U2329 (N_2329,In_1617,In_1468);
or U2330 (N_2330,In_323,In_1795);
xnor U2331 (N_2331,In_1936,In_1342);
nor U2332 (N_2332,In_219,In_781);
nor U2333 (N_2333,In_760,In_1166);
and U2334 (N_2334,In_1459,In_980);
or U2335 (N_2335,In_1928,In_566);
or U2336 (N_2336,In_1346,In_1954);
and U2337 (N_2337,In_1741,In_871);
xor U2338 (N_2338,In_1580,In_1829);
and U2339 (N_2339,In_401,In_1858);
or U2340 (N_2340,In_1025,In_1301);
or U2341 (N_2341,In_454,In_1596);
or U2342 (N_2342,In_929,In_665);
and U2343 (N_2343,In_1446,In_344);
nor U2344 (N_2344,In_1218,In_1466);
xor U2345 (N_2345,In_427,In_523);
nand U2346 (N_2346,In_52,In_756);
nor U2347 (N_2347,In_1157,In_1015);
and U2348 (N_2348,In_603,In_1449);
nand U2349 (N_2349,In_879,In_423);
nand U2350 (N_2350,In_1335,In_855);
nor U2351 (N_2351,In_890,In_1685);
or U2352 (N_2352,In_451,In_1275);
or U2353 (N_2353,In_1144,In_1046);
or U2354 (N_2354,In_166,In_1734);
nand U2355 (N_2355,In_1236,In_1058);
or U2356 (N_2356,In_518,In_1870);
xnor U2357 (N_2357,In_1459,In_669);
nand U2358 (N_2358,In_1724,In_1911);
or U2359 (N_2359,In_505,In_1925);
nor U2360 (N_2360,In_630,In_220);
or U2361 (N_2361,In_1602,In_1661);
nand U2362 (N_2362,In_859,In_867);
and U2363 (N_2363,In_637,In_306);
xor U2364 (N_2364,In_1396,In_815);
xor U2365 (N_2365,In_940,In_751);
and U2366 (N_2366,In_1724,In_715);
or U2367 (N_2367,In_1489,In_1636);
nand U2368 (N_2368,In_919,In_1127);
or U2369 (N_2369,In_1577,In_251);
nor U2370 (N_2370,In_955,In_1079);
or U2371 (N_2371,In_898,In_1235);
and U2372 (N_2372,In_763,In_1412);
and U2373 (N_2373,In_1101,In_1536);
or U2374 (N_2374,In_1856,In_379);
nand U2375 (N_2375,In_343,In_1323);
nand U2376 (N_2376,In_1446,In_1636);
or U2377 (N_2377,In_1163,In_306);
nor U2378 (N_2378,In_51,In_1652);
nand U2379 (N_2379,In_1629,In_1276);
and U2380 (N_2380,In_1249,In_1023);
and U2381 (N_2381,In_945,In_461);
or U2382 (N_2382,In_1901,In_1167);
or U2383 (N_2383,In_1156,In_1827);
nor U2384 (N_2384,In_707,In_46);
nor U2385 (N_2385,In_834,In_1910);
or U2386 (N_2386,In_297,In_1196);
xor U2387 (N_2387,In_259,In_1493);
nor U2388 (N_2388,In_1237,In_114);
nor U2389 (N_2389,In_95,In_1297);
and U2390 (N_2390,In_1752,In_77);
nand U2391 (N_2391,In_1251,In_923);
nor U2392 (N_2392,In_714,In_980);
nand U2393 (N_2393,In_1611,In_1450);
and U2394 (N_2394,In_810,In_689);
nand U2395 (N_2395,In_761,In_399);
nor U2396 (N_2396,In_931,In_208);
and U2397 (N_2397,In_1850,In_241);
xor U2398 (N_2398,In_163,In_851);
or U2399 (N_2399,In_1821,In_1061);
nand U2400 (N_2400,In_1269,In_1030);
or U2401 (N_2401,In_1418,In_1469);
and U2402 (N_2402,In_1483,In_401);
xor U2403 (N_2403,In_133,In_1286);
nand U2404 (N_2404,In_515,In_421);
and U2405 (N_2405,In_866,In_1178);
and U2406 (N_2406,In_1536,In_1909);
and U2407 (N_2407,In_1823,In_1194);
nand U2408 (N_2408,In_689,In_170);
nand U2409 (N_2409,In_805,In_1540);
nor U2410 (N_2410,In_1206,In_291);
or U2411 (N_2411,In_634,In_1693);
nor U2412 (N_2412,In_1669,In_1604);
nor U2413 (N_2413,In_385,In_1702);
nand U2414 (N_2414,In_1045,In_1054);
nor U2415 (N_2415,In_749,In_1735);
nand U2416 (N_2416,In_1888,In_929);
nand U2417 (N_2417,In_1244,In_503);
or U2418 (N_2418,In_1542,In_1776);
xnor U2419 (N_2419,In_131,In_1169);
or U2420 (N_2420,In_390,In_938);
nand U2421 (N_2421,In_121,In_1441);
or U2422 (N_2422,In_782,In_1433);
and U2423 (N_2423,In_663,In_78);
nor U2424 (N_2424,In_440,In_489);
and U2425 (N_2425,In_1455,In_500);
nand U2426 (N_2426,In_1803,In_1577);
or U2427 (N_2427,In_1444,In_959);
nand U2428 (N_2428,In_1982,In_584);
nor U2429 (N_2429,In_1061,In_1263);
and U2430 (N_2430,In_1833,In_1312);
or U2431 (N_2431,In_506,In_219);
nor U2432 (N_2432,In_283,In_640);
or U2433 (N_2433,In_436,In_473);
or U2434 (N_2434,In_743,In_1004);
and U2435 (N_2435,In_248,In_1282);
xor U2436 (N_2436,In_1261,In_102);
nor U2437 (N_2437,In_904,In_378);
and U2438 (N_2438,In_1935,In_727);
or U2439 (N_2439,In_143,In_489);
nand U2440 (N_2440,In_307,In_153);
and U2441 (N_2441,In_1684,In_1402);
nor U2442 (N_2442,In_510,In_1731);
nand U2443 (N_2443,In_791,In_239);
or U2444 (N_2444,In_1672,In_1342);
and U2445 (N_2445,In_149,In_1186);
nor U2446 (N_2446,In_692,In_26);
nor U2447 (N_2447,In_475,In_1396);
and U2448 (N_2448,In_1701,In_894);
nand U2449 (N_2449,In_448,In_1838);
and U2450 (N_2450,In_1026,In_1662);
and U2451 (N_2451,In_1689,In_250);
and U2452 (N_2452,In_1319,In_1569);
and U2453 (N_2453,In_1392,In_864);
or U2454 (N_2454,In_784,In_468);
nand U2455 (N_2455,In_390,In_702);
nand U2456 (N_2456,In_1275,In_1779);
nand U2457 (N_2457,In_1521,In_1540);
nand U2458 (N_2458,In_152,In_1777);
or U2459 (N_2459,In_667,In_1932);
and U2460 (N_2460,In_820,In_300);
nor U2461 (N_2461,In_674,In_478);
and U2462 (N_2462,In_278,In_1376);
nor U2463 (N_2463,In_275,In_902);
nand U2464 (N_2464,In_672,In_633);
nor U2465 (N_2465,In_1821,In_1594);
and U2466 (N_2466,In_1466,In_1777);
or U2467 (N_2467,In_996,In_689);
and U2468 (N_2468,In_758,In_702);
nor U2469 (N_2469,In_217,In_1637);
or U2470 (N_2470,In_1076,In_1248);
nand U2471 (N_2471,In_1873,In_1052);
or U2472 (N_2472,In_1951,In_460);
nand U2473 (N_2473,In_1405,In_657);
or U2474 (N_2474,In_559,In_1403);
nor U2475 (N_2475,In_1322,In_1012);
nand U2476 (N_2476,In_758,In_93);
nand U2477 (N_2477,In_1629,In_360);
and U2478 (N_2478,In_839,In_289);
and U2479 (N_2479,In_704,In_336);
and U2480 (N_2480,In_1642,In_1008);
or U2481 (N_2481,In_1534,In_758);
nand U2482 (N_2482,In_1891,In_1690);
nand U2483 (N_2483,In_111,In_1568);
nand U2484 (N_2484,In_99,In_1419);
or U2485 (N_2485,In_1359,In_266);
nor U2486 (N_2486,In_1783,In_355);
xnor U2487 (N_2487,In_969,In_333);
nor U2488 (N_2488,In_762,In_1516);
nor U2489 (N_2489,In_1532,In_837);
and U2490 (N_2490,In_369,In_803);
nor U2491 (N_2491,In_1735,In_1945);
or U2492 (N_2492,In_73,In_647);
nor U2493 (N_2493,In_794,In_399);
or U2494 (N_2494,In_363,In_1299);
nand U2495 (N_2495,In_1996,In_1112);
or U2496 (N_2496,In_260,In_1140);
nand U2497 (N_2497,In_163,In_1476);
and U2498 (N_2498,In_628,In_1382);
and U2499 (N_2499,In_1712,In_1021);
or U2500 (N_2500,In_1026,In_116);
or U2501 (N_2501,In_409,In_1770);
and U2502 (N_2502,In_454,In_92);
nand U2503 (N_2503,In_130,In_1069);
nand U2504 (N_2504,In_1628,In_1895);
nand U2505 (N_2505,In_540,In_557);
nand U2506 (N_2506,In_271,In_740);
nor U2507 (N_2507,In_497,In_706);
nand U2508 (N_2508,In_1384,In_315);
or U2509 (N_2509,In_1863,In_516);
nor U2510 (N_2510,In_988,In_952);
nand U2511 (N_2511,In_620,In_43);
and U2512 (N_2512,In_319,In_803);
nor U2513 (N_2513,In_1298,In_1376);
nor U2514 (N_2514,In_693,In_177);
or U2515 (N_2515,In_735,In_1490);
and U2516 (N_2516,In_1339,In_866);
nor U2517 (N_2517,In_1948,In_1966);
nand U2518 (N_2518,In_645,In_816);
nand U2519 (N_2519,In_321,In_1238);
nand U2520 (N_2520,In_1493,In_73);
nand U2521 (N_2521,In_304,In_638);
xor U2522 (N_2522,In_515,In_655);
xnor U2523 (N_2523,In_700,In_941);
and U2524 (N_2524,In_1072,In_1082);
nand U2525 (N_2525,In_1613,In_1981);
or U2526 (N_2526,In_1255,In_1414);
xor U2527 (N_2527,In_189,In_1481);
xnor U2528 (N_2528,In_940,In_272);
or U2529 (N_2529,In_1987,In_148);
or U2530 (N_2530,In_1776,In_1880);
and U2531 (N_2531,In_1074,In_1647);
nand U2532 (N_2532,In_509,In_1276);
nor U2533 (N_2533,In_1618,In_353);
nor U2534 (N_2534,In_230,In_1517);
and U2535 (N_2535,In_835,In_1193);
and U2536 (N_2536,In_1968,In_88);
and U2537 (N_2537,In_57,In_1707);
or U2538 (N_2538,In_1034,In_59);
and U2539 (N_2539,In_1791,In_1818);
nor U2540 (N_2540,In_1314,In_1392);
or U2541 (N_2541,In_1198,In_755);
nor U2542 (N_2542,In_810,In_1183);
nand U2543 (N_2543,In_756,In_888);
nor U2544 (N_2544,In_1451,In_918);
nor U2545 (N_2545,In_412,In_1190);
and U2546 (N_2546,In_802,In_209);
or U2547 (N_2547,In_85,In_961);
and U2548 (N_2548,In_1236,In_984);
xnor U2549 (N_2549,In_1438,In_1978);
nor U2550 (N_2550,In_1236,In_1122);
nor U2551 (N_2551,In_149,In_1150);
nand U2552 (N_2552,In_600,In_675);
and U2553 (N_2553,In_412,In_917);
or U2554 (N_2554,In_954,In_196);
nor U2555 (N_2555,In_887,In_1476);
and U2556 (N_2556,In_1428,In_314);
or U2557 (N_2557,In_6,In_675);
and U2558 (N_2558,In_1520,In_888);
nor U2559 (N_2559,In_1985,In_709);
or U2560 (N_2560,In_315,In_1655);
nor U2561 (N_2561,In_166,In_853);
or U2562 (N_2562,In_802,In_452);
or U2563 (N_2563,In_1175,In_1798);
nor U2564 (N_2564,In_732,In_844);
or U2565 (N_2565,In_1144,In_1179);
nor U2566 (N_2566,In_1529,In_142);
nor U2567 (N_2567,In_1400,In_1720);
nand U2568 (N_2568,In_1146,In_581);
nand U2569 (N_2569,In_1118,In_940);
nor U2570 (N_2570,In_815,In_881);
nand U2571 (N_2571,In_382,In_1848);
or U2572 (N_2572,In_1941,In_870);
or U2573 (N_2573,In_194,In_988);
or U2574 (N_2574,In_1067,In_447);
or U2575 (N_2575,In_1491,In_532);
nand U2576 (N_2576,In_1813,In_1517);
nand U2577 (N_2577,In_510,In_1453);
or U2578 (N_2578,In_703,In_246);
nor U2579 (N_2579,In_569,In_882);
nor U2580 (N_2580,In_861,In_966);
xnor U2581 (N_2581,In_1245,In_1256);
nand U2582 (N_2582,In_1965,In_397);
nand U2583 (N_2583,In_859,In_1441);
and U2584 (N_2584,In_1220,In_1314);
nand U2585 (N_2585,In_548,In_1688);
and U2586 (N_2586,In_816,In_1012);
or U2587 (N_2587,In_684,In_1161);
xnor U2588 (N_2588,In_782,In_1864);
nand U2589 (N_2589,In_1546,In_1834);
nand U2590 (N_2590,In_350,In_1547);
and U2591 (N_2591,In_1056,In_1778);
xnor U2592 (N_2592,In_1984,In_305);
nand U2593 (N_2593,In_218,In_1670);
nand U2594 (N_2594,In_1894,In_1778);
nor U2595 (N_2595,In_1114,In_1261);
nor U2596 (N_2596,In_532,In_187);
and U2597 (N_2597,In_1195,In_45);
nand U2598 (N_2598,In_1535,In_1219);
or U2599 (N_2599,In_37,In_571);
and U2600 (N_2600,In_74,In_137);
and U2601 (N_2601,In_1597,In_78);
and U2602 (N_2602,In_733,In_1248);
and U2603 (N_2603,In_802,In_1144);
xor U2604 (N_2604,In_1848,In_1323);
nand U2605 (N_2605,In_955,In_984);
xor U2606 (N_2606,In_817,In_1281);
nor U2607 (N_2607,In_1649,In_1440);
or U2608 (N_2608,In_100,In_218);
and U2609 (N_2609,In_370,In_1677);
nor U2610 (N_2610,In_570,In_258);
and U2611 (N_2611,In_435,In_1102);
and U2612 (N_2612,In_1855,In_1223);
nand U2613 (N_2613,In_1787,In_1903);
and U2614 (N_2614,In_215,In_536);
nor U2615 (N_2615,In_309,In_1292);
xor U2616 (N_2616,In_22,In_1923);
nand U2617 (N_2617,In_764,In_1708);
and U2618 (N_2618,In_1711,In_1360);
nor U2619 (N_2619,In_512,In_473);
and U2620 (N_2620,In_1573,In_1646);
or U2621 (N_2621,In_1420,In_596);
or U2622 (N_2622,In_738,In_869);
nand U2623 (N_2623,In_1746,In_895);
and U2624 (N_2624,In_1325,In_1127);
nand U2625 (N_2625,In_281,In_1552);
or U2626 (N_2626,In_1503,In_1266);
nand U2627 (N_2627,In_1314,In_909);
or U2628 (N_2628,In_215,In_1070);
and U2629 (N_2629,In_1356,In_381);
or U2630 (N_2630,In_1400,In_110);
and U2631 (N_2631,In_1271,In_1112);
or U2632 (N_2632,In_588,In_630);
nor U2633 (N_2633,In_1216,In_153);
nor U2634 (N_2634,In_1426,In_869);
nor U2635 (N_2635,In_591,In_846);
and U2636 (N_2636,In_355,In_170);
nand U2637 (N_2637,In_1095,In_1674);
and U2638 (N_2638,In_948,In_231);
xnor U2639 (N_2639,In_1206,In_289);
or U2640 (N_2640,In_1497,In_669);
nor U2641 (N_2641,In_1730,In_163);
or U2642 (N_2642,In_157,In_1339);
nor U2643 (N_2643,In_754,In_307);
nor U2644 (N_2644,In_1813,In_1416);
or U2645 (N_2645,In_851,In_1302);
xor U2646 (N_2646,In_1375,In_339);
nor U2647 (N_2647,In_848,In_799);
nor U2648 (N_2648,In_1725,In_292);
nor U2649 (N_2649,In_349,In_1139);
nor U2650 (N_2650,In_1559,In_60);
nand U2651 (N_2651,In_747,In_1712);
nor U2652 (N_2652,In_477,In_436);
nor U2653 (N_2653,In_212,In_951);
nor U2654 (N_2654,In_1819,In_630);
or U2655 (N_2655,In_866,In_1972);
nand U2656 (N_2656,In_959,In_1067);
and U2657 (N_2657,In_1407,In_698);
nand U2658 (N_2658,In_843,In_1039);
and U2659 (N_2659,In_337,In_1715);
and U2660 (N_2660,In_508,In_1202);
nand U2661 (N_2661,In_1683,In_284);
and U2662 (N_2662,In_792,In_1167);
nor U2663 (N_2663,In_1984,In_691);
nand U2664 (N_2664,In_1032,In_252);
nand U2665 (N_2665,In_1682,In_45);
nor U2666 (N_2666,In_642,In_1420);
nand U2667 (N_2667,In_1990,In_1823);
and U2668 (N_2668,In_289,In_1560);
nor U2669 (N_2669,In_723,In_1796);
nand U2670 (N_2670,In_1224,In_1718);
or U2671 (N_2671,In_803,In_1213);
nand U2672 (N_2672,In_484,In_181);
xor U2673 (N_2673,In_662,In_1951);
nand U2674 (N_2674,In_699,In_139);
nor U2675 (N_2675,In_683,In_429);
nand U2676 (N_2676,In_654,In_1828);
or U2677 (N_2677,In_1968,In_51);
nor U2678 (N_2678,In_49,In_78);
and U2679 (N_2679,In_1605,In_1487);
xnor U2680 (N_2680,In_287,In_1913);
or U2681 (N_2681,In_509,In_1824);
nor U2682 (N_2682,In_962,In_1880);
and U2683 (N_2683,In_1986,In_1004);
xor U2684 (N_2684,In_891,In_395);
and U2685 (N_2685,In_1187,In_1224);
nor U2686 (N_2686,In_1047,In_1066);
and U2687 (N_2687,In_908,In_119);
nor U2688 (N_2688,In_835,In_785);
or U2689 (N_2689,In_801,In_859);
or U2690 (N_2690,In_606,In_1840);
nor U2691 (N_2691,In_533,In_1387);
nor U2692 (N_2692,In_130,In_611);
or U2693 (N_2693,In_1123,In_1501);
nand U2694 (N_2694,In_1126,In_891);
or U2695 (N_2695,In_343,In_594);
or U2696 (N_2696,In_1532,In_449);
or U2697 (N_2697,In_1127,In_1400);
nor U2698 (N_2698,In_701,In_538);
or U2699 (N_2699,In_236,In_627);
nand U2700 (N_2700,In_224,In_234);
nand U2701 (N_2701,In_784,In_101);
or U2702 (N_2702,In_507,In_318);
or U2703 (N_2703,In_1541,In_333);
nor U2704 (N_2704,In_292,In_985);
nor U2705 (N_2705,In_1186,In_1021);
nand U2706 (N_2706,In_1302,In_1119);
or U2707 (N_2707,In_1786,In_596);
or U2708 (N_2708,In_1734,In_660);
nand U2709 (N_2709,In_1882,In_514);
nand U2710 (N_2710,In_1541,In_1550);
and U2711 (N_2711,In_253,In_821);
and U2712 (N_2712,In_246,In_575);
nand U2713 (N_2713,In_137,In_1592);
nor U2714 (N_2714,In_1299,In_1564);
nand U2715 (N_2715,In_297,In_1243);
or U2716 (N_2716,In_604,In_189);
and U2717 (N_2717,In_187,In_1038);
and U2718 (N_2718,In_756,In_1710);
or U2719 (N_2719,In_1541,In_38);
or U2720 (N_2720,In_627,In_240);
or U2721 (N_2721,In_1462,In_615);
or U2722 (N_2722,In_143,In_1520);
or U2723 (N_2723,In_588,In_1098);
or U2724 (N_2724,In_1533,In_367);
or U2725 (N_2725,In_1525,In_503);
nor U2726 (N_2726,In_1540,In_1539);
nor U2727 (N_2727,In_921,In_1121);
nor U2728 (N_2728,In_272,In_544);
and U2729 (N_2729,In_558,In_1463);
or U2730 (N_2730,In_362,In_940);
or U2731 (N_2731,In_124,In_1087);
nand U2732 (N_2732,In_1898,In_1938);
xor U2733 (N_2733,In_1389,In_1154);
nand U2734 (N_2734,In_1124,In_1661);
and U2735 (N_2735,In_1438,In_70);
nor U2736 (N_2736,In_1697,In_1195);
nand U2737 (N_2737,In_1916,In_270);
nor U2738 (N_2738,In_1043,In_1590);
or U2739 (N_2739,In_1867,In_1899);
and U2740 (N_2740,In_215,In_809);
xor U2741 (N_2741,In_1851,In_1161);
nand U2742 (N_2742,In_798,In_1456);
and U2743 (N_2743,In_777,In_1235);
nor U2744 (N_2744,In_336,In_842);
and U2745 (N_2745,In_15,In_812);
and U2746 (N_2746,In_220,In_1312);
nor U2747 (N_2747,In_1136,In_775);
or U2748 (N_2748,In_746,In_1992);
nor U2749 (N_2749,In_1171,In_47);
and U2750 (N_2750,In_1013,In_466);
nand U2751 (N_2751,In_1478,In_1172);
and U2752 (N_2752,In_56,In_1068);
nand U2753 (N_2753,In_1046,In_74);
or U2754 (N_2754,In_589,In_1484);
and U2755 (N_2755,In_1935,In_1861);
nor U2756 (N_2756,In_670,In_244);
and U2757 (N_2757,In_1877,In_1497);
and U2758 (N_2758,In_91,In_212);
nand U2759 (N_2759,In_1534,In_239);
nor U2760 (N_2760,In_43,In_655);
or U2761 (N_2761,In_405,In_404);
and U2762 (N_2762,In_1161,In_1158);
nand U2763 (N_2763,In_461,In_443);
nand U2764 (N_2764,In_61,In_1092);
nor U2765 (N_2765,In_1971,In_1563);
nor U2766 (N_2766,In_520,In_405);
nor U2767 (N_2767,In_1664,In_63);
and U2768 (N_2768,In_409,In_34);
and U2769 (N_2769,In_1904,In_1765);
xnor U2770 (N_2770,In_106,In_1574);
or U2771 (N_2771,In_1930,In_993);
xnor U2772 (N_2772,In_1554,In_48);
and U2773 (N_2773,In_1037,In_442);
nand U2774 (N_2774,In_1481,In_732);
and U2775 (N_2775,In_672,In_4);
or U2776 (N_2776,In_1588,In_1434);
nand U2777 (N_2777,In_717,In_934);
nor U2778 (N_2778,In_1446,In_924);
nand U2779 (N_2779,In_255,In_1796);
or U2780 (N_2780,In_391,In_1343);
and U2781 (N_2781,In_1279,In_1771);
or U2782 (N_2782,In_1374,In_181);
and U2783 (N_2783,In_1279,In_767);
nor U2784 (N_2784,In_1732,In_1675);
nand U2785 (N_2785,In_188,In_744);
nor U2786 (N_2786,In_1190,In_278);
or U2787 (N_2787,In_378,In_1676);
or U2788 (N_2788,In_1355,In_1256);
xnor U2789 (N_2789,In_807,In_1468);
nor U2790 (N_2790,In_52,In_251);
xor U2791 (N_2791,In_851,In_1882);
nor U2792 (N_2792,In_232,In_875);
and U2793 (N_2793,In_117,In_1689);
nor U2794 (N_2794,In_1084,In_440);
nor U2795 (N_2795,In_852,In_1517);
or U2796 (N_2796,In_775,In_1838);
and U2797 (N_2797,In_967,In_197);
xnor U2798 (N_2798,In_84,In_80);
nand U2799 (N_2799,In_427,In_261);
nand U2800 (N_2800,In_274,In_1019);
nor U2801 (N_2801,In_565,In_999);
or U2802 (N_2802,In_671,In_1455);
nand U2803 (N_2803,In_384,In_1332);
nor U2804 (N_2804,In_179,In_519);
nor U2805 (N_2805,In_1759,In_348);
xnor U2806 (N_2806,In_1860,In_428);
or U2807 (N_2807,In_877,In_280);
xor U2808 (N_2808,In_654,In_1670);
or U2809 (N_2809,In_1049,In_802);
nand U2810 (N_2810,In_1879,In_1428);
nand U2811 (N_2811,In_1097,In_1390);
nand U2812 (N_2812,In_1724,In_1926);
and U2813 (N_2813,In_1893,In_1197);
and U2814 (N_2814,In_759,In_1936);
and U2815 (N_2815,In_1539,In_1171);
nor U2816 (N_2816,In_1555,In_1019);
and U2817 (N_2817,In_993,In_1449);
or U2818 (N_2818,In_1978,In_277);
nor U2819 (N_2819,In_1,In_437);
or U2820 (N_2820,In_1261,In_38);
and U2821 (N_2821,In_283,In_1513);
nor U2822 (N_2822,In_606,In_1605);
nand U2823 (N_2823,In_172,In_873);
or U2824 (N_2824,In_1494,In_867);
nor U2825 (N_2825,In_693,In_1597);
xor U2826 (N_2826,In_736,In_833);
nand U2827 (N_2827,In_768,In_650);
or U2828 (N_2828,In_792,In_1019);
nand U2829 (N_2829,In_73,In_566);
nand U2830 (N_2830,In_423,In_563);
or U2831 (N_2831,In_1094,In_858);
nor U2832 (N_2832,In_1618,In_1218);
or U2833 (N_2833,In_1292,In_1);
or U2834 (N_2834,In_1794,In_1612);
or U2835 (N_2835,In_1874,In_875);
or U2836 (N_2836,In_1142,In_1299);
nor U2837 (N_2837,In_11,In_185);
and U2838 (N_2838,In_1684,In_331);
nor U2839 (N_2839,In_1656,In_624);
xnor U2840 (N_2840,In_1214,In_987);
nand U2841 (N_2841,In_1119,In_844);
and U2842 (N_2842,In_1143,In_1103);
nor U2843 (N_2843,In_242,In_678);
or U2844 (N_2844,In_635,In_414);
and U2845 (N_2845,In_329,In_852);
or U2846 (N_2846,In_911,In_1537);
nand U2847 (N_2847,In_1536,In_1282);
or U2848 (N_2848,In_82,In_655);
nor U2849 (N_2849,In_1098,In_627);
nor U2850 (N_2850,In_1197,In_896);
nand U2851 (N_2851,In_542,In_1060);
nand U2852 (N_2852,In_1467,In_906);
xnor U2853 (N_2853,In_163,In_723);
or U2854 (N_2854,In_994,In_695);
nor U2855 (N_2855,In_1339,In_854);
nor U2856 (N_2856,In_1976,In_1476);
and U2857 (N_2857,In_863,In_1074);
or U2858 (N_2858,In_968,In_1169);
nand U2859 (N_2859,In_157,In_849);
and U2860 (N_2860,In_563,In_1018);
nand U2861 (N_2861,In_397,In_1915);
nand U2862 (N_2862,In_1968,In_718);
nand U2863 (N_2863,In_1396,In_670);
and U2864 (N_2864,In_396,In_1662);
nor U2865 (N_2865,In_1460,In_1793);
and U2866 (N_2866,In_182,In_1119);
or U2867 (N_2867,In_461,In_1617);
and U2868 (N_2868,In_678,In_273);
nand U2869 (N_2869,In_27,In_201);
or U2870 (N_2870,In_296,In_770);
nand U2871 (N_2871,In_731,In_164);
or U2872 (N_2872,In_235,In_564);
xnor U2873 (N_2873,In_1362,In_1251);
and U2874 (N_2874,In_1395,In_1757);
or U2875 (N_2875,In_368,In_1013);
nor U2876 (N_2876,In_1861,In_1290);
nand U2877 (N_2877,In_577,In_1702);
or U2878 (N_2878,In_771,In_808);
xnor U2879 (N_2879,In_270,In_260);
nor U2880 (N_2880,In_333,In_966);
nor U2881 (N_2881,In_1253,In_1404);
and U2882 (N_2882,In_314,In_714);
nand U2883 (N_2883,In_1082,In_328);
xor U2884 (N_2884,In_1968,In_1999);
and U2885 (N_2885,In_495,In_1712);
or U2886 (N_2886,In_441,In_720);
and U2887 (N_2887,In_477,In_1660);
nand U2888 (N_2888,In_1798,In_276);
and U2889 (N_2889,In_1421,In_839);
and U2890 (N_2890,In_1181,In_76);
or U2891 (N_2891,In_1971,In_611);
and U2892 (N_2892,In_960,In_1530);
nand U2893 (N_2893,In_1738,In_1632);
and U2894 (N_2894,In_126,In_1910);
and U2895 (N_2895,In_854,In_1690);
nor U2896 (N_2896,In_1228,In_1);
xnor U2897 (N_2897,In_1281,In_1698);
and U2898 (N_2898,In_902,In_859);
nor U2899 (N_2899,In_909,In_800);
nand U2900 (N_2900,In_1484,In_972);
and U2901 (N_2901,In_1294,In_616);
nand U2902 (N_2902,In_1770,In_1409);
and U2903 (N_2903,In_1061,In_358);
xnor U2904 (N_2904,In_1659,In_729);
xor U2905 (N_2905,In_1337,In_543);
and U2906 (N_2906,In_338,In_633);
nand U2907 (N_2907,In_194,In_1695);
nor U2908 (N_2908,In_729,In_340);
nand U2909 (N_2909,In_1334,In_38);
and U2910 (N_2910,In_1353,In_787);
and U2911 (N_2911,In_800,In_1006);
and U2912 (N_2912,In_606,In_1690);
xor U2913 (N_2913,In_1253,In_0);
nand U2914 (N_2914,In_165,In_15);
and U2915 (N_2915,In_828,In_1767);
and U2916 (N_2916,In_317,In_320);
nand U2917 (N_2917,In_19,In_182);
nor U2918 (N_2918,In_1819,In_1416);
nand U2919 (N_2919,In_1564,In_1492);
and U2920 (N_2920,In_1012,In_1284);
or U2921 (N_2921,In_1417,In_654);
or U2922 (N_2922,In_242,In_1995);
nand U2923 (N_2923,In_1661,In_1234);
and U2924 (N_2924,In_1738,In_1981);
and U2925 (N_2925,In_1620,In_585);
and U2926 (N_2926,In_1351,In_1683);
and U2927 (N_2927,In_642,In_805);
nor U2928 (N_2928,In_1040,In_1617);
nor U2929 (N_2929,In_1098,In_1440);
nand U2930 (N_2930,In_1820,In_1742);
and U2931 (N_2931,In_1352,In_1443);
or U2932 (N_2932,In_470,In_1424);
or U2933 (N_2933,In_1371,In_417);
or U2934 (N_2934,In_1856,In_1946);
nor U2935 (N_2935,In_454,In_741);
and U2936 (N_2936,In_1546,In_771);
or U2937 (N_2937,In_474,In_1420);
or U2938 (N_2938,In_252,In_1495);
nand U2939 (N_2939,In_845,In_851);
or U2940 (N_2940,In_545,In_155);
and U2941 (N_2941,In_1929,In_958);
and U2942 (N_2942,In_1671,In_320);
and U2943 (N_2943,In_771,In_1205);
and U2944 (N_2944,In_315,In_126);
and U2945 (N_2945,In_1925,In_833);
xor U2946 (N_2946,In_1666,In_847);
nor U2947 (N_2947,In_490,In_224);
nor U2948 (N_2948,In_1926,In_1562);
nand U2949 (N_2949,In_391,In_186);
or U2950 (N_2950,In_1271,In_1461);
xor U2951 (N_2951,In_924,In_770);
nor U2952 (N_2952,In_354,In_1355);
nor U2953 (N_2953,In_1166,In_836);
xnor U2954 (N_2954,In_761,In_841);
and U2955 (N_2955,In_197,In_107);
nor U2956 (N_2956,In_1380,In_1162);
and U2957 (N_2957,In_1965,In_832);
and U2958 (N_2958,In_995,In_1222);
nand U2959 (N_2959,In_668,In_1853);
xor U2960 (N_2960,In_1456,In_1916);
nand U2961 (N_2961,In_403,In_1306);
nor U2962 (N_2962,In_185,In_14);
or U2963 (N_2963,In_342,In_619);
nand U2964 (N_2964,In_1950,In_700);
nor U2965 (N_2965,In_1584,In_1438);
nand U2966 (N_2966,In_1820,In_1061);
or U2967 (N_2967,In_279,In_313);
and U2968 (N_2968,In_1014,In_314);
nor U2969 (N_2969,In_921,In_240);
nand U2970 (N_2970,In_1568,In_398);
nand U2971 (N_2971,In_1722,In_1325);
and U2972 (N_2972,In_932,In_151);
or U2973 (N_2973,In_979,In_1968);
nand U2974 (N_2974,In_1652,In_1501);
and U2975 (N_2975,In_801,In_1066);
or U2976 (N_2976,In_1411,In_136);
nand U2977 (N_2977,In_1305,In_1657);
and U2978 (N_2978,In_97,In_910);
xnor U2979 (N_2979,In_333,In_1011);
nor U2980 (N_2980,In_336,In_1032);
and U2981 (N_2981,In_1946,In_1159);
xor U2982 (N_2982,In_512,In_55);
xnor U2983 (N_2983,In_1070,In_1317);
xor U2984 (N_2984,In_1230,In_1101);
nand U2985 (N_2985,In_1789,In_1488);
and U2986 (N_2986,In_1380,In_950);
or U2987 (N_2987,In_352,In_1027);
and U2988 (N_2988,In_1119,In_161);
nand U2989 (N_2989,In_980,In_1412);
nor U2990 (N_2990,In_1720,In_1944);
and U2991 (N_2991,In_358,In_1625);
or U2992 (N_2992,In_174,In_682);
or U2993 (N_2993,In_190,In_1808);
or U2994 (N_2994,In_417,In_837);
xnor U2995 (N_2995,In_73,In_1165);
nand U2996 (N_2996,In_1031,In_1033);
or U2997 (N_2997,In_1645,In_1466);
and U2998 (N_2998,In_1216,In_1279);
or U2999 (N_2999,In_284,In_1422);
xor U3000 (N_3000,In_1467,In_1123);
and U3001 (N_3001,In_1293,In_1540);
or U3002 (N_3002,In_1724,In_557);
xor U3003 (N_3003,In_721,In_133);
nand U3004 (N_3004,In_1871,In_1134);
and U3005 (N_3005,In_1455,In_1197);
or U3006 (N_3006,In_904,In_1914);
nand U3007 (N_3007,In_927,In_225);
nand U3008 (N_3008,In_767,In_318);
nand U3009 (N_3009,In_228,In_884);
nand U3010 (N_3010,In_266,In_1579);
nand U3011 (N_3011,In_1525,In_441);
xnor U3012 (N_3012,In_954,In_845);
nand U3013 (N_3013,In_950,In_1570);
nor U3014 (N_3014,In_1813,In_924);
and U3015 (N_3015,In_1894,In_1699);
nor U3016 (N_3016,In_1951,In_361);
or U3017 (N_3017,In_1521,In_1428);
nor U3018 (N_3018,In_800,In_980);
and U3019 (N_3019,In_1705,In_242);
or U3020 (N_3020,In_442,In_761);
nor U3021 (N_3021,In_97,In_1209);
and U3022 (N_3022,In_1900,In_1802);
or U3023 (N_3023,In_1770,In_1939);
nor U3024 (N_3024,In_1343,In_1358);
or U3025 (N_3025,In_473,In_1842);
nand U3026 (N_3026,In_1695,In_1026);
or U3027 (N_3027,In_91,In_1129);
nor U3028 (N_3028,In_1485,In_1624);
xor U3029 (N_3029,In_700,In_109);
nand U3030 (N_3030,In_362,In_961);
nor U3031 (N_3031,In_986,In_1809);
and U3032 (N_3032,In_1410,In_173);
nand U3033 (N_3033,In_1714,In_1103);
nor U3034 (N_3034,In_1196,In_1916);
nand U3035 (N_3035,In_963,In_7);
nand U3036 (N_3036,In_1724,In_1554);
and U3037 (N_3037,In_203,In_1910);
xor U3038 (N_3038,In_1933,In_751);
or U3039 (N_3039,In_1179,In_107);
or U3040 (N_3040,In_479,In_1062);
or U3041 (N_3041,In_1057,In_1326);
nor U3042 (N_3042,In_1904,In_1876);
nand U3043 (N_3043,In_923,In_1940);
and U3044 (N_3044,In_1185,In_204);
xor U3045 (N_3045,In_550,In_1266);
xor U3046 (N_3046,In_20,In_286);
nand U3047 (N_3047,In_1651,In_555);
xor U3048 (N_3048,In_1612,In_1026);
nor U3049 (N_3049,In_1331,In_385);
and U3050 (N_3050,In_820,In_1736);
xnor U3051 (N_3051,In_238,In_1547);
nor U3052 (N_3052,In_1621,In_656);
nor U3053 (N_3053,In_1129,In_1047);
nand U3054 (N_3054,In_1434,In_932);
or U3055 (N_3055,In_1143,In_325);
and U3056 (N_3056,In_1869,In_1536);
nor U3057 (N_3057,In_781,In_1074);
nand U3058 (N_3058,In_955,In_147);
or U3059 (N_3059,In_955,In_1619);
nand U3060 (N_3060,In_112,In_717);
and U3061 (N_3061,In_1433,In_1567);
xor U3062 (N_3062,In_699,In_219);
nor U3063 (N_3063,In_1990,In_1559);
nand U3064 (N_3064,In_1475,In_979);
nor U3065 (N_3065,In_1626,In_1685);
and U3066 (N_3066,In_995,In_1269);
nand U3067 (N_3067,In_1030,In_1348);
and U3068 (N_3068,In_1493,In_1258);
xor U3069 (N_3069,In_274,In_1956);
xor U3070 (N_3070,In_166,In_488);
or U3071 (N_3071,In_1438,In_1907);
or U3072 (N_3072,In_297,In_182);
and U3073 (N_3073,In_1138,In_623);
xor U3074 (N_3074,In_769,In_1469);
and U3075 (N_3075,In_502,In_960);
and U3076 (N_3076,In_787,In_1299);
or U3077 (N_3077,In_1434,In_510);
nand U3078 (N_3078,In_370,In_1980);
and U3079 (N_3079,In_778,In_1073);
nor U3080 (N_3080,In_208,In_1419);
and U3081 (N_3081,In_815,In_726);
nand U3082 (N_3082,In_318,In_783);
and U3083 (N_3083,In_18,In_489);
nand U3084 (N_3084,In_579,In_1109);
nand U3085 (N_3085,In_137,In_1503);
nand U3086 (N_3086,In_275,In_249);
nor U3087 (N_3087,In_530,In_287);
nor U3088 (N_3088,In_1126,In_885);
nor U3089 (N_3089,In_814,In_958);
and U3090 (N_3090,In_827,In_473);
or U3091 (N_3091,In_610,In_1649);
xnor U3092 (N_3092,In_469,In_1919);
and U3093 (N_3093,In_990,In_1114);
and U3094 (N_3094,In_545,In_1454);
and U3095 (N_3095,In_679,In_739);
nand U3096 (N_3096,In_1105,In_594);
nor U3097 (N_3097,In_1005,In_838);
or U3098 (N_3098,In_1786,In_343);
nand U3099 (N_3099,In_881,In_1049);
nand U3100 (N_3100,In_806,In_1455);
or U3101 (N_3101,In_1246,In_1230);
nand U3102 (N_3102,In_1471,In_1304);
and U3103 (N_3103,In_736,In_1701);
nand U3104 (N_3104,In_935,In_1222);
nor U3105 (N_3105,In_1839,In_810);
and U3106 (N_3106,In_496,In_1585);
nor U3107 (N_3107,In_1396,In_1515);
and U3108 (N_3108,In_1193,In_1797);
and U3109 (N_3109,In_1212,In_88);
and U3110 (N_3110,In_891,In_1756);
and U3111 (N_3111,In_239,In_1628);
or U3112 (N_3112,In_690,In_1995);
xnor U3113 (N_3113,In_1398,In_1598);
or U3114 (N_3114,In_682,In_673);
nor U3115 (N_3115,In_1901,In_708);
nand U3116 (N_3116,In_1433,In_778);
nand U3117 (N_3117,In_1930,In_667);
and U3118 (N_3118,In_1271,In_590);
nor U3119 (N_3119,In_1778,In_1544);
nand U3120 (N_3120,In_798,In_1896);
nand U3121 (N_3121,In_1613,In_1336);
nor U3122 (N_3122,In_1059,In_1133);
nor U3123 (N_3123,In_617,In_1017);
nand U3124 (N_3124,In_1970,In_1288);
nor U3125 (N_3125,In_52,In_1226);
nor U3126 (N_3126,In_774,In_1805);
nand U3127 (N_3127,In_1183,In_1906);
nand U3128 (N_3128,In_1371,In_1833);
or U3129 (N_3129,In_272,In_1609);
xor U3130 (N_3130,In_1700,In_1667);
nor U3131 (N_3131,In_1950,In_1274);
nand U3132 (N_3132,In_1105,In_1708);
nor U3133 (N_3133,In_1914,In_857);
nor U3134 (N_3134,In_1171,In_720);
or U3135 (N_3135,In_650,In_1395);
and U3136 (N_3136,In_1094,In_273);
nor U3137 (N_3137,In_1926,In_1452);
and U3138 (N_3138,In_114,In_1556);
nor U3139 (N_3139,In_307,In_1526);
nor U3140 (N_3140,In_1549,In_890);
and U3141 (N_3141,In_1608,In_1792);
or U3142 (N_3142,In_1128,In_1641);
nor U3143 (N_3143,In_1292,In_1345);
xnor U3144 (N_3144,In_1434,In_955);
nor U3145 (N_3145,In_943,In_1420);
nor U3146 (N_3146,In_1512,In_1100);
xnor U3147 (N_3147,In_1862,In_869);
nor U3148 (N_3148,In_1037,In_409);
xor U3149 (N_3149,In_1843,In_204);
or U3150 (N_3150,In_150,In_705);
or U3151 (N_3151,In_1225,In_741);
and U3152 (N_3152,In_541,In_132);
and U3153 (N_3153,In_1281,In_543);
and U3154 (N_3154,In_1869,In_16);
nand U3155 (N_3155,In_1084,In_1203);
nand U3156 (N_3156,In_206,In_1177);
or U3157 (N_3157,In_561,In_888);
or U3158 (N_3158,In_1842,In_1340);
nand U3159 (N_3159,In_224,In_1501);
xor U3160 (N_3160,In_1604,In_284);
nand U3161 (N_3161,In_1430,In_1814);
nand U3162 (N_3162,In_1116,In_1951);
and U3163 (N_3163,In_731,In_1505);
and U3164 (N_3164,In_1113,In_1897);
nor U3165 (N_3165,In_1119,In_1858);
or U3166 (N_3166,In_1041,In_1504);
nor U3167 (N_3167,In_792,In_1127);
nor U3168 (N_3168,In_56,In_1165);
nand U3169 (N_3169,In_129,In_1381);
xnor U3170 (N_3170,In_777,In_57);
xnor U3171 (N_3171,In_1294,In_195);
and U3172 (N_3172,In_1450,In_367);
nor U3173 (N_3173,In_286,In_83);
nor U3174 (N_3174,In_1529,In_365);
and U3175 (N_3175,In_1438,In_1896);
nand U3176 (N_3176,In_824,In_589);
xor U3177 (N_3177,In_689,In_1949);
nand U3178 (N_3178,In_316,In_1052);
or U3179 (N_3179,In_672,In_646);
or U3180 (N_3180,In_115,In_1236);
nor U3181 (N_3181,In_1038,In_1414);
nand U3182 (N_3182,In_1351,In_210);
or U3183 (N_3183,In_1128,In_1961);
and U3184 (N_3184,In_1034,In_1258);
nor U3185 (N_3185,In_1505,In_447);
and U3186 (N_3186,In_1565,In_621);
and U3187 (N_3187,In_406,In_315);
or U3188 (N_3188,In_1410,In_564);
xnor U3189 (N_3189,In_190,In_93);
or U3190 (N_3190,In_377,In_923);
nor U3191 (N_3191,In_428,In_249);
nand U3192 (N_3192,In_570,In_1552);
nor U3193 (N_3193,In_339,In_781);
nand U3194 (N_3194,In_1206,In_1490);
nor U3195 (N_3195,In_583,In_937);
and U3196 (N_3196,In_956,In_1872);
nor U3197 (N_3197,In_1335,In_625);
and U3198 (N_3198,In_858,In_1828);
xnor U3199 (N_3199,In_340,In_836);
and U3200 (N_3200,In_1119,In_238);
or U3201 (N_3201,In_903,In_1170);
nor U3202 (N_3202,In_156,In_368);
xnor U3203 (N_3203,In_1836,In_7);
nor U3204 (N_3204,In_1448,In_566);
or U3205 (N_3205,In_1018,In_1757);
and U3206 (N_3206,In_248,In_463);
nor U3207 (N_3207,In_116,In_1011);
or U3208 (N_3208,In_438,In_1514);
xnor U3209 (N_3209,In_308,In_1507);
and U3210 (N_3210,In_1094,In_974);
or U3211 (N_3211,In_1139,In_447);
or U3212 (N_3212,In_89,In_594);
or U3213 (N_3213,In_551,In_948);
xor U3214 (N_3214,In_1828,In_1646);
or U3215 (N_3215,In_1025,In_1700);
and U3216 (N_3216,In_494,In_1516);
xnor U3217 (N_3217,In_123,In_528);
xnor U3218 (N_3218,In_956,In_1932);
nor U3219 (N_3219,In_700,In_565);
nand U3220 (N_3220,In_1754,In_518);
or U3221 (N_3221,In_1645,In_196);
or U3222 (N_3222,In_1484,In_577);
nand U3223 (N_3223,In_1395,In_1643);
nand U3224 (N_3224,In_1186,In_700);
xnor U3225 (N_3225,In_1715,In_1932);
nor U3226 (N_3226,In_490,In_1610);
or U3227 (N_3227,In_298,In_326);
nor U3228 (N_3228,In_225,In_1066);
nand U3229 (N_3229,In_1402,In_856);
nor U3230 (N_3230,In_1849,In_1343);
and U3231 (N_3231,In_1014,In_1523);
nand U3232 (N_3232,In_1594,In_1347);
nand U3233 (N_3233,In_804,In_1905);
xnor U3234 (N_3234,In_1163,In_1375);
xnor U3235 (N_3235,In_981,In_1387);
and U3236 (N_3236,In_1632,In_471);
and U3237 (N_3237,In_483,In_210);
and U3238 (N_3238,In_1331,In_47);
xor U3239 (N_3239,In_1727,In_776);
nor U3240 (N_3240,In_933,In_1066);
nor U3241 (N_3241,In_1687,In_1029);
and U3242 (N_3242,In_217,In_1070);
and U3243 (N_3243,In_195,In_1068);
nand U3244 (N_3244,In_1744,In_1368);
nand U3245 (N_3245,In_1141,In_582);
nand U3246 (N_3246,In_221,In_502);
nor U3247 (N_3247,In_208,In_439);
nand U3248 (N_3248,In_1501,In_1811);
nor U3249 (N_3249,In_1695,In_474);
nor U3250 (N_3250,In_1905,In_452);
and U3251 (N_3251,In_1188,In_424);
and U3252 (N_3252,In_1466,In_440);
and U3253 (N_3253,In_1711,In_1497);
and U3254 (N_3254,In_1645,In_866);
xor U3255 (N_3255,In_1676,In_969);
or U3256 (N_3256,In_1122,In_1106);
and U3257 (N_3257,In_760,In_394);
or U3258 (N_3258,In_365,In_1468);
or U3259 (N_3259,In_1893,In_1275);
and U3260 (N_3260,In_830,In_934);
nand U3261 (N_3261,In_471,In_38);
xnor U3262 (N_3262,In_1797,In_27);
nand U3263 (N_3263,In_363,In_687);
xnor U3264 (N_3264,In_1598,In_446);
or U3265 (N_3265,In_1905,In_1151);
nor U3266 (N_3266,In_1327,In_470);
or U3267 (N_3267,In_1791,In_1571);
and U3268 (N_3268,In_825,In_1539);
nand U3269 (N_3269,In_459,In_680);
or U3270 (N_3270,In_846,In_834);
nor U3271 (N_3271,In_1157,In_1610);
nand U3272 (N_3272,In_537,In_129);
or U3273 (N_3273,In_431,In_1471);
or U3274 (N_3274,In_699,In_1024);
xor U3275 (N_3275,In_1874,In_938);
nand U3276 (N_3276,In_564,In_1493);
nor U3277 (N_3277,In_23,In_1832);
xnor U3278 (N_3278,In_1543,In_537);
and U3279 (N_3279,In_1388,In_1451);
nand U3280 (N_3280,In_90,In_190);
or U3281 (N_3281,In_641,In_785);
or U3282 (N_3282,In_740,In_813);
or U3283 (N_3283,In_990,In_748);
nor U3284 (N_3284,In_1323,In_559);
or U3285 (N_3285,In_1883,In_1956);
or U3286 (N_3286,In_596,In_609);
or U3287 (N_3287,In_1487,In_76);
or U3288 (N_3288,In_88,In_35);
xor U3289 (N_3289,In_1348,In_1442);
xnor U3290 (N_3290,In_1918,In_1159);
nand U3291 (N_3291,In_1553,In_362);
or U3292 (N_3292,In_881,In_918);
nor U3293 (N_3293,In_616,In_1424);
or U3294 (N_3294,In_819,In_171);
and U3295 (N_3295,In_1774,In_135);
nor U3296 (N_3296,In_1586,In_1765);
or U3297 (N_3297,In_1081,In_779);
or U3298 (N_3298,In_1411,In_1094);
or U3299 (N_3299,In_490,In_1066);
nor U3300 (N_3300,In_923,In_1674);
nand U3301 (N_3301,In_53,In_525);
or U3302 (N_3302,In_473,In_750);
and U3303 (N_3303,In_523,In_1268);
nor U3304 (N_3304,In_1157,In_1568);
and U3305 (N_3305,In_1567,In_1346);
nor U3306 (N_3306,In_136,In_1731);
and U3307 (N_3307,In_973,In_448);
or U3308 (N_3308,In_926,In_1087);
and U3309 (N_3309,In_263,In_1341);
nand U3310 (N_3310,In_2,In_1597);
or U3311 (N_3311,In_1092,In_1636);
or U3312 (N_3312,In_1415,In_1870);
and U3313 (N_3313,In_317,In_606);
nor U3314 (N_3314,In_1071,In_186);
nor U3315 (N_3315,In_1201,In_1205);
or U3316 (N_3316,In_483,In_1620);
and U3317 (N_3317,In_335,In_1466);
or U3318 (N_3318,In_673,In_1817);
nand U3319 (N_3319,In_643,In_761);
nand U3320 (N_3320,In_301,In_1491);
nor U3321 (N_3321,In_119,In_1142);
xnor U3322 (N_3322,In_1895,In_1658);
nor U3323 (N_3323,In_1370,In_773);
nand U3324 (N_3324,In_340,In_606);
and U3325 (N_3325,In_1588,In_1840);
nand U3326 (N_3326,In_194,In_1346);
nand U3327 (N_3327,In_1783,In_498);
nor U3328 (N_3328,In_275,In_1991);
xnor U3329 (N_3329,In_818,In_1332);
or U3330 (N_3330,In_1276,In_1782);
and U3331 (N_3331,In_1571,In_409);
nand U3332 (N_3332,In_413,In_94);
nor U3333 (N_3333,In_1396,In_1340);
or U3334 (N_3334,In_769,In_1750);
nand U3335 (N_3335,In_818,In_791);
or U3336 (N_3336,In_971,In_1195);
nor U3337 (N_3337,In_1307,In_729);
nand U3338 (N_3338,In_1422,In_758);
nor U3339 (N_3339,In_318,In_888);
nor U3340 (N_3340,In_1032,In_1003);
xnor U3341 (N_3341,In_755,In_608);
nor U3342 (N_3342,In_648,In_1669);
nor U3343 (N_3343,In_1817,In_801);
nand U3344 (N_3344,In_424,In_927);
and U3345 (N_3345,In_1150,In_1183);
xnor U3346 (N_3346,In_1652,In_871);
and U3347 (N_3347,In_671,In_524);
nand U3348 (N_3348,In_718,In_1727);
nand U3349 (N_3349,In_1016,In_663);
nor U3350 (N_3350,In_1328,In_542);
xnor U3351 (N_3351,In_447,In_1532);
or U3352 (N_3352,In_473,In_1544);
or U3353 (N_3353,In_629,In_1408);
and U3354 (N_3354,In_1314,In_459);
and U3355 (N_3355,In_1698,In_964);
and U3356 (N_3356,In_549,In_1561);
or U3357 (N_3357,In_1696,In_1173);
nand U3358 (N_3358,In_1056,In_1647);
or U3359 (N_3359,In_929,In_558);
or U3360 (N_3360,In_792,In_1586);
and U3361 (N_3361,In_1256,In_1440);
nor U3362 (N_3362,In_802,In_1826);
nor U3363 (N_3363,In_1649,In_1634);
xor U3364 (N_3364,In_1289,In_1005);
nand U3365 (N_3365,In_765,In_569);
or U3366 (N_3366,In_1466,In_950);
xor U3367 (N_3367,In_211,In_1497);
nand U3368 (N_3368,In_1271,In_267);
nand U3369 (N_3369,In_1326,In_44);
nor U3370 (N_3370,In_1484,In_985);
and U3371 (N_3371,In_946,In_1971);
and U3372 (N_3372,In_1547,In_808);
and U3373 (N_3373,In_28,In_160);
nand U3374 (N_3374,In_339,In_164);
or U3375 (N_3375,In_1425,In_878);
nand U3376 (N_3376,In_352,In_1145);
nand U3377 (N_3377,In_32,In_278);
and U3378 (N_3378,In_1988,In_1978);
and U3379 (N_3379,In_153,In_98);
xnor U3380 (N_3380,In_1634,In_1737);
and U3381 (N_3381,In_692,In_1141);
nand U3382 (N_3382,In_1197,In_646);
and U3383 (N_3383,In_705,In_1917);
nand U3384 (N_3384,In_232,In_51);
and U3385 (N_3385,In_567,In_1583);
nor U3386 (N_3386,In_437,In_1827);
nor U3387 (N_3387,In_621,In_763);
and U3388 (N_3388,In_834,In_980);
and U3389 (N_3389,In_1328,In_1582);
and U3390 (N_3390,In_1573,In_1099);
or U3391 (N_3391,In_215,In_508);
or U3392 (N_3392,In_1225,In_1729);
and U3393 (N_3393,In_924,In_1443);
nand U3394 (N_3394,In_1118,In_400);
or U3395 (N_3395,In_29,In_1524);
nor U3396 (N_3396,In_239,In_1788);
nand U3397 (N_3397,In_21,In_1962);
and U3398 (N_3398,In_1366,In_1184);
nor U3399 (N_3399,In_619,In_1785);
nor U3400 (N_3400,In_706,In_1657);
nand U3401 (N_3401,In_684,In_1565);
nor U3402 (N_3402,In_1133,In_1775);
and U3403 (N_3403,In_384,In_1711);
nand U3404 (N_3404,In_926,In_1920);
nand U3405 (N_3405,In_1029,In_821);
or U3406 (N_3406,In_616,In_783);
and U3407 (N_3407,In_819,In_232);
nor U3408 (N_3408,In_429,In_718);
nor U3409 (N_3409,In_1454,In_409);
nand U3410 (N_3410,In_66,In_1071);
nand U3411 (N_3411,In_30,In_1265);
nor U3412 (N_3412,In_1283,In_1478);
and U3413 (N_3413,In_272,In_265);
nand U3414 (N_3414,In_1965,In_1876);
nor U3415 (N_3415,In_852,In_276);
nor U3416 (N_3416,In_1269,In_690);
nor U3417 (N_3417,In_443,In_560);
and U3418 (N_3418,In_755,In_1642);
or U3419 (N_3419,In_285,In_522);
nor U3420 (N_3420,In_424,In_811);
nor U3421 (N_3421,In_1796,In_738);
or U3422 (N_3422,In_340,In_1353);
nand U3423 (N_3423,In_1764,In_1528);
nand U3424 (N_3424,In_1439,In_992);
xnor U3425 (N_3425,In_539,In_1589);
nor U3426 (N_3426,In_1529,In_79);
nand U3427 (N_3427,In_1202,In_1508);
xnor U3428 (N_3428,In_65,In_1202);
xor U3429 (N_3429,In_668,In_915);
or U3430 (N_3430,In_1534,In_1657);
nor U3431 (N_3431,In_1465,In_1925);
xnor U3432 (N_3432,In_1448,In_1826);
nand U3433 (N_3433,In_560,In_1385);
or U3434 (N_3434,In_1110,In_1802);
nand U3435 (N_3435,In_402,In_327);
nor U3436 (N_3436,In_119,In_213);
and U3437 (N_3437,In_697,In_1874);
nor U3438 (N_3438,In_1307,In_1405);
nor U3439 (N_3439,In_38,In_1947);
nand U3440 (N_3440,In_1244,In_1424);
nand U3441 (N_3441,In_1134,In_1459);
nor U3442 (N_3442,In_648,In_75);
or U3443 (N_3443,In_1564,In_1842);
or U3444 (N_3444,In_749,In_865);
nand U3445 (N_3445,In_1160,In_1790);
and U3446 (N_3446,In_715,In_239);
nand U3447 (N_3447,In_859,In_1693);
or U3448 (N_3448,In_1304,In_1351);
nor U3449 (N_3449,In_1156,In_1654);
or U3450 (N_3450,In_195,In_692);
and U3451 (N_3451,In_1911,In_24);
or U3452 (N_3452,In_177,In_1458);
xnor U3453 (N_3453,In_1444,In_869);
nor U3454 (N_3454,In_1429,In_1982);
and U3455 (N_3455,In_1462,In_1773);
and U3456 (N_3456,In_1147,In_1415);
xnor U3457 (N_3457,In_1839,In_570);
or U3458 (N_3458,In_1585,In_269);
or U3459 (N_3459,In_1643,In_325);
and U3460 (N_3460,In_1031,In_1939);
or U3461 (N_3461,In_1156,In_896);
and U3462 (N_3462,In_1128,In_380);
or U3463 (N_3463,In_22,In_1030);
xnor U3464 (N_3464,In_1946,In_57);
nor U3465 (N_3465,In_1525,In_725);
or U3466 (N_3466,In_1998,In_1986);
nand U3467 (N_3467,In_402,In_812);
xor U3468 (N_3468,In_196,In_1063);
and U3469 (N_3469,In_250,In_1711);
or U3470 (N_3470,In_1526,In_1036);
nand U3471 (N_3471,In_1180,In_1041);
and U3472 (N_3472,In_598,In_783);
nor U3473 (N_3473,In_1196,In_38);
and U3474 (N_3474,In_329,In_31);
or U3475 (N_3475,In_556,In_1225);
or U3476 (N_3476,In_1576,In_622);
and U3477 (N_3477,In_972,In_1875);
xor U3478 (N_3478,In_97,In_878);
nand U3479 (N_3479,In_19,In_370);
xor U3480 (N_3480,In_97,In_1456);
nor U3481 (N_3481,In_868,In_1963);
and U3482 (N_3482,In_1084,In_1589);
nor U3483 (N_3483,In_1932,In_1339);
xnor U3484 (N_3484,In_824,In_722);
and U3485 (N_3485,In_897,In_1601);
and U3486 (N_3486,In_1203,In_557);
nand U3487 (N_3487,In_1721,In_994);
nor U3488 (N_3488,In_862,In_1294);
or U3489 (N_3489,In_765,In_467);
or U3490 (N_3490,In_24,In_21);
nand U3491 (N_3491,In_1125,In_1706);
nand U3492 (N_3492,In_1940,In_1202);
or U3493 (N_3493,In_561,In_965);
nand U3494 (N_3494,In_219,In_1676);
nor U3495 (N_3495,In_802,In_604);
nor U3496 (N_3496,In_584,In_1738);
or U3497 (N_3497,In_1051,In_1367);
nand U3498 (N_3498,In_1015,In_393);
and U3499 (N_3499,In_337,In_724);
or U3500 (N_3500,In_12,In_1126);
xnor U3501 (N_3501,In_1442,In_938);
and U3502 (N_3502,In_610,In_1957);
nor U3503 (N_3503,In_453,In_1529);
xor U3504 (N_3504,In_1263,In_806);
or U3505 (N_3505,In_299,In_941);
nand U3506 (N_3506,In_822,In_1970);
nand U3507 (N_3507,In_24,In_1915);
or U3508 (N_3508,In_396,In_1308);
nor U3509 (N_3509,In_1573,In_1143);
nand U3510 (N_3510,In_826,In_833);
nor U3511 (N_3511,In_1044,In_474);
and U3512 (N_3512,In_1561,In_564);
xor U3513 (N_3513,In_1505,In_140);
nor U3514 (N_3514,In_1786,In_1511);
or U3515 (N_3515,In_1489,In_1433);
or U3516 (N_3516,In_774,In_233);
nand U3517 (N_3517,In_1468,In_654);
nor U3518 (N_3518,In_1482,In_1645);
or U3519 (N_3519,In_514,In_1449);
nand U3520 (N_3520,In_64,In_799);
nor U3521 (N_3521,In_846,In_1833);
xor U3522 (N_3522,In_647,In_753);
nor U3523 (N_3523,In_1723,In_216);
and U3524 (N_3524,In_1624,In_551);
and U3525 (N_3525,In_1437,In_277);
nand U3526 (N_3526,In_1610,In_1778);
or U3527 (N_3527,In_1777,In_892);
or U3528 (N_3528,In_1622,In_3);
or U3529 (N_3529,In_691,In_57);
nand U3530 (N_3530,In_1728,In_352);
nor U3531 (N_3531,In_43,In_636);
nand U3532 (N_3532,In_98,In_531);
and U3533 (N_3533,In_406,In_760);
nand U3534 (N_3534,In_178,In_606);
or U3535 (N_3535,In_314,In_1368);
and U3536 (N_3536,In_1353,In_240);
or U3537 (N_3537,In_492,In_1027);
and U3538 (N_3538,In_1975,In_1129);
and U3539 (N_3539,In_32,In_376);
and U3540 (N_3540,In_127,In_328);
and U3541 (N_3541,In_1204,In_1168);
or U3542 (N_3542,In_832,In_34);
nand U3543 (N_3543,In_309,In_132);
and U3544 (N_3544,In_1618,In_1396);
and U3545 (N_3545,In_1132,In_1512);
and U3546 (N_3546,In_428,In_363);
xor U3547 (N_3547,In_184,In_589);
nor U3548 (N_3548,In_535,In_1285);
and U3549 (N_3549,In_108,In_1927);
and U3550 (N_3550,In_643,In_1433);
and U3551 (N_3551,In_1567,In_491);
nand U3552 (N_3552,In_196,In_1577);
or U3553 (N_3553,In_449,In_1293);
and U3554 (N_3554,In_69,In_1167);
nand U3555 (N_3555,In_1459,In_902);
and U3556 (N_3556,In_681,In_1688);
nor U3557 (N_3557,In_1077,In_817);
nand U3558 (N_3558,In_1719,In_1838);
nand U3559 (N_3559,In_188,In_1048);
nand U3560 (N_3560,In_1470,In_676);
and U3561 (N_3561,In_186,In_138);
nand U3562 (N_3562,In_723,In_788);
nand U3563 (N_3563,In_196,In_1235);
and U3564 (N_3564,In_45,In_470);
nand U3565 (N_3565,In_1283,In_1341);
nor U3566 (N_3566,In_887,In_455);
nor U3567 (N_3567,In_1628,In_1811);
and U3568 (N_3568,In_1760,In_1500);
or U3569 (N_3569,In_1241,In_403);
xnor U3570 (N_3570,In_1546,In_1960);
or U3571 (N_3571,In_1589,In_974);
or U3572 (N_3572,In_1727,In_1792);
or U3573 (N_3573,In_60,In_773);
or U3574 (N_3574,In_97,In_68);
or U3575 (N_3575,In_288,In_1458);
or U3576 (N_3576,In_794,In_1570);
and U3577 (N_3577,In_33,In_1802);
nor U3578 (N_3578,In_505,In_431);
and U3579 (N_3579,In_500,In_422);
or U3580 (N_3580,In_740,In_1483);
nor U3581 (N_3581,In_1923,In_828);
xor U3582 (N_3582,In_9,In_391);
nand U3583 (N_3583,In_286,In_668);
and U3584 (N_3584,In_363,In_980);
nand U3585 (N_3585,In_253,In_1468);
nor U3586 (N_3586,In_1668,In_161);
nor U3587 (N_3587,In_512,In_1712);
xor U3588 (N_3588,In_1773,In_431);
and U3589 (N_3589,In_1682,In_185);
nor U3590 (N_3590,In_1861,In_1011);
or U3591 (N_3591,In_957,In_1261);
or U3592 (N_3592,In_491,In_1657);
nand U3593 (N_3593,In_73,In_435);
or U3594 (N_3594,In_1266,In_1846);
or U3595 (N_3595,In_1813,In_1240);
nor U3596 (N_3596,In_2,In_892);
nor U3597 (N_3597,In_892,In_1473);
nor U3598 (N_3598,In_282,In_1223);
or U3599 (N_3599,In_1122,In_1713);
nand U3600 (N_3600,In_1506,In_802);
nor U3601 (N_3601,In_1892,In_1456);
nand U3602 (N_3602,In_1155,In_868);
nand U3603 (N_3603,In_9,In_262);
nor U3604 (N_3604,In_222,In_77);
nor U3605 (N_3605,In_1890,In_650);
nand U3606 (N_3606,In_1627,In_1710);
nand U3607 (N_3607,In_1859,In_1323);
nor U3608 (N_3608,In_371,In_1254);
and U3609 (N_3609,In_918,In_1299);
nand U3610 (N_3610,In_1058,In_315);
nor U3611 (N_3611,In_1602,In_183);
nand U3612 (N_3612,In_800,In_1728);
and U3613 (N_3613,In_1310,In_897);
nand U3614 (N_3614,In_1365,In_1645);
nand U3615 (N_3615,In_219,In_1526);
xor U3616 (N_3616,In_1798,In_1326);
or U3617 (N_3617,In_41,In_167);
or U3618 (N_3618,In_895,In_783);
nand U3619 (N_3619,In_402,In_1098);
and U3620 (N_3620,In_1956,In_1607);
and U3621 (N_3621,In_424,In_1292);
or U3622 (N_3622,In_1620,In_1286);
and U3623 (N_3623,In_1582,In_737);
nor U3624 (N_3624,In_1575,In_1570);
nor U3625 (N_3625,In_376,In_803);
xnor U3626 (N_3626,In_915,In_822);
nor U3627 (N_3627,In_692,In_1781);
or U3628 (N_3628,In_1771,In_545);
nand U3629 (N_3629,In_673,In_348);
or U3630 (N_3630,In_540,In_325);
or U3631 (N_3631,In_1373,In_891);
nand U3632 (N_3632,In_1667,In_187);
or U3633 (N_3633,In_1094,In_1232);
xnor U3634 (N_3634,In_998,In_528);
nor U3635 (N_3635,In_1948,In_746);
nor U3636 (N_3636,In_459,In_1163);
nand U3637 (N_3637,In_417,In_818);
nor U3638 (N_3638,In_1925,In_255);
nand U3639 (N_3639,In_1525,In_1921);
nand U3640 (N_3640,In_739,In_1884);
nand U3641 (N_3641,In_1369,In_1804);
and U3642 (N_3642,In_380,In_0);
or U3643 (N_3643,In_1238,In_1260);
or U3644 (N_3644,In_426,In_1915);
or U3645 (N_3645,In_463,In_443);
or U3646 (N_3646,In_502,In_1706);
nand U3647 (N_3647,In_1621,In_223);
and U3648 (N_3648,In_159,In_8);
or U3649 (N_3649,In_1019,In_1899);
xnor U3650 (N_3650,In_1824,In_431);
or U3651 (N_3651,In_555,In_793);
nor U3652 (N_3652,In_1924,In_1739);
or U3653 (N_3653,In_239,In_1698);
xor U3654 (N_3654,In_1657,In_1310);
or U3655 (N_3655,In_1143,In_1278);
nor U3656 (N_3656,In_996,In_1321);
nor U3657 (N_3657,In_1405,In_1662);
and U3658 (N_3658,In_1289,In_961);
or U3659 (N_3659,In_1036,In_1008);
or U3660 (N_3660,In_1716,In_1339);
or U3661 (N_3661,In_473,In_91);
nand U3662 (N_3662,In_1369,In_1483);
nand U3663 (N_3663,In_1971,In_1159);
xnor U3664 (N_3664,In_1461,In_7);
nand U3665 (N_3665,In_66,In_657);
nor U3666 (N_3666,In_1967,In_907);
nand U3667 (N_3667,In_1151,In_1476);
nand U3668 (N_3668,In_712,In_1867);
and U3669 (N_3669,In_1114,In_589);
nand U3670 (N_3670,In_1412,In_1678);
nand U3671 (N_3671,In_1071,In_1750);
or U3672 (N_3672,In_1815,In_1715);
and U3673 (N_3673,In_951,In_1897);
or U3674 (N_3674,In_963,In_722);
nand U3675 (N_3675,In_426,In_1154);
and U3676 (N_3676,In_660,In_173);
nor U3677 (N_3677,In_638,In_1250);
nand U3678 (N_3678,In_381,In_855);
nand U3679 (N_3679,In_928,In_1657);
nand U3680 (N_3680,In_590,In_557);
and U3681 (N_3681,In_1198,In_362);
nand U3682 (N_3682,In_689,In_535);
nor U3683 (N_3683,In_1512,In_994);
nand U3684 (N_3684,In_1751,In_522);
nand U3685 (N_3685,In_276,In_358);
nand U3686 (N_3686,In_1060,In_1751);
or U3687 (N_3687,In_1664,In_1146);
nand U3688 (N_3688,In_1016,In_793);
xor U3689 (N_3689,In_1271,In_375);
and U3690 (N_3690,In_1975,In_796);
xnor U3691 (N_3691,In_215,In_435);
and U3692 (N_3692,In_274,In_1507);
and U3693 (N_3693,In_1303,In_954);
and U3694 (N_3694,In_1396,In_205);
and U3695 (N_3695,In_565,In_857);
or U3696 (N_3696,In_281,In_1973);
nand U3697 (N_3697,In_1325,In_1017);
or U3698 (N_3698,In_532,In_38);
or U3699 (N_3699,In_929,In_524);
or U3700 (N_3700,In_982,In_155);
nor U3701 (N_3701,In_1502,In_236);
and U3702 (N_3702,In_1061,In_1200);
nand U3703 (N_3703,In_1370,In_797);
xor U3704 (N_3704,In_1057,In_1411);
nand U3705 (N_3705,In_82,In_1382);
and U3706 (N_3706,In_1920,In_975);
xnor U3707 (N_3707,In_461,In_663);
nand U3708 (N_3708,In_1909,In_1715);
or U3709 (N_3709,In_1172,In_553);
nand U3710 (N_3710,In_1957,In_1750);
nand U3711 (N_3711,In_26,In_1254);
nand U3712 (N_3712,In_631,In_109);
or U3713 (N_3713,In_1245,In_1634);
xor U3714 (N_3714,In_256,In_34);
or U3715 (N_3715,In_1988,In_565);
nor U3716 (N_3716,In_1966,In_311);
or U3717 (N_3717,In_689,In_443);
and U3718 (N_3718,In_752,In_171);
or U3719 (N_3719,In_829,In_270);
and U3720 (N_3720,In_1455,In_727);
or U3721 (N_3721,In_303,In_16);
nand U3722 (N_3722,In_64,In_1180);
and U3723 (N_3723,In_549,In_693);
or U3724 (N_3724,In_207,In_12);
nand U3725 (N_3725,In_646,In_635);
xor U3726 (N_3726,In_1578,In_1428);
or U3727 (N_3727,In_1700,In_1914);
nor U3728 (N_3728,In_1493,In_417);
nand U3729 (N_3729,In_1164,In_294);
nor U3730 (N_3730,In_450,In_515);
nand U3731 (N_3731,In_236,In_1651);
nand U3732 (N_3732,In_145,In_1287);
nand U3733 (N_3733,In_1248,In_654);
nand U3734 (N_3734,In_834,In_932);
nor U3735 (N_3735,In_891,In_1318);
or U3736 (N_3736,In_1766,In_47);
nand U3737 (N_3737,In_1253,In_753);
nor U3738 (N_3738,In_1043,In_435);
and U3739 (N_3739,In_385,In_1279);
and U3740 (N_3740,In_556,In_534);
or U3741 (N_3741,In_1353,In_368);
nand U3742 (N_3742,In_1695,In_1400);
or U3743 (N_3743,In_1363,In_804);
nor U3744 (N_3744,In_1236,In_372);
xor U3745 (N_3745,In_447,In_477);
or U3746 (N_3746,In_1936,In_18);
and U3747 (N_3747,In_1942,In_1652);
or U3748 (N_3748,In_88,In_1179);
or U3749 (N_3749,In_150,In_729);
nor U3750 (N_3750,In_52,In_361);
and U3751 (N_3751,In_84,In_244);
or U3752 (N_3752,In_1573,In_517);
or U3753 (N_3753,In_272,In_1651);
or U3754 (N_3754,In_1948,In_149);
or U3755 (N_3755,In_559,In_349);
xnor U3756 (N_3756,In_1214,In_163);
nor U3757 (N_3757,In_1290,In_1196);
and U3758 (N_3758,In_1390,In_1917);
xnor U3759 (N_3759,In_669,In_207);
nor U3760 (N_3760,In_1750,In_475);
or U3761 (N_3761,In_1149,In_1786);
xor U3762 (N_3762,In_863,In_1558);
and U3763 (N_3763,In_1148,In_1697);
nand U3764 (N_3764,In_1169,In_1518);
nor U3765 (N_3765,In_1880,In_1672);
nand U3766 (N_3766,In_356,In_799);
nor U3767 (N_3767,In_1378,In_1184);
xnor U3768 (N_3768,In_1708,In_1637);
and U3769 (N_3769,In_1555,In_941);
and U3770 (N_3770,In_790,In_665);
or U3771 (N_3771,In_1296,In_472);
xnor U3772 (N_3772,In_1484,In_1528);
nand U3773 (N_3773,In_1872,In_412);
and U3774 (N_3774,In_1699,In_1814);
xnor U3775 (N_3775,In_273,In_1941);
nand U3776 (N_3776,In_467,In_1171);
or U3777 (N_3777,In_119,In_132);
nand U3778 (N_3778,In_1278,In_1403);
xnor U3779 (N_3779,In_1336,In_947);
xnor U3780 (N_3780,In_831,In_1505);
nor U3781 (N_3781,In_1347,In_1212);
nand U3782 (N_3782,In_1183,In_216);
and U3783 (N_3783,In_888,In_1231);
or U3784 (N_3784,In_1059,In_200);
xor U3785 (N_3785,In_886,In_1126);
nor U3786 (N_3786,In_371,In_489);
or U3787 (N_3787,In_938,In_1301);
nand U3788 (N_3788,In_1825,In_1808);
or U3789 (N_3789,In_1908,In_817);
and U3790 (N_3790,In_1372,In_855);
nor U3791 (N_3791,In_793,In_1355);
nand U3792 (N_3792,In_64,In_717);
nand U3793 (N_3793,In_1066,In_47);
or U3794 (N_3794,In_1481,In_20);
and U3795 (N_3795,In_1202,In_545);
nand U3796 (N_3796,In_1604,In_623);
or U3797 (N_3797,In_305,In_1641);
and U3798 (N_3798,In_210,In_621);
and U3799 (N_3799,In_832,In_79);
nor U3800 (N_3800,In_146,In_1331);
nor U3801 (N_3801,In_221,In_832);
and U3802 (N_3802,In_436,In_1501);
nand U3803 (N_3803,In_1005,In_1846);
nand U3804 (N_3804,In_1344,In_1843);
nor U3805 (N_3805,In_72,In_1348);
nand U3806 (N_3806,In_767,In_1067);
nor U3807 (N_3807,In_1312,In_612);
or U3808 (N_3808,In_1718,In_19);
nand U3809 (N_3809,In_591,In_739);
nand U3810 (N_3810,In_842,In_953);
and U3811 (N_3811,In_54,In_1174);
nor U3812 (N_3812,In_278,In_28);
and U3813 (N_3813,In_34,In_1950);
and U3814 (N_3814,In_131,In_1659);
and U3815 (N_3815,In_1740,In_1367);
nand U3816 (N_3816,In_164,In_1412);
or U3817 (N_3817,In_1488,In_1360);
nand U3818 (N_3818,In_931,In_754);
nor U3819 (N_3819,In_548,In_924);
xnor U3820 (N_3820,In_705,In_1245);
xnor U3821 (N_3821,In_430,In_1699);
and U3822 (N_3822,In_868,In_167);
or U3823 (N_3823,In_790,In_152);
nand U3824 (N_3824,In_880,In_1114);
or U3825 (N_3825,In_717,In_1370);
or U3826 (N_3826,In_1216,In_899);
and U3827 (N_3827,In_51,In_1358);
or U3828 (N_3828,In_80,In_219);
nand U3829 (N_3829,In_492,In_1493);
and U3830 (N_3830,In_1135,In_763);
and U3831 (N_3831,In_1196,In_1546);
or U3832 (N_3832,In_940,In_168);
xor U3833 (N_3833,In_347,In_1218);
nor U3834 (N_3834,In_265,In_1943);
and U3835 (N_3835,In_904,In_36);
nand U3836 (N_3836,In_464,In_1835);
and U3837 (N_3837,In_491,In_692);
nand U3838 (N_3838,In_644,In_1066);
nor U3839 (N_3839,In_219,In_692);
and U3840 (N_3840,In_1488,In_322);
or U3841 (N_3841,In_566,In_299);
nor U3842 (N_3842,In_822,In_1418);
and U3843 (N_3843,In_1525,In_978);
or U3844 (N_3844,In_413,In_391);
or U3845 (N_3845,In_1720,In_1306);
or U3846 (N_3846,In_35,In_579);
or U3847 (N_3847,In_325,In_1259);
and U3848 (N_3848,In_1902,In_1080);
nor U3849 (N_3849,In_349,In_211);
nor U3850 (N_3850,In_467,In_1218);
or U3851 (N_3851,In_1168,In_1573);
nor U3852 (N_3852,In_108,In_1736);
or U3853 (N_3853,In_1546,In_302);
nand U3854 (N_3854,In_1963,In_764);
or U3855 (N_3855,In_1998,In_1923);
nand U3856 (N_3856,In_1500,In_1529);
and U3857 (N_3857,In_801,In_1268);
or U3858 (N_3858,In_341,In_1751);
or U3859 (N_3859,In_913,In_1662);
or U3860 (N_3860,In_1815,In_829);
and U3861 (N_3861,In_1271,In_608);
xnor U3862 (N_3862,In_1495,In_99);
and U3863 (N_3863,In_1732,In_1218);
nand U3864 (N_3864,In_952,In_13);
nor U3865 (N_3865,In_1745,In_1209);
nand U3866 (N_3866,In_1113,In_889);
or U3867 (N_3867,In_1799,In_379);
nand U3868 (N_3868,In_786,In_1162);
and U3869 (N_3869,In_797,In_1619);
nor U3870 (N_3870,In_169,In_102);
and U3871 (N_3871,In_1576,In_1229);
or U3872 (N_3872,In_1488,In_105);
nor U3873 (N_3873,In_403,In_343);
or U3874 (N_3874,In_535,In_782);
nor U3875 (N_3875,In_168,In_353);
nor U3876 (N_3876,In_376,In_1162);
nand U3877 (N_3877,In_1135,In_486);
or U3878 (N_3878,In_190,In_1421);
nand U3879 (N_3879,In_1310,In_1273);
and U3880 (N_3880,In_1992,In_447);
nand U3881 (N_3881,In_597,In_111);
or U3882 (N_3882,In_26,In_780);
nor U3883 (N_3883,In_944,In_1432);
nor U3884 (N_3884,In_1804,In_1816);
nor U3885 (N_3885,In_1085,In_1243);
nand U3886 (N_3886,In_1548,In_551);
nand U3887 (N_3887,In_1461,In_1533);
or U3888 (N_3888,In_853,In_1549);
xnor U3889 (N_3889,In_32,In_1201);
or U3890 (N_3890,In_387,In_1326);
nor U3891 (N_3891,In_763,In_855);
nand U3892 (N_3892,In_1512,In_149);
nor U3893 (N_3893,In_1423,In_1067);
nor U3894 (N_3894,In_177,In_1846);
nor U3895 (N_3895,In_1039,In_1212);
nand U3896 (N_3896,In_86,In_1274);
and U3897 (N_3897,In_411,In_805);
nor U3898 (N_3898,In_849,In_1440);
nor U3899 (N_3899,In_1829,In_1253);
or U3900 (N_3900,In_1959,In_484);
or U3901 (N_3901,In_1917,In_659);
nor U3902 (N_3902,In_1814,In_1086);
nor U3903 (N_3903,In_1137,In_54);
and U3904 (N_3904,In_1051,In_540);
and U3905 (N_3905,In_941,In_1580);
nand U3906 (N_3906,In_582,In_181);
or U3907 (N_3907,In_1031,In_928);
nand U3908 (N_3908,In_1159,In_512);
and U3909 (N_3909,In_464,In_1931);
and U3910 (N_3910,In_1956,In_841);
or U3911 (N_3911,In_776,In_65);
nand U3912 (N_3912,In_1691,In_790);
nand U3913 (N_3913,In_187,In_1862);
nand U3914 (N_3914,In_1576,In_1675);
or U3915 (N_3915,In_689,In_1146);
and U3916 (N_3916,In_551,In_151);
or U3917 (N_3917,In_1695,In_1892);
nand U3918 (N_3918,In_1292,In_704);
nand U3919 (N_3919,In_86,In_628);
and U3920 (N_3920,In_1748,In_499);
nand U3921 (N_3921,In_1119,In_36);
and U3922 (N_3922,In_712,In_1723);
nand U3923 (N_3923,In_206,In_1555);
and U3924 (N_3924,In_1760,In_1868);
and U3925 (N_3925,In_84,In_265);
nor U3926 (N_3926,In_107,In_1982);
and U3927 (N_3927,In_1606,In_1411);
and U3928 (N_3928,In_869,In_916);
or U3929 (N_3929,In_1929,In_219);
and U3930 (N_3930,In_76,In_1678);
nand U3931 (N_3931,In_1867,In_439);
nor U3932 (N_3932,In_548,In_90);
nand U3933 (N_3933,In_732,In_501);
or U3934 (N_3934,In_221,In_303);
and U3935 (N_3935,In_324,In_1900);
or U3936 (N_3936,In_376,In_613);
and U3937 (N_3937,In_1176,In_402);
nor U3938 (N_3938,In_1993,In_592);
nand U3939 (N_3939,In_646,In_676);
or U3940 (N_3940,In_1150,In_989);
nor U3941 (N_3941,In_1397,In_28);
nor U3942 (N_3942,In_359,In_1079);
xor U3943 (N_3943,In_913,In_232);
and U3944 (N_3944,In_727,In_1783);
and U3945 (N_3945,In_1048,In_703);
nor U3946 (N_3946,In_1118,In_964);
nand U3947 (N_3947,In_1389,In_1245);
and U3948 (N_3948,In_1701,In_1466);
or U3949 (N_3949,In_1597,In_503);
or U3950 (N_3950,In_681,In_692);
nor U3951 (N_3951,In_317,In_241);
nor U3952 (N_3952,In_770,In_508);
nand U3953 (N_3953,In_1641,In_732);
and U3954 (N_3954,In_1066,In_1717);
nor U3955 (N_3955,In_1181,In_100);
xor U3956 (N_3956,In_1360,In_1216);
and U3957 (N_3957,In_1740,In_1904);
or U3958 (N_3958,In_1290,In_214);
nand U3959 (N_3959,In_663,In_1163);
nor U3960 (N_3960,In_1534,In_1271);
or U3961 (N_3961,In_1441,In_1774);
or U3962 (N_3962,In_983,In_1842);
or U3963 (N_3963,In_1500,In_1979);
and U3964 (N_3964,In_602,In_1667);
nand U3965 (N_3965,In_784,In_1561);
or U3966 (N_3966,In_1515,In_1120);
or U3967 (N_3967,In_419,In_909);
nand U3968 (N_3968,In_427,In_152);
nor U3969 (N_3969,In_1108,In_462);
or U3970 (N_3970,In_1488,In_976);
nand U3971 (N_3971,In_1480,In_1944);
or U3972 (N_3972,In_1181,In_309);
nand U3973 (N_3973,In_499,In_1369);
or U3974 (N_3974,In_1108,In_1842);
nor U3975 (N_3975,In_1674,In_1907);
nand U3976 (N_3976,In_910,In_181);
nand U3977 (N_3977,In_281,In_811);
nor U3978 (N_3978,In_804,In_934);
xor U3979 (N_3979,In_922,In_1744);
xnor U3980 (N_3980,In_1433,In_168);
nor U3981 (N_3981,In_508,In_1147);
nor U3982 (N_3982,In_1164,In_90);
nand U3983 (N_3983,In_983,In_452);
nor U3984 (N_3984,In_445,In_1475);
xor U3985 (N_3985,In_703,In_701);
nor U3986 (N_3986,In_754,In_1812);
and U3987 (N_3987,In_1626,In_1581);
nand U3988 (N_3988,In_51,In_1936);
nor U3989 (N_3989,In_1736,In_1539);
xor U3990 (N_3990,In_354,In_946);
nor U3991 (N_3991,In_1707,In_452);
or U3992 (N_3992,In_1242,In_1542);
and U3993 (N_3993,In_769,In_1907);
nor U3994 (N_3994,In_889,In_1580);
or U3995 (N_3995,In_498,In_1196);
nand U3996 (N_3996,In_618,In_1251);
and U3997 (N_3997,In_1872,In_1569);
or U3998 (N_3998,In_1759,In_448);
nand U3999 (N_3999,In_844,In_873);
nor U4000 (N_4000,In_596,In_1074);
nand U4001 (N_4001,In_1858,In_697);
nor U4002 (N_4002,In_611,In_693);
nand U4003 (N_4003,In_295,In_1053);
and U4004 (N_4004,In_338,In_132);
nor U4005 (N_4005,In_305,In_1123);
xnor U4006 (N_4006,In_225,In_840);
and U4007 (N_4007,In_1007,In_227);
nand U4008 (N_4008,In_493,In_458);
or U4009 (N_4009,In_1328,In_139);
nor U4010 (N_4010,In_766,In_325);
nand U4011 (N_4011,In_1581,In_1318);
or U4012 (N_4012,In_1979,In_465);
and U4013 (N_4013,In_431,In_1606);
and U4014 (N_4014,In_54,In_478);
and U4015 (N_4015,In_650,In_1884);
or U4016 (N_4016,In_1200,In_1895);
xor U4017 (N_4017,In_1820,In_1517);
nand U4018 (N_4018,In_1543,In_1075);
nand U4019 (N_4019,In_785,In_1695);
and U4020 (N_4020,In_1936,In_678);
nand U4021 (N_4021,In_1509,In_1016);
and U4022 (N_4022,In_1923,In_404);
xnor U4023 (N_4023,In_131,In_337);
and U4024 (N_4024,In_431,In_188);
nor U4025 (N_4025,In_636,In_1370);
or U4026 (N_4026,In_1362,In_1886);
nand U4027 (N_4027,In_1516,In_402);
nor U4028 (N_4028,In_534,In_397);
nand U4029 (N_4029,In_1455,In_559);
nand U4030 (N_4030,In_1347,In_918);
nand U4031 (N_4031,In_676,In_279);
or U4032 (N_4032,In_768,In_556);
nor U4033 (N_4033,In_1215,In_1195);
or U4034 (N_4034,In_1462,In_139);
or U4035 (N_4035,In_614,In_1503);
and U4036 (N_4036,In_861,In_1851);
or U4037 (N_4037,In_912,In_701);
nor U4038 (N_4038,In_1755,In_1709);
or U4039 (N_4039,In_142,In_1724);
and U4040 (N_4040,In_863,In_1541);
xor U4041 (N_4041,In_902,In_1378);
nand U4042 (N_4042,In_540,In_1832);
nand U4043 (N_4043,In_738,In_171);
nand U4044 (N_4044,In_1988,In_1558);
nor U4045 (N_4045,In_758,In_1474);
or U4046 (N_4046,In_1313,In_570);
or U4047 (N_4047,In_1545,In_1076);
nand U4048 (N_4048,In_1261,In_1406);
or U4049 (N_4049,In_796,In_98);
and U4050 (N_4050,In_583,In_1942);
and U4051 (N_4051,In_856,In_601);
and U4052 (N_4052,In_233,In_1223);
and U4053 (N_4053,In_439,In_152);
or U4054 (N_4054,In_725,In_440);
or U4055 (N_4055,In_1529,In_301);
nor U4056 (N_4056,In_361,In_61);
and U4057 (N_4057,In_1882,In_633);
xnor U4058 (N_4058,In_929,In_33);
and U4059 (N_4059,In_896,In_994);
nor U4060 (N_4060,In_1797,In_1224);
and U4061 (N_4061,In_174,In_817);
nand U4062 (N_4062,In_1087,In_718);
nand U4063 (N_4063,In_766,In_526);
nand U4064 (N_4064,In_1923,In_1573);
or U4065 (N_4065,In_847,In_48);
nand U4066 (N_4066,In_1850,In_1508);
nand U4067 (N_4067,In_461,In_195);
or U4068 (N_4068,In_923,In_1140);
and U4069 (N_4069,In_444,In_459);
or U4070 (N_4070,In_1960,In_1144);
xor U4071 (N_4071,In_829,In_1327);
nor U4072 (N_4072,In_239,In_588);
nand U4073 (N_4073,In_1444,In_1508);
xor U4074 (N_4074,In_682,In_1918);
or U4075 (N_4075,In_654,In_358);
nand U4076 (N_4076,In_1217,In_1341);
nor U4077 (N_4077,In_1256,In_683);
and U4078 (N_4078,In_980,In_1196);
nand U4079 (N_4079,In_1788,In_449);
or U4080 (N_4080,In_583,In_25);
nand U4081 (N_4081,In_296,In_1445);
nor U4082 (N_4082,In_1374,In_687);
nor U4083 (N_4083,In_1995,In_683);
nor U4084 (N_4084,In_409,In_1882);
xnor U4085 (N_4085,In_448,In_1781);
nand U4086 (N_4086,In_923,In_292);
xnor U4087 (N_4087,In_464,In_208);
and U4088 (N_4088,In_212,In_1079);
nor U4089 (N_4089,In_1529,In_59);
and U4090 (N_4090,In_851,In_661);
nor U4091 (N_4091,In_804,In_1469);
and U4092 (N_4092,In_568,In_1063);
nor U4093 (N_4093,In_1775,In_1232);
nor U4094 (N_4094,In_1577,In_1239);
and U4095 (N_4095,In_879,In_1570);
or U4096 (N_4096,In_946,In_217);
nand U4097 (N_4097,In_1144,In_785);
xnor U4098 (N_4098,In_820,In_235);
nand U4099 (N_4099,In_518,In_700);
and U4100 (N_4100,In_763,In_1140);
xor U4101 (N_4101,In_1342,In_874);
nor U4102 (N_4102,In_1735,In_466);
nor U4103 (N_4103,In_973,In_1872);
and U4104 (N_4104,In_1662,In_1378);
and U4105 (N_4105,In_597,In_1449);
and U4106 (N_4106,In_1019,In_371);
and U4107 (N_4107,In_1493,In_36);
and U4108 (N_4108,In_1186,In_1822);
nand U4109 (N_4109,In_622,In_1267);
or U4110 (N_4110,In_1719,In_346);
and U4111 (N_4111,In_1457,In_96);
nor U4112 (N_4112,In_502,In_146);
nor U4113 (N_4113,In_1288,In_1781);
and U4114 (N_4114,In_88,In_606);
nand U4115 (N_4115,In_502,In_1218);
or U4116 (N_4116,In_567,In_1261);
nor U4117 (N_4117,In_742,In_1369);
nand U4118 (N_4118,In_1295,In_1929);
nor U4119 (N_4119,In_646,In_779);
or U4120 (N_4120,In_267,In_623);
nor U4121 (N_4121,In_109,In_1834);
or U4122 (N_4122,In_914,In_1902);
xnor U4123 (N_4123,In_1042,In_1337);
nor U4124 (N_4124,In_739,In_1274);
xnor U4125 (N_4125,In_985,In_1061);
and U4126 (N_4126,In_564,In_93);
and U4127 (N_4127,In_1983,In_358);
nand U4128 (N_4128,In_1420,In_1071);
or U4129 (N_4129,In_1458,In_1252);
nand U4130 (N_4130,In_1046,In_111);
and U4131 (N_4131,In_1830,In_696);
or U4132 (N_4132,In_741,In_1988);
nor U4133 (N_4133,In_59,In_498);
and U4134 (N_4134,In_1342,In_1457);
nand U4135 (N_4135,In_115,In_1363);
nand U4136 (N_4136,In_500,In_195);
or U4137 (N_4137,In_1418,In_887);
or U4138 (N_4138,In_1688,In_1043);
or U4139 (N_4139,In_1735,In_608);
or U4140 (N_4140,In_134,In_1341);
and U4141 (N_4141,In_634,In_80);
nand U4142 (N_4142,In_726,In_971);
nor U4143 (N_4143,In_1878,In_1536);
or U4144 (N_4144,In_1874,In_544);
xnor U4145 (N_4145,In_1993,In_191);
nand U4146 (N_4146,In_405,In_796);
nand U4147 (N_4147,In_1218,In_1137);
nor U4148 (N_4148,In_964,In_454);
and U4149 (N_4149,In_1928,In_33);
and U4150 (N_4150,In_366,In_1987);
and U4151 (N_4151,In_1531,In_1845);
or U4152 (N_4152,In_840,In_160);
and U4153 (N_4153,In_1314,In_1589);
and U4154 (N_4154,In_304,In_457);
nand U4155 (N_4155,In_851,In_914);
nor U4156 (N_4156,In_1809,In_342);
nand U4157 (N_4157,In_1865,In_1581);
nand U4158 (N_4158,In_848,In_122);
nor U4159 (N_4159,In_1030,In_635);
nor U4160 (N_4160,In_205,In_928);
and U4161 (N_4161,In_1910,In_920);
and U4162 (N_4162,In_470,In_498);
or U4163 (N_4163,In_1055,In_1199);
and U4164 (N_4164,In_1198,In_133);
and U4165 (N_4165,In_509,In_1831);
xnor U4166 (N_4166,In_1363,In_1656);
and U4167 (N_4167,In_1388,In_1692);
nand U4168 (N_4168,In_380,In_1780);
nand U4169 (N_4169,In_1891,In_1928);
nor U4170 (N_4170,In_1615,In_1373);
nand U4171 (N_4171,In_1651,In_1105);
xnor U4172 (N_4172,In_1845,In_1134);
and U4173 (N_4173,In_761,In_1318);
or U4174 (N_4174,In_633,In_1866);
nor U4175 (N_4175,In_1661,In_435);
nand U4176 (N_4176,In_1272,In_1047);
nor U4177 (N_4177,In_1304,In_966);
and U4178 (N_4178,In_1524,In_593);
nand U4179 (N_4179,In_839,In_960);
nand U4180 (N_4180,In_1293,In_1949);
or U4181 (N_4181,In_134,In_1611);
or U4182 (N_4182,In_671,In_455);
nor U4183 (N_4183,In_1437,In_734);
or U4184 (N_4184,In_516,In_1952);
nor U4185 (N_4185,In_82,In_708);
or U4186 (N_4186,In_732,In_1315);
nor U4187 (N_4187,In_597,In_1940);
or U4188 (N_4188,In_1595,In_789);
or U4189 (N_4189,In_1435,In_1174);
and U4190 (N_4190,In_53,In_1434);
nand U4191 (N_4191,In_736,In_708);
nand U4192 (N_4192,In_976,In_1832);
or U4193 (N_4193,In_1583,In_1331);
xnor U4194 (N_4194,In_1152,In_1993);
nor U4195 (N_4195,In_219,In_1338);
nand U4196 (N_4196,In_194,In_49);
nor U4197 (N_4197,In_1559,In_341);
or U4198 (N_4198,In_75,In_1962);
and U4199 (N_4199,In_25,In_1371);
nand U4200 (N_4200,In_448,In_1106);
and U4201 (N_4201,In_251,In_461);
nand U4202 (N_4202,In_1229,In_112);
or U4203 (N_4203,In_1550,In_1181);
and U4204 (N_4204,In_251,In_1980);
nor U4205 (N_4205,In_1380,In_555);
or U4206 (N_4206,In_1524,In_1975);
nor U4207 (N_4207,In_1332,In_1090);
and U4208 (N_4208,In_1437,In_171);
nor U4209 (N_4209,In_1377,In_687);
or U4210 (N_4210,In_888,In_1024);
nor U4211 (N_4211,In_84,In_1534);
and U4212 (N_4212,In_1481,In_1283);
nor U4213 (N_4213,In_1278,In_1093);
xor U4214 (N_4214,In_1561,In_1792);
nand U4215 (N_4215,In_1699,In_108);
or U4216 (N_4216,In_1654,In_1123);
nand U4217 (N_4217,In_116,In_1308);
nand U4218 (N_4218,In_515,In_451);
or U4219 (N_4219,In_1614,In_1539);
nor U4220 (N_4220,In_1689,In_1284);
nor U4221 (N_4221,In_217,In_959);
or U4222 (N_4222,In_1289,In_1073);
or U4223 (N_4223,In_1894,In_785);
or U4224 (N_4224,In_17,In_1817);
or U4225 (N_4225,In_1165,In_310);
and U4226 (N_4226,In_904,In_978);
nor U4227 (N_4227,In_385,In_1856);
or U4228 (N_4228,In_883,In_604);
nand U4229 (N_4229,In_1106,In_75);
nor U4230 (N_4230,In_453,In_367);
or U4231 (N_4231,In_1963,In_1725);
nor U4232 (N_4232,In_1122,In_984);
or U4233 (N_4233,In_1457,In_1876);
and U4234 (N_4234,In_1614,In_1817);
nor U4235 (N_4235,In_708,In_865);
nor U4236 (N_4236,In_1355,In_1511);
nand U4237 (N_4237,In_891,In_516);
xor U4238 (N_4238,In_579,In_113);
or U4239 (N_4239,In_241,In_1838);
nor U4240 (N_4240,In_1638,In_1009);
xor U4241 (N_4241,In_1172,In_1444);
or U4242 (N_4242,In_562,In_1498);
and U4243 (N_4243,In_1404,In_667);
and U4244 (N_4244,In_122,In_1798);
nand U4245 (N_4245,In_307,In_1873);
or U4246 (N_4246,In_1678,In_1698);
or U4247 (N_4247,In_158,In_889);
nor U4248 (N_4248,In_631,In_289);
and U4249 (N_4249,In_1436,In_594);
nand U4250 (N_4250,In_375,In_703);
or U4251 (N_4251,In_357,In_652);
nor U4252 (N_4252,In_1383,In_51);
or U4253 (N_4253,In_205,In_134);
nand U4254 (N_4254,In_937,In_1802);
nor U4255 (N_4255,In_841,In_241);
or U4256 (N_4256,In_810,In_56);
or U4257 (N_4257,In_1874,In_1701);
and U4258 (N_4258,In_548,In_1415);
and U4259 (N_4259,In_387,In_1322);
nor U4260 (N_4260,In_541,In_1742);
nor U4261 (N_4261,In_1607,In_1719);
nand U4262 (N_4262,In_1009,In_945);
nor U4263 (N_4263,In_773,In_1436);
nor U4264 (N_4264,In_1471,In_963);
nor U4265 (N_4265,In_283,In_904);
nor U4266 (N_4266,In_216,In_1835);
nor U4267 (N_4267,In_1149,In_1395);
and U4268 (N_4268,In_1927,In_745);
or U4269 (N_4269,In_1350,In_900);
and U4270 (N_4270,In_1058,In_1466);
xor U4271 (N_4271,In_1881,In_21);
nor U4272 (N_4272,In_727,In_1232);
and U4273 (N_4273,In_981,In_1658);
and U4274 (N_4274,In_1863,In_157);
nor U4275 (N_4275,In_1940,In_1626);
or U4276 (N_4276,In_1831,In_1436);
xor U4277 (N_4277,In_915,In_861);
or U4278 (N_4278,In_1318,In_1826);
or U4279 (N_4279,In_1143,In_73);
and U4280 (N_4280,In_1763,In_605);
nand U4281 (N_4281,In_467,In_1908);
or U4282 (N_4282,In_1842,In_927);
or U4283 (N_4283,In_681,In_1071);
nor U4284 (N_4284,In_1712,In_1127);
nor U4285 (N_4285,In_634,In_1779);
nand U4286 (N_4286,In_1556,In_775);
nor U4287 (N_4287,In_444,In_102);
and U4288 (N_4288,In_404,In_551);
or U4289 (N_4289,In_1332,In_775);
nor U4290 (N_4290,In_543,In_1837);
or U4291 (N_4291,In_1241,In_92);
nor U4292 (N_4292,In_1368,In_371);
or U4293 (N_4293,In_1762,In_1946);
nand U4294 (N_4294,In_37,In_1940);
or U4295 (N_4295,In_1349,In_976);
or U4296 (N_4296,In_327,In_1139);
nand U4297 (N_4297,In_1304,In_413);
and U4298 (N_4298,In_949,In_897);
or U4299 (N_4299,In_902,In_377);
nand U4300 (N_4300,In_1070,In_1220);
or U4301 (N_4301,In_741,In_1339);
nor U4302 (N_4302,In_98,In_895);
nand U4303 (N_4303,In_460,In_1024);
or U4304 (N_4304,In_762,In_1403);
and U4305 (N_4305,In_246,In_312);
nand U4306 (N_4306,In_1281,In_640);
and U4307 (N_4307,In_1279,In_412);
xor U4308 (N_4308,In_1524,In_425);
and U4309 (N_4309,In_796,In_1266);
nor U4310 (N_4310,In_1647,In_406);
nor U4311 (N_4311,In_1788,In_503);
nand U4312 (N_4312,In_145,In_1865);
or U4313 (N_4313,In_383,In_1374);
xnor U4314 (N_4314,In_1592,In_1762);
nand U4315 (N_4315,In_538,In_1877);
xor U4316 (N_4316,In_275,In_93);
or U4317 (N_4317,In_913,In_1817);
nand U4318 (N_4318,In_1568,In_645);
nand U4319 (N_4319,In_1257,In_535);
and U4320 (N_4320,In_365,In_1838);
xor U4321 (N_4321,In_78,In_1992);
or U4322 (N_4322,In_1010,In_1987);
nor U4323 (N_4323,In_1467,In_1984);
nor U4324 (N_4324,In_1774,In_1734);
nand U4325 (N_4325,In_367,In_499);
nor U4326 (N_4326,In_1786,In_1175);
or U4327 (N_4327,In_480,In_1629);
nor U4328 (N_4328,In_1385,In_1151);
nor U4329 (N_4329,In_1477,In_1654);
or U4330 (N_4330,In_121,In_568);
nor U4331 (N_4331,In_435,In_1078);
xnor U4332 (N_4332,In_841,In_614);
nand U4333 (N_4333,In_1404,In_957);
nand U4334 (N_4334,In_1011,In_1765);
nand U4335 (N_4335,In_842,In_873);
and U4336 (N_4336,In_1221,In_1416);
xnor U4337 (N_4337,In_1817,In_1260);
nand U4338 (N_4338,In_1562,In_851);
nor U4339 (N_4339,In_1708,In_738);
and U4340 (N_4340,In_997,In_1094);
nand U4341 (N_4341,In_118,In_1583);
nand U4342 (N_4342,In_251,In_1181);
nor U4343 (N_4343,In_520,In_124);
and U4344 (N_4344,In_1526,In_1281);
nor U4345 (N_4345,In_1645,In_1805);
and U4346 (N_4346,In_931,In_841);
and U4347 (N_4347,In_729,In_1448);
and U4348 (N_4348,In_1168,In_1023);
nand U4349 (N_4349,In_218,In_82);
and U4350 (N_4350,In_300,In_1133);
or U4351 (N_4351,In_327,In_1361);
or U4352 (N_4352,In_1553,In_1232);
nor U4353 (N_4353,In_1876,In_982);
nand U4354 (N_4354,In_39,In_3);
and U4355 (N_4355,In_248,In_407);
nor U4356 (N_4356,In_672,In_975);
and U4357 (N_4357,In_7,In_1113);
and U4358 (N_4358,In_137,In_1020);
xor U4359 (N_4359,In_318,In_1564);
and U4360 (N_4360,In_1491,In_1899);
nand U4361 (N_4361,In_331,In_1411);
and U4362 (N_4362,In_1702,In_1604);
or U4363 (N_4363,In_610,In_1374);
nand U4364 (N_4364,In_769,In_1564);
nand U4365 (N_4365,In_730,In_1272);
nor U4366 (N_4366,In_1232,In_1923);
xnor U4367 (N_4367,In_916,In_1293);
nor U4368 (N_4368,In_854,In_1371);
nor U4369 (N_4369,In_1859,In_731);
nor U4370 (N_4370,In_579,In_627);
or U4371 (N_4371,In_977,In_1121);
and U4372 (N_4372,In_1516,In_308);
xnor U4373 (N_4373,In_1138,In_625);
and U4374 (N_4374,In_560,In_708);
and U4375 (N_4375,In_1952,In_1116);
nor U4376 (N_4376,In_1729,In_1766);
nor U4377 (N_4377,In_1151,In_1508);
nand U4378 (N_4378,In_111,In_1167);
or U4379 (N_4379,In_1132,In_660);
nor U4380 (N_4380,In_415,In_861);
nand U4381 (N_4381,In_929,In_1933);
and U4382 (N_4382,In_78,In_1562);
or U4383 (N_4383,In_125,In_1172);
nand U4384 (N_4384,In_1068,In_925);
and U4385 (N_4385,In_1138,In_1332);
nor U4386 (N_4386,In_670,In_585);
or U4387 (N_4387,In_21,In_1720);
nand U4388 (N_4388,In_1275,In_1654);
nor U4389 (N_4389,In_1656,In_1924);
nor U4390 (N_4390,In_680,In_1555);
and U4391 (N_4391,In_264,In_440);
and U4392 (N_4392,In_1815,In_1686);
nor U4393 (N_4393,In_732,In_1621);
and U4394 (N_4394,In_1673,In_646);
nor U4395 (N_4395,In_195,In_859);
nand U4396 (N_4396,In_31,In_452);
or U4397 (N_4397,In_430,In_1284);
xor U4398 (N_4398,In_76,In_1069);
nor U4399 (N_4399,In_1496,In_1161);
xor U4400 (N_4400,In_766,In_906);
nor U4401 (N_4401,In_179,In_1479);
nand U4402 (N_4402,In_1506,In_29);
and U4403 (N_4403,In_1996,In_772);
or U4404 (N_4404,In_591,In_1769);
or U4405 (N_4405,In_1493,In_215);
nor U4406 (N_4406,In_1096,In_1711);
xnor U4407 (N_4407,In_1284,In_586);
nor U4408 (N_4408,In_345,In_860);
or U4409 (N_4409,In_70,In_1972);
nand U4410 (N_4410,In_1495,In_573);
or U4411 (N_4411,In_1155,In_1688);
nor U4412 (N_4412,In_1522,In_835);
nor U4413 (N_4413,In_865,In_440);
nor U4414 (N_4414,In_677,In_153);
nand U4415 (N_4415,In_1690,In_712);
nor U4416 (N_4416,In_1257,In_1463);
and U4417 (N_4417,In_814,In_1589);
nand U4418 (N_4418,In_252,In_1314);
nor U4419 (N_4419,In_83,In_1425);
nor U4420 (N_4420,In_361,In_389);
and U4421 (N_4421,In_645,In_895);
and U4422 (N_4422,In_218,In_1797);
nor U4423 (N_4423,In_1325,In_1798);
xnor U4424 (N_4424,In_1681,In_693);
nor U4425 (N_4425,In_950,In_1405);
xor U4426 (N_4426,In_1255,In_1625);
nand U4427 (N_4427,In_1931,In_1864);
nor U4428 (N_4428,In_993,In_392);
xnor U4429 (N_4429,In_578,In_1635);
nor U4430 (N_4430,In_1614,In_1033);
nor U4431 (N_4431,In_1740,In_967);
or U4432 (N_4432,In_147,In_1703);
and U4433 (N_4433,In_275,In_813);
nand U4434 (N_4434,In_827,In_1523);
and U4435 (N_4435,In_1302,In_713);
nand U4436 (N_4436,In_895,In_875);
nand U4437 (N_4437,In_604,In_1629);
nand U4438 (N_4438,In_31,In_965);
nand U4439 (N_4439,In_1991,In_404);
or U4440 (N_4440,In_935,In_180);
or U4441 (N_4441,In_1740,In_692);
nor U4442 (N_4442,In_1483,In_983);
or U4443 (N_4443,In_1513,In_957);
nand U4444 (N_4444,In_152,In_40);
and U4445 (N_4445,In_1038,In_1326);
nand U4446 (N_4446,In_595,In_975);
or U4447 (N_4447,In_1453,In_204);
or U4448 (N_4448,In_1103,In_64);
nor U4449 (N_4449,In_884,In_860);
nor U4450 (N_4450,In_629,In_960);
and U4451 (N_4451,In_1870,In_1077);
nand U4452 (N_4452,In_1431,In_390);
and U4453 (N_4453,In_547,In_484);
and U4454 (N_4454,In_1464,In_1796);
xnor U4455 (N_4455,In_1283,In_274);
and U4456 (N_4456,In_537,In_42);
nand U4457 (N_4457,In_1018,In_663);
and U4458 (N_4458,In_596,In_1040);
and U4459 (N_4459,In_1390,In_127);
and U4460 (N_4460,In_1806,In_226);
and U4461 (N_4461,In_1053,In_161);
xor U4462 (N_4462,In_1687,In_578);
and U4463 (N_4463,In_396,In_1179);
nand U4464 (N_4464,In_1930,In_705);
or U4465 (N_4465,In_973,In_1052);
or U4466 (N_4466,In_729,In_1440);
nor U4467 (N_4467,In_1928,In_1205);
xor U4468 (N_4468,In_1420,In_1316);
or U4469 (N_4469,In_1335,In_350);
nor U4470 (N_4470,In_80,In_172);
and U4471 (N_4471,In_429,In_875);
or U4472 (N_4472,In_411,In_1993);
nor U4473 (N_4473,In_1706,In_11);
and U4474 (N_4474,In_718,In_207);
nand U4475 (N_4475,In_401,In_1959);
or U4476 (N_4476,In_484,In_1008);
xnor U4477 (N_4477,In_198,In_1593);
nand U4478 (N_4478,In_824,In_1210);
and U4479 (N_4479,In_1643,In_1247);
nor U4480 (N_4480,In_36,In_1971);
and U4481 (N_4481,In_1945,In_1689);
and U4482 (N_4482,In_1415,In_256);
and U4483 (N_4483,In_366,In_1741);
and U4484 (N_4484,In_176,In_50);
xnor U4485 (N_4485,In_328,In_1407);
and U4486 (N_4486,In_1067,In_1057);
nand U4487 (N_4487,In_1418,In_1508);
and U4488 (N_4488,In_1132,In_1289);
or U4489 (N_4489,In_1603,In_297);
and U4490 (N_4490,In_569,In_861);
nand U4491 (N_4491,In_1909,In_1071);
nor U4492 (N_4492,In_309,In_1598);
nor U4493 (N_4493,In_1454,In_1417);
nand U4494 (N_4494,In_587,In_223);
xnor U4495 (N_4495,In_423,In_829);
or U4496 (N_4496,In_1067,In_593);
or U4497 (N_4497,In_1781,In_797);
nand U4498 (N_4498,In_183,In_322);
nand U4499 (N_4499,In_396,In_786);
xnor U4500 (N_4500,In_994,In_469);
xnor U4501 (N_4501,In_418,In_1018);
nor U4502 (N_4502,In_1325,In_261);
nor U4503 (N_4503,In_1960,In_512);
or U4504 (N_4504,In_1559,In_1584);
or U4505 (N_4505,In_74,In_786);
nand U4506 (N_4506,In_1481,In_1307);
nand U4507 (N_4507,In_772,In_822);
nand U4508 (N_4508,In_1459,In_493);
nand U4509 (N_4509,In_1657,In_446);
and U4510 (N_4510,In_12,In_1412);
nand U4511 (N_4511,In_56,In_220);
nor U4512 (N_4512,In_793,In_1581);
nor U4513 (N_4513,In_1378,In_618);
nand U4514 (N_4514,In_95,In_1599);
xnor U4515 (N_4515,In_759,In_1164);
nand U4516 (N_4516,In_40,In_1277);
nor U4517 (N_4517,In_1935,In_1708);
nand U4518 (N_4518,In_223,In_1391);
nor U4519 (N_4519,In_825,In_1368);
nor U4520 (N_4520,In_1608,In_915);
and U4521 (N_4521,In_1337,In_13);
nand U4522 (N_4522,In_1110,In_1601);
nor U4523 (N_4523,In_1413,In_1183);
and U4524 (N_4524,In_1450,In_1209);
or U4525 (N_4525,In_1430,In_937);
or U4526 (N_4526,In_1035,In_1472);
xnor U4527 (N_4527,In_1280,In_248);
nor U4528 (N_4528,In_140,In_1464);
nor U4529 (N_4529,In_555,In_1978);
nand U4530 (N_4530,In_1108,In_1266);
and U4531 (N_4531,In_1366,In_641);
or U4532 (N_4532,In_1599,In_86);
nand U4533 (N_4533,In_544,In_620);
or U4534 (N_4534,In_703,In_615);
nand U4535 (N_4535,In_49,In_120);
xor U4536 (N_4536,In_1884,In_1431);
nor U4537 (N_4537,In_1126,In_876);
nand U4538 (N_4538,In_265,In_1922);
or U4539 (N_4539,In_1224,In_1324);
nand U4540 (N_4540,In_1173,In_495);
and U4541 (N_4541,In_1349,In_715);
nand U4542 (N_4542,In_1249,In_1505);
and U4543 (N_4543,In_65,In_1123);
and U4544 (N_4544,In_1550,In_144);
or U4545 (N_4545,In_504,In_781);
nand U4546 (N_4546,In_309,In_741);
or U4547 (N_4547,In_1018,In_1781);
or U4548 (N_4548,In_188,In_1055);
or U4549 (N_4549,In_1189,In_1237);
nand U4550 (N_4550,In_94,In_1758);
and U4551 (N_4551,In_752,In_105);
nand U4552 (N_4552,In_375,In_68);
nand U4553 (N_4553,In_229,In_1708);
and U4554 (N_4554,In_650,In_207);
or U4555 (N_4555,In_265,In_1335);
or U4556 (N_4556,In_1047,In_421);
and U4557 (N_4557,In_34,In_263);
or U4558 (N_4558,In_1319,In_430);
and U4559 (N_4559,In_346,In_994);
and U4560 (N_4560,In_774,In_361);
xnor U4561 (N_4561,In_8,In_97);
nor U4562 (N_4562,In_528,In_1816);
and U4563 (N_4563,In_1601,In_397);
and U4564 (N_4564,In_476,In_1369);
and U4565 (N_4565,In_1948,In_18);
and U4566 (N_4566,In_184,In_911);
and U4567 (N_4567,In_112,In_1339);
nor U4568 (N_4568,In_1706,In_1380);
or U4569 (N_4569,In_1015,In_641);
xor U4570 (N_4570,In_1455,In_581);
nor U4571 (N_4571,In_1331,In_1322);
and U4572 (N_4572,In_720,In_71);
nor U4573 (N_4573,In_1646,In_1928);
xnor U4574 (N_4574,In_1849,In_548);
nor U4575 (N_4575,In_118,In_1197);
or U4576 (N_4576,In_912,In_1063);
nor U4577 (N_4577,In_471,In_327);
or U4578 (N_4578,In_697,In_1305);
and U4579 (N_4579,In_1790,In_1546);
nand U4580 (N_4580,In_115,In_578);
and U4581 (N_4581,In_1810,In_1412);
nand U4582 (N_4582,In_793,In_724);
or U4583 (N_4583,In_1160,In_1409);
xor U4584 (N_4584,In_1338,In_1320);
and U4585 (N_4585,In_293,In_1448);
nor U4586 (N_4586,In_871,In_1815);
nor U4587 (N_4587,In_832,In_1538);
nor U4588 (N_4588,In_1007,In_134);
nand U4589 (N_4589,In_132,In_1348);
nor U4590 (N_4590,In_1022,In_550);
nor U4591 (N_4591,In_913,In_1044);
and U4592 (N_4592,In_404,In_1870);
and U4593 (N_4593,In_1579,In_1494);
nor U4594 (N_4594,In_1181,In_542);
or U4595 (N_4595,In_1881,In_1812);
and U4596 (N_4596,In_1188,In_1043);
or U4597 (N_4597,In_968,In_1996);
and U4598 (N_4598,In_1083,In_1876);
nand U4599 (N_4599,In_1062,In_739);
or U4600 (N_4600,In_443,In_1452);
or U4601 (N_4601,In_1963,In_1116);
nand U4602 (N_4602,In_951,In_30);
nor U4603 (N_4603,In_1779,In_612);
nand U4604 (N_4604,In_1029,In_507);
and U4605 (N_4605,In_1816,In_1978);
and U4606 (N_4606,In_125,In_579);
and U4607 (N_4607,In_392,In_1292);
and U4608 (N_4608,In_648,In_878);
and U4609 (N_4609,In_1609,In_824);
xor U4610 (N_4610,In_1596,In_1989);
or U4611 (N_4611,In_1005,In_1347);
or U4612 (N_4612,In_1750,In_960);
nand U4613 (N_4613,In_918,In_1319);
xnor U4614 (N_4614,In_1621,In_954);
nand U4615 (N_4615,In_1812,In_1016);
and U4616 (N_4616,In_1831,In_528);
xor U4617 (N_4617,In_1840,In_775);
or U4618 (N_4618,In_886,In_111);
nand U4619 (N_4619,In_445,In_1216);
and U4620 (N_4620,In_557,In_1779);
nor U4621 (N_4621,In_1914,In_1746);
or U4622 (N_4622,In_1575,In_823);
nor U4623 (N_4623,In_760,In_745);
and U4624 (N_4624,In_834,In_1467);
or U4625 (N_4625,In_102,In_865);
xor U4626 (N_4626,In_1284,In_1104);
nor U4627 (N_4627,In_818,In_1473);
nor U4628 (N_4628,In_608,In_537);
or U4629 (N_4629,In_1517,In_1493);
or U4630 (N_4630,In_1250,In_1788);
and U4631 (N_4631,In_1793,In_1707);
xnor U4632 (N_4632,In_1057,In_1514);
xnor U4633 (N_4633,In_662,In_1204);
and U4634 (N_4634,In_1637,In_279);
nand U4635 (N_4635,In_125,In_1091);
and U4636 (N_4636,In_1580,In_915);
nand U4637 (N_4637,In_822,In_1604);
and U4638 (N_4638,In_992,In_289);
xor U4639 (N_4639,In_1619,In_711);
nor U4640 (N_4640,In_1353,In_957);
or U4641 (N_4641,In_1495,In_763);
nand U4642 (N_4642,In_965,In_184);
nor U4643 (N_4643,In_758,In_907);
and U4644 (N_4644,In_483,In_1042);
or U4645 (N_4645,In_523,In_1773);
and U4646 (N_4646,In_259,In_268);
nand U4647 (N_4647,In_1953,In_1692);
and U4648 (N_4648,In_1683,In_170);
and U4649 (N_4649,In_970,In_135);
or U4650 (N_4650,In_976,In_490);
xnor U4651 (N_4651,In_929,In_1033);
nand U4652 (N_4652,In_238,In_1857);
nor U4653 (N_4653,In_174,In_1832);
or U4654 (N_4654,In_1994,In_311);
and U4655 (N_4655,In_1376,In_1694);
nand U4656 (N_4656,In_158,In_1407);
nor U4657 (N_4657,In_668,In_236);
xnor U4658 (N_4658,In_1632,In_1042);
or U4659 (N_4659,In_1472,In_983);
or U4660 (N_4660,In_1164,In_835);
nor U4661 (N_4661,In_763,In_1005);
and U4662 (N_4662,In_1160,In_1997);
nand U4663 (N_4663,In_230,In_1956);
and U4664 (N_4664,In_1268,In_271);
xnor U4665 (N_4665,In_448,In_1229);
nor U4666 (N_4666,In_540,In_165);
or U4667 (N_4667,In_1787,In_1618);
xnor U4668 (N_4668,In_337,In_1702);
and U4669 (N_4669,In_1000,In_1635);
nand U4670 (N_4670,In_747,In_1413);
and U4671 (N_4671,In_1660,In_937);
xor U4672 (N_4672,In_1145,In_1982);
or U4673 (N_4673,In_1622,In_754);
or U4674 (N_4674,In_595,In_1194);
nand U4675 (N_4675,In_906,In_392);
nand U4676 (N_4676,In_1404,In_972);
nand U4677 (N_4677,In_1375,In_509);
and U4678 (N_4678,In_623,In_309);
or U4679 (N_4679,In_1928,In_1406);
and U4680 (N_4680,In_1010,In_1379);
or U4681 (N_4681,In_562,In_479);
or U4682 (N_4682,In_196,In_603);
nor U4683 (N_4683,In_617,In_1557);
and U4684 (N_4684,In_1829,In_625);
xnor U4685 (N_4685,In_1577,In_951);
xor U4686 (N_4686,In_1019,In_474);
xnor U4687 (N_4687,In_1397,In_1579);
and U4688 (N_4688,In_1374,In_901);
nand U4689 (N_4689,In_238,In_126);
and U4690 (N_4690,In_1098,In_795);
nand U4691 (N_4691,In_149,In_643);
and U4692 (N_4692,In_1224,In_1375);
nor U4693 (N_4693,In_681,In_1941);
nor U4694 (N_4694,In_1285,In_1692);
and U4695 (N_4695,In_27,In_550);
nor U4696 (N_4696,In_1186,In_1462);
or U4697 (N_4697,In_382,In_860);
or U4698 (N_4698,In_538,In_1309);
xor U4699 (N_4699,In_963,In_196);
and U4700 (N_4700,In_1099,In_540);
nand U4701 (N_4701,In_1611,In_893);
or U4702 (N_4702,In_1025,In_811);
nor U4703 (N_4703,In_1868,In_1634);
or U4704 (N_4704,In_328,In_189);
xor U4705 (N_4705,In_1972,In_824);
nor U4706 (N_4706,In_841,In_1169);
or U4707 (N_4707,In_1052,In_341);
or U4708 (N_4708,In_1219,In_1077);
or U4709 (N_4709,In_1028,In_1835);
nand U4710 (N_4710,In_1200,In_564);
nor U4711 (N_4711,In_1640,In_111);
nand U4712 (N_4712,In_1633,In_404);
nor U4713 (N_4713,In_988,In_1280);
nor U4714 (N_4714,In_1544,In_508);
or U4715 (N_4715,In_7,In_19);
nand U4716 (N_4716,In_1939,In_1159);
or U4717 (N_4717,In_1937,In_1873);
nand U4718 (N_4718,In_1710,In_1759);
nor U4719 (N_4719,In_1493,In_1929);
and U4720 (N_4720,In_760,In_721);
or U4721 (N_4721,In_456,In_965);
or U4722 (N_4722,In_1747,In_799);
nand U4723 (N_4723,In_364,In_323);
nor U4724 (N_4724,In_400,In_1120);
and U4725 (N_4725,In_1576,In_1821);
nor U4726 (N_4726,In_1436,In_1350);
or U4727 (N_4727,In_1113,In_1118);
and U4728 (N_4728,In_1740,In_1907);
and U4729 (N_4729,In_670,In_766);
nor U4730 (N_4730,In_893,In_58);
and U4731 (N_4731,In_207,In_529);
nand U4732 (N_4732,In_913,In_1535);
xor U4733 (N_4733,In_370,In_1173);
and U4734 (N_4734,In_1342,In_1117);
nand U4735 (N_4735,In_905,In_1573);
or U4736 (N_4736,In_200,In_970);
nor U4737 (N_4737,In_1403,In_1127);
nor U4738 (N_4738,In_1644,In_1233);
nor U4739 (N_4739,In_1625,In_1279);
or U4740 (N_4740,In_1818,In_1136);
nor U4741 (N_4741,In_185,In_736);
and U4742 (N_4742,In_738,In_1916);
or U4743 (N_4743,In_59,In_1303);
or U4744 (N_4744,In_888,In_709);
or U4745 (N_4745,In_810,In_726);
or U4746 (N_4746,In_54,In_469);
and U4747 (N_4747,In_1743,In_1354);
nor U4748 (N_4748,In_1215,In_1063);
and U4749 (N_4749,In_324,In_225);
or U4750 (N_4750,In_1720,In_1742);
or U4751 (N_4751,In_1232,In_652);
nor U4752 (N_4752,In_731,In_1529);
nor U4753 (N_4753,In_808,In_1919);
nor U4754 (N_4754,In_1956,In_910);
nor U4755 (N_4755,In_1415,In_732);
or U4756 (N_4756,In_1831,In_442);
or U4757 (N_4757,In_1069,In_1571);
and U4758 (N_4758,In_392,In_1037);
and U4759 (N_4759,In_1378,In_1866);
xor U4760 (N_4760,In_864,In_481);
nor U4761 (N_4761,In_1837,In_1233);
and U4762 (N_4762,In_766,In_1618);
nor U4763 (N_4763,In_836,In_1470);
nand U4764 (N_4764,In_91,In_1789);
or U4765 (N_4765,In_410,In_372);
xnor U4766 (N_4766,In_1391,In_188);
and U4767 (N_4767,In_726,In_1010);
and U4768 (N_4768,In_245,In_1150);
and U4769 (N_4769,In_628,In_400);
or U4770 (N_4770,In_947,In_231);
nor U4771 (N_4771,In_439,In_1793);
or U4772 (N_4772,In_1487,In_527);
nand U4773 (N_4773,In_947,In_948);
or U4774 (N_4774,In_615,In_839);
nand U4775 (N_4775,In_1831,In_953);
and U4776 (N_4776,In_1913,In_714);
nand U4777 (N_4777,In_148,In_57);
nand U4778 (N_4778,In_281,In_949);
and U4779 (N_4779,In_804,In_298);
or U4780 (N_4780,In_700,In_1609);
nand U4781 (N_4781,In_1311,In_1182);
nor U4782 (N_4782,In_1512,In_1210);
nand U4783 (N_4783,In_628,In_1461);
nor U4784 (N_4784,In_246,In_1299);
and U4785 (N_4785,In_905,In_1787);
xor U4786 (N_4786,In_1027,In_648);
or U4787 (N_4787,In_666,In_701);
or U4788 (N_4788,In_1434,In_446);
nor U4789 (N_4789,In_447,In_1369);
nor U4790 (N_4790,In_1466,In_1287);
xnor U4791 (N_4791,In_113,In_139);
nand U4792 (N_4792,In_1938,In_1407);
and U4793 (N_4793,In_350,In_1183);
and U4794 (N_4794,In_1163,In_411);
nand U4795 (N_4795,In_1300,In_1386);
nand U4796 (N_4796,In_1221,In_15);
xor U4797 (N_4797,In_1282,In_884);
nand U4798 (N_4798,In_1497,In_370);
and U4799 (N_4799,In_930,In_1025);
nor U4800 (N_4800,In_683,In_1993);
nor U4801 (N_4801,In_519,In_98);
nor U4802 (N_4802,In_1098,In_1186);
and U4803 (N_4803,In_1033,In_429);
nor U4804 (N_4804,In_1184,In_999);
and U4805 (N_4805,In_777,In_178);
and U4806 (N_4806,In_1814,In_25);
nand U4807 (N_4807,In_808,In_299);
or U4808 (N_4808,In_1605,In_1038);
nand U4809 (N_4809,In_11,In_1214);
nand U4810 (N_4810,In_996,In_200);
and U4811 (N_4811,In_1498,In_1603);
or U4812 (N_4812,In_727,In_1861);
xnor U4813 (N_4813,In_1774,In_79);
and U4814 (N_4814,In_1883,In_727);
and U4815 (N_4815,In_1102,In_1377);
nor U4816 (N_4816,In_1988,In_160);
or U4817 (N_4817,In_954,In_231);
xnor U4818 (N_4818,In_10,In_1917);
nor U4819 (N_4819,In_1846,In_953);
and U4820 (N_4820,In_881,In_272);
nor U4821 (N_4821,In_768,In_1306);
xnor U4822 (N_4822,In_1352,In_652);
nor U4823 (N_4823,In_1023,In_628);
xnor U4824 (N_4824,In_1951,In_1700);
or U4825 (N_4825,In_957,In_74);
nand U4826 (N_4826,In_250,In_853);
nor U4827 (N_4827,In_1570,In_142);
nor U4828 (N_4828,In_56,In_991);
nand U4829 (N_4829,In_658,In_1067);
or U4830 (N_4830,In_572,In_1422);
nand U4831 (N_4831,In_1601,In_704);
nor U4832 (N_4832,In_637,In_1808);
nand U4833 (N_4833,In_133,In_153);
nand U4834 (N_4834,In_764,In_1440);
or U4835 (N_4835,In_1378,In_932);
or U4836 (N_4836,In_7,In_1066);
or U4837 (N_4837,In_1124,In_184);
xnor U4838 (N_4838,In_801,In_600);
and U4839 (N_4839,In_1550,In_1397);
and U4840 (N_4840,In_293,In_1551);
nor U4841 (N_4841,In_19,In_1408);
or U4842 (N_4842,In_1093,In_1376);
xor U4843 (N_4843,In_819,In_1752);
nor U4844 (N_4844,In_872,In_89);
or U4845 (N_4845,In_1752,In_1252);
nand U4846 (N_4846,In_1630,In_1641);
nor U4847 (N_4847,In_1100,In_264);
nand U4848 (N_4848,In_1108,In_1820);
or U4849 (N_4849,In_416,In_1944);
or U4850 (N_4850,In_1526,In_1411);
or U4851 (N_4851,In_1998,In_1991);
nor U4852 (N_4852,In_1563,In_670);
and U4853 (N_4853,In_1819,In_24);
nand U4854 (N_4854,In_1690,In_126);
and U4855 (N_4855,In_1048,In_1498);
nand U4856 (N_4856,In_1254,In_1143);
and U4857 (N_4857,In_424,In_1839);
and U4858 (N_4858,In_685,In_1419);
and U4859 (N_4859,In_1436,In_73);
xor U4860 (N_4860,In_635,In_1072);
and U4861 (N_4861,In_1447,In_759);
nor U4862 (N_4862,In_939,In_1642);
xor U4863 (N_4863,In_280,In_1635);
nor U4864 (N_4864,In_1407,In_1484);
and U4865 (N_4865,In_1471,In_866);
nand U4866 (N_4866,In_293,In_903);
nor U4867 (N_4867,In_1407,In_1007);
xnor U4868 (N_4868,In_1410,In_1062);
and U4869 (N_4869,In_1090,In_1306);
and U4870 (N_4870,In_689,In_1124);
nor U4871 (N_4871,In_1922,In_1779);
nand U4872 (N_4872,In_1192,In_290);
and U4873 (N_4873,In_1235,In_125);
nor U4874 (N_4874,In_1689,In_936);
nand U4875 (N_4875,In_1954,In_226);
nand U4876 (N_4876,In_971,In_1591);
nor U4877 (N_4877,In_587,In_1581);
nand U4878 (N_4878,In_688,In_1371);
nand U4879 (N_4879,In_256,In_73);
or U4880 (N_4880,In_1723,In_1612);
or U4881 (N_4881,In_187,In_136);
and U4882 (N_4882,In_982,In_442);
nor U4883 (N_4883,In_1832,In_1029);
nand U4884 (N_4884,In_1843,In_1360);
nor U4885 (N_4885,In_252,In_1145);
nand U4886 (N_4886,In_604,In_1690);
xor U4887 (N_4887,In_1772,In_756);
nand U4888 (N_4888,In_206,In_1289);
xnor U4889 (N_4889,In_554,In_1375);
nand U4890 (N_4890,In_1590,In_873);
or U4891 (N_4891,In_244,In_1934);
and U4892 (N_4892,In_1845,In_1143);
nand U4893 (N_4893,In_1757,In_95);
nand U4894 (N_4894,In_420,In_1754);
nand U4895 (N_4895,In_144,In_1496);
or U4896 (N_4896,In_1093,In_1378);
and U4897 (N_4897,In_1017,In_409);
or U4898 (N_4898,In_154,In_1237);
or U4899 (N_4899,In_847,In_352);
nand U4900 (N_4900,In_311,In_1657);
xnor U4901 (N_4901,In_263,In_1649);
nor U4902 (N_4902,In_1450,In_490);
nor U4903 (N_4903,In_522,In_572);
or U4904 (N_4904,In_395,In_1152);
or U4905 (N_4905,In_1196,In_1071);
nor U4906 (N_4906,In_864,In_1459);
or U4907 (N_4907,In_11,In_1428);
nor U4908 (N_4908,In_579,In_1625);
and U4909 (N_4909,In_180,In_1628);
nand U4910 (N_4910,In_965,In_66);
nand U4911 (N_4911,In_960,In_229);
nand U4912 (N_4912,In_1107,In_1250);
or U4913 (N_4913,In_1269,In_281);
or U4914 (N_4914,In_1909,In_1455);
nand U4915 (N_4915,In_846,In_1286);
and U4916 (N_4916,In_908,In_846);
nor U4917 (N_4917,In_1405,In_1460);
nor U4918 (N_4918,In_902,In_1181);
nor U4919 (N_4919,In_1038,In_1015);
nand U4920 (N_4920,In_550,In_20);
and U4921 (N_4921,In_220,In_1086);
xnor U4922 (N_4922,In_6,In_746);
nand U4923 (N_4923,In_0,In_1286);
nor U4924 (N_4924,In_1442,In_613);
or U4925 (N_4925,In_250,In_241);
nor U4926 (N_4926,In_460,In_1851);
or U4927 (N_4927,In_340,In_963);
or U4928 (N_4928,In_1285,In_99);
nor U4929 (N_4929,In_494,In_863);
nand U4930 (N_4930,In_1317,In_897);
and U4931 (N_4931,In_1713,In_1578);
and U4932 (N_4932,In_84,In_782);
nand U4933 (N_4933,In_230,In_303);
or U4934 (N_4934,In_1723,In_940);
and U4935 (N_4935,In_1663,In_1312);
or U4936 (N_4936,In_752,In_575);
nand U4937 (N_4937,In_4,In_1378);
and U4938 (N_4938,In_889,In_502);
and U4939 (N_4939,In_1456,In_140);
or U4940 (N_4940,In_631,In_305);
or U4941 (N_4941,In_394,In_491);
and U4942 (N_4942,In_858,In_143);
or U4943 (N_4943,In_1295,In_36);
or U4944 (N_4944,In_1143,In_917);
xor U4945 (N_4945,In_747,In_522);
nor U4946 (N_4946,In_805,In_1575);
nand U4947 (N_4947,In_803,In_870);
and U4948 (N_4948,In_1296,In_834);
and U4949 (N_4949,In_43,In_714);
nor U4950 (N_4950,In_391,In_1099);
nand U4951 (N_4951,In_208,In_1940);
xnor U4952 (N_4952,In_965,In_371);
nand U4953 (N_4953,In_272,In_1248);
nand U4954 (N_4954,In_1064,In_1099);
nor U4955 (N_4955,In_60,In_818);
nand U4956 (N_4956,In_1212,In_1155);
and U4957 (N_4957,In_1248,In_261);
xnor U4958 (N_4958,In_1523,In_626);
nor U4959 (N_4959,In_56,In_1316);
xor U4960 (N_4960,In_1249,In_1674);
or U4961 (N_4961,In_1682,In_370);
xnor U4962 (N_4962,In_1396,In_154);
nand U4963 (N_4963,In_1206,In_1477);
and U4964 (N_4964,In_1315,In_1628);
xnor U4965 (N_4965,In_195,In_726);
and U4966 (N_4966,In_654,In_1093);
xor U4967 (N_4967,In_1776,In_8);
and U4968 (N_4968,In_902,In_161);
nor U4969 (N_4969,In_801,In_1468);
nand U4970 (N_4970,In_63,In_1493);
nor U4971 (N_4971,In_1425,In_1610);
nand U4972 (N_4972,In_358,In_134);
nand U4973 (N_4973,In_1185,In_639);
nand U4974 (N_4974,In_142,In_206);
and U4975 (N_4975,In_53,In_432);
or U4976 (N_4976,In_1188,In_902);
and U4977 (N_4977,In_526,In_301);
nand U4978 (N_4978,In_1200,In_816);
nand U4979 (N_4979,In_170,In_848);
or U4980 (N_4980,In_376,In_599);
nand U4981 (N_4981,In_1489,In_1428);
nor U4982 (N_4982,In_1433,In_786);
or U4983 (N_4983,In_1731,In_1677);
and U4984 (N_4984,In_744,In_1718);
and U4985 (N_4985,In_1822,In_425);
xnor U4986 (N_4986,In_1016,In_800);
nand U4987 (N_4987,In_1292,In_1514);
or U4988 (N_4988,In_1754,In_41);
or U4989 (N_4989,In_1905,In_182);
nor U4990 (N_4990,In_384,In_381);
nand U4991 (N_4991,In_1772,In_1361);
nor U4992 (N_4992,In_1296,In_364);
nand U4993 (N_4993,In_154,In_1285);
and U4994 (N_4994,In_567,In_24);
and U4995 (N_4995,In_213,In_137);
or U4996 (N_4996,In_670,In_281);
xor U4997 (N_4997,In_1008,In_1401);
nand U4998 (N_4998,In_729,In_211);
or U4999 (N_4999,In_200,In_1956);
nand U5000 (N_5000,N_3269,N_2687);
or U5001 (N_5001,N_4654,N_3571);
nand U5002 (N_5002,N_1221,N_2831);
and U5003 (N_5003,N_3899,N_765);
or U5004 (N_5004,N_756,N_1042);
nand U5005 (N_5005,N_3740,N_3719);
nor U5006 (N_5006,N_4191,N_259);
or U5007 (N_5007,N_4621,N_263);
or U5008 (N_5008,N_1264,N_335);
or U5009 (N_5009,N_2828,N_4125);
nor U5010 (N_5010,N_3757,N_115);
nand U5011 (N_5011,N_2055,N_685);
nand U5012 (N_5012,N_1251,N_1223);
nand U5013 (N_5013,N_4607,N_2827);
nor U5014 (N_5014,N_879,N_2583);
nand U5015 (N_5015,N_470,N_4674);
or U5016 (N_5016,N_971,N_4578);
nand U5017 (N_5017,N_4019,N_2532);
nor U5018 (N_5018,N_2764,N_327);
and U5019 (N_5019,N_4758,N_3940);
nand U5020 (N_5020,N_4404,N_3287);
nor U5021 (N_5021,N_2013,N_1517);
and U5022 (N_5022,N_2578,N_862);
or U5023 (N_5023,N_1879,N_715);
or U5024 (N_5024,N_3540,N_890);
and U5025 (N_5025,N_4165,N_3822);
nor U5026 (N_5026,N_3453,N_197);
and U5027 (N_5027,N_4056,N_53);
nor U5028 (N_5028,N_2354,N_4310);
nor U5029 (N_5029,N_1790,N_176);
or U5030 (N_5030,N_4440,N_846);
and U5031 (N_5031,N_1808,N_2962);
nor U5032 (N_5032,N_1319,N_4737);
nand U5033 (N_5033,N_1300,N_4907);
and U5034 (N_5034,N_189,N_3624);
nor U5035 (N_5035,N_4114,N_2032);
xnor U5036 (N_5036,N_4452,N_3946);
nand U5037 (N_5037,N_2692,N_814);
xor U5038 (N_5038,N_1035,N_641);
nor U5039 (N_5039,N_491,N_4086);
or U5040 (N_5040,N_3234,N_3629);
nand U5041 (N_5041,N_4435,N_3444);
nand U5042 (N_5042,N_2915,N_3779);
xor U5043 (N_5043,N_26,N_3794);
nor U5044 (N_5044,N_2627,N_747);
nand U5045 (N_5045,N_1586,N_2907);
nor U5046 (N_5046,N_1148,N_520);
and U5047 (N_5047,N_1579,N_4096);
and U5048 (N_5048,N_4969,N_1490);
nor U5049 (N_5049,N_4542,N_365);
or U5050 (N_5050,N_2768,N_1479);
nor U5051 (N_5051,N_3374,N_1342);
or U5052 (N_5052,N_4927,N_4162);
and U5053 (N_5053,N_4210,N_1603);
and U5054 (N_5054,N_1701,N_4324);
and U5055 (N_5055,N_656,N_2664);
nand U5056 (N_5056,N_3448,N_2806);
nor U5057 (N_5057,N_2665,N_3416);
nand U5058 (N_5058,N_4460,N_615);
nand U5059 (N_5059,N_212,N_3782);
nor U5060 (N_5060,N_1537,N_1581);
nor U5061 (N_5061,N_2037,N_3766);
and U5062 (N_5062,N_2990,N_2909);
or U5063 (N_5063,N_3456,N_4519);
or U5064 (N_5064,N_1591,N_3233);
nand U5065 (N_5065,N_2501,N_4020);
and U5066 (N_5066,N_1937,N_3531);
or U5067 (N_5067,N_4691,N_749);
or U5068 (N_5068,N_1767,N_2486);
nand U5069 (N_5069,N_2033,N_4084);
nor U5070 (N_5070,N_4928,N_2191);
and U5071 (N_5071,N_233,N_2411);
and U5072 (N_5072,N_891,N_1661);
and U5073 (N_5073,N_4805,N_1002);
and U5074 (N_5074,N_1670,N_213);
or U5075 (N_5075,N_497,N_2181);
or U5076 (N_5076,N_1774,N_1644);
nand U5077 (N_5077,N_2548,N_1078);
or U5078 (N_5078,N_983,N_1668);
nor U5079 (N_5079,N_1157,N_2622);
nor U5080 (N_5080,N_2799,N_4611);
nand U5081 (N_5081,N_2413,N_193);
nor U5082 (N_5082,N_3969,N_4494);
or U5083 (N_5083,N_2313,N_2149);
and U5084 (N_5084,N_4391,N_2816);
and U5085 (N_5085,N_583,N_3783);
and U5086 (N_5086,N_3631,N_1919);
nand U5087 (N_5087,N_1830,N_1032);
nor U5088 (N_5088,N_1017,N_707);
and U5089 (N_5089,N_3599,N_11);
nand U5090 (N_5090,N_3149,N_2763);
nor U5091 (N_5091,N_141,N_2320);
and U5092 (N_5092,N_1468,N_1832);
nor U5093 (N_5093,N_959,N_4793);
nor U5094 (N_5094,N_1665,N_4095);
nand U5095 (N_5095,N_2557,N_2285);
nor U5096 (N_5096,N_618,N_4597);
and U5097 (N_5097,N_3710,N_3851);
nor U5098 (N_5098,N_1008,N_2446);
and U5099 (N_5099,N_1461,N_3076);
or U5100 (N_5100,N_3016,N_4827);
nor U5101 (N_5101,N_4221,N_4294);
xnor U5102 (N_5102,N_4033,N_4733);
xnor U5103 (N_5103,N_3220,N_3956);
or U5104 (N_5104,N_4650,N_4574);
nor U5105 (N_5105,N_2155,N_2228);
or U5106 (N_5106,N_2043,N_444);
nand U5107 (N_5107,N_4302,N_3472);
xnor U5108 (N_5108,N_3840,N_1142);
nor U5109 (N_5109,N_4980,N_801);
or U5110 (N_5110,N_4756,N_1676);
or U5111 (N_5111,N_1706,N_2840);
or U5112 (N_5112,N_1496,N_4340);
nor U5113 (N_5113,N_3742,N_2061);
or U5114 (N_5114,N_2637,N_3979);
nand U5115 (N_5115,N_892,N_3700);
nor U5116 (N_5116,N_4577,N_1134);
nand U5117 (N_5117,N_3194,N_413);
and U5118 (N_5118,N_2537,N_4040);
or U5119 (N_5119,N_3084,N_1215);
or U5120 (N_5120,N_1420,N_4591);
nor U5121 (N_5121,N_3141,N_1269);
and U5122 (N_5122,N_2914,N_226);
nor U5123 (N_5123,N_27,N_4216);
xor U5124 (N_5124,N_3341,N_3195);
or U5125 (N_5125,N_4858,N_3254);
or U5126 (N_5126,N_3587,N_3106);
nor U5127 (N_5127,N_2882,N_2607);
and U5128 (N_5128,N_2940,N_4012);
or U5129 (N_5129,N_0,N_3803);
and U5130 (N_5130,N_3484,N_4497);
nor U5131 (N_5131,N_2267,N_1716);
nor U5132 (N_5132,N_3704,N_2345);
nor U5133 (N_5133,N_4192,N_3662);
xor U5134 (N_5134,N_1241,N_4026);
nand U5135 (N_5135,N_3775,N_3047);
or U5136 (N_5136,N_87,N_4748);
nand U5137 (N_5137,N_3862,N_4580);
nor U5138 (N_5138,N_4380,N_4146);
or U5139 (N_5139,N_929,N_1677);
xnor U5140 (N_5140,N_952,N_2098);
and U5141 (N_5141,N_2384,N_1837);
nor U5142 (N_5142,N_663,N_4878);
nand U5143 (N_5143,N_2776,N_4762);
or U5144 (N_5144,N_2897,N_1120);
nor U5145 (N_5145,N_2208,N_1273);
nand U5146 (N_5146,N_3365,N_645);
or U5147 (N_5147,N_1130,N_3980);
and U5148 (N_5148,N_2654,N_4979);
and U5149 (N_5149,N_4054,N_4799);
nand U5150 (N_5150,N_1355,N_1006);
nand U5151 (N_5151,N_4724,N_555);
or U5152 (N_5152,N_2551,N_4124);
nor U5153 (N_5153,N_3402,N_3485);
nor U5154 (N_5154,N_4803,N_2732);
and U5155 (N_5155,N_2959,N_1266);
and U5156 (N_5156,N_1759,N_1763);
nor U5157 (N_5157,N_78,N_4958);
and U5158 (N_5158,N_390,N_4899);
nand U5159 (N_5159,N_2142,N_2030);
and U5160 (N_5160,N_4744,N_3666);
nor U5161 (N_5161,N_2131,N_4475);
nand U5162 (N_5162,N_54,N_4840);
nor U5163 (N_5163,N_690,N_2024);
nand U5164 (N_5164,N_1481,N_3277);
nand U5165 (N_5165,N_4070,N_525);
or U5166 (N_5166,N_3375,N_1527);
and U5167 (N_5167,N_295,N_4353);
xnor U5168 (N_5168,N_705,N_1073);
and U5169 (N_5169,N_3814,N_2456);
nor U5170 (N_5170,N_2618,N_4952);
and U5171 (N_5171,N_1548,N_3860);
and U5172 (N_5172,N_2021,N_3983);
nand U5173 (N_5173,N_1252,N_4912);
or U5174 (N_5174,N_1923,N_381);
and U5175 (N_5175,N_4203,N_791);
nand U5176 (N_5176,N_4428,N_4182);
or U5177 (N_5177,N_4579,N_1904);
nor U5178 (N_5178,N_1782,N_2182);
nand U5179 (N_5179,N_3808,N_2430);
and U5180 (N_5180,N_2552,N_313);
and U5181 (N_5181,N_1641,N_2334);
nor U5182 (N_5182,N_4627,N_4815);
nor U5183 (N_5183,N_3907,N_4141);
xor U5184 (N_5184,N_2054,N_551);
and U5185 (N_5185,N_3210,N_235);
and U5186 (N_5186,N_4856,N_1526);
or U5187 (N_5187,N_4777,N_1839);
or U5188 (N_5188,N_4971,N_4743);
xnor U5189 (N_5189,N_2025,N_2502);
xor U5190 (N_5190,N_1039,N_3502);
nand U5191 (N_5191,N_2358,N_2388);
nor U5192 (N_5192,N_1056,N_1528);
nor U5193 (N_5193,N_4480,N_1399);
and U5194 (N_5194,N_3255,N_691);
and U5195 (N_5195,N_2613,N_2489);
and U5196 (N_5196,N_3155,N_3861);
or U5197 (N_5197,N_4249,N_1369);
and U5198 (N_5198,N_2729,N_3103);
xnor U5199 (N_5199,N_261,N_18);
or U5200 (N_5200,N_772,N_150);
nor U5201 (N_5201,N_4385,N_2516);
nor U5202 (N_5202,N_793,N_4469);
and U5203 (N_5203,N_650,N_4386);
and U5204 (N_5204,N_4648,N_2623);
and U5205 (N_5205,N_3207,N_1942);
xnor U5206 (N_5206,N_1571,N_3809);
nand U5207 (N_5207,N_2937,N_4853);
and U5208 (N_5208,N_2066,N_2185);
and U5209 (N_5209,N_2350,N_1324);
nor U5210 (N_5210,N_4595,N_4568);
nand U5211 (N_5211,N_1088,N_3584);
or U5212 (N_5212,N_3268,N_3503);
nor U5213 (N_5213,N_2461,N_4438);
nor U5214 (N_5214,N_348,N_302);
nand U5215 (N_5215,N_3401,N_2808);
or U5216 (N_5216,N_4430,N_4166);
nand U5217 (N_5217,N_2370,N_158);
and U5218 (N_5218,N_52,N_2368);
nand U5219 (N_5219,N_1080,N_3098);
nor U5220 (N_5220,N_1689,N_825);
and U5221 (N_5221,N_1636,N_72);
nand U5222 (N_5222,N_532,N_3323);
and U5223 (N_5223,N_2600,N_1866);
or U5224 (N_5224,N_2148,N_3945);
xnor U5225 (N_5225,N_1272,N_626);
nand U5226 (N_5226,N_4936,N_4420);
nor U5227 (N_5227,N_3392,N_3483);
and U5228 (N_5228,N_1805,N_4807);
nand U5229 (N_5229,N_119,N_3048);
and U5230 (N_5230,N_2609,N_4305);
nor U5231 (N_5231,N_2097,N_3475);
or U5232 (N_5232,N_1060,N_2567);
or U5233 (N_5233,N_2304,N_1344);
or U5234 (N_5234,N_75,N_1564);
nor U5235 (N_5235,N_3586,N_1705);
or U5236 (N_5236,N_2193,N_1351);
nor U5237 (N_5237,N_4254,N_184);
or U5238 (N_5238,N_1519,N_1557);
and U5239 (N_5239,N_3542,N_3145);
nand U5240 (N_5240,N_2553,N_3867);
and U5241 (N_5241,N_3964,N_4226);
nor U5242 (N_5242,N_1389,N_522);
nand U5243 (N_5243,N_1589,N_1655);
nor U5244 (N_5244,N_3085,N_2893);
and U5245 (N_5245,N_4194,N_3957);
and U5246 (N_5246,N_3651,N_3912);
nor U5247 (N_5247,N_4620,N_4987);
and U5248 (N_5248,N_831,N_2283);
or U5249 (N_5249,N_4163,N_2722);
and U5250 (N_5250,N_4325,N_1093);
nand U5251 (N_5251,N_4372,N_3797);
or U5252 (N_5252,N_800,N_3683);
or U5253 (N_5253,N_769,N_806);
xor U5254 (N_5254,N_4399,N_1491);
xor U5255 (N_5255,N_1509,N_2500);
or U5256 (N_5256,N_1973,N_3967);
nor U5257 (N_5257,N_2412,N_4334);
xnor U5258 (N_5258,N_3516,N_301);
xnor U5259 (N_5259,N_3590,N_2984);
nand U5260 (N_5260,N_2906,N_2956);
nor U5261 (N_5261,N_1849,N_3603);
and U5262 (N_5262,N_2256,N_1723);
and U5263 (N_5263,N_3099,N_4161);
or U5264 (N_5264,N_544,N_220);
and U5265 (N_5265,N_3682,N_3425);
nor U5266 (N_5266,N_4456,N_2524);
and U5267 (N_5267,N_3110,N_2617);
nor U5268 (N_5268,N_3183,N_576);
and U5269 (N_5269,N_592,N_504);
xor U5270 (N_5270,N_2439,N_1529);
or U5271 (N_5271,N_1694,N_731);
nor U5272 (N_5272,N_3299,N_1753);
nand U5273 (N_5273,N_4295,N_4562);
or U5274 (N_5274,N_1307,N_1218);
nor U5275 (N_5275,N_1431,N_2257);
or U5276 (N_5276,N_3904,N_4132);
nand U5277 (N_5277,N_1840,N_662);
and U5278 (N_5278,N_936,N_646);
nor U5279 (N_5279,N_94,N_4929);
or U5280 (N_5280,N_540,N_3345);
or U5281 (N_5281,N_1722,N_1859);
nand U5282 (N_5282,N_2641,N_1531);
and U5283 (N_5283,N_989,N_148);
nand U5284 (N_5284,N_2428,N_38);
nor U5285 (N_5285,N_4660,N_4407);
nor U5286 (N_5286,N_2895,N_4575);
or U5287 (N_5287,N_1929,N_1725);
nor U5288 (N_5288,N_1608,N_4930);
or U5289 (N_5289,N_223,N_2450);
nand U5290 (N_5290,N_2601,N_4964);
nand U5291 (N_5291,N_2137,N_909);
or U5292 (N_5292,N_1822,N_4989);
nor U5293 (N_5293,N_356,N_2473);
and U5294 (N_5294,N_3131,N_3870);
and U5295 (N_5295,N_1204,N_374);
or U5296 (N_5296,N_968,N_192);
nand U5297 (N_5297,N_3019,N_590);
or U5298 (N_5298,N_1762,N_276);
and U5299 (N_5299,N_807,N_4122);
nor U5300 (N_5300,N_1971,N_4247);
nor U5301 (N_5301,N_2154,N_2344);
xor U5302 (N_5302,N_669,N_3674);
nand U5303 (N_5303,N_369,N_2514);
xnor U5304 (N_5304,N_910,N_4222);
nor U5305 (N_5305,N_2086,N_1930);
and U5306 (N_5306,N_3937,N_3333);
nor U5307 (N_5307,N_681,N_2935);
nand U5308 (N_5308,N_1729,N_3158);
nor U5309 (N_5309,N_673,N_4066);
nor U5310 (N_5310,N_1543,N_4496);
and U5311 (N_5311,N_4833,N_818);
xor U5312 (N_5312,N_3184,N_1792);
or U5313 (N_5313,N_1547,N_2420);
xnor U5314 (N_5314,N_1749,N_172);
and U5315 (N_5315,N_821,N_3060);
and U5316 (N_5316,N_346,N_1402);
nand U5317 (N_5317,N_4649,N_1077);
nand U5318 (N_5318,N_4903,N_4327);
or U5319 (N_5319,N_1024,N_3817);
xor U5320 (N_5320,N_1189,N_4999);
and U5321 (N_5321,N_3944,N_2530);
nand U5322 (N_5322,N_4035,N_1760);
and U5323 (N_5323,N_251,N_3720);
nand U5324 (N_5324,N_73,N_1615);
nand U5325 (N_5325,N_1202,N_4937);
and U5326 (N_5326,N_2821,N_3072);
or U5327 (N_5327,N_1754,N_3216);
nand U5328 (N_5328,N_1957,N_3335);
xor U5329 (N_5329,N_225,N_2253);
nor U5330 (N_5330,N_2792,N_2386);
or U5331 (N_5331,N_489,N_2157);
or U5332 (N_5332,N_1124,N_3021);
and U5333 (N_5333,N_1275,N_2046);
and U5334 (N_5334,N_90,N_4272);
nand U5335 (N_5335,N_914,N_1566);
nor U5336 (N_5336,N_2168,N_1208);
and U5337 (N_5337,N_4373,N_1649);
xor U5338 (N_5338,N_55,N_49);
nor U5339 (N_5339,N_2885,N_667);
or U5340 (N_5340,N_3768,N_1478);
and U5341 (N_5341,N_1188,N_2478);
nor U5342 (N_5342,N_399,N_4439);
nand U5343 (N_5343,N_1881,N_2487);
and U5344 (N_5344,N_1746,N_4094);
and U5345 (N_5345,N_2710,N_516);
or U5346 (N_5346,N_992,N_4961);
nor U5347 (N_5347,N_3627,N_4945);
and U5348 (N_5348,N_4291,N_4424);
nor U5349 (N_5349,N_3736,N_2198);
and U5350 (N_5350,N_970,N_3798);
nor U5351 (N_5351,N_4730,N_431);
nand U5352 (N_5352,N_3534,N_252);
nor U5353 (N_5353,N_737,N_229);
nand U5354 (N_5354,N_3310,N_2515);
xor U5355 (N_5355,N_4230,N_598);
nor U5356 (N_5356,N_363,N_1857);
or U5357 (N_5357,N_2049,N_3143);
nor U5358 (N_5358,N_3741,N_4766);
and U5359 (N_5359,N_2919,N_377);
or U5360 (N_5360,N_2499,N_2340);
nand U5361 (N_5361,N_4479,N_773);
nor U5362 (N_5362,N_3726,N_1633);
xnor U5363 (N_5363,N_4449,N_1287);
nor U5364 (N_5364,N_1294,N_3621);
nor U5365 (N_5365,N_445,N_4278);
or U5366 (N_5366,N_4136,N_2911);
and U5367 (N_5367,N_4594,N_2277);
and U5368 (N_5368,N_573,N_1632);
nor U5369 (N_5369,N_1736,N_2878);
or U5370 (N_5370,N_955,N_1087);
nor U5371 (N_5371,N_4336,N_4018);
nand U5372 (N_5372,N_398,N_304);
or U5373 (N_5373,N_2569,N_3230);
or U5374 (N_5374,N_3007,N_3306);
nand U5375 (N_5375,N_3154,N_1781);
or U5376 (N_5376,N_768,N_3319);
and U5377 (N_5377,N_135,N_3977);
nand U5378 (N_5378,N_4919,N_559);
and U5379 (N_5379,N_1520,N_4118);
xor U5380 (N_5380,N_2513,N_2682);
and U5381 (N_5381,N_3272,N_4689);
nor U5382 (N_5382,N_4872,N_1820);
nor U5383 (N_5383,N_312,N_3898);
and U5384 (N_5384,N_897,N_4843);
nor U5385 (N_5385,N_1824,N_4003);
nor U5386 (N_5386,N_298,N_3396);
and U5387 (N_5387,N_4371,N_4786);
nor U5388 (N_5388,N_4553,N_1101);
and U5389 (N_5389,N_542,N_2635);
nand U5390 (N_5390,N_3369,N_1841);
nand U5391 (N_5391,N_4729,N_3015);
and U5392 (N_5392,N_1426,N_1681);
nand U5393 (N_5393,N_3811,N_2643);
or U5394 (N_5394,N_736,N_1972);
nand U5395 (N_5395,N_597,N_3812);
or U5396 (N_5396,N_774,N_2031);
nand U5397 (N_5397,N_4024,N_2785);
nand U5398 (N_5398,N_1623,N_4817);
nand U5399 (N_5399,N_3632,N_25);
or U5400 (N_5400,N_3819,N_1889);
nand U5401 (N_5401,N_2251,N_2881);
nor U5402 (N_5402,N_4663,N_4721);
nand U5403 (N_5403,N_4457,N_1220);
nand U5404 (N_5404,N_3156,N_4264);
nor U5405 (N_5405,N_2987,N_687);
nand U5406 (N_5406,N_426,N_2357);
nand U5407 (N_5407,N_1821,N_809);
nor U5408 (N_5408,N_4156,N_4117);
or U5409 (N_5409,N_2734,N_4376);
nand U5410 (N_5410,N_4069,N_1277);
nand U5411 (N_5411,N_1766,N_627);
nor U5412 (N_5412,N_2760,N_3340);
nand U5413 (N_5413,N_487,N_682);
and U5414 (N_5414,N_3971,N_3707);
and U5415 (N_5415,N_1439,N_1176);
nand U5416 (N_5416,N_165,N_282);
and U5417 (N_5417,N_2559,N_149);
and U5418 (N_5418,N_3687,N_1046);
nand U5419 (N_5419,N_2332,N_1651);
or U5420 (N_5420,N_255,N_2109);
nand U5421 (N_5421,N_142,N_2402);
or U5422 (N_5422,N_917,N_2452);
xor U5423 (N_5423,N_3780,N_240);
nor U5424 (N_5424,N_4426,N_3070);
nor U5425 (N_5425,N_560,N_3031);
xor U5426 (N_5426,N_3724,N_3857);
nand U5427 (N_5427,N_4665,N_314);
xor U5428 (N_5428,N_616,N_4462);
and U5429 (N_5429,N_3238,N_2014);
nand U5430 (N_5430,N_296,N_2661);
or U5431 (N_5431,N_2765,N_4911);
or U5432 (N_5432,N_3303,N_4888);
and U5433 (N_5433,N_535,N_404);
and U5434 (N_5434,N_808,N_878);
or U5435 (N_5435,N_4842,N_56);
nor U5436 (N_5436,N_2406,N_280);
and U5437 (N_5437,N_1909,N_2300);
or U5438 (N_5438,N_2606,N_2852);
nor U5439 (N_5439,N_2586,N_2705);
or U5440 (N_5440,N_3579,N_3816);
and U5441 (N_5441,N_657,N_2711);
and U5442 (N_5442,N_4005,N_3002);
nand U5443 (N_5443,N_3479,N_3445);
nand U5444 (N_5444,N_3294,N_3136);
xor U5445 (N_5445,N_1379,N_2761);
or U5446 (N_5446,N_1020,N_4696);
and U5447 (N_5447,N_941,N_257);
nor U5448 (N_5448,N_612,N_4783);
nor U5449 (N_5449,N_3591,N_2465);
xnor U5450 (N_5450,N_2671,N_3180);
and U5451 (N_5451,N_4101,N_1406);
nor U5452 (N_5452,N_3725,N_2346);
nand U5453 (N_5453,N_3615,N_3382);
or U5454 (N_5454,N_2988,N_2020);
or U5455 (N_5455,N_3745,N_4516);
nand U5456 (N_5456,N_4677,N_2697);
nand U5457 (N_5457,N_2407,N_688);
nand U5458 (N_5458,N_723,N_2669);
nand U5459 (N_5459,N_126,N_1952);
nand U5460 (N_5460,N_2405,N_3077);
or U5461 (N_5461,N_3829,N_600);
or U5462 (N_5462,N_557,N_473);
nor U5463 (N_5463,N_4281,N_1068);
nor U5464 (N_5464,N_2124,N_4431);
or U5465 (N_5465,N_2477,N_655);
nand U5466 (N_5466,N_4751,N_1397);
nor U5467 (N_5467,N_1550,N_4869);
and U5468 (N_5468,N_4021,N_2158);
nand U5469 (N_5469,N_2645,N_2504);
nor U5470 (N_5470,N_2490,N_3372);
or U5471 (N_5471,N_4686,N_1788);
nor U5472 (N_5472,N_2337,N_3337);
and U5473 (N_5473,N_4234,N_322);
nor U5474 (N_5474,N_4251,N_1235);
nor U5475 (N_5475,N_713,N_3185);
and U5476 (N_5476,N_2783,N_3827);
nand U5477 (N_5477,N_2180,N_3985);
nor U5478 (N_5478,N_287,N_994);
nand U5479 (N_5479,N_1475,N_4918);
and U5480 (N_5480,N_3787,N_4300);
nor U5481 (N_5481,N_3873,N_4395);
and U5482 (N_5482,N_1422,N_3188);
nor U5483 (N_5483,N_3711,N_2209);
nand U5484 (N_5484,N_1113,N_2485);
and U5485 (N_5485,N_4513,N_4285);
xor U5486 (N_5486,N_3146,N_2296);
nor U5487 (N_5487,N_3377,N_961);
nand U5488 (N_5488,N_2562,N_2996);
and U5489 (N_5489,N_3746,N_2943);
xor U5490 (N_5490,N_2292,N_977);
and U5491 (N_5491,N_432,N_3801);
xor U5492 (N_5492,N_243,N_4603);
nand U5493 (N_5493,N_1198,N_2232);
or U5494 (N_5494,N_594,N_2653);
or U5495 (N_5495,N_3581,N_3054);
and U5496 (N_5496,N_4983,N_916);
and U5497 (N_5497,N_4616,N_3252);
and U5498 (N_5498,N_3880,N_4659);
xnor U5499 (N_5499,N_1114,N_1675);
xor U5500 (N_5500,N_3610,N_3352);
or U5501 (N_5501,N_3789,N_3496);
nor U5502 (N_5502,N_1184,N_1748);
and U5503 (N_5503,N_1048,N_3022);
and U5504 (N_5504,N_751,N_2858);
and U5505 (N_5505,N_3555,N_693);
or U5506 (N_5506,N_4592,N_1780);
or U5507 (N_5507,N_3030,N_4064);
nor U5508 (N_5508,N_4240,N_3909);
or U5509 (N_5509,N_60,N_4544);
nand U5510 (N_5510,N_2162,N_3212);
or U5511 (N_5511,N_493,N_2493);
nor U5512 (N_5512,N_4408,N_869);
and U5513 (N_5513,N_2901,N_112);
or U5514 (N_5514,N_2132,N_4501);
nand U5515 (N_5515,N_4304,N_3291);
nand U5516 (N_5516,N_4666,N_930);
nor U5517 (N_5517,N_3832,N_2077);
nor U5518 (N_5518,N_4115,N_649);
nor U5519 (N_5519,N_4850,N_3421);
and U5520 (N_5520,N_2712,N_2983);
nor U5521 (N_5521,N_394,N_4922);
and U5522 (N_5522,N_1352,N_2812);
or U5523 (N_5523,N_4409,N_2028);
and U5524 (N_5524,N_2856,N_2690);
and U5525 (N_5525,N_1278,N_58);
xor U5526 (N_5526,N_3122,N_1842);
nand U5527 (N_5527,N_29,N_250);
nor U5528 (N_5528,N_2241,N_4341);
nor U5529 (N_5529,N_3083,N_3737);
and U5530 (N_5530,N_4362,N_1447);
or U5531 (N_5531,N_2503,N_2945);
and U5532 (N_5532,N_4382,N_4032);
and U5533 (N_5533,N_2947,N_2992);
or U5534 (N_5534,N_2480,N_827);
nor U5535 (N_5535,N_3092,N_4867);
xor U5536 (N_5536,N_4991,N_2318);
nand U5537 (N_5537,N_2464,N_3850);
nor U5538 (N_5538,N_3750,N_474);
nor U5539 (N_5539,N_3138,N_4631);
nor U5540 (N_5540,N_4746,N_4641);
and U5541 (N_5541,N_3288,N_2924);
and U5542 (N_5542,N_3955,N_47);
nor U5543 (N_5543,N_3614,N_2991);
and U5544 (N_5544,N_1247,N_3600);
and U5545 (N_5545,N_3691,N_3973);
and U5546 (N_5546,N_785,N_1454);
and U5547 (N_5547,N_81,N_1110);
and U5548 (N_5548,N_4676,N_1695);
or U5549 (N_5549,N_3404,N_2795);
nand U5550 (N_5550,N_2787,N_3815);
and U5551 (N_5551,N_2593,N_2753);
nor U5552 (N_5552,N_3244,N_1819);
or U5553 (N_5553,N_3876,N_2353);
or U5554 (N_5554,N_334,N_4109);
nor U5555 (N_5555,N_4195,N_4551);
nor U5556 (N_5556,N_4121,N_2560);
nand U5557 (N_5557,N_1552,N_2355);
or U5558 (N_5558,N_3813,N_4819);
or U5559 (N_5559,N_1348,N_3929);
and U5560 (N_5560,N_4255,N_4184);
and U5561 (N_5561,N_4896,N_610);
nor U5562 (N_5562,N_4736,N_4901);
or U5563 (N_5563,N_434,N_3588);
and U5564 (N_5564,N_4453,N_4968);
xnor U5565 (N_5565,N_817,N_461);
nand U5566 (N_5566,N_1932,N_4477);
nand U5567 (N_5567,N_964,N_3253);
nor U5568 (N_5568,N_2976,N_811);
and U5569 (N_5569,N_1688,N_3082);
and U5570 (N_5570,N_1321,N_367);
nor U5571 (N_5571,N_4492,N_620);
nor U5572 (N_5572,N_3660,N_900);
and U5573 (N_5573,N_1876,N_1980);
nand U5574 (N_5574,N_860,N_86);
or U5575 (N_5575,N_2325,N_2261);
and U5576 (N_5576,N_2394,N_380);
and U5577 (N_5577,N_3838,N_4068);
xnor U5578 (N_5578,N_1569,N_2335);
and U5579 (N_5579,N_1535,N_730);
xnor U5580 (N_5580,N_2400,N_582);
nand U5581 (N_5581,N_3762,N_3573);
nand U5582 (N_5582,N_1410,N_3981);
or U5583 (N_5583,N_3894,N_3576);
or U5584 (N_5584,N_2434,N_2542);
or U5585 (N_5585,N_3856,N_4227);
and U5586 (N_5586,N_1939,N_3518);
nand U5587 (N_5587,N_2571,N_4149);
and U5588 (N_5588,N_3714,N_4831);
and U5589 (N_5589,N_948,N_3892);
xnor U5590 (N_5590,N_4486,N_2244);
and U5591 (N_5591,N_1357,N_1826);
or U5592 (N_5592,N_1469,N_2543);
or U5593 (N_5593,N_4732,N_3931);
nand U5594 (N_5594,N_2696,N_3258);
nand U5595 (N_5595,N_1099,N_1684);
xor U5596 (N_5596,N_3150,N_2004);
nor U5597 (N_5597,N_1126,N_4589);
nand U5598 (N_5598,N_3437,N_1000);
nor U5599 (N_5599,N_841,N_4681);
or U5600 (N_5600,N_1950,N_2800);
nand U5601 (N_5601,N_940,N_1690);
nand U5602 (N_5602,N_2259,N_4455);
nor U5603 (N_5603,N_702,N_4555);
nand U5604 (N_5604,N_1427,N_4406);
and U5605 (N_5605,N_315,N_2550);
and U5606 (N_5606,N_1495,N_1238);
xor U5607 (N_5607,N_2746,N_3703);
nor U5608 (N_5608,N_3645,N_4013);
or U5609 (N_5609,N_2519,N_1456);
or U5610 (N_5610,N_1714,N_4345);
nor U5611 (N_5611,N_3457,N_4413);
or U5612 (N_5612,N_3129,N_3101);
xnor U5613 (N_5613,N_1914,N_3367);
nor U5614 (N_5614,N_4262,N_1333);
or U5615 (N_5615,N_1128,N_4990);
nand U5616 (N_5616,N_2016,N_4976);
and U5617 (N_5617,N_3875,N_3593);
or U5618 (N_5618,N_3917,N_4996);
or U5619 (N_5619,N_4367,N_1462);
nand U5620 (N_5620,N_3261,N_922);
or U5621 (N_5621,N_1570,N_351);
nand U5622 (N_5622,N_1164,N_77);
nor U5623 (N_5623,N_4702,N_2592);
and U5624 (N_5624,N_2539,N_2419);
and U5625 (N_5625,N_3059,N_659);
nor U5626 (N_5626,N_4214,N_2052);
nor U5627 (N_5627,N_4105,N_4206);
and U5628 (N_5628,N_3293,N_3539);
nand U5629 (N_5629,N_4865,N_1804);
and U5630 (N_5630,N_873,N_2683);
nand U5631 (N_5631,N_981,N_3301);
nand U5632 (N_5632,N_2989,N_1525);
nand U5633 (N_5633,N_4606,N_2979);
nand U5634 (N_5634,N_57,N_4351);
nor U5635 (N_5635,N_1390,N_76);
nor U5636 (N_5636,N_2777,N_3492);
nand U5637 (N_5637,N_2842,N_1330);
and U5638 (N_5638,N_2404,N_3249);
or U5639 (N_5639,N_195,N_4127);
or U5640 (N_5640,N_472,N_3089);
nor U5641 (N_5641,N_3130,N_2647);
and U5642 (N_5642,N_3500,N_926);
and U5643 (N_5643,N_1827,N_3498);
nor U5644 (N_5644,N_4835,N_4466);
nand U5645 (N_5645,N_134,N_3357);
nand U5646 (N_5646,N_4967,N_3203);
nand U5647 (N_5647,N_757,N_2604);
and U5648 (N_5648,N_120,N_3609);
and U5649 (N_5649,N_1563,N_4312);
and U5650 (N_5650,N_4828,N_1775);
nor U5651 (N_5651,N_2491,N_1979);
nor U5652 (N_5652,N_3232,N_2873);
nor U5653 (N_5653,N_395,N_3830);
nand U5654 (N_5654,N_2297,N_4427);
and U5655 (N_5655,N_2196,N_571);
or U5656 (N_5656,N_614,N_1236);
nand U5657 (N_5657,N_3936,N_1734);
nand U5658 (N_5658,N_1429,N_1415);
nor U5659 (N_5659,N_1288,N_3749);
and U5660 (N_5660,N_4178,N_775);
nand U5661 (N_5661,N_1997,N_1726);
or U5662 (N_5662,N_2214,N_1865);
or U5663 (N_5663,N_4642,N_3752);
nand U5664 (N_5664,N_1817,N_1358);
nand U5665 (N_5665,N_847,N_2362);
xor U5666 (N_5666,N_2040,N_701);
nand U5667 (N_5667,N_3686,N_622);
or U5668 (N_5668,N_4583,N_4314);
or U5669 (N_5669,N_1067,N_3428);
nor U5670 (N_5670,N_2508,N_3635);
xor U5671 (N_5671,N_661,N_1281);
or U5672 (N_5672,N_4914,N_819);
xnor U5673 (N_5673,N_2742,N_4925);
and U5674 (N_5674,N_74,N_3735);
or U5675 (N_5675,N_254,N_1445);
nor U5676 (N_5676,N_932,N_4712);
nand U5677 (N_5677,N_1231,N_1850);
and U5678 (N_5678,N_2823,N_1737);
or U5679 (N_5679,N_127,N_1409);
or U5680 (N_5680,N_1401,N_4891);
or U5681 (N_5681,N_3664,N_587);
or U5682 (N_5682,N_3784,N_105);
or U5683 (N_5683,N_2201,N_3908);
nand U5684 (N_5684,N_536,N_689);
and U5685 (N_5685,N_4953,N_2850);
and U5686 (N_5686,N_717,N_2273);
nand U5687 (N_5687,N_3463,N_1064);
or U5688 (N_5688,N_1750,N_2786);
and U5689 (N_5689,N_4522,N_2248);
and U5690 (N_5690,N_3458,N_4993);
or U5691 (N_5691,N_305,N_490);
nor U5692 (N_5692,N_2679,N_3987);
nand U5693 (N_5693,N_3537,N_4811);
nand U5694 (N_5694,N_4349,N_2851);
nand U5695 (N_5695,N_4232,N_1951);
nand U5696 (N_5696,N_2752,N_1104);
nand U5697 (N_5697,N_1335,N_4852);
nand U5698 (N_5698,N_2939,N_658);
or U5699 (N_5699,N_1800,N_998);
nand U5700 (N_5700,N_1105,N_2321);
nor U5701 (N_5701,N_4784,N_4207);
and U5702 (N_5702,N_41,N_1034);
and U5703 (N_5703,N_1811,N_3992);
or U5704 (N_5704,N_786,N_2662);
nand U5705 (N_5705,N_2751,N_4363);
nand U5706 (N_5706,N_3302,N_2074);
nor U5707 (N_5707,N_2718,N_1908);
nand U5708 (N_5708,N_427,N_795);
and U5709 (N_5709,N_4379,N_1186);
nor U5710 (N_5710,N_4097,N_907);
and U5711 (N_5711,N_1743,N_1616);
or U5712 (N_5712,N_3434,N_1796);
and U5713 (N_5713,N_4458,N_908);
nor U5714 (N_5714,N_95,N_3001);
and U5715 (N_5715,N_3693,N_248);
xor U5716 (N_5716,N_741,N_440);
and U5717 (N_5717,N_4061,N_1313);
nor U5718 (N_5718,N_4714,N_996);
or U5719 (N_5719,N_1449,N_2212);
and U5720 (N_5720,N_4800,N_2757);
nand U5721 (N_5721,N_1707,N_85);
nand U5722 (N_5722,N_3821,N_1210);
nor U5723 (N_5723,N_4419,N_3094);
nor U5724 (N_5724,N_2007,N_2950);
nand U5725 (N_5725,N_3597,N_1337);
or U5726 (N_5726,N_2372,N_1228);
or U5727 (N_5727,N_2660,N_586);
nand U5728 (N_5728,N_2068,N_4267);
nand U5729 (N_5729,N_1147,N_4653);
nand U5730 (N_5730,N_3467,N_1136);
or U5731 (N_5731,N_761,N_1648);
and U5732 (N_5732,N_3105,N_1693);
or U5733 (N_5733,N_3834,N_4299);
nand U5734 (N_5734,N_1372,N_1201);
xor U5735 (N_5735,N_4009,N_1769);
xnor U5736 (N_5736,N_4079,N_3311);
or U5737 (N_5737,N_2269,N_450);
and U5738 (N_5738,N_2134,N_3558);
nor U5739 (N_5739,N_4506,N_3991);
xor U5740 (N_5740,N_2846,N_2565);
or U5741 (N_5741,N_1474,N_4771);
xor U5742 (N_5742,N_3659,N_1158);
or U5743 (N_5743,N_1065,N_4790);
nor U5744 (N_5744,N_1991,N_2190);
nand U5745 (N_5745,N_3895,N_4429);
nor U5746 (N_5746,N_1424,N_1671);
xor U5747 (N_5747,N_3777,N_4639);
or U5748 (N_5748,N_425,N_2417);
xnor U5749 (N_5749,N_310,N_3761);
or U5750 (N_5750,N_1868,N_1386);
and U5751 (N_5751,N_4504,N_1948);
nand U5752 (N_5752,N_3889,N_2997);
nor U5753 (N_5753,N_1985,N_4383);
and U5754 (N_5754,N_2903,N_4339);
xor U5755 (N_5755,N_1757,N_2608);
nand U5756 (N_5756,N_3028,N_2708);
or U5757 (N_5757,N_3366,N_2570);
nor U5758 (N_5758,N_110,N_1216);
nor U5759 (N_5759,N_872,N_2233);
nand U5760 (N_5760,N_3474,N_2121);
and U5761 (N_5761,N_2955,N_3116);
nor U5762 (N_5762,N_2245,N_1869);
xnor U5763 (N_5763,N_2649,N_2472);
or U5764 (N_5764,N_1191,N_2739);
xor U5765 (N_5765,N_1453,N_843);
nand U5766 (N_5766,N_3698,N_696);
nand U5767 (N_5767,N_1448,N_319);
and U5768 (N_5768,N_4031,N_492);
nand U5769 (N_5769,N_2965,N_2782);
xnor U5770 (N_5770,N_4527,N_281);
nor U5771 (N_5771,N_4242,N_3247);
nor U5772 (N_5772,N_2611,N_4375);
nor U5773 (N_5773,N_4767,N_1637);
xor U5774 (N_5774,N_3117,N_1556);
or U5775 (N_5775,N_3037,N_330);
nand U5776 (N_5776,N_1200,N_595);
and U5777 (N_5777,N_4701,N_4180);
and U5778 (N_5778,N_3257,N_4416);
nand U5779 (N_5779,N_1504,N_3673);
nor U5780 (N_5780,N_4433,N_3442);
nor U5781 (N_5781,N_2582,N_3179);
and U5782 (N_5782,N_2738,N_558);
and U5783 (N_5783,N_2681,N_3701);
nand U5784 (N_5784,N_1970,N_320);
nor U5785 (N_5785,N_4089,N_3706);
xnor U5786 (N_5786,N_1298,N_2819);
or U5787 (N_5787,N_161,N_810);
nand U5788 (N_5788,N_4798,N_4401);
or U5789 (N_5789,N_1855,N_3743);
or U5790 (N_5790,N_4643,N_2366);
nor U5791 (N_5791,N_2085,N_1996);
nor U5792 (N_5792,N_1106,N_480);
or U5793 (N_5793,N_871,N_1727);
nand U5794 (N_5794,N_2964,N_3665);
nor U5795 (N_5795,N_4112,N_4498);
and U5796 (N_5796,N_1450,N_4770);
nand U5797 (N_5797,N_99,N_564);
and U5798 (N_5798,N_3669,N_4683);
or U5799 (N_5799,N_1183,N_1473);
nand U5800 (N_5800,N_905,N_4742);
and U5801 (N_5801,N_2392,N_4241);
nor U5802 (N_5802,N_2048,N_1883);
or U5803 (N_5803,N_606,N_3915);
and U5804 (N_5804,N_4,N_835);
nand U5805 (N_5805,N_3032,N_4248);
and U5806 (N_5806,N_3962,N_514);
and U5807 (N_5807,N_294,N_3135);
and U5808 (N_5808,N_4738,N_4753);
nor U5809 (N_5809,N_4849,N_4881);
nand U5810 (N_5810,N_3174,N_3035);
nand U5811 (N_5811,N_1901,N_529);
nand U5812 (N_5812,N_4050,N_3260);
nor U5813 (N_5813,N_3582,N_783);
and U5814 (N_5814,N_3043,N_4845);
and U5815 (N_5815,N_1656,N_4731);
or U5816 (N_5816,N_3661,N_2000);
nor U5817 (N_5817,N_2899,N_771);
or U5818 (N_5818,N_1323,N_788);
nor U5819 (N_5819,N_2106,N_2274);
nor U5820 (N_5820,N_1590,N_143);
or U5821 (N_5821,N_838,N_2371);
xor U5822 (N_5822,N_4038,N_4396);
or U5823 (N_5823,N_4754,N_1451);
and U5824 (N_5824,N_2348,N_4100);
or U5825 (N_5825,N_919,N_3676);
nand U5826 (N_5826,N_1091,N_506);
nor U5827 (N_5827,N_4014,N_4211);
nor U5828 (N_5828,N_1360,N_4049);
or U5829 (N_5829,N_1935,N_986);
nor U5830 (N_5830,N_3217,N_4451);
or U5831 (N_5831,N_1925,N_2603);
and U5832 (N_5832,N_326,N_3221);
nand U5833 (N_5833,N_3239,N_1823);
or U5834 (N_5834,N_2869,N_1057);
nor U5835 (N_5835,N_4675,N_758);
and U5836 (N_5836,N_4781,N_2985);
xor U5837 (N_5837,N_3109,N_1540);
or U5838 (N_5838,N_2468,N_415);
and U5839 (N_5839,N_3429,N_4158);
and U5840 (N_5840,N_2838,N_3888);
and U5841 (N_5841,N_343,N_1193);
xnor U5842 (N_5842,N_4046,N_325);
and U5843 (N_5843,N_3902,N_154);
nand U5844 (N_5844,N_4776,N_3452);
and U5845 (N_5845,N_3884,N_4157);
and U5846 (N_5846,N_3430,N_4864);
or U5847 (N_5847,N_3267,N_3694);
nor U5848 (N_5848,N_3755,N_183);
nand U5849 (N_5849,N_1284,N_3381);
xor U5850 (N_5850,N_861,N_1650);
nand U5851 (N_5851,N_1507,N_1467);
nor U5852 (N_5852,N_4787,N_1893);
nand U5853 (N_5853,N_3229,N_2150);
nand U5854 (N_5854,N_4212,N_2589);
nor U5855 (N_5855,N_1030,N_1617);
or U5856 (N_5856,N_311,N_2202);
nand U5857 (N_5857,N_4632,N_4129);
nor U5858 (N_5858,N_1594,N_3911);
or U5859 (N_5859,N_2811,N_1384);
nand U5860 (N_5860,N_1408,N_3450);
nor U5861 (N_5861,N_830,N_1692);
and U5862 (N_5862,N_4077,N_3006);
or U5863 (N_5863,N_4286,N_3270);
and U5864 (N_5864,N_2735,N_4662);
and U5865 (N_5865,N_4685,N_1249);
nand U5866 (N_5866,N_4365,N_4092);
nand U5867 (N_5867,N_3246,N_4369);
nand U5868 (N_5868,N_2794,N_1559);
or U5869 (N_5869,N_2584,N_1019);
and U5870 (N_5870,N_874,N_1974);
and U5871 (N_5871,N_1995,N_2216);
and U5872 (N_5872,N_3171,N_3702);
nand U5873 (N_5873,N_852,N_2308);
or U5874 (N_5874,N_4520,N_949);
nor U5875 (N_5875,N_554,N_933);
and U5876 (N_5876,N_2949,N_4876);
nor U5877 (N_5877,N_1463,N_4785);
nand U5878 (N_5878,N_2636,N_3494);
and U5879 (N_5879,N_3334,N_3577);
or U5880 (N_5880,N_4684,N_3634);
nor U5881 (N_5881,N_4599,N_1915);
nand U5882 (N_5882,N_328,N_2576);
nor U5883 (N_5883,N_4087,N_1992);
nor U5884 (N_5884,N_1392,N_4393);
nor U5885 (N_5885,N_3709,N_2079);
nor U5886 (N_5886,N_3295,N_3390);
nor U5887 (N_5887,N_762,N_3296);
nor U5888 (N_5888,N_4252,N_4797);
or U5889 (N_5889,N_1041,N_4671);
and U5890 (N_5890,N_3713,N_4320);
or U5891 (N_5891,N_1667,N_3486);
and U5892 (N_5892,N_2804,N_2129);
or U5893 (N_5893,N_3841,N_2597);
and U5894 (N_5894,N_589,N_3874);
xor U5895 (N_5895,N_2818,N_1375);
nor U5896 (N_5896,N_1314,N_1261);
nand U5897 (N_5897,N_4582,N_4189);
and U5898 (N_5898,N_2925,N_1488);
or U5899 (N_5899,N_633,N_3641);
nor U5900 (N_5900,N_4188,N_4143);
nand U5901 (N_5901,N_820,N_2381);
or U5902 (N_5902,N_2280,N_200);
nand U5903 (N_5903,N_103,N_738);
and U5904 (N_5904,N_1789,N_2507);
nor U5905 (N_5905,N_3201,N_2247);
nor U5906 (N_5906,N_837,N_4741);
nor U5907 (N_5907,N_2186,N_782);
nor U5908 (N_5908,N_3871,N_2380);
nor U5909 (N_5909,N_2509,N_1040);
nand U5910 (N_5910,N_889,N_4584);
and U5911 (N_5911,N_1012,N_1377);
nand U5912 (N_5912,N_2210,N_221);
nand U5913 (N_5913,N_306,N_1887);
or U5914 (N_5914,N_1332,N_1374);
or U5915 (N_5915,N_2737,N_609);
or U5916 (N_5916,N_4823,N_4564);
or U5917 (N_5917,N_3459,N_842);
and U5918 (N_5918,N_4509,N_4319);
and U5919 (N_5919,N_2391,N_152);
nor U5920 (N_5920,N_4998,N_14);
xor U5921 (N_5921,N_1365,N_4769);
or U5922 (N_5922,N_2271,N_3013);
and U5923 (N_5923,N_4388,N_3469);
nand U5924 (N_5924,N_3753,N_2177);
nand U5925 (N_5925,N_2460,N_4202);
nand U5926 (N_5926,N_796,N_4126);
nand U5927 (N_5927,N_2923,N_279);
nand U5928 (N_5928,N_2429,N_714);
nand U5929 (N_5929,N_4636,N_1607);
nand U5930 (N_5930,N_4532,N_3137);
nand U5931 (N_5931,N_3209,N_269);
nor U5932 (N_5932,N_4004,N_3852);
nand U5933 (N_5933,N_2815,N_3653);
and U5934 (N_5934,N_3667,N_447);
nor U5935 (N_5935,N_979,N_4713);
or U5936 (N_5936,N_2934,N_2172);
nor U5937 (N_5937,N_3356,N_4090);
and U5938 (N_5938,N_2715,N_2270);
and U5939 (N_5939,N_4008,N_1404);
and U5940 (N_5940,N_375,N_3513);
and U5941 (N_5941,N_3901,N_3276);
nand U5942 (N_5942,N_3400,N_608);
xnor U5943 (N_5943,N_4055,N_1654);
or U5944 (N_5944,N_2122,N_3938);
nor U5945 (N_5945,N_4160,N_4634);
nor U5946 (N_5946,N_3080,N_2217);
and U5947 (N_5947,N_1118,N_2326);
xor U5948 (N_5948,N_503,N_635);
or U5949 (N_5949,N_3243,N_2047);
nor U5950 (N_5950,N_3869,N_67);
and U5951 (N_5951,N_3039,N_34);
or U5952 (N_5952,N_3994,N_3471);
xnor U5953 (N_5953,N_9,N_3204);
nand U5954 (N_5954,N_2316,N_4860);
or U5955 (N_5955,N_753,N_1685);
nand U5956 (N_5956,N_1156,N_4402);
nand U5957 (N_5957,N_1015,N_1732);
and U5958 (N_5958,N_3885,N_2234);
or U5959 (N_5959,N_316,N_3914);
nand U5960 (N_5960,N_2063,N_523);
or U5961 (N_5961,N_2284,N_3968);
or U5962 (N_5962,N_3930,N_3050);
nand U5963 (N_5963,N_1483,N_3435);
and U5964 (N_5964,N_4119,N_1079);
xor U5965 (N_5965,N_4330,N_718);
nor U5966 (N_5966,N_3045,N_4994);
xnor U5967 (N_5967,N_2807,N_288);
or U5968 (N_5968,N_37,N_1835);
nor U5969 (N_5969,N_2704,N_1809);
nor U5970 (N_5970,N_3681,N_2449);
nor U5971 (N_5971,N_802,N_1924);
nor U5972 (N_5972,N_829,N_895);
and U5973 (N_5973,N_2883,N_2699);
or U5974 (N_5974,N_4058,N_3005);
and U5975 (N_5975,N_2276,N_1553);
or U5976 (N_5976,N_511,N_3623);
nand U5977 (N_5977,N_2069,N_1686);
nor U5978 (N_5978,N_2264,N_3868);
or U5979 (N_5979,N_2103,N_4208);
or U5980 (N_5980,N_4057,N_3536);
and U5981 (N_5981,N_3383,N_546);
nor U5982 (N_5982,N_901,N_2237);
or U5983 (N_5983,N_4900,N_755);
nor U5984 (N_5984,N_3308,N_556);
and U5985 (N_5985,N_3616,N_2759);
nand U5986 (N_5986,N_3617,N_4000);
nor U5987 (N_5987,N_3626,N_1250);
or U5988 (N_5988,N_2754,N_2327);
nand U5989 (N_5989,N_4443,N_1578);
or U5990 (N_5990,N_601,N_3169);
and U5991 (N_5991,N_2698,N_3102);
and U5992 (N_5992,N_1621,N_1669);
or U5993 (N_5993,N_4355,N_4710);
nor U5994 (N_5994,N_4507,N_116);
nand U5995 (N_5995,N_1248,N_2861);
or U5996 (N_5996,N_4465,N_3197);
nand U5997 (N_5997,N_4481,N_4082);
or U5998 (N_5998,N_3280,N_2390);
or U5999 (N_5999,N_2774,N_3568);
xor U6000 (N_6000,N_157,N_4280);
and U6001 (N_6001,N_1969,N_2798);
or U6002 (N_6002,N_2820,N_4224);
nor U6003 (N_6003,N_3763,N_924);
nand U6004 (N_6004,N_2306,N_1145);
or U6005 (N_6005,N_1306,N_4768);
nor U6006 (N_6006,N_400,N_4028);
or U6007 (N_6007,N_3769,N_3517);
and U6008 (N_6008,N_3920,N_4102);
nor U6009 (N_6009,N_3650,N_2338);
or U6010 (N_6010,N_3081,N_3118);
nand U6011 (N_6011,N_4045,N_2772);
xor U6012 (N_6012,N_496,N_3115);
xnor U6013 (N_6013,N_2463,N_1764);
nor U6014 (N_6014,N_3391,N_2497);
nand U6015 (N_6015,N_2226,N_2029);
nor U6016 (N_6016,N_4658,N_3818);
and U6017 (N_6017,N_1712,N_4331);
xor U6018 (N_6018,N_3040,N_1022);
nor U6019 (N_6019,N_4403,N_1072);
or U6020 (N_6020,N_211,N_210);
or U6021 (N_6021,N_3387,N_3849);
or U6022 (N_6022,N_4318,N_2295);
and U6023 (N_6023,N_3023,N_1920);
xor U6024 (N_6024,N_2139,N_4570);
and U6025 (N_6025,N_4110,N_2771);
or U6026 (N_6026,N_1103,N_3881);
nor U6027 (N_6027,N_3176,N_2072);
xnor U6028 (N_6028,N_2230,N_1159);
nand U6029 (N_6029,N_4609,N_384);
and U6030 (N_6030,N_324,N_2409);
nand U6031 (N_6031,N_4957,N_208);
or U6032 (N_6032,N_2791,N_4493);
nor U6033 (N_6033,N_2633,N_3836);
nor U6034 (N_6034,N_4932,N_3567);
xor U6035 (N_6035,N_4871,N_853);
nand U6036 (N_6036,N_1354,N_2929);
or U6037 (N_6037,N_265,N_1587);
or U6038 (N_6038,N_3426,N_877);
and U6039 (N_6039,N_3927,N_4411);
and U6040 (N_6040,N_3984,N_4332);
xor U6041 (N_6041,N_2866,N_2026);
xnor U6042 (N_6042,N_4213,N_163);
or U6043 (N_6043,N_4277,N_2015);
or U6044 (N_6044,N_3134,N_236);
nand U6045 (N_6045,N_3211,N_438);
nand U6046 (N_6046,N_4450,N_2263);
nor U6047 (N_6047,N_1260,N_1212);
nor U6048 (N_6048,N_3727,N_2009);
or U6049 (N_6049,N_1738,N_3422);
nand U6050 (N_6050,N_4680,N_4904);
nor U6051 (N_6051,N_4540,N_336);
and U6052 (N_6052,N_4487,N_884);
and U6053 (N_6053,N_1112,N_1163);
or U6054 (N_6054,N_297,N_1976);
nor U6055 (N_6055,N_3104,N_1501);
or U6056 (N_6056,N_1791,N_4346);
nor U6057 (N_6057,N_3073,N_458);
nor U6058 (N_6058,N_500,N_3592);
and U6059 (N_6059,N_1018,N_4778);
nor U6060 (N_6060,N_2088,N_4605);
or U6061 (N_6061,N_2178,N_2522);
and U6062 (N_6062,N_102,N_946);
or U6063 (N_6063,N_2666,N_3300);
and U6064 (N_6064,N_3202,N_3893);
nand U6065 (N_6065,N_4317,N_613);
nor U6066 (N_6066,N_2147,N_2206);
nor U6067 (N_6067,N_1432,N_2453);
or U6068 (N_6068,N_71,N_942);
and U6069 (N_6069,N_4489,N_1393);
nor U6070 (N_6070,N_3793,N_3760);
or U6071 (N_6071,N_178,N_4001);
nor U6072 (N_6072,N_1958,N_1076);
and U6073 (N_6073,N_1583,N_3866);
or U6074 (N_6074,N_4854,N_2652);
and U6075 (N_6075,N_156,N_666);
nand U6076 (N_6076,N_2960,N_227);
or U6077 (N_6077,N_876,N_2467);
or U6078 (N_6078,N_1666,N_1978);
or U6079 (N_6079,N_129,N_1853);
or U6080 (N_6080,N_2755,N_3389);
nor U6081 (N_6081,N_923,N_1895);
nand U6082 (N_6082,N_2287,N_3096);
and U6083 (N_6083,N_4760,N_4261);
nor U6084 (N_6084,N_1512,N_1524);
nor U6085 (N_6085,N_2549,N_2323);
nor U6086 (N_6086,N_3482,N_2998);
xor U6087 (N_6087,N_1897,N_1534);
or U6088 (N_6088,N_3918,N_833);
or U6089 (N_6089,N_23,N_3107);
or U6090 (N_6090,N_3563,N_92);
nand U6091 (N_6091,N_3044,N_1874);
nor U6092 (N_6092,N_237,N_144);
xnor U6093 (N_6093,N_3785,N_2741);
nor U6094 (N_6094,N_1464,N_2056);
nor U6095 (N_6095,N_2126,N_3585);
nor U6096 (N_6096,N_1366,N_2416);
and U6097 (N_6097,N_2442,N_2254);
nor U6098 (N_6098,N_3640,N_3312);
nor U6099 (N_6099,N_1625,N_965);
nand U6100 (N_6100,N_230,N_1917);
and U6101 (N_6101,N_2192,N_191);
and U6102 (N_6102,N_4392,N_2138);
nor U6103 (N_6103,N_1003,N_3684);
nand U6104 (N_6104,N_1168,N_4530);
or U6105 (N_6105,N_4343,N_947);
nor U6106 (N_6106,N_4818,N_4935);
xor U6107 (N_6107,N_3863,N_4011);
nand U6108 (N_6108,N_1628,N_1949);
and U6109 (N_6109,N_3004,N_903);
nor U6110 (N_6110,N_2946,N_683);
and U6111 (N_6111,N_1884,N_4588);
nor U6112 (N_6112,N_3289,N_813);
and U6113 (N_6113,N_1334,N_1047);
or U6114 (N_6114,N_1794,N_262);
and U6115 (N_6115,N_1132,N_2036);
nand U6116 (N_6116,N_1858,N_1051);
or U6117 (N_6117,N_3522,N_3436);
nor U6118 (N_6118,N_624,N_2926);
and U6119 (N_6119,N_3304,N_3067);
nand U6120 (N_6120,N_1271,N_4946);
and U6121 (N_6121,N_199,N_1797);
nor U6122 (N_6122,N_4523,N_4834);
nand U6123 (N_6123,N_437,N_4656);
or U6124 (N_6124,N_4552,N_2528);
nor U6125 (N_6125,N_2680,N_2676);
nor U6126 (N_6126,N_3088,N_2488);
or U6127 (N_6127,N_145,N_2011);
or U6128 (N_6128,N_1739,N_4688);
nand U6129 (N_6129,N_2598,N_61);
or U6130 (N_6130,N_3941,N_359);
xor U6131 (N_6131,N_3410,N_3636);
nand U6132 (N_6132,N_3854,N_4984);
or U6133 (N_6133,N_3820,N_2171);
nand U6134 (N_6134,N_712,N_3464);
and U6135 (N_6135,N_3061,N_902);
nand U6136 (N_6136,N_341,N_4511);
nor U6137 (N_6137,N_391,N_834);
and U6138 (N_6138,N_3493,N_1169);
or U6139 (N_6139,N_1940,N_1492);
and U6140 (N_6140,N_778,N_1229);
xor U6141 (N_6141,N_547,N_371);
and U6142 (N_6142,N_2176,N_2045);
nand U6143 (N_6143,N_2322,N_3153);
nor U6144 (N_6144,N_2349,N_4296);
xnor U6145 (N_6145,N_1329,N_4761);
or U6146 (N_6146,N_4694,N_1891);
and U6147 (N_6147,N_1477,N_2969);
nor U6148 (N_6148,N_277,N_4895);
nor U6149 (N_6149,N_4333,N_2369);
or U6150 (N_6150,N_2612,N_764);
nand U6151 (N_6151,N_194,N_253);
nand U6152 (N_6152,N_3358,N_1458);
nand U6153 (N_6153,N_2832,N_3990);
nand U6154 (N_6154,N_870,N_2886);
and U6155 (N_6155,N_4025,N_3398);
nand U6156 (N_6156,N_815,N_1482);
and U6157 (N_6157,N_1845,N_1873);
nor U6158 (N_6158,N_2303,N_4716);
and U6159 (N_6159,N_160,N_4525);
xor U6160 (N_6160,N_3119,N_2376);
nand U6161 (N_6161,N_2331,N_3688);
nor U6162 (N_6162,N_2972,N_2620);
or U6163 (N_6163,N_4897,N_4950);
nor U6164 (N_6164,N_1038,N_3637);
xor U6165 (N_6165,N_2781,N_4941);
nand U6166 (N_6166,N_2275,N_209);
nor U6167 (N_6167,N_2075,N_4954);
nor U6168 (N_6168,N_3433,N_4723);
xnor U6169 (N_6169,N_1982,N_2540);
xnor U6170 (N_6170,N_50,N_2942);
nor U6171 (N_6171,N_4866,N_468);
and U6172 (N_6172,N_2890,N_794);
or U6173 (N_6173,N_1715,N_1597);
and U6174 (N_6174,N_2723,N_2538);
nand U6175 (N_6175,N_537,N_3695);
nand U6176 (N_6176,N_951,N_4175);
or U6177 (N_6177,N_1353,N_3388);
nor U6178 (N_6178,N_925,N_1702);
nor U6179 (N_6179,N_1983,N_1214);
nor U6180 (N_6180,N_867,N_893);
nand U6181 (N_6181,N_1143,N_1799);
nand U6182 (N_6182,N_804,N_3068);
or U6183 (N_6183,N_2833,N_409);
and U6184 (N_6184,N_2022,N_4476);
nand U6185 (N_6185,N_1510,N_3512);
and U6186 (N_6186,N_2136,N_2476);
and U6187 (N_6187,N_214,N_4661);
and U6188 (N_6188,N_4921,N_3953);
or U6189 (N_6189,N_2561,N_1683);
nand U6190 (N_6190,N_3142,N_4036);
and U6191 (N_6191,N_3842,N_2789);
or U6192 (N_6192,N_151,N_4265);
nor U6193 (N_6193,N_2780,N_3583);
xor U6194 (N_6194,N_566,N_3510);
nand U6195 (N_6195,N_3339,N_3501);
and U6196 (N_6196,N_3839,N_2145);
or U6197 (N_6197,N_4471,N_17);
xor U6198 (N_6198,N_2492,N_234);
and U6199 (N_6199,N_424,N_3314);
xnor U6200 (N_6200,N_3733,N_2352);
or U6201 (N_6201,N_2822,N_1139);
or U6202 (N_6202,N_973,N_4644);
and U6203 (N_6203,N_2803,N_3844);
nor U6204 (N_6204,N_2581,N_1836);
and U6205 (N_6205,N_1918,N_2053);
or U6206 (N_6206,N_4137,N_3251);
nor U6207 (N_6207,N_1023,N_4626);
xor U6208 (N_6208,N_4780,N_4750);
nor U6209 (N_6209,N_2511,N_4851);
and U6210 (N_6210,N_2,N_787);
xnor U6211 (N_6211,N_3996,N_4545);
nor U6212 (N_6212,N_106,N_4699);
nor U6213 (N_6213,N_4541,N_3690);
and U6214 (N_6214,N_4104,N_2591);
nor U6215 (N_6215,N_2169,N_1455);
or U6216 (N_6216,N_2038,N_824);
nor U6217 (N_6217,N_370,N_665);
or U6218 (N_6218,N_1998,N_2658);
and U6219 (N_6219,N_3379,N_4531);
and U6220 (N_6220,N_1844,N_3896);
xor U6221 (N_6221,N_3853,N_1194);
nor U6222 (N_6222,N_3263,N_3455);
and U6223 (N_6223,N_4861,N_3327);
nand U6224 (N_6224,N_3320,N_2330);
nor U6225 (N_6225,N_2222,N_3805);
nand U6226 (N_6226,N_848,N_4601);
and U6227 (N_6227,N_3316,N_155);
nand U6228 (N_6228,N_1911,N_4276);
nor U6229 (N_6229,N_4687,N_3497);
nand U6230 (N_6230,N_4228,N_2342);
or U6231 (N_6231,N_4902,N_3923);
or U6232 (N_6232,N_4802,N_1962);
nor U6233 (N_6233,N_1311,N_1538);
nand U6234 (N_6234,N_2204,N_3647);
nand U6235 (N_6235,N_1741,N_1771);
nand U6236 (N_6236,N_2484,N_716);
nand U6237 (N_6237,N_3679,N_875);
or U6238 (N_6238,N_4791,N_2187);
nand U6239 (N_6239,N_1806,N_1703);
nand U6240 (N_6240,N_3245,N_4361);
nand U6241 (N_6241,N_2227,N_636);
nor U6242 (N_6242,N_4123,N_3186);
and U6243 (N_6243,N_2717,N_1831);
nand U6244 (N_6244,N_4062,N_990);
xnor U6245 (N_6245,N_1787,N_1931);
nor U6246 (N_6246,N_3066,N_704);
and U6247 (N_6247,N_412,N_1523);
nor U6248 (N_6248,N_4233,N_3362);
and U6249 (N_6249,N_4910,N_911);
and U6250 (N_6250,N_3190,N_2558);
nand U6251 (N_6251,N_3652,N_978);
nand U6252 (N_6252,N_4405,N_2314);
nor U6253 (N_6253,N_4533,N_4268);
xor U6254 (N_6254,N_82,N_677);
and U6255 (N_6255,N_3406,N_4782);
nand U6256 (N_6256,N_648,N_4311);
and U6257 (N_6257,N_4467,N_1867);
nand U6258 (N_6258,N_686,N_832);
nor U6259 (N_6259,N_4947,N_4108);
or U6260 (N_6260,N_1555,N_1802);
and U6261 (N_6261,N_2932,N_984);
xnor U6262 (N_6262,N_4892,N_3313);
or U6263 (N_6263,N_3575,N_1532);
nand U6264 (N_6264,N_1133,N_1443);
nor U6265 (N_6265,N_179,N_1010);
nor U6266 (N_6266,N_108,N_3326);
nor U6267 (N_6267,N_1549,N_1009);
or U6268 (N_6268,N_2849,N_2301);
xor U6269 (N_6269,N_1416,N_238);
and U6270 (N_6270,N_4647,N_1166);
nor U6271 (N_6271,N_1336,N_1779);
nand U6272 (N_6272,N_4657,N_3511);
nor U6273 (N_6273,N_1493,N_2498);
nor U6274 (N_6274,N_1745,N_3882);
and U6275 (N_6275,N_2494,N_1711);
and U6276 (N_6276,N_885,N_483);
and U6277 (N_6277,N_477,N_1127);
or U6278 (N_6278,N_3405,N_3241);
and U6279 (N_6279,N_3172,N_858);
xnor U6280 (N_6280,N_4640,N_2720);
nand U6281 (N_6281,N_3151,N_1237);
or U6282 (N_6282,N_1933,N_397);
nand U6283 (N_6283,N_2957,N_1192);
xnor U6284 (N_6284,N_2311,N_4245);
and U6285 (N_6285,N_1902,N_2481);
xnor U6286 (N_6286,N_3826,N_967);
and U6287 (N_6287,N_4347,N_1007);
xnor U6288 (N_6288,N_2512,N_2383);
or U6289 (N_6289,N_1363,N_46);
nor U6290 (N_6290,N_224,N_3950);
xor U6291 (N_6291,N_1339,N_1489);
nor U6292 (N_6292,N_2398,N_1777);
or U6293 (N_6293,N_1572,N_231);
nor U6294 (N_6294,N_3525,N_446);
and U6295 (N_6295,N_1302,N_1177);
and U6296 (N_6296,N_4502,N_1052);
and U6297 (N_6297,N_3148,N_1310);
or U6298 (N_6298,N_3461,N_1089);
nand U6299 (N_6299,N_4931,N_1364);
nand U6300 (N_6300,N_651,N_70);
nor U6301 (N_6301,N_2418,N_4259);
nand U6302 (N_6302,N_4966,N_3124);
nand U6303 (N_6303,N_3910,N_1383);
nor U6304 (N_6304,N_4986,N_2272);
xnor U6305 (N_6305,N_3934,N_3646);
or U6306 (N_6306,N_286,N_1744);
nor U6307 (N_6307,N_1875,N_389);
and U6308 (N_6308,N_2286,N_1282);
nand U6309 (N_6309,N_4600,N_1013);
xnor U6310 (N_6310,N_4814,N_1213);
nor U6311 (N_6311,N_3633,N_3165);
or U6312 (N_6312,N_2100,N_845);
and U6313 (N_6313,N_3064,N_4772);
nor U6314 (N_6314,N_3281,N_1916);
and U6315 (N_6315,N_784,N_2123);
xnor U6316 (N_6316,N_1577,N_3630);
nor U6317 (N_6317,N_4563,N_980);
nor U6318 (N_6318,N_4549,N_4887);
and U6319 (N_6319,N_4154,N_3018);
nor U6320 (N_6320,N_2012,N_1913);
nand U6321 (N_6321,N_637,N_4612);
or U6322 (N_6322,N_2001,N_2133);
nand U6323 (N_6323,N_740,N_1435);
xnor U6324 (N_6324,N_4812,N_3499);
or U6325 (N_6325,N_1631,N_2317);
and U6326 (N_6326,N_1936,N_4219);
and U6327 (N_6327,N_746,N_1246);
nand U6328 (N_6328,N_3113,N_2422);
and U6329 (N_6329,N_937,N_3530);
and U6330 (N_6330,N_1446,N_2520);
nand U6331 (N_6331,N_1152,N_459);
or U6332 (N_6332,N_1053,N_1614);
nor U6333 (N_6333,N_3226,N_2140);
nor U6334 (N_6334,N_1430,N_268);
and U6335 (N_6335,N_3978,N_2691);
and U6336 (N_6336,N_887,N_652);
xnor U6337 (N_6337,N_2778,N_4974);
nor U6338 (N_6338,N_565,N_1405);
xor U6339 (N_6339,N_318,N_1146);
and U6340 (N_6340,N_4470,N_3325);
nor U6341 (N_6341,N_3928,N_3505);
nor U6342 (N_6342,N_4765,N_4326);
nor U6343 (N_6343,N_4690,N_3601);
and U6344 (N_6344,N_2078,N_2246);
nand U6345 (N_6345,N_1086,N_3227);
nor U6346 (N_6346,N_799,N_457);
and U6347 (N_6347,N_383,N_4081);
or U6348 (N_6348,N_244,N_2880);
xnor U6349 (N_6349,N_3491,N_410);
xnor U6350 (N_6350,N_4495,N_131);
xor U6351 (N_6351,N_3348,N_1276);
or U6352 (N_6352,N_1417,N_1662);
nand U6353 (N_6353,N_4836,N_2005);
nand U6354 (N_6354,N_4432,N_2262);
nand U6355 (N_6355,N_1240,N_3132);
or U6356 (N_6356,N_4445,N_171);
nand U6357 (N_6357,N_3413,N_836);
and U6358 (N_6358,N_4655,N_1986);
or U6359 (N_6359,N_4204,N_3432);
or U6360 (N_6360,N_3264,N_345);
nand U6361 (N_6361,N_664,N_2910);
or U6362 (N_6362,N_3748,N_162);
xnor U6363 (N_6363,N_2117,N_190);
or U6364 (N_6364,N_1516,N_3622);
nor U6365 (N_6365,N_3173,N_1315);
or U6366 (N_6366,N_3781,N_1601);
nand U6367 (N_6367,N_4628,N_4002);
and U6368 (N_6368,N_1137,N_42);
nor U6369 (N_6369,N_944,N_4099);
nor U6370 (N_6370,N_1498,N_1029);
nand U6371 (N_6371,N_241,N_3086);
nand U6372 (N_6372,N_1317,N_2870);
nor U6373 (N_6373,N_118,N_1618);
and U6374 (N_6374,N_4488,N_1768);
nand U6375 (N_6375,N_2999,N_4360);
nor U6376 (N_6376,N_2670,N_2229);
and U6377 (N_6377,N_2090,N_4181);
or U6378 (N_6378,N_3657,N_2646);
or U6379 (N_6379,N_101,N_1226);
or U6380 (N_6380,N_1465,N_4825);
nand U6381 (N_6381,N_3608,N_4855);
or U6382 (N_6382,N_4521,N_2810);
nor U6383 (N_6383,N_43,N_4328);
nand U6384 (N_6384,N_215,N_1322);
xnor U6385 (N_6385,N_1539,N_3935);
nand U6386 (N_6386,N_2836,N_113);
nand U6387 (N_6387,N_2266,N_1622);
and U6388 (N_6388,N_4107,N_3166);
or U6389 (N_6389,N_4164,N_3409);
or U6390 (N_6390,N_3997,N_2431);
nor U6391 (N_6391,N_1170,N_2888);
and U6392 (N_6392,N_1503,N_1021);
nor U6393 (N_6393,N_4863,N_2564);
nand U6394 (N_6394,N_744,N_3790);
nor U6395 (N_6395,N_4637,N_588);
xor U6396 (N_6396,N_228,N_4586);
nor U6397 (N_6397,N_1343,N_2164);
nand U6398 (N_6398,N_4250,N_2039);
and U6399 (N_6399,N_3580,N_337);
nor U6400 (N_6400,N_4585,N_4988);
nand U6401 (N_6401,N_3556,N_4279);
nor U6402 (N_6402,N_4059,N_1513);
or U6403 (N_6403,N_1638,N_632);
nor U6404 (N_6404,N_2767,N_3317);
and U6405 (N_6405,N_2496,N_196);
and U6406 (N_6406,N_2689,N_407);
nand U6407 (N_6407,N_549,N_4491);
and U6408 (N_6408,N_1291,N_1442);
or U6409 (N_6409,N_4548,N_2291);
or U6410 (N_6410,N_4321,N_2459);
or U6411 (N_6411,N_1151,N_3236);
xor U6412 (N_6412,N_868,N_3123);
nand U6413 (N_6413,N_2930,N_3140);
nor U6414 (N_6414,N_4437,N_1733);
and U6415 (N_6415,N_2677,N_4053);
nand U6416 (N_6416,N_3877,N_3473);
nor U6417 (N_6417,N_117,N_2740);
or U6418 (N_6418,N_1412,N_174);
nor U6419 (N_6419,N_1639,N_4478);
and U6420 (N_6420,N_3925,N_780);
nand U6421 (N_6421,N_1338,N_2135);
and U6422 (N_6422,N_4400,N_3806);
nand U6423 (N_6423,N_3,N_2091);
and U6424 (N_6424,N_4960,N_816);
or U6425 (N_6425,N_792,N_3481);
or U6426 (N_6426,N_1233,N_3214);
xnor U6427 (N_6427,N_2339,N_2747);
nor U6428 (N_6428,N_3776,N_2748);
xor U6429 (N_6429,N_20,N_3170);
xor U6430 (N_6430,N_1906,N_676);
nand U6431 (N_6431,N_1829,N_4173);
or U6432 (N_6432,N_4421,N_2060);
and U6433 (N_6433,N_3298,N_2104);
nand U6434 (N_6434,N_3731,N_4253);
nand U6435 (N_6435,N_307,N_2215);
and U6436 (N_6436,N_4503,N_3206);
nor U6437 (N_6437,N_3613,N_4307);
and U6438 (N_6438,N_486,N_4015);
nor U6439 (N_6439,N_40,N_2195);
and U6440 (N_6440,N_4283,N_671);
or U6441 (N_6441,N_605,N_4071);
or U6442 (N_6442,N_1899,N_1921);
nand U6443 (N_6443,N_3017,N_3810);
nor U6444 (N_6444,N_849,N_4841);
nor U6445 (N_6445,N_4029,N_3128);
nand U6446 (N_6446,N_2638,N_732);
nor U6447 (N_6447,N_1293,N_1558);
and U6448 (N_6448,N_488,N_1784);
nand U6449 (N_6449,N_4951,N_36);
or U6450 (N_6450,N_2700,N_1165);
nor U6451 (N_6451,N_247,N_1634);
nand U6452 (N_6452,N_3734,N_3087);
nor U6453 (N_6453,N_1244,N_577);
xor U6454 (N_6454,N_4709,N_912);
or U6455 (N_6455,N_4972,N_2745);
and U6456 (N_6456,N_4859,N_3765);
nand U6457 (N_6457,N_130,N_4943);
or U6458 (N_6458,N_3193,N_2517);
nand U6459 (N_6459,N_2743,N_4223);
xnor U6460 (N_6460,N_3949,N_347);
xnor U6461 (N_6461,N_1206,N_2399);
or U6462 (N_6462,N_3774,N_509);
nand U6463 (N_6463,N_2845,N_4394);
nor U6464 (N_6464,N_3786,N_2615);
and U6465 (N_6465,N_1055,N_2309);
xnor U6466 (N_6466,N_4134,N_1773);
and U6467 (N_6467,N_1011,N_2876);
and U6468 (N_6468,N_4364,N_181);
and U6469 (N_6469,N_2424,N_3181);
nor U6470 (N_6470,N_4745,N_1141);
or U6471 (N_6471,N_729,N_1852);
and U6472 (N_6472,N_1848,N_2414);
nor U6473 (N_6473,N_411,N_3546);
and U6474 (N_6474,N_3125,N_1425);
and U6475 (N_6475,N_3057,N_3282);
and U6476 (N_6476,N_66,N_1928);
or U6477 (N_6477,N_3112,N_1219);
nor U6478 (N_6478,N_4920,N_1441);
nor U6479 (N_6479,N_4235,N_4366);
or U6480 (N_6480,N_3551,N_3027);
xor U6481 (N_6481,N_3926,N_2769);
nor U6482 (N_6482,N_2707,N_2110);
nor U6483 (N_6483,N_4944,N_2203);
and U6484 (N_6484,N_2443,N_481);
nor U6485 (N_6485,N_4890,N_4187);
and U6486 (N_6486,N_939,N_3845);
and U6487 (N_6487,N_4567,N_3053);
xnor U6488 (N_6488,N_2116,N_303);
xnor U6489 (N_6489,N_611,N_2220);
nor U6490 (N_6490,N_1599,N_654);
nor U6491 (N_6491,N_3349,N_1090);
or U6492 (N_6492,N_2382,N_4536);
and U6493 (N_6493,N_935,N_855);
nand U6494 (N_6494,N_863,N_1783);
nand U6495 (N_6495,N_4167,N_3480);
nor U6496 (N_6496,N_1533,N_4030);
and U6497 (N_6497,N_1515,N_4284);
or U6498 (N_6498,N_1346,N_2994);
nand U6499 (N_6499,N_3602,N_3696);
nor U6500 (N_6500,N_2268,N_4560);
xor U6501 (N_6501,N_1259,N_3034);
nor U6502 (N_6502,N_1843,N_4415);
and U6503 (N_6503,N_2290,N_2594);
or U6504 (N_6504,N_1673,N_3376);
or U6505 (N_6505,N_3976,N_2779);
nor U6506 (N_6506,N_748,N_4801);
or U6507 (N_6507,N_943,N_1660);
nand U6508 (N_6508,N_1761,N_4201);
nand U6509 (N_6509,N_1297,N_1304);
xor U6510 (N_6510,N_3605,N_2017);
or U6511 (N_6511,N_1115,N_2260);
nand U6512 (N_6512,N_1604,N_3164);
nand U6513 (N_6513,N_906,N_2451);
nor U6514 (N_6514,N_494,N_894);
nor U6515 (N_6515,N_3026,N_3939);
nand U6516 (N_6516,N_4569,N_2249);
or U6517 (N_6517,N_443,N_3677);
nor U6518 (N_6518,N_4474,N_534);
and U6519 (N_6519,N_1394,N_1049);
or U6520 (N_6520,N_3948,N_2235);
nand U6521 (N_6521,N_2278,N_568);
or U6522 (N_6522,N_187,N_640);
nor U6523 (N_6523,N_4007,N_3900);
nand U6524 (N_6524,N_2351,N_4598);
nor U6525 (N_6525,N_2684,N_1256);
or U6526 (N_6526,N_4418,N_4414);
nand U6527 (N_6527,N_1965,N_1283);
nand U6528 (N_6528,N_4959,N_2454);
and U6529 (N_6529,N_2678,N_1630);
xor U6530 (N_6530,N_1232,N_3589);
nand U6531 (N_6531,N_4153,N_4422);
or U6532 (N_6532,N_2374,N_3891);
nor U6533 (N_6533,N_2385,N_3965);
or U6534 (N_6534,N_2333,N_4652);
or U6535 (N_6535,N_2982,N_1111);
or U6536 (N_6536,N_4926,N_4229);
nand U6537 (N_6537,N_3205,N_1485);
or U6538 (N_6538,N_1207,N_4794);
or U6539 (N_6539,N_218,N_4995);
and U6540 (N_6540,N_2058,N_4698);
and U6541 (N_6541,N_2793,N_3049);
nor U6542 (N_6542,N_2396,N_2282);
nor U6543 (N_6543,N_300,N_2986);
or U6544 (N_6544,N_505,N_1989);
nor U6545 (N_6545,N_4271,N_3932);
nor U6546 (N_6546,N_1963,N_1699);
nand U6547 (N_6547,N_4447,N_4697);
nor U6548 (N_6548,N_2588,N_4830);
nand U6549 (N_6549,N_4218,N_1036);
nand U6550 (N_6550,N_2084,N_1100);
or U6551 (N_6551,N_4006,N_1645);
or U6552 (N_6552,N_3835,N_2573);
nor U6553 (N_6553,N_3778,N_3344);
nor U6554 (N_6554,N_405,N_3329);
nand U6555 (N_6555,N_570,N_3611);
or U6556 (N_6556,N_4282,N_1345);
xor U6557 (N_6557,N_1144,N_1575);
xnor U6558 (N_6558,N_2995,N_1098);
or U6559 (N_6559,N_2980,N_1814);
nor U6560 (N_6560,N_3121,N_4217);
and U6561 (N_6561,N_1347,N_580);
nor U6562 (N_6562,N_3275,N_2656);
and U6563 (N_6563,N_2908,N_4368);
and U6564 (N_6564,N_4826,N_2064);
or U6565 (N_6565,N_2621,N_2614);
nand U6566 (N_6566,N_2624,N_3843);
nand U6567 (N_6567,N_3477,N_3476);
nor U6568 (N_6568,N_3259,N_3330);
and U6569 (N_6569,N_1502,N_4728);
xor U6570 (N_6570,N_379,N_2367);
nand U6571 (N_6571,N_2648,N_4348);
or U6572 (N_6572,N_4615,N_2329);
nor U6573 (N_6573,N_2531,N_519);
nand U6574 (N_6574,N_1205,N_2628);
nor U6575 (N_6575,N_4288,N_3025);
xor U6576 (N_6576,N_4463,N_2427);
nor U6577 (N_6577,N_1653,N_3466);
and U6578 (N_6578,N_3570,N_1303);
xor U6579 (N_6579,N_4412,N_1663);
and U6580 (N_6580,N_1234,N_1295);
and U6581 (N_6581,N_4338,N_4645);
and U6582 (N_6582,N_3353,N_3465);
nand U6583 (N_6583,N_4176,N_742);
nand U6584 (N_6584,N_4485,N_3069);
and U6585 (N_6585,N_1107,N_1254);
nor U6586 (N_6586,N_3058,N_1546);
xor U6587 (N_6587,N_1828,N_2146);
or U6588 (N_6588,N_4749,N_4538);
nor U6589 (N_6589,N_4434,N_822);
or U6590 (N_6590,N_3462,N_1149);
nand U6591 (N_6591,N_1943,N_1898);
or U6592 (N_6592,N_4808,N_1071);
nor U6593 (N_6593,N_1742,N_4442);
nand U6594 (N_6594,N_4581,N_1679);
nor U6595 (N_6595,N_703,N_376);
and U6596 (N_6596,N_812,N_159);
nor U6597 (N_6597,N_881,N_3559);
xnor U6598 (N_6598,N_3160,N_2457);
nor U6599 (N_6599,N_1955,N_3751);
and U6600 (N_6600,N_1885,N_1239);
xor U6601 (N_6601,N_2483,N_1178);
xor U6602 (N_6602,N_4047,N_619);
nor U6603 (N_6603,N_4231,N_64);
nand U6604 (N_6604,N_2928,N_864);
nand U6605 (N_6605,N_4596,N_2805);
nor U6606 (N_6606,N_2378,N_1698);
or U6607 (N_6607,N_3438,N_2790);
and U6608 (N_6608,N_1864,N_526);
nand U6609 (N_6609,N_1135,N_2087);
nor U6610 (N_6610,N_420,N_3200);
or U6611 (N_6611,N_4963,N_4804);
nor U6612 (N_6612,N_2008,N_4292);
and U6613 (N_6613,N_3346,N_2898);
and U6614 (N_6614,N_4679,N_2113);
and U6615 (N_6615,N_1584,N_4120);
or U6616 (N_6616,N_1005,N_275);
and U6617 (N_6617,N_1062,N_2685);
xnor U6618 (N_6618,N_2587,N_4788);
or U6619 (N_6619,N_3208,N_3256);
and U6620 (N_6620,N_4992,N_3393);
nand U6621 (N_6621,N_1717,N_2572);
or U6622 (N_6622,N_4973,N_2479);
or U6623 (N_6623,N_222,N_2730);
or U6624 (N_6624,N_435,N_292);
nor U6625 (N_6625,N_107,N_4557);
or U6626 (N_6626,N_2936,N_1102);
nor U6627 (N_6627,N_3959,N_1265);
or U6628 (N_6628,N_2871,N_456);
nand U6629 (N_6629,N_349,N_4824);
and U6630 (N_6630,N_1263,N_3533);
or U6631 (N_6631,N_3758,N_1044);
or U6632 (N_6632,N_2387,N_2605);
and U6633 (N_6633,N_4938,N_4917);
nand U6634 (N_6634,N_1657,N_596);
nor U6635 (N_6635,N_2541,N_340);
or U6636 (N_6636,N_1097,N_828);
nor U6637 (N_6637,N_423,N_4239);
nand U6638 (N_6638,N_169,N_1437);
nor U6639 (N_6639,N_2341,N_797);
and U6640 (N_6640,N_545,N_759);
nor U6641 (N_6641,N_309,N_138);
nand U6642 (N_6642,N_4719,N_4410);
and U6643 (N_6643,N_264,N_4358);
and U6644 (N_6644,N_3847,N_754);
and U6645 (N_6645,N_643,N_567);
nand U6646 (N_6646,N_3628,N_2373);
and U6647 (N_6647,N_1961,N_1640);
xor U6648 (N_6648,N_3671,N_1719);
or U6649 (N_6649,N_3225,N_1747);
or U6650 (N_6650,N_321,N_2107);
and U6651 (N_6651,N_724,N_403);
or U6652 (N_6652,N_3554,N_1816);
nor U6653 (N_6653,N_1894,N_1376);
and U6654 (N_6654,N_2667,N_3689);
nand U6655 (N_6655,N_2574,N_2279);
and U6656 (N_6656,N_3897,N_217);
nor U6657 (N_6657,N_2954,N_4726);
or U6658 (N_6658,N_1765,N_239);
nand U6659 (N_6659,N_3460,N_2525);
nand U6660 (N_6660,N_2829,N_3451);
nor U6661 (N_6661,N_840,N_4243);
or U6662 (N_6662,N_109,N_4444);
nor U6663 (N_6663,N_464,N_4725);
nor U6664 (N_6664,N_4106,N_4908);
nand U6665 (N_6665,N_350,N_2616);
nor U6666 (N_6666,N_362,N_4774);
nand U6667 (N_6667,N_2801,N_958);
and U6668 (N_6668,N_3359,N_3520);
nor U6669 (N_6669,N_4186,N_2293);
and U6670 (N_6670,N_3529,N_242);
nand U6671 (N_6671,N_3447,N_355);
or U6672 (N_6672,N_4236,N_2188);
or U6673 (N_6673,N_1854,N_2073);
nor U6674 (N_6674,N_1185,N_599);
or U6675 (N_6675,N_1349,N_2948);
or U6676 (N_6676,N_2458,N_1350);
nand U6677 (N_6677,N_4608,N_4838);
and U6678 (N_6678,N_3952,N_4752);
nand U6679 (N_6679,N_3848,N_4695);
or U6680 (N_6680,N_1861,N_2634);
nand U6681 (N_6681,N_2448,N_4322);
nor U6682 (N_6682,N_1946,N_332);
nor U6683 (N_6683,N_2343,N_4140);
nor U6684 (N_6684,N_3872,N_789);
and U6685 (N_6685,N_3126,N_921);
nor U6686 (N_6686,N_1187,N_3240);
or U6687 (N_6687,N_2521,N_1487);
nor U6688 (N_6688,N_1262,N_4155);
and U6689 (N_6689,N_4571,N_3544);
nor U6690 (N_6690,N_3468,N_4734);
nand U6691 (N_6691,N_2545,N_3739);
nand U6692 (N_6692,N_2963,N_2784);
xnor U6693 (N_6693,N_1061,N_1434);
nand U6694 (N_6694,N_3823,N_3515);
or U6695 (N_6695,N_3903,N_575);
nor U6696 (N_6696,N_3446,N_591);
nand U6697 (N_6697,N_2211,N_3771);
or U6698 (N_6698,N_2941,N_3307);
or U6699 (N_6699,N_1696,N_1058);
nor U6700 (N_6700,N_2703,N_4537);
xnor U6701 (N_6701,N_3161,N_2904);
nor U6702 (N_6702,N_4975,N_1308);
or U6703 (N_6703,N_515,N_1801);
or U6704 (N_6704,N_4193,N_1004);
and U6705 (N_6705,N_2365,N_3993);
nor U6706 (N_6706,N_401,N_4940);
or U6707 (N_6707,N_1600,N_1438);
xnor U6708 (N_6708,N_1785,N_2590);
nor U6709 (N_6709,N_3010,N_1016);
nor U6710 (N_6710,N_743,N_3552);
nand U6711 (N_6711,N_3824,N_2953);
nand U6712 (N_6712,N_4934,N_12);
nor U6713 (N_6713,N_2931,N_454);
nor U6714 (N_6714,N_1175,N_3309);
nand U6715 (N_6715,N_2128,N_1735);
nor U6716 (N_6716,N_2526,N_1270);
nor U6717 (N_6717,N_3770,N_4209);
or U6718 (N_6718,N_1400,N_3519);
nor U6719 (N_6719,N_1459,N_2281);
and U6720 (N_6720,N_1751,N_2651);
nor U6721 (N_6721,N_4832,N_1);
nand U6722 (N_6722,N_3380,N_2130);
or U6723 (N_6723,N_2105,N_122);
nand U6724 (N_6724,N_2631,N_4461);
nor U6725 (N_6725,N_482,N_3297);
or U6726 (N_6726,N_3565,N_2817);
nor U6727 (N_6727,N_2770,N_2762);
and U6728 (N_6728,N_581,N_1045);
or U6729 (N_6729,N_2555,N_4316);
and U6730 (N_6730,N_2867,N_3144);
or U6731 (N_6731,N_4417,N_2663);
or U6732 (N_6732,N_4468,N_3942);
nand U6733 (N_6733,N_776,N_3759);
nand U6734 (N_6734,N_512,N_2425);
xnor U6735 (N_6735,N_2243,N_4673);
nand U6736 (N_6736,N_3139,N_3807);
or U6737 (N_6737,N_2070,N_4128);
or U6738 (N_6738,N_4613,N_2223);
nand U6739 (N_6739,N_4256,N_1423);
nand U6740 (N_6740,N_272,N_1856);
nand U6741 (N_6741,N_177,N_628);
nor U6742 (N_6742,N_3831,N_4130);
xor U6743 (N_6743,N_4113,N_3538);
and U6744 (N_6744,N_3024,N_1731);
nand U6745 (N_6745,N_4075,N_4517);
xnor U6746 (N_6746,N_4651,N_3315);
nor U6747 (N_6747,N_1752,N_4505);
nand U6748 (N_6748,N_4133,N_2059);
nand U6749 (N_6749,N_4977,N_2853);
nand U6750 (N_6750,N_1966,N_3561);
or U6751 (N_6751,N_1643,N_4244);
and U6752 (N_6752,N_4622,N_3638);
nor U6753 (N_6753,N_3242,N_2673);
and U6754 (N_6754,N_2120,N_408);
nor U6755 (N_6755,N_4848,N_33);
nand U6756 (N_6756,N_518,N_527);
nor U6757 (N_6757,N_4547,N_1279);
and U6758 (N_6758,N_2444,N_1514);
nand U6759 (N_6759,N_4027,N_982);
or U6760 (N_6760,N_623,N_888);
and U6761 (N_6761,N_2221,N_694);
and U6762 (N_6762,N_1981,N_3182);
or U6763 (N_6763,N_4423,N_1059);
nand U6764 (N_6764,N_267,N_1092);
and U6765 (N_6765,N_2076,N_2035);
nor U6766 (N_6766,N_455,N_1652);
xnor U6767 (N_6767,N_3656,N_84);
or U6768 (N_6768,N_2265,N_2102);
nor U6769 (N_6769,N_278,N_1545);
nor U6770 (N_6770,N_1941,N_803);
nor U6771 (N_6771,N_1083,N_1309);
and U6772 (N_6772,N_2389,N_2184);
nand U6773 (N_6773,N_3224,N_2042);
nor U6774 (N_6774,N_4610,N_3399);
or U6775 (N_6775,N_1154,N_2108);
and U6776 (N_6776,N_2239,N_4775);
nand U6777 (N_6777,N_4329,N_2258);
and U6778 (N_6778,N_3441,N_4370);
nand U6779 (N_6779,N_1691,N_1253);
or U6780 (N_6780,N_1905,N_4664);
and U6781 (N_6781,N_1312,N_3111);
xor U6782 (N_6782,N_4602,N_1522);
nand U6783 (N_6783,N_3248,N_1834);
nor U6784 (N_6784,N_100,N_354);
or U6785 (N_6785,N_1195,N_2835);
and U6786 (N_6786,N_1624,N_4882);
and U6787 (N_6787,N_953,N_3705);
nand U6788 (N_6788,N_1325,N_1440);
nand U6789 (N_6789,N_4170,N_2596);
xnor U6790 (N_6790,N_1290,N_4258);
or U6791 (N_6791,N_4915,N_3454);
and U6792 (N_6792,N_3363,N_517);
nor U6793 (N_6793,N_1211,N_2860);
nor U6794 (N_6794,N_1756,N_1672);
and U6795 (N_6795,N_4667,N_2166);
or U6796 (N_6796,N_4715,N_3639);
or U6797 (N_6797,N_604,N_3014);
and U6798 (N_6798,N_4526,N_1947);
nor U6799 (N_6799,N_4981,N_2153);
nor U6800 (N_6800,N_1122,N_3846);
nor U6801 (N_6801,N_1833,N_1812);
or U6802 (N_6802,N_826,N_4387);
nor U6803 (N_6803,N_1460,N_3859);
and U6804 (N_6804,N_89,N_1318);
or U6805 (N_6805,N_3865,N_1838);
nand U6806 (N_6806,N_1900,N_4955);
nand U6807 (N_6807,N_3419,N_3091);
or U6808 (N_6808,N_972,N_2887);
or U6809 (N_6809,N_3079,N_4200);
nand U6810 (N_6810,N_3553,N_4023);
nand U6811 (N_6811,N_4060,N_1179);
nor U6812 (N_6812,N_698,N_4266);
xnor U6813 (N_6813,N_4169,N_593);
nand U6814 (N_6814,N_569,N_2288);
or U6815 (N_6815,N_617,N_4356);
nor U6816 (N_6816,N_3192,N_2595);
nand U6817 (N_6817,N_1267,N_2554);
nand U6818 (N_6818,N_4529,N_4880);
and U6819 (N_6819,N_4078,N_3672);
and U6820 (N_6820,N_3384,N_4238);
nor U6821 (N_6821,N_4572,N_3403);
or U6822 (N_6822,N_2205,N_4246);
nand U6823 (N_6823,N_4985,N_201);
xnor U6824 (N_6824,N_3478,N_2006);
nand U6825 (N_6825,N_2529,N_882);
nor U6826 (N_6826,N_1224,N_572);
xor U6827 (N_6827,N_4561,N_4682);
or U6828 (N_6828,N_3360,N_164);
or U6829 (N_6829,N_3933,N_4846);
nand U6830 (N_6830,N_1230,N_1368);
nor U6831 (N_6831,N_2706,N_4747);
or U6832 (N_6832,N_2978,N_678);
nor U6833 (N_6833,N_1444,N_2933);
and U6834 (N_6834,N_1605,N_2726);
nor U6835 (N_6835,N_2534,N_2951);
nand U6836 (N_6836,N_2580,N_2518);
nand U6837 (N_6837,N_317,N_4287);
and U6838 (N_6838,N_2970,N_3147);
nand U6839 (N_6839,N_3986,N_3879);
nor U6840 (N_6840,N_3654,N_3802);
or U6841 (N_6841,N_2065,N_2917);
nor U6842 (N_6842,N_1094,N_2151);
and U6843 (N_6843,N_1629,N_3385);
and U6844 (N_6844,N_476,N_584);
nor U6845 (N_6845,N_308,N_232);
nor U6846 (N_6846,N_552,N_945);
nand U6847 (N_6847,N_3618,N_4543);
nor U6848 (N_6848,N_3833,N_3729);
and U6849 (N_6849,N_2912,N_4116);
xor U6850 (N_6850,N_4795,N_3071);
nand U6851 (N_6851,N_1203,N_854);
nor U6852 (N_6852,N_2826,N_3215);
nand U6853 (N_6853,N_4374,N_711);
nor U6854 (N_6854,N_501,N_3338);
and U6855 (N_6855,N_1258,N_1466);
and U6856 (N_6856,N_3528,N_3773);
nor U6857 (N_6857,N_299,N_137);
and U6858 (N_6858,N_2905,N_1718);
xor U6859 (N_6859,N_1975,N_393);
and U6860 (N_6860,N_4335,N_3550);
and U6861 (N_6861,N_4301,N_4604);
and U6862 (N_6862,N_4906,N_4809);
and U6863 (N_6863,N_634,N_2395);
nor U6864 (N_6864,N_125,N_3487);
nand U6865 (N_6865,N_1082,N_1328);
nor U6866 (N_6866,N_2099,N_4398);
nor U6867 (N_6867,N_607,N_721);
or U6868 (N_6868,N_485,N_3495);
nand U6869 (N_6869,N_1209,N_4074);
nand U6870 (N_6870,N_1506,N_2544);
or U6871 (N_6871,N_96,N_4297);
nor U6872 (N_6872,N_4534,N_3090);
or U6873 (N_6873,N_960,N_3423);
and U6874 (N_6874,N_733,N_4757);
or U6875 (N_6875,N_3078,N_3560);
and U6876 (N_6876,N_1758,N_3065);
nor U6877 (N_6877,N_3038,N_8);
nand U6878 (N_6878,N_507,N_1627);
xnor U6879 (N_6879,N_1391,N_3625);
nor U6880 (N_6880,N_3995,N_502);
or U6881 (N_6881,N_726,N_2475);
and U6882 (N_6882,N_1161,N_2347);
nor U6883 (N_6883,N_1697,N_19);
or U6884 (N_6884,N_3919,N_2579);
or U6885 (N_6885,N_2027,N_3564);
and U6886 (N_6886,N_1411,N_3361);
nand U6887 (N_6887,N_3285,N_4135);
and U6888 (N_6888,N_3738,N_245);
xor U6889 (N_6889,N_4875,N_4198);
or U6890 (N_6890,N_3342,N_3052);
nand U6891 (N_6891,N_1380,N_4722);
nor U6892 (N_6892,N_3506,N_1541);
nand U6893 (N_6893,N_1580,N_3321);
xor U6894 (N_6894,N_1117,N_1903);
nand U6895 (N_6895,N_1500,N_2175);
and U6896 (N_6896,N_4197,N_219);
or U6897 (N_6897,N_3157,N_3825);
nor U6898 (N_6898,N_471,N_2733);
or U6899 (N_6899,N_3187,N_2563);
xor U6900 (N_6900,N_2179,N_3490);
or U6901 (N_6901,N_1243,N_2938);
or U6902 (N_6902,N_153,N_4514);
nor U6903 (N_6903,N_1371,N_1647);
xnor U6904 (N_6904,N_2112,N_3235);
nor U6905 (N_6905,N_3878,N_79);
nand U6906 (N_6906,N_3056,N_3041);
xnor U6907 (N_6907,N_4573,N_539);
or U6908 (N_6908,N_2644,N_993);
and U6909 (N_6909,N_2927,N_4720);
or U6910 (N_6910,N_850,N_2640);
or U6911 (N_6911,N_3371,N_3982);
or U6912 (N_6912,N_2189,N_3427);
or U6913 (N_6913,N_857,N_3178);
and U6914 (N_6914,N_4779,N_2441);
nor U6915 (N_6915,N_216,N_2546);
nand U6916 (N_6916,N_3095,N_4717);
and U6917 (N_6917,N_1860,N_1626);
or U6918 (N_6918,N_4727,N_2813);
or U6919 (N_6919,N_2165,N_3998);
nand U6920 (N_6920,N_4459,N_466);
nand U6921 (N_6921,N_3274,N_2672);
nand U6922 (N_6922,N_2863,N_3008);
xor U6923 (N_6923,N_2336,N_4323);
xnor U6924 (N_6924,N_578,N_1561);
or U6925 (N_6925,N_1642,N_3887);
nor U6926 (N_6926,N_402,N_3508);
or U6927 (N_6927,N_1511,N_289);
xnor U6928 (N_6928,N_3648,N_2432);
nand U6929 (N_6929,N_2750,N_3595);
xnor U6930 (N_6930,N_10,N_1418);
and U6931 (N_6931,N_1910,N_1054);
nor U6932 (N_6932,N_1542,N_1069);
and U6933 (N_6933,N_3250,N_4692);
and U6934 (N_6934,N_3728,N_2825);
nand U6935 (N_6935,N_1387,N_4472);
or U6936 (N_6936,N_4446,N_2225);
nor U6937 (N_6937,N_421,N_1150);
nor U6938 (N_6938,N_1680,N_4565);
nor U6939 (N_6939,N_2119,N_35);
or U6940 (N_6940,N_2101,N_886);
or U6941 (N_6941,N_4381,N_1602);
nand U6942 (N_6942,N_2377,N_4144);
nor U6943 (N_6943,N_1428,N_1953);
nand U6944 (N_6944,N_4508,N_3747);
or U6945 (N_6945,N_4257,N_2874);
nor U6946 (N_6946,N_3292,N_2403);
and U6947 (N_6947,N_4923,N_3127);
nor U6948 (N_6948,N_1674,N_2695);
nor U6949 (N_6949,N_621,N_167);
or U6950 (N_6950,N_4933,N_2163);
xnor U6951 (N_6951,N_4705,N_3449);
nor U6952 (N_6952,N_7,N_3265);
or U6953 (N_6953,N_2659,N_4225);
nor U6954 (N_6954,N_69,N_3218);
nand U6955 (N_6955,N_1862,N_991);
nand U6956 (N_6956,N_1026,N_205);
nand U6957 (N_6957,N_533,N_2141);
nand U6958 (N_6958,N_3177,N_2125);
xnor U6959 (N_6959,N_1922,N_898);
nand U6960 (N_6960,N_4886,N_452);
xnor U6961 (N_6961,N_2194,N_508);
nor U6962 (N_6962,N_4490,N_2018);
or U6963 (N_6963,N_2756,N_4270);
and U6964 (N_6964,N_781,N_1907);
nor U6965 (N_6965,N_2859,N_915);
or U6966 (N_6966,N_3507,N_865);
and U6967 (N_6967,N_4623,N_357);
nand U6968 (N_6968,N_68,N_188);
or U6969 (N_6969,N_3414,N_2082);
or U6970 (N_6970,N_3642,N_3924);
nand U6971 (N_6971,N_1994,N_114);
nor U6972 (N_6972,N_1066,N_1382);
or U6973 (N_6973,N_6,N_2843);
nor U6974 (N_6974,N_4810,N_3578);
and U6975 (N_6975,N_745,N_839);
and U6976 (N_6976,N_3524,N_3424);
and U6977 (N_6977,N_2426,N_3350);
and U6978 (N_6978,N_2824,N_2802);
nor U6979 (N_6979,N_927,N_1967);
xnor U6980 (N_6980,N_767,N_1070);
nand U6981 (N_6981,N_4816,N_16);
nand U6982 (N_6982,N_2455,N_4755);
nand U6983 (N_6983,N_1934,N_2916);
and U6984 (N_6984,N_1728,N_2397);
nor U6985 (N_6985,N_3569,N_1912);
nand U6986 (N_6986,N_4576,N_1174);
nor U6987 (N_6987,N_2721,N_4042);
nand U6988 (N_6988,N_1296,N_392);
and U6989 (N_6989,N_182,N_763);
and U6990 (N_6990,N_2505,N_3386);
nand U6991 (N_6991,N_1938,N_1197);
and U6992 (N_6992,N_2630,N_4073);
and U6993 (N_6993,N_4822,N_4017);
nor U6994 (N_6994,N_4344,N_553);
and U6995 (N_6995,N_2920,N_1398);
xnor U6996 (N_6996,N_2872,N_1530);
and U6997 (N_6997,N_1886,N_1988);
and U6998 (N_6998,N_185,N_4829);
nand U6999 (N_6999,N_1063,N_4484);
or U7000 (N_7000,N_1108,N_2536);
and U7001 (N_7001,N_204,N_4308);
nand U7002 (N_7002,N_2324,N_4293);
nor U7003 (N_7003,N_3535,N_1217);
xor U7004 (N_7004,N_2152,N_198);
nand U7005 (N_7005,N_2393,N_823);
and U7006 (N_7006,N_2071,N_498);
nand U7007 (N_7007,N_4263,N_4147);
nor U7008 (N_7008,N_4274,N_266);
nand U7009 (N_7009,N_4065,N_13);
xor U7010 (N_7010,N_1772,N_2289);
nand U7011 (N_7011,N_880,N_2255);
and U7012 (N_7012,N_3033,N_1081);
nand U7013 (N_7013,N_2363,N_4614);
nor U7014 (N_7014,N_4773,N_4205);
nand U7015 (N_7015,N_528,N_2642);
nand U7016 (N_7016,N_469,N_1222);
nor U7017 (N_7017,N_4313,N_2547);
or U7018 (N_7018,N_4500,N_3972);
nor U7019 (N_7019,N_256,N_1340);
nor U7020 (N_7020,N_128,N_1658);
nand U7021 (N_7021,N_2298,N_1378);
and U7022 (N_7022,N_4982,N_417);
and U7023 (N_7023,N_4179,N_603);
and U7024 (N_7024,N_2921,N_1327);
nand U7025 (N_7025,N_3855,N_3523);
or U7026 (N_7026,N_1359,N_132);
nand U7027 (N_7027,N_3012,N_988);
xnor U7028 (N_7028,N_3283,N_4518);
and U7029 (N_7029,N_3063,N_4948);
or U7030 (N_7030,N_3488,N_4260);
or U7031 (N_7031,N_679,N_1803);
or U7032 (N_7032,N_2143,N_140);
nand U7033 (N_7033,N_3418,N_1172);
and U7034 (N_7034,N_2889,N_4044);
and U7035 (N_7035,N_2902,N_1320);
nor U7036 (N_7036,N_4796,N_2159);
or U7037 (N_7037,N_530,N_30);
xnor U7038 (N_7038,N_2083,N_1494);
xnor U7039 (N_7039,N_2438,N_4735);
and U7040 (N_7040,N_3228,N_3799);
nand U7041 (N_7041,N_675,N_4700);
or U7042 (N_7042,N_3572,N_3411);
nand U7043 (N_7043,N_2713,N_997);
xor U7044 (N_7044,N_3557,N_3351);
and U7045 (N_7045,N_4706,N_1596);
or U7046 (N_7046,N_3440,N_1611);
and U7047 (N_7047,N_342,N_3042);
nor U7048 (N_7048,N_4150,N_720);
and U7049 (N_7049,N_39,N_995);
or U7050 (N_7050,N_4131,N_2701);
or U7051 (N_7051,N_4898,N_4949);
nor U7052 (N_7052,N_91,N_3905);
or U7053 (N_7053,N_48,N_270);
nand U7054 (N_7054,N_2092,N_1999);
nor U7055 (N_7055,N_2127,N_4624);
xnor U7056 (N_7056,N_4885,N_2668);
xor U7057 (N_7057,N_3644,N_3266);
nor U7058 (N_7058,N_644,N_1585);
nand U7059 (N_7059,N_574,N_4550);
nor U7060 (N_7060,N_2892,N_170);
or U7061 (N_7061,N_2993,N_2328);
nand U7062 (N_7062,N_1508,N_538);
or U7063 (N_7063,N_1871,N_3722);
or U7064 (N_7064,N_388,N_4378);
nand U7065 (N_7065,N_3431,N_2568);
xnor U7066 (N_7066,N_3612,N_4889);
nand U7067 (N_7067,N_2862,N_166);
or U7068 (N_7068,N_3198,N_139);
or U7069 (N_7069,N_4139,N_1292);
nor U7070 (N_7070,N_3966,N_3347);
xnor U7071 (N_7071,N_2144,N_859);
nand U7072 (N_7072,N_475,N_4554);
nand U7073 (N_7073,N_4792,N_3947);
nand U7074 (N_7074,N_104,N_3549);
and U7075 (N_7075,N_4962,N_2575);
nor U7076 (N_7076,N_4764,N_2410);
and U7077 (N_7077,N_3527,N_3545);
and U7078 (N_7078,N_3020,N_1593);
or U7079 (N_7079,N_3800,N_1870);
or U7080 (N_7080,N_2809,N_1095);
nand U7081 (N_7081,N_4151,N_3721);
nand U7082 (N_7082,N_1190,N_1274);
nand U7083 (N_7083,N_2305,N_2966);
or U7084 (N_7084,N_3332,N_1245);
nand U7085 (N_7085,N_3093,N_3685);
and U7086 (N_7086,N_3598,N_3643);
and U7087 (N_7087,N_3951,N_670);
or U7088 (N_7088,N_2535,N_2814);
nand U7089 (N_7089,N_3231,N_2625);
and U7090 (N_7090,N_80,N_1776);
xnor U7091 (N_7091,N_1452,N_290);
xnor U7092 (N_7092,N_1155,N_3009);
and U7093 (N_7093,N_2958,N_3886);
nand U7094 (N_7094,N_3697,N_3331);
and U7095 (N_7095,N_63,N_750);
and U7096 (N_7096,N_1014,N_1620);
and U7097 (N_7097,N_3133,N_1268);
or U7098 (N_7098,N_2639,N_777);
nand U7099 (N_7099,N_1740,N_531);
nand U7100 (N_7100,N_2632,N_98);
nand U7101 (N_7101,N_1896,N_433);
and U7102 (N_7102,N_2731,N_88);
or U7103 (N_7103,N_249,N_4617);
nor U7104 (N_7104,N_1825,N_3715);
nand U7105 (N_7105,N_3343,N_124);
nand U7106 (N_7106,N_2973,N_4718);
or U7107 (N_7107,N_1316,N_3355);
xor U7108 (N_7108,N_1880,N_674);
nor U7109 (N_7109,N_2307,N_414);
and U7110 (N_7110,N_2944,N_709);
nor U7111 (N_7111,N_1574,N_358);
or U7112 (N_7112,N_962,N_478);
or U7113 (N_7113,N_4354,N_1568);
and U7114 (N_7114,N_585,N_24);
xnor U7115 (N_7115,N_4633,N_1028);
and U7116 (N_7116,N_4315,N_3219);
nand U7117 (N_7117,N_83,N_904);
nor U7118 (N_7118,N_28,N_1199);
nand U7119 (N_7119,N_3732,N_1565);
or U7120 (N_7120,N_3412,N_2242);
and U7121 (N_7121,N_1480,N_2240);
or U7122 (N_7122,N_2875,N_331);
nand U7123 (N_7123,N_3114,N_3574);
nor U7124 (N_7124,N_1367,N_2865);
nand U7125 (N_7125,N_4357,N_779);
and U7126 (N_7126,N_3318,N_4556);
xnor U7127 (N_7127,N_928,N_1131);
nand U7128 (N_7128,N_3322,N_2839);
nor U7129 (N_7129,N_4635,N_372);
nand U7130 (N_7130,N_2218,N_4048);
or U7131 (N_7131,N_2023,N_1255);
or U7132 (N_7132,N_4273,N_660);
nand U7133 (N_7133,N_1878,N_4884);
and U7134 (N_7134,N_387,N_918);
nor U7135 (N_7135,N_2470,N_856);
nand U7136 (N_7136,N_2466,N_1659);
xor U7137 (N_7137,N_2364,N_1121);
or U7138 (N_7138,N_1968,N_3890);
or U7139 (N_7139,N_3804,N_1285);
and U7140 (N_7140,N_1227,N_4821);
nor U7141 (N_7141,N_562,N_175);
xnor U7142 (N_7142,N_3943,N_896);
xnor U7143 (N_7143,N_883,N_462);
nand U7144 (N_7144,N_1786,N_805);
and U7145 (N_7145,N_3378,N_97);
and U7146 (N_7146,N_2650,N_1793);
nor U7147 (N_7147,N_1289,N_353);
or U7148 (N_7148,N_4103,N_602);
nand U7149 (N_7149,N_430,N_1612);
and U7150 (N_7150,N_2114,N_1419);
and U7151 (N_7151,N_1700,N_561);
nor U7152 (N_7152,N_2224,N_4668);
nor U7153 (N_7153,N_3514,N_1085);
nand U7154 (N_7154,N_1567,N_4873);
and U7155 (N_7155,N_3906,N_442);
or U7156 (N_7156,N_2469,N_1499);
and U7157 (N_7157,N_3604,N_32);
nand U7158 (N_7158,N_31,N_3489);
nor U7159 (N_7159,N_4499,N_4098);
nor U7160 (N_7160,N_722,N_3223);
nand U7161 (N_7161,N_15,N_2952);
nand U7162 (N_7162,N_2702,N_934);
and U7163 (N_7163,N_4759,N_4711);
nor U7164 (N_7164,N_406,N_2961);
nand U7165 (N_7165,N_3754,N_2854);
nand U7166 (N_7166,N_422,N_706);
xnor U7167 (N_7167,N_4083,N_3961);
and U7168 (N_7168,N_1182,N_4384);
nor U7169 (N_7169,N_2156,N_323);
or U7170 (N_7170,N_543,N_3547);
and U7171 (N_7171,N_931,N_1180);
or U7172 (N_7172,N_734,N_2050);
and U7173 (N_7173,N_3532,N_4010);
and U7174 (N_7174,N_291,N_2967);
nand U7175 (N_7175,N_3960,N_366);
xor U7176 (N_7176,N_3792,N_2051);
nand U7177 (N_7177,N_1709,N_735);
nand U7178 (N_7178,N_1471,N_2510);
nand U7179 (N_7179,N_642,N_4837);
or U7180 (N_7180,N_1119,N_524);
or U7181 (N_7181,N_2968,N_4425);
xnor U7182 (N_7182,N_2118,N_44);
or U7183 (N_7183,N_4171,N_1153);
xnor U7184 (N_7184,N_2577,N_4763);
or U7185 (N_7185,N_3029,N_1031);
or U7186 (N_7186,N_4883,N_4559);
and U7187 (N_7187,N_2981,N_2495);
and U7188 (N_7188,N_22,N_4539);
nor U7189 (N_7189,N_1720,N_2977);
or U7190 (N_7190,N_913,N_1280);
or U7191 (N_7191,N_4965,N_4275);
nand U7192 (N_7192,N_3175,N_360);
nor U7193 (N_7193,N_21,N_416);
nor U7194 (N_7194,N_513,N_2095);
and U7195 (N_7195,N_4619,N_4039);
and U7196 (N_7196,N_4051,N_2094);
and U7197 (N_7197,N_699,N_3470);
nand U7198 (N_7198,N_352,N_4558);
and U7199 (N_7199,N_2174,N_692);
or U7200 (N_7200,N_3199,N_2067);
and U7201 (N_7201,N_668,N_4215);
and U7202 (N_7202,N_3958,N_338);
or U7203 (N_7203,N_3368,N_1421);
nand U7204 (N_7204,N_441,N_4566);
and U7205 (N_7205,N_449,N_1518);
nand U7206 (N_7206,N_639,N_2161);
and U7207 (N_7207,N_4390,N_4111);
nand U7208 (N_7208,N_448,N_3913);
nor U7209 (N_7209,N_3336,N_3788);
or U7210 (N_7210,N_260,N_4309);
and U7211 (N_7211,N_4220,N_4813);
nor U7212 (N_7212,N_1927,N_2830);
and U7213 (N_7213,N_246,N_1872);
nand U7214 (N_7214,N_1687,N_1770);
nor U7215 (N_7215,N_2207,N_4337);
nor U7216 (N_7216,N_1882,N_2884);
nor U7217 (N_7217,N_1457,N_2375);
or U7218 (N_7218,N_2864,N_1635);
and U7219 (N_7219,N_579,N_4043);
xnor U7220 (N_7220,N_180,N_2626);
or U7221 (N_7221,N_521,N_3562);
and U7222 (N_7222,N_4877,N_1708);
nor U7223 (N_7223,N_708,N_2003);
and U7224 (N_7224,N_2361,N_3397);
or U7225 (N_7225,N_59,N_1551);
nand U7226 (N_7226,N_382,N_3699);
nand U7227 (N_7227,N_3837,N_1807);
nand U7228 (N_7228,N_4857,N_4473);
and U7229 (N_7229,N_4483,N_2714);
nor U7230 (N_7230,N_451,N_1778);
or U7231 (N_7231,N_3364,N_638);
nand U7232 (N_7232,N_3168,N_3286);
or U7233 (N_7233,N_1181,N_3883);
and U7234 (N_7234,N_2971,N_1954);
or U7235 (N_7235,N_1582,N_725);
nor U7236 (N_7236,N_3526,N_3011);
or U7237 (N_7237,N_1476,N_4352);
or U7238 (N_7238,N_4708,N_2440);
nor U7239 (N_7239,N_3278,N_3213);
nand U7240 (N_7240,N_4298,N_3521);
nor U7241 (N_7241,N_3305,N_1301);
xnor U7242 (N_7242,N_2199,N_3772);
and U7243 (N_7243,N_2315,N_3828);
and U7244 (N_7244,N_2173,N_2167);
nand U7245 (N_7245,N_1598,N_2857);
nand U7246 (N_7246,N_146,N_3271);
nand U7247 (N_7247,N_1433,N_3764);
xor U7248 (N_7248,N_1505,N_2629);
nand U7249 (N_7249,N_2974,N_1138);
or U7250 (N_7250,N_1001,N_1025);
nand U7251 (N_7251,N_2093,N_3543);
and U7252 (N_7252,N_4970,N_1096);
or U7253 (N_7253,N_4646,N_2688);
and U7254 (N_7254,N_203,N_3262);
nor U7255 (N_7255,N_2766,N_4359);
or U7256 (N_7256,N_1810,N_3692);
nor U7257 (N_7257,N_4629,N_4034);
nor U7258 (N_7258,N_1984,N_1592);
and U7259 (N_7259,N_4893,N_4303);
or U7260 (N_7260,N_3407,N_1678);
or U7261 (N_7261,N_4587,N_3420);
and U7262 (N_7262,N_284,N_45);
and U7263 (N_7263,N_1050,N_1385);
and U7264 (N_7264,N_3963,N_2081);
nor U7265 (N_7265,N_1167,N_2719);
nand U7266 (N_7266,N_2788,N_938);
or U7267 (N_7267,N_3167,N_1043);
nand U7268 (N_7268,N_4091,N_2506);
xnor U7269 (N_7269,N_976,N_65);
or U7270 (N_7270,N_1926,N_2922);
nor U7271 (N_7271,N_4067,N_2360);
nor U7272 (N_7272,N_3108,N_653);
nor U7273 (N_7273,N_1977,N_2447);
nand U7274 (N_7274,N_3795,N_4839);
or U7275 (N_7275,N_3191,N_2115);
nand U7276 (N_7276,N_3290,N_93);
or U7277 (N_7277,N_4290,N_1109);
nand U7278 (N_7278,N_2877,N_4956);
nand U7279 (N_7279,N_1381,N_3370);
nand U7280 (N_7280,N_770,N_364);
nand U7281 (N_7281,N_4350,N_168);
and U7282 (N_7282,N_4546,N_133);
and U7283 (N_7283,N_2675,N_969);
or U7284 (N_7284,N_3723,N_2057);
nor U7285 (N_7285,N_766,N_710);
nand U7286 (N_7286,N_4448,N_2379);
nand U7287 (N_7287,N_4183,N_3237);
nor U7288 (N_7288,N_2471,N_4016);
xor U7289 (N_7289,N_920,N_1356);
and U7290 (N_7290,N_1407,N_2610);
and U7291 (N_7291,N_3606,N_1160);
nor U7292 (N_7292,N_465,N_1863);
nor U7293 (N_7293,N_3678,N_739);
nand U7294 (N_7294,N_4185,N_510);
nor U7295 (N_7295,N_2894,N_51);
nand U7296 (N_7296,N_2716,N_1536);
or U7297 (N_7297,N_2356,N_1846);
and U7298 (N_7298,N_2421,N_4535);
nor U7299 (N_7299,N_2044,N_4142);
or U7300 (N_7300,N_1521,N_3655);
and U7301 (N_7301,N_647,N_541);
nor U7302 (N_7302,N_1497,N_1713);
or U7303 (N_7303,N_1305,N_987);
nand U7304 (N_7304,N_378,N_1472);
nor U7305 (N_7305,N_2302,N_4145);
nand U7306 (N_7306,N_62,N_2796);
or U7307 (N_7307,N_1877,N_625);
and U7308 (N_7308,N_1560,N_4844);
nand U7309 (N_7309,N_630,N_4847);
nor U7310 (N_7310,N_2359,N_1964);
nand U7311 (N_7311,N_368,N_1562);
or U7312 (N_7312,N_3858,N_975);
nand U7313 (N_7313,N_719,N_4997);
xor U7314 (N_7314,N_173,N_1361);
nor U7315 (N_7315,N_2062,N_4524);
xor U7316 (N_7316,N_1125,N_3395);
nor U7317 (N_7317,N_3120,N_4052);
and U7318 (N_7318,N_4678,N_2758);
nand U7319 (N_7319,N_3439,N_3999);
or U7320 (N_7320,N_1173,N_2775);
xor U7321 (N_7321,N_629,N_2619);
and U7322 (N_7322,N_136,N_3324);
nor U7323 (N_7323,N_2462,N_2019);
and U7324 (N_7324,N_2436,N_3767);
nor U7325 (N_7325,N_3373,N_3055);
or U7326 (N_7326,N_1890,N_4905);
and U7327 (N_7327,N_3675,N_2847);
nand U7328 (N_7328,N_3415,N_4528);
nor U7329 (N_7329,N_1484,N_2837);
or U7330 (N_7330,N_2727,N_2566);
nor U7331 (N_7331,N_1993,N_3864);
and U7332 (N_7332,N_3619,N_3921);
xor U7333 (N_7333,N_2445,N_957);
nor U7334 (N_7334,N_2913,N_1373);
or U7335 (N_7335,N_1956,N_2844);
and U7336 (N_7336,N_3712,N_1847);
xor U7337 (N_7337,N_1990,N_1242);
nand U7338 (N_7338,N_2749,N_3152);
or U7339 (N_7339,N_1140,N_1646);
or U7340 (N_7340,N_4389,N_1664);
and U7341 (N_7341,N_2319,N_3159);
nand U7342 (N_7342,N_4820,N_467);
nand U7343 (N_7343,N_1162,N_460);
xor U7344 (N_7344,N_2010,N_2655);
nand U7345 (N_7345,N_550,N_1171);
nor U7346 (N_7346,N_1987,N_123);
and U7347 (N_7347,N_4237,N_4088);
and U7348 (N_7348,N_2401,N_1554);
and U7349 (N_7349,N_1037,N_844);
nand U7350 (N_7350,N_4177,N_631);
or U7351 (N_7351,N_1944,N_798);
and U7352 (N_7352,N_1286,N_484);
nand U7353 (N_7353,N_974,N_2423);
or U7354 (N_7354,N_2896,N_3988);
nand U7355 (N_7355,N_4874,N_4693);
or U7356 (N_7356,N_453,N_1331);
and U7357 (N_7357,N_1123,N_985);
nor U7358 (N_7358,N_2686,N_4669);
nand U7359 (N_7359,N_2868,N_851);
xnor U7360 (N_7360,N_548,N_3062);
nor U7361 (N_7361,N_5,N_2252);
nor U7362 (N_7362,N_2602,N_4510);
or U7363 (N_7363,N_3954,N_697);
nor U7364 (N_7364,N_1129,N_3989);
nand U7365 (N_7365,N_2657,N_4482);
and U7366 (N_7366,N_1613,N_2408);
and U7367 (N_7367,N_695,N_4913);
nand U7368 (N_7368,N_479,N_1544);
nor U7369 (N_7369,N_121,N_3730);
or U7370 (N_7370,N_2034,N_4063);
nor U7371 (N_7371,N_293,N_3354);
xnor U7372 (N_7372,N_1892,N_4093);
nor U7373 (N_7373,N_1721,N_3658);
and U7374 (N_7374,N_2736,N_361);
nand U7375 (N_7375,N_3000,N_344);
or U7376 (N_7376,N_2527,N_2674);
or U7377 (N_7377,N_4377,N_3922);
nor U7378 (N_7378,N_3916,N_2002);
nand U7379 (N_7379,N_4625,N_3100);
and U7380 (N_7380,N_1710,N_1610);
nor U7381 (N_7381,N_1116,N_2724);
xnor U7382 (N_7382,N_1959,N_4894);
and U7383 (N_7383,N_3620,N_436);
and U7384 (N_7384,N_4172,N_1396);
nor U7385 (N_7385,N_4515,N_4638);
and U7386 (N_7386,N_4041,N_684);
and U7387 (N_7387,N_4512,N_1682);
nand U7388 (N_7388,N_2523,N_954);
or U7389 (N_7389,N_2855,N_2918);
or U7390 (N_7390,N_2080,N_2236);
nand U7391 (N_7391,N_4740,N_463);
nand U7392 (N_7392,N_700,N_1299);
nor U7393 (N_7393,N_1027,N_386);
nor U7394 (N_7394,N_4916,N_4593);
nand U7395 (N_7395,N_1362,N_3796);
and U7396 (N_7396,N_2693,N_1403);
or U7397 (N_7397,N_3003,N_3718);
nor U7398 (N_7398,N_1704,N_1960);
nand U7399 (N_7399,N_3717,N_4454);
nor U7400 (N_7400,N_3566,N_2834);
xnor U7401 (N_7401,N_4037,N_3970);
nand U7402 (N_7402,N_1815,N_499);
nor U7403 (N_7403,N_2200,N_3504);
nand U7404 (N_7404,N_4862,N_2299);
nor U7405 (N_7405,N_2797,N_4806);
nand U7406 (N_7406,N_2900,N_4939);
and U7407 (N_7407,N_2435,N_3668);
or U7408 (N_7408,N_1074,N_1724);
nor U7409 (N_7409,N_966,N_1395);
and U7410 (N_7410,N_4168,N_2183);
nand U7411 (N_7411,N_2533,N_4152);
and U7412 (N_7412,N_206,N_396);
and U7413 (N_7413,N_4924,N_4196);
or U7414 (N_7414,N_3974,N_4138);
and U7415 (N_7415,N_418,N_2089);
and U7416 (N_7416,N_563,N_1730);
and U7417 (N_7417,N_1436,N_2437);
xor U7418 (N_7418,N_3607,N_1606);
and U7419 (N_7419,N_373,N_2096);
nor U7420 (N_7420,N_2891,N_274);
nor U7421 (N_7421,N_4909,N_950);
nor U7422 (N_7422,N_3394,N_4148);
nor U7423 (N_7423,N_4707,N_3594);
nor U7424 (N_7424,N_4590,N_2879);
nor U7425 (N_7425,N_3649,N_2219);
nor U7426 (N_7426,N_4076,N_1413);
nand U7427 (N_7427,N_3756,N_790);
nand U7428 (N_7428,N_2310,N_2474);
and U7429 (N_7429,N_866,N_3716);
or U7430 (N_7430,N_2556,N_495);
and U7431 (N_7431,N_1609,N_4868);
or U7432 (N_7432,N_2725,N_1084);
or U7433 (N_7433,N_3196,N_3074);
nand U7434 (N_7434,N_760,N_3548);
or U7435 (N_7435,N_1818,N_4789);
xnor U7436 (N_7436,N_429,N_2728);
or U7437 (N_7437,N_1075,N_3075);
nand U7438 (N_7438,N_2231,N_1851);
nand U7439 (N_7439,N_1225,N_2433);
and U7440 (N_7440,N_3046,N_1755);
nor U7441 (N_7441,N_3541,N_419);
and U7442 (N_7442,N_3708,N_3791);
nor U7443 (N_7443,N_728,N_2709);
and U7444 (N_7444,N_4704,N_1888);
xnor U7445 (N_7445,N_2585,N_2250);
or U7446 (N_7446,N_1341,N_111);
and U7447 (N_7447,N_4618,N_899);
xnor U7448 (N_7448,N_271,N_1576);
or U7449 (N_7449,N_4306,N_1795);
and U7450 (N_7450,N_3162,N_339);
nand U7451 (N_7451,N_4879,N_3443);
nor U7452 (N_7452,N_4199,N_956);
or U7453 (N_7453,N_1470,N_3097);
and U7454 (N_7454,N_4289,N_4630);
nor U7455 (N_7455,N_2312,N_4670);
nor U7456 (N_7456,N_3051,N_2841);
nand U7457 (N_7457,N_999,N_2170);
nand U7458 (N_7458,N_1033,N_1813);
xnor U7459 (N_7459,N_2213,N_4739);
or U7460 (N_7460,N_4703,N_1326);
nand U7461 (N_7461,N_4870,N_2238);
and U7462 (N_7462,N_1257,N_3670);
or U7463 (N_7463,N_4342,N_202);
nor U7464 (N_7464,N_258,N_1573);
and U7465 (N_7465,N_4022,N_3279);
or U7466 (N_7466,N_3596,N_4942);
or U7467 (N_7467,N_752,N_3509);
and U7468 (N_7468,N_329,N_4464);
nand U7469 (N_7469,N_2111,N_4085);
xnor U7470 (N_7470,N_2694,N_3163);
nor U7471 (N_7471,N_3680,N_2848);
nor U7472 (N_7472,N_4672,N_147);
or U7473 (N_7473,N_1945,N_186);
or U7474 (N_7474,N_3273,N_3744);
or U7475 (N_7475,N_4080,N_207);
and U7476 (N_7476,N_2415,N_672);
or U7477 (N_7477,N_1486,N_3284);
nor U7478 (N_7478,N_285,N_1414);
and U7479 (N_7479,N_2599,N_283);
xnor U7480 (N_7480,N_3417,N_273);
or U7481 (N_7481,N_1370,N_2197);
nor U7482 (N_7482,N_2482,N_428);
nor U7483 (N_7483,N_4190,N_1196);
xor U7484 (N_7484,N_3189,N_3036);
nand U7485 (N_7485,N_2975,N_4978);
and U7486 (N_7486,N_4072,N_727);
nor U7487 (N_7487,N_3328,N_1588);
nand U7488 (N_7488,N_3408,N_3975);
or U7489 (N_7489,N_4174,N_2160);
and U7490 (N_7490,N_4159,N_4397);
nor U7491 (N_7491,N_4441,N_4269);
nand U7492 (N_7492,N_2294,N_1595);
nand U7493 (N_7493,N_1388,N_439);
and U7494 (N_7494,N_2773,N_4436);
nor U7495 (N_7495,N_1798,N_1619);
nand U7496 (N_7496,N_385,N_963);
nor U7497 (N_7497,N_3663,N_2744);
nor U7498 (N_7498,N_333,N_2041);
xnor U7499 (N_7499,N_3222,N_680);
and U7500 (N_7500,N_3803,N_4274);
nand U7501 (N_7501,N_1707,N_2260);
nand U7502 (N_7502,N_1966,N_2533);
xor U7503 (N_7503,N_365,N_3875);
and U7504 (N_7504,N_1949,N_335);
and U7505 (N_7505,N_1870,N_18);
nor U7506 (N_7506,N_2163,N_336);
nand U7507 (N_7507,N_2128,N_2559);
and U7508 (N_7508,N_2114,N_3166);
nand U7509 (N_7509,N_85,N_4465);
nand U7510 (N_7510,N_1903,N_402);
or U7511 (N_7511,N_1003,N_2003);
nand U7512 (N_7512,N_3945,N_1212);
nor U7513 (N_7513,N_644,N_4694);
and U7514 (N_7514,N_1493,N_2273);
nor U7515 (N_7515,N_4354,N_429);
nor U7516 (N_7516,N_4026,N_3540);
nand U7517 (N_7517,N_2006,N_868);
and U7518 (N_7518,N_3306,N_3639);
and U7519 (N_7519,N_1200,N_3522);
nand U7520 (N_7520,N_4472,N_3323);
nand U7521 (N_7521,N_436,N_3640);
nor U7522 (N_7522,N_143,N_1847);
nor U7523 (N_7523,N_2268,N_3136);
or U7524 (N_7524,N_929,N_916);
nor U7525 (N_7525,N_1750,N_2723);
and U7526 (N_7526,N_4145,N_1969);
and U7527 (N_7527,N_2753,N_4971);
xnor U7528 (N_7528,N_1552,N_4208);
xor U7529 (N_7529,N_1175,N_715);
nor U7530 (N_7530,N_1354,N_1234);
and U7531 (N_7531,N_3416,N_587);
nand U7532 (N_7532,N_3719,N_451);
xor U7533 (N_7533,N_4249,N_3836);
and U7534 (N_7534,N_3498,N_792);
nand U7535 (N_7535,N_1155,N_1957);
nor U7536 (N_7536,N_4664,N_4227);
or U7537 (N_7537,N_4147,N_1162);
or U7538 (N_7538,N_2514,N_2309);
or U7539 (N_7539,N_2290,N_814);
or U7540 (N_7540,N_4549,N_4339);
xnor U7541 (N_7541,N_3286,N_362);
and U7542 (N_7542,N_4477,N_3644);
xnor U7543 (N_7543,N_655,N_948);
or U7544 (N_7544,N_2983,N_914);
or U7545 (N_7545,N_4986,N_1930);
nor U7546 (N_7546,N_1929,N_857);
or U7547 (N_7547,N_3706,N_121);
nor U7548 (N_7548,N_1982,N_1033);
nand U7549 (N_7549,N_2640,N_531);
and U7550 (N_7550,N_1529,N_4029);
or U7551 (N_7551,N_4820,N_1574);
nand U7552 (N_7552,N_3941,N_4339);
or U7553 (N_7553,N_2066,N_906);
and U7554 (N_7554,N_655,N_2333);
nand U7555 (N_7555,N_2704,N_216);
nor U7556 (N_7556,N_3129,N_3808);
nand U7557 (N_7557,N_3691,N_716);
or U7558 (N_7558,N_1215,N_2061);
and U7559 (N_7559,N_2692,N_3652);
and U7560 (N_7560,N_1185,N_3443);
and U7561 (N_7561,N_4762,N_1983);
nand U7562 (N_7562,N_3376,N_3039);
xnor U7563 (N_7563,N_4878,N_4124);
and U7564 (N_7564,N_255,N_2737);
nand U7565 (N_7565,N_2802,N_3579);
and U7566 (N_7566,N_65,N_4883);
nand U7567 (N_7567,N_2997,N_1746);
nand U7568 (N_7568,N_1229,N_2343);
nand U7569 (N_7569,N_4884,N_3941);
nor U7570 (N_7570,N_4890,N_1762);
nor U7571 (N_7571,N_4350,N_1134);
and U7572 (N_7572,N_1533,N_4243);
xor U7573 (N_7573,N_1377,N_1906);
nand U7574 (N_7574,N_243,N_1498);
nand U7575 (N_7575,N_1665,N_1270);
nor U7576 (N_7576,N_3778,N_1909);
or U7577 (N_7577,N_1925,N_4015);
xnor U7578 (N_7578,N_4502,N_445);
or U7579 (N_7579,N_4807,N_3575);
and U7580 (N_7580,N_2868,N_2263);
and U7581 (N_7581,N_1,N_1409);
nor U7582 (N_7582,N_363,N_3542);
nand U7583 (N_7583,N_4622,N_103);
nand U7584 (N_7584,N_3164,N_2390);
and U7585 (N_7585,N_3469,N_3695);
nand U7586 (N_7586,N_2413,N_2004);
xnor U7587 (N_7587,N_4876,N_406);
or U7588 (N_7588,N_2555,N_4191);
nor U7589 (N_7589,N_3952,N_3461);
and U7590 (N_7590,N_666,N_956);
nor U7591 (N_7591,N_3646,N_1376);
and U7592 (N_7592,N_2956,N_2777);
nor U7593 (N_7593,N_4390,N_4726);
and U7594 (N_7594,N_263,N_4856);
nand U7595 (N_7595,N_658,N_1492);
or U7596 (N_7596,N_2641,N_4337);
and U7597 (N_7597,N_2899,N_673);
nand U7598 (N_7598,N_2903,N_358);
nor U7599 (N_7599,N_2886,N_983);
xor U7600 (N_7600,N_4663,N_2804);
nor U7601 (N_7601,N_2251,N_469);
or U7602 (N_7602,N_1820,N_260);
nand U7603 (N_7603,N_825,N_2997);
nor U7604 (N_7604,N_1811,N_4717);
and U7605 (N_7605,N_4008,N_4512);
nor U7606 (N_7606,N_4121,N_3068);
nand U7607 (N_7607,N_2573,N_569);
xor U7608 (N_7608,N_4233,N_3408);
or U7609 (N_7609,N_2145,N_658);
nor U7610 (N_7610,N_3078,N_158);
and U7611 (N_7611,N_4219,N_2258);
nor U7612 (N_7612,N_954,N_120);
or U7613 (N_7613,N_2001,N_1164);
or U7614 (N_7614,N_4695,N_1900);
xor U7615 (N_7615,N_4051,N_905);
or U7616 (N_7616,N_4862,N_308);
or U7617 (N_7617,N_2078,N_4396);
nand U7618 (N_7618,N_2073,N_3808);
nor U7619 (N_7619,N_1997,N_1263);
or U7620 (N_7620,N_3847,N_1829);
or U7621 (N_7621,N_343,N_2287);
or U7622 (N_7622,N_4951,N_2949);
and U7623 (N_7623,N_2884,N_1960);
nand U7624 (N_7624,N_2457,N_4098);
nand U7625 (N_7625,N_2444,N_1776);
nand U7626 (N_7626,N_1284,N_2099);
or U7627 (N_7627,N_1295,N_1014);
xor U7628 (N_7628,N_2154,N_4655);
xor U7629 (N_7629,N_1206,N_1753);
nand U7630 (N_7630,N_1099,N_1010);
nand U7631 (N_7631,N_3480,N_4663);
or U7632 (N_7632,N_2782,N_319);
xnor U7633 (N_7633,N_4438,N_3642);
and U7634 (N_7634,N_3360,N_3472);
nand U7635 (N_7635,N_3844,N_3522);
nor U7636 (N_7636,N_2517,N_3286);
xor U7637 (N_7637,N_595,N_4244);
nand U7638 (N_7638,N_1405,N_1469);
and U7639 (N_7639,N_838,N_3798);
and U7640 (N_7640,N_4843,N_1282);
or U7641 (N_7641,N_4315,N_1618);
nor U7642 (N_7642,N_1007,N_4684);
and U7643 (N_7643,N_601,N_2090);
nor U7644 (N_7644,N_3301,N_707);
or U7645 (N_7645,N_3297,N_4525);
nor U7646 (N_7646,N_4469,N_910);
xnor U7647 (N_7647,N_2141,N_1904);
or U7648 (N_7648,N_991,N_2941);
nor U7649 (N_7649,N_4161,N_4393);
nand U7650 (N_7650,N_2899,N_3147);
or U7651 (N_7651,N_4789,N_1617);
and U7652 (N_7652,N_141,N_4311);
nand U7653 (N_7653,N_693,N_3043);
and U7654 (N_7654,N_1711,N_3346);
nand U7655 (N_7655,N_3885,N_1828);
and U7656 (N_7656,N_3964,N_4800);
nand U7657 (N_7657,N_3613,N_4948);
nor U7658 (N_7658,N_803,N_4265);
nand U7659 (N_7659,N_2588,N_815);
nand U7660 (N_7660,N_4454,N_2715);
nand U7661 (N_7661,N_4437,N_3097);
nor U7662 (N_7662,N_3239,N_545);
and U7663 (N_7663,N_1525,N_2246);
nor U7664 (N_7664,N_3652,N_827);
nor U7665 (N_7665,N_277,N_1038);
or U7666 (N_7666,N_1454,N_446);
nor U7667 (N_7667,N_1684,N_2719);
xor U7668 (N_7668,N_83,N_4983);
nor U7669 (N_7669,N_2665,N_4179);
xnor U7670 (N_7670,N_4409,N_3841);
nand U7671 (N_7671,N_1757,N_4973);
and U7672 (N_7672,N_2389,N_2645);
and U7673 (N_7673,N_4656,N_1668);
nand U7674 (N_7674,N_490,N_2896);
and U7675 (N_7675,N_748,N_2257);
nor U7676 (N_7676,N_4776,N_4418);
and U7677 (N_7677,N_572,N_509);
and U7678 (N_7678,N_2065,N_3009);
and U7679 (N_7679,N_4605,N_925);
nand U7680 (N_7680,N_1696,N_3745);
nor U7681 (N_7681,N_1378,N_3093);
nor U7682 (N_7682,N_1572,N_1427);
and U7683 (N_7683,N_2344,N_3656);
xnor U7684 (N_7684,N_3625,N_2317);
and U7685 (N_7685,N_1293,N_2358);
xor U7686 (N_7686,N_227,N_2845);
nand U7687 (N_7687,N_3854,N_212);
nand U7688 (N_7688,N_1139,N_3402);
nor U7689 (N_7689,N_11,N_3103);
and U7690 (N_7690,N_4917,N_2786);
and U7691 (N_7691,N_3,N_1314);
nor U7692 (N_7692,N_3521,N_3985);
xnor U7693 (N_7693,N_2326,N_576);
xor U7694 (N_7694,N_4966,N_337);
nand U7695 (N_7695,N_4212,N_889);
or U7696 (N_7696,N_3753,N_3692);
and U7697 (N_7697,N_4716,N_1466);
and U7698 (N_7698,N_1493,N_4144);
and U7699 (N_7699,N_1285,N_4313);
nor U7700 (N_7700,N_1671,N_3326);
or U7701 (N_7701,N_3702,N_3920);
xnor U7702 (N_7702,N_382,N_2257);
nand U7703 (N_7703,N_4339,N_4866);
nand U7704 (N_7704,N_2347,N_4921);
and U7705 (N_7705,N_2053,N_4397);
and U7706 (N_7706,N_4368,N_3439);
nor U7707 (N_7707,N_3977,N_3644);
or U7708 (N_7708,N_3400,N_3977);
or U7709 (N_7709,N_2016,N_1619);
and U7710 (N_7710,N_2461,N_3478);
and U7711 (N_7711,N_1472,N_140);
and U7712 (N_7712,N_915,N_1806);
or U7713 (N_7713,N_1643,N_2561);
or U7714 (N_7714,N_4993,N_272);
or U7715 (N_7715,N_2396,N_3359);
and U7716 (N_7716,N_99,N_4779);
nand U7717 (N_7717,N_2605,N_4721);
and U7718 (N_7718,N_258,N_2304);
or U7719 (N_7719,N_4299,N_3160);
and U7720 (N_7720,N_683,N_979);
nor U7721 (N_7721,N_951,N_1705);
and U7722 (N_7722,N_2486,N_2456);
nor U7723 (N_7723,N_3922,N_1530);
xor U7724 (N_7724,N_4939,N_3411);
nor U7725 (N_7725,N_2110,N_3787);
and U7726 (N_7726,N_2905,N_281);
or U7727 (N_7727,N_2234,N_4772);
nor U7728 (N_7728,N_2273,N_3661);
and U7729 (N_7729,N_3668,N_1012);
nand U7730 (N_7730,N_3670,N_477);
nor U7731 (N_7731,N_1398,N_3178);
nor U7732 (N_7732,N_4458,N_1534);
nand U7733 (N_7733,N_4482,N_509);
and U7734 (N_7734,N_4631,N_2558);
and U7735 (N_7735,N_2584,N_3293);
xor U7736 (N_7736,N_4289,N_2586);
nand U7737 (N_7737,N_3404,N_2395);
nand U7738 (N_7738,N_4192,N_1615);
xnor U7739 (N_7739,N_683,N_3888);
nor U7740 (N_7740,N_1493,N_694);
or U7741 (N_7741,N_4957,N_926);
nand U7742 (N_7742,N_1738,N_980);
xor U7743 (N_7743,N_2854,N_445);
nand U7744 (N_7744,N_2599,N_39);
xor U7745 (N_7745,N_1562,N_2879);
xor U7746 (N_7746,N_3953,N_342);
nand U7747 (N_7747,N_2367,N_2509);
nor U7748 (N_7748,N_1921,N_827);
and U7749 (N_7749,N_3154,N_4452);
xnor U7750 (N_7750,N_4362,N_961);
and U7751 (N_7751,N_2564,N_2744);
and U7752 (N_7752,N_413,N_62);
and U7753 (N_7753,N_4470,N_2225);
or U7754 (N_7754,N_4244,N_860);
or U7755 (N_7755,N_3996,N_1604);
xnor U7756 (N_7756,N_4545,N_2373);
nand U7757 (N_7757,N_4433,N_2518);
and U7758 (N_7758,N_4189,N_2480);
nor U7759 (N_7759,N_1346,N_1328);
and U7760 (N_7760,N_4951,N_2469);
and U7761 (N_7761,N_3447,N_1637);
nor U7762 (N_7762,N_1928,N_3129);
nor U7763 (N_7763,N_529,N_4587);
xnor U7764 (N_7764,N_1892,N_1385);
nor U7765 (N_7765,N_2954,N_1782);
nand U7766 (N_7766,N_3660,N_4890);
xor U7767 (N_7767,N_2159,N_2032);
nor U7768 (N_7768,N_4261,N_696);
xnor U7769 (N_7769,N_2245,N_3229);
nand U7770 (N_7770,N_4346,N_752);
nor U7771 (N_7771,N_4250,N_2080);
nand U7772 (N_7772,N_2209,N_856);
nor U7773 (N_7773,N_1677,N_406);
or U7774 (N_7774,N_388,N_3939);
and U7775 (N_7775,N_103,N_1750);
nand U7776 (N_7776,N_3168,N_356);
nor U7777 (N_7777,N_1797,N_2872);
or U7778 (N_7778,N_97,N_3853);
nand U7779 (N_7779,N_4471,N_4358);
xnor U7780 (N_7780,N_1993,N_2374);
and U7781 (N_7781,N_4343,N_4158);
nand U7782 (N_7782,N_2300,N_4246);
or U7783 (N_7783,N_1779,N_76);
or U7784 (N_7784,N_1683,N_4944);
or U7785 (N_7785,N_290,N_3498);
nor U7786 (N_7786,N_1275,N_4133);
xor U7787 (N_7787,N_3443,N_4435);
nor U7788 (N_7788,N_3093,N_2577);
or U7789 (N_7789,N_4668,N_925);
and U7790 (N_7790,N_3282,N_2816);
or U7791 (N_7791,N_2336,N_1781);
or U7792 (N_7792,N_930,N_4870);
or U7793 (N_7793,N_2114,N_1446);
nand U7794 (N_7794,N_405,N_1927);
or U7795 (N_7795,N_2687,N_4805);
and U7796 (N_7796,N_1722,N_4813);
and U7797 (N_7797,N_4628,N_1261);
nand U7798 (N_7798,N_2784,N_1961);
nor U7799 (N_7799,N_2486,N_691);
nand U7800 (N_7800,N_1114,N_2137);
and U7801 (N_7801,N_3506,N_3624);
and U7802 (N_7802,N_3985,N_4667);
or U7803 (N_7803,N_4588,N_1255);
nor U7804 (N_7804,N_373,N_775);
and U7805 (N_7805,N_711,N_105);
or U7806 (N_7806,N_4571,N_2061);
and U7807 (N_7807,N_1248,N_1276);
or U7808 (N_7808,N_2355,N_1532);
or U7809 (N_7809,N_1032,N_4574);
nand U7810 (N_7810,N_1890,N_3418);
nor U7811 (N_7811,N_1069,N_2752);
nor U7812 (N_7812,N_1458,N_4928);
or U7813 (N_7813,N_2360,N_2982);
nand U7814 (N_7814,N_296,N_4419);
nor U7815 (N_7815,N_1658,N_529);
nand U7816 (N_7816,N_2318,N_4366);
nor U7817 (N_7817,N_743,N_1886);
and U7818 (N_7818,N_2421,N_1262);
nand U7819 (N_7819,N_2459,N_863);
nand U7820 (N_7820,N_2341,N_3546);
and U7821 (N_7821,N_4344,N_3337);
and U7822 (N_7822,N_3048,N_459);
and U7823 (N_7823,N_1211,N_4394);
nor U7824 (N_7824,N_4082,N_2402);
and U7825 (N_7825,N_1031,N_2472);
and U7826 (N_7826,N_4814,N_1747);
xnor U7827 (N_7827,N_2770,N_4871);
or U7828 (N_7828,N_1738,N_647);
and U7829 (N_7829,N_4041,N_4202);
xor U7830 (N_7830,N_272,N_2432);
nand U7831 (N_7831,N_1195,N_1486);
and U7832 (N_7832,N_490,N_1863);
or U7833 (N_7833,N_3361,N_4315);
or U7834 (N_7834,N_1813,N_4075);
and U7835 (N_7835,N_78,N_2617);
xnor U7836 (N_7836,N_1481,N_3635);
or U7837 (N_7837,N_1970,N_1034);
and U7838 (N_7838,N_204,N_2783);
nand U7839 (N_7839,N_3729,N_3982);
nand U7840 (N_7840,N_4388,N_3446);
or U7841 (N_7841,N_3312,N_592);
or U7842 (N_7842,N_3446,N_3107);
nand U7843 (N_7843,N_3544,N_1911);
nand U7844 (N_7844,N_1431,N_345);
and U7845 (N_7845,N_4759,N_3039);
nand U7846 (N_7846,N_1453,N_3516);
nor U7847 (N_7847,N_3288,N_2190);
nor U7848 (N_7848,N_3355,N_3379);
nand U7849 (N_7849,N_1239,N_831);
and U7850 (N_7850,N_1891,N_4392);
nor U7851 (N_7851,N_4599,N_1157);
and U7852 (N_7852,N_305,N_2607);
or U7853 (N_7853,N_1620,N_1492);
or U7854 (N_7854,N_1285,N_3598);
and U7855 (N_7855,N_1901,N_3793);
nor U7856 (N_7856,N_4134,N_1996);
xnor U7857 (N_7857,N_233,N_27);
and U7858 (N_7858,N_1708,N_4190);
nand U7859 (N_7859,N_4365,N_3690);
or U7860 (N_7860,N_3615,N_4714);
and U7861 (N_7861,N_4372,N_2343);
nor U7862 (N_7862,N_4511,N_1889);
or U7863 (N_7863,N_3607,N_2295);
nor U7864 (N_7864,N_4804,N_3027);
nor U7865 (N_7865,N_1599,N_4332);
and U7866 (N_7866,N_502,N_172);
xor U7867 (N_7867,N_4634,N_2981);
nand U7868 (N_7868,N_2863,N_3925);
or U7869 (N_7869,N_4876,N_2791);
or U7870 (N_7870,N_4472,N_3633);
and U7871 (N_7871,N_4236,N_2487);
or U7872 (N_7872,N_4099,N_1719);
xor U7873 (N_7873,N_2233,N_1488);
nand U7874 (N_7874,N_2676,N_458);
nand U7875 (N_7875,N_4014,N_4108);
nand U7876 (N_7876,N_138,N_2596);
or U7877 (N_7877,N_245,N_2500);
and U7878 (N_7878,N_917,N_4829);
or U7879 (N_7879,N_1811,N_1552);
nand U7880 (N_7880,N_3193,N_2376);
nand U7881 (N_7881,N_4116,N_2240);
or U7882 (N_7882,N_4888,N_1140);
or U7883 (N_7883,N_4276,N_3671);
nor U7884 (N_7884,N_1412,N_2572);
and U7885 (N_7885,N_2947,N_4902);
nor U7886 (N_7886,N_3692,N_2283);
nand U7887 (N_7887,N_1050,N_1875);
nand U7888 (N_7888,N_3716,N_2979);
nor U7889 (N_7889,N_55,N_1044);
and U7890 (N_7890,N_2102,N_4909);
or U7891 (N_7891,N_3128,N_2529);
nand U7892 (N_7892,N_4299,N_2650);
nor U7893 (N_7893,N_379,N_4564);
or U7894 (N_7894,N_1364,N_3913);
nor U7895 (N_7895,N_4185,N_4803);
nor U7896 (N_7896,N_1002,N_4318);
nand U7897 (N_7897,N_4316,N_2397);
and U7898 (N_7898,N_829,N_4022);
xnor U7899 (N_7899,N_3107,N_3720);
xnor U7900 (N_7900,N_4475,N_406);
and U7901 (N_7901,N_1517,N_2708);
nand U7902 (N_7902,N_1616,N_682);
or U7903 (N_7903,N_2280,N_523);
xnor U7904 (N_7904,N_395,N_4903);
nand U7905 (N_7905,N_3288,N_1935);
or U7906 (N_7906,N_2584,N_3678);
nor U7907 (N_7907,N_2690,N_3518);
nand U7908 (N_7908,N_4971,N_3641);
and U7909 (N_7909,N_1051,N_4440);
or U7910 (N_7910,N_2541,N_2074);
nor U7911 (N_7911,N_1854,N_4304);
nor U7912 (N_7912,N_4155,N_954);
or U7913 (N_7913,N_1285,N_3982);
nand U7914 (N_7914,N_4545,N_1331);
nand U7915 (N_7915,N_1888,N_3088);
and U7916 (N_7916,N_1698,N_1721);
xor U7917 (N_7917,N_2798,N_1453);
nand U7918 (N_7918,N_948,N_1861);
nand U7919 (N_7919,N_1604,N_2793);
nand U7920 (N_7920,N_4099,N_2976);
nand U7921 (N_7921,N_899,N_2054);
nor U7922 (N_7922,N_2959,N_4930);
and U7923 (N_7923,N_980,N_2882);
or U7924 (N_7924,N_1143,N_4068);
nand U7925 (N_7925,N_85,N_2520);
nand U7926 (N_7926,N_3248,N_1721);
nand U7927 (N_7927,N_1669,N_3915);
or U7928 (N_7928,N_4918,N_1866);
nor U7929 (N_7929,N_2448,N_3537);
or U7930 (N_7930,N_3322,N_1258);
or U7931 (N_7931,N_156,N_4364);
or U7932 (N_7932,N_2549,N_2925);
nand U7933 (N_7933,N_2466,N_2432);
nor U7934 (N_7934,N_3593,N_2651);
nor U7935 (N_7935,N_3299,N_485);
nand U7936 (N_7936,N_1867,N_2408);
nor U7937 (N_7937,N_4568,N_3078);
or U7938 (N_7938,N_1888,N_442);
nor U7939 (N_7939,N_547,N_3627);
nand U7940 (N_7940,N_4915,N_4801);
nand U7941 (N_7941,N_446,N_403);
or U7942 (N_7942,N_716,N_2321);
xnor U7943 (N_7943,N_4750,N_4720);
nor U7944 (N_7944,N_791,N_729);
or U7945 (N_7945,N_1812,N_3480);
nand U7946 (N_7946,N_974,N_989);
or U7947 (N_7947,N_715,N_1109);
nand U7948 (N_7948,N_4262,N_861);
xnor U7949 (N_7949,N_4529,N_1638);
nand U7950 (N_7950,N_4872,N_857);
and U7951 (N_7951,N_3966,N_478);
nand U7952 (N_7952,N_1049,N_4665);
nor U7953 (N_7953,N_1933,N_3454);
or U7954 (N_7954,N_1562,N_2652);
nor U7955 (N_7955,N_1896,N_1427);
nand U7956 (N_7956,N_2516,N_328);
nand U7957 (N_7957,N_347,N_735);
nor U7958 (N_7958,N_2723,N_2666);
and U7959 (N_7959,N_922,N_517);
nor U7960 (N_7960,N_1965,N_1792);
nand U7961 (N_7961,N_4585,N_1756);
and U7962 (N_7962,N_2369,N_3556);
nand U7963 (N_7963,N_400,N_1981);
nand U7964 (N_7964,N_364,N_1981);
nor U7965 (N_7965,N_4066,N_985);
and U7966 (N_7966,N_1106,N_1509);
xor U7967 (N_7967,N_1802,N_2506);
or U7968 (N_7968,N_2149,N_2103);
and U7969 (N_7969,N_3442,N_4442);
and U7970 (N_7970,N_639,N_4032);
and U7971 (N_7971,N_2798,N_2199);
nor U7972 (N_7972,N_1708,N_2530);
xor U7973 (N_7973,N_4103,N_1705);
or U7974 (N_7974,N_1601,N_2775);
or U7975 (N_7975,N_4483,N_655);
xor U7976 (N_7976,N_2140,N_3534);
or U7977 (N_7977,N_4467,N_1457);
or U7978 (N_7978,N_2668,N_1917);
or U7979 (N_7979,N_465,N_922);
nand U7980 (N_7980,N_2969,N_365);
xor U7981 (N_7981,N_3590,N_1907);
nor U7982 (N_7982,N_3073,N_4966);
nor U7983 (N_7983,N_3053,N_246);
or U7984 (N_7984,N_2270,N_3046);
and U7985 (N_7985,N_3384,N_4099);
and U7986 (N_7986,N_4200,N_4817);
and U7987 (N_7987,N_2565,N_1355);
or U7988 (N_7988,N_2629,N_3241);
nor U7989 (N_7989,N_2456,N_4106);
nand U7990 (N_7990,N_3065,N_1126);
or U7991 (N_7991,N_1236,N_3915);
and U7992 (N_7992,N_2153,N_4312);
or U7993 (N_7993,N_4012,N_341);
nand U7994 (N_7994,N_2218,N_1870);
or U7995 (N_7995,N_1899,N_2032);
nor U7996 (N_7996,N_4199,N_3317);
or U7997 (N_7997,N_599,N_4235);
xor U7998 (N_7998,N_611,N_2084);
and U7999 (N_7999,N_4224,N_141);
or U8000 (N_8000,N_3641,N_2997);
nor U8001 (N_8001,N_1357,N_1232);
nor U8002 (N_8002,N_913,N_3446);
nor U8003 (N_8003,N_948,N_2357);
nor U8004 (N_8004,N_1108,N_4349);
xor U8005 (N_8005,N_2341,N_3292);
xor U8006 (N_8006,N_1433,N_2611);
nor U8007 (N_8007,N_2796,N_4840);
and U8008 (N_8008,N_2511,N_255);
nand U8009 (N_8009,N_14,N_1020);
and U8010 (N_8010,N_2381,N_4570);
or U8011 (N_8011,N_2636,N_1926);
or U8012 (N_8012,N_3575,N_3783);
and U8013 (N_8013,N_4477,N_3135);
or U8014 (N_8014,N_985,N_1838);
nand U8015 (N_8015,N_2458,N_904);
or U8016 (N_8016,N_1293,N_3687);
and U8017 (N_8017,N_441,N_4311);
or U8018 (N_8018,N_715,N_4686);
nor U8019 (N_8019,N_1183,N_274);
xor U8020 (N_8020,N_2098,N_975);
nor U8021 (N_8021,N_3690,N_4761);
nor U8022 (N_8022,N_2068,N_1318);
and U8023 (N_8023,N_1332,N_3036);
nor U8024 (N_8024,N_807,N_1091);
nand U8025 (N_8025,N_3369,N_1087);
or U8026 (N_8026,N_4249,N_3139);
or U8027 (N_8027,N_4211,N_3136);
and U8028 (N_8028,N_4482,N_2433);
and U8029 (N_8029,N_798,N_2119);
and U8030 (N_8030,N_260,N_230);
nand U8031 (N_8031,N_1064,N_3137);
and U8032 (N_8032,N_3354,N_990);
xor U8033 (N_8033,N_4656,N_3428);
and U8034 (N_8034,N_1944,N_2239);
xnor U8035 (N_8035,N_4904,N_717);
nor U8036 (N_8036,N_3248,N_4003);
or U8037 (N_8037,N_2887,N_3081);
nand U8038 (N_8038,N_2909,N_3665);
and U8039 (N_8039,N_3505,N_4803);
xor U8040 (N_8040,N_4051,N_4850);
and U8041 (N_8041,N_3342,N_164);
nor U8042 (N_8042,N_2995,N_3337);
or U8043 (N_8043,N_4255,N_202);
xor U8044 (N_8044,N_1016,N_75);
nor U8045 (N_8045,N_942,N_4879);
and U8046 (N_8046,N_3196,N_4213);
nor U8047 (N_8047,N_4564,N_33);
nor U8048 (N_8048,N_4863,N_143);
and U8049 (N_8049,N_1312,N_1059);
or U8050 (N_8050,N_4434,N_706);
or U8051 (N_8051,N_3026,N_1480);
nand U8052 (N_8052,N_4386,N_1980);
and U8053 (N_8053,N_1815,N_346);
or U8054 (N_8054,N_1342,N_3022);
and U8055 (N_8055,N_647,N_4703);
nand U8056 (N_8056,N_4085,N_4995);
nand U8057 (N_8057,N_1082,N_3636);
nor U8058 (N_8058,N_4198,N_2753);
xnor U8059 (N_8059,N_1956,N_4169);
nor U8060 (N_8060,N_4142,N_3638);
or U8061 (N_8061,N_3478,N_978);
nor U8062 (N_8062,N_2826,N_177);
or U8063 (N_8063,N_4521,N_522);
nor U8064 (N_8064,N_3885,N_2131);
nand U8065 (N_8065,N_3099,N_11);
or U8066 (N_8066,N_975,N_4868);
nor U8067 (N_8067,N_2685,N_1105);
nand U8068 (N_8068,N_2742,N_1204);
nand U8069 (N_8069,N_3344,N_4668);
nor U8070 (N_8070,N_1066,N_2418);
xor U8071 (N_8071,N_1209,N_4112);
nor U8072 (N_8072,N_1454,N_3275);
nor U8073 (N_8073,N_2665,N_4823);
nor U8074 (N_8074,N_4879,N_1758);
nand U8075 (N_8075,N_4880,N_3522);
or U8076 (N_8076,N_2451,N_1732);
or U8077 (N_8077,N_237,N_4477);
nand U8078 (N_8078,N_4251,N_3145);
nand U8079 (N_8079,N_173,N_3687);
or U8080 (N_8080,N_418,N_1033);
xnor U8081 (N_8081,N_689,N_2600);
and U8082 (N_8082,N_684,N_2663);
and U8083 (N_8083,N_4126,N_1591);
nor U8084 (N_8084,N_4341,N_859);
or U8085 (N_8085,N_2726,N_1656);
or U8086 (N_8086,N_2977,N_2353);
nand U8087 (N_8087,N_1732,N_3898);
or U8088 (N_8088,N_428,N_3290);
or U8089 (N_8089,N_3000,N_4838);
xnor U8090 (N_8090,N_997,N_4669);
or U8091 (N_8091,N_4995,N_1107);
nor U8092 (N_8092,N_1332,N_1068);
or U8093 (N_8093,N_2145,N_1909);
or U8094 (N_8094,N_4231,N_3433);
nand U8095 (N_8095,N_1729,N_3695);
or U8096 (N_8096,N_1434,N_3148);
or U8097 (N_8097,N_3730,N_1310);
nand U8098 (N_8098,N_848,N_3031);
and U8099 (N_8099,N_4893,N_2446);
xor U8100 (N_8100,N_972,N_4461);
nand U8101 (N_8101,N_413,N_3597);
nor U8102 (N_8102,N_4238,N_4104);
nand U8103 (N_8103,N_41,N_3095);
nand U8104 (N_8104,N_1694,N_1154);
and U8105 (N_8105,N_4473,N_4366);
nand U8106 (N_8106,N_4296,N_1092);
nand U8107 (N_8107,N_1231,N_4738);
or U8108 (N_8108,N_1880,N_298);
and U8109 (N_8109,N_378,N_4984);
or U8110 (N_8110,N_3728,N_124);
and U8111 (N_8111,N_4829,N_1658);
or U8112 (N_8112,N_835,N_1027);
nand U8113 (N_8113,N_612,N_2458);
nand U8114 (N_8114,N_2996,N_1009);
or U8115 (N_8115,N_620,N_173);
nor U8116 (N_8116,N_3725,N_4561);
nor U8117 (N_8117,N_393,N_2734);
nor U8118 (N_8118,N_4052,N_1223);
nor U8119 (N_8119,N_3673,N_4456);
or U8120 (N_8120,N_2843,N_958);
nand U8121 (N_8121,N_1829,N_1429);
and U8122 (N_8122,N_3494,N_4887);
or U8123 (N_8123,N_524,N_2037);
nand U8124 (N_8124,N_3144,N_1204);
xor U8125 (N_8125,N_3494,N_3859);
nand U8126 (N_8126,N_2094,N_564);
nand U8127 (N_8127,N_539,N_2206);
or U8128 (N_8128,N_2334,N_748);
and U8129 (N_8129,N_984,N_430);
nor U8130 (N_8130,N_980,N_4669);
nor U8131 (N_8131,N_3011,N_1630);
nor U8132 (N_8132,N_2115,N_4841);
nor U8133 (N_8133,N_4141,N_1415);
or U8134 (N_8134,N_3857,N_2343);
xor U8135 (N_8135,N_3498,N_4515);
and U8136 (N_8136,N_1702,N_1418);
nand U8137 (N_8137,N_353,N_3748);
and U8138 (N_8138,N_2499,N_3728);
nor U8139 (N_8139,N_3749,N_4787);
nand U8140 (N_8140,N_4697,N_4402);
and U8141 (N_8141,N_709,N_1955);
or U8142 (N_8142,N_3729,N_1322);
xor U8143 (N_8143,N_1984,N_1362);
nor U8144 (N_8144,N_2105,N_2650);
nand U8145 (N_8145,N_4237,N_653);
or U8146 (N_8146,N_3086,N_4736);
or U8147 (N_8147,N_367,N_2697);
nand U8148 (N_8148,N_3414,N_2814);
nor U8149 (N_8149,N_3358,N_3478);
xor U8150 (N_8150,N_3702,N_3329);
nor U8151 (N_8151,N_1220,N_3477);
or U8152 (N_8152,N_4466,N_4879);
nor U8153 (N_8153,N_4436,N_1260);
and U8154 (N_8154,N_767,N_1444);
nor U8155 (N_8155,N_478,N_2125);
nand U8156 (N_8156,N_4428,N_2834);
and U8157 (N_8157,N_3799,N_1774);
and U8158 (N_8158,N_2293,N_4464);
or U8159 (N_8159,N_2540,N_4791);
and U8160 (N_8160,N_737,N_4678);
nand U8161 (N_8161,N_4419,N_4999);
nor U8162 (N_8162,N_2494,N_4965);
or U8163 (N_8163,N_3089,N_512);
nand U8164 (N_8164,N_2241,N_1815);
and U8165 (N_8165,N_4904,N_55);
nand U8166 (N_8166,N_1751,N_4904);
nor U8167 (N_8167,N_2390,N_997);
nand U8168 (N_8168,N_2872,N_2167);
xor U8169 (N_8169,N_3743,N_3940);
and U8170 (N_8170,N_4228,N_3961);
nor U8171 (N_8171,N_3904,N_846);
nor U8172 (N_8172,N_3818,N_2945);
nand U8173 (N_8173,N_4015,N_2334);
and U8174 (N_8174,N_506,N_2719);
xnor U8175 (N_8175,N_3366,N_679);
or U8176 (N_8176,N_2561,N_4475);
and U8177 (N_8177,N_4492,N_4656);
nand U8178 (N_8178,N_3240,N_1221);
and U8179 (N_8179,N_271,N_1532);
nand U8180 (N_8180,N_1398,N_2342);
or U8181 (N_8181,N_4746,N_228);
nor U8182 (N_8182,N_2043,N_1484);
nor U8183 (N_8183,N_3545,N_4293);
or U8184 (N_8184,N_2502,N_2011);
or U8185 (N_8185,N_1405,N_3710);
nand U8186 (N_8186,N_1641,N_580);
or U8187 (N_8187,N_2836,N_157);
nand U8188 (N_8188,N_3247,N_3219);
and U8189 (N_8189,N_1686,N_1249);
nor U8190 (N_8190,N_200,N_2875);
nand U8191 (N_8191,N_4639,N_417);
xnor U8192 (N_8192,N_4780,N_4511);
nor U8193 (N_8193,N_4537,N_2591);
nand U8194 (N_8194,N_2173,N_3045);
nand U8195 (N_8195,N_2718,N_1482);
nor U8196 (N_8196,N_927,N_1784);
or U8197 (N_8197,N_1691,N_4212);
and U8198 (N_8198,N_1022,N_867);
or U8199 (N_8199,N_1447,N_4980);
nand U8200 (N_8200,N_4979,N_2357);
nor U8201 (N_8201,N_4876,N_1881);
nor U8202 (N_8202,N_2730,N_4976);
or U8203 (N_8203,N_2600,N_3449);
nand U8204 (N_8204,N_2925,N_1099);
nor U8205 (N_8205,N_2841,N_1167);
or U8206 (N_8206,N_2616,N_4732);
and U8207 (N_8207,N_4481,N_1892);
nand U8208 (N_8208,N_495,N_1565);
nand U8209 (N_8209,N_1452,N_651);
xnor U8210 (N_8210,N_1587,N_4273);
xor U8211 (N_8211,N_819,N_3874);
nor U8212 (N_8212,N_1597,N_2230);
and U8213 (N_8213,N_3599,N_4136);
and U8214 (N_8214,N_2089,N_4286);
nand U8215 (N_8215,N_3601,N_542);
and U8216 (N_8216,N_3204,N_4396);
nand U8217 (N_8217,N_3130,N_4660);
nor U8218 (N_8218,N_1883,N_3708);
nor U8219 (N_8219,N_2597,N_3151);
nand U8220 (N_8220,N_3347,N_2980);
nor U8221 (N_8221,N_3744,N_3007);
nor U8222 (N_8222,N_2140,N_3406);
nor U8223 (N_8223,N_3385,N_3051);
and U8224 (N_8224,N_4405,N_2311);
nor U8225 (N_8225,N_1595,N_1551);
or U8226 (N_8226,N_25,N_175);
and U8227 (N_8227,N_3931,N_3851);
nand U8228 (N_8228,N_577,N_3429);
and U8229 (N_8229,N_993,N_4772);
and U8230 (N_8230,N_247,N_4955);
and U8231 (N_8231,N_3435,N_4180);
xnor U8232 (N_8232,N_3571,N_453);
nand U8233 (N_8233,N_823,N_3229);
nand U8234 (N_8234,N_3219,N_4440);
xnor U8235 (N_8235,N_3913,N_401);
or U8236 (N_8236,N_2622,N_2791);
nor U8237 (N_8237,N_189,N_2121);
nand U8238 (N_8238,N_3376,N_3658);
and U8239 (N_8239,N_4013,N_4781);
nand U8240 (N_8240,N_2826,N_3805);
nor U8241 (N_8241,N_3894,N_86);
or U8242 (N_8242,N_89,N_4765);
or U8243 (N_8243,N_4613,N_1364);
nand U8244 (N_8244,N_3075,N_150);
nand U8245 (N_8245,N_4901,N_4651);
and U8246 (N_8246,N_2940,N_1945);
and U8247 (N_8247,N_4647,N_1549);
xor U8248 (N_8248,N_3307,N_3442);
and U8249 (N_8249,N_1579,N_523);
xor U8250 (N_8250,N_4829,N_1034);
nand U8251 (N_8251,N_890,N_641);
nand U8252 (N_8252,N_2955,N_3417);
nor U8253 (N_8253,N_2443,N_4299);
nand U8254 (N_8254,N_796,N_3825);
xor U8255 (N_8255,N_653,N_4899);
and U8256 (N_8256,N_4466,N_3020);
and U8257 (N_8257,N_4876,N_3056);
nor U8258 (N_8258,N_4729,N_3979);
nand U8259 (N_8259,N_2251,N_1330);
xor U8260 (N_8260,N_3739,N_1512);
nand U8261 (N_8261,N_3467,N_4058);
nand U8262 (N_8262,N_1808,N_3405);
or U8263 (N_8263,N_4159,N_775);
and U8264 (N_8264,N_1211,N_4455);
or U8265 (N_8265,N_1744,N_2609);
nor U8266 (N_8266,N_3505,N_18);
and U8267 (N_8267,N_1172,N_2251);
nor U8268 (N_8268,N_3370,N_2164);
and U8269 (N_8269,N_4293,N_2713);
nor U8270 (N_8270,N_1618,N_3593);
nor U8271 (N_8271,N_52,N_162);
or U8272 (N_8272,N_3265,N_1366);
and U8273 (N_8273,N_1723,N_1661);
nand U8274 (N_8274,N_450,N_1730);
nor U8275 (N_8275,N_4973,N_3058);
and U8276 (N_8276,N_1383,N_3396);
nand U8277 (N_8277,N_2835,N_2688);
and U8278 (N_8278,N_2079,N_1542);
and U8279 (N_8279,N_972,N_3469);
nand U8280 (N_8280,N_2063,N_4841);
nor U8281 (N_8281,N_1884,N_4266);
or U8282 (N_8282,N_1186,N_3367);
or U8283 (N_8283,N_1365,N_3602);
or U8284 (N_8284,N_3267,N_2370);
or U8285 (N_8285,N_1626,N_3240);
nor U8286 (N_8286,N_3995,N_1181);
and U8287 (N_8287,N_545,N_2971);
nand U8288 (N_8288,N_634,N_1424);
nor U8289 (N_8289,N_2809,N_4965);
nor U8290 (N_8290,N_2165,N_3481);
xnor U8291 (N_8291,N_2101,N_1528);
nand U8292 (N_8292,N_554,N_2242);
and U8293 (N_8293,N_448,N_2595);
and U8294 (N_8294,N_1624,N_845);
and U8295 (N_8295,N_3390,N_3782);
nor U8296 (N_8296,N_4848,N_2683);
nor U8297 (N_8297,N_215,N_4562);
nand U8298 (N_8298,N_1907,N_2880);
or U8299 (N_8299,N_4020,N_1113);
nand U8300 (N_8300,N_2633,N_3252);
nand U8301 (N_8301,N_4822,N_4516);
or U8302 (N_8302,N_793,N_4269);
nor U8303 (N_8303,N_3095,N_4455);
nor U8304 (N_8304,N_3237,N_1934);
xor U8305 (N_8305,N_3088,N_1540);
or U8306 (N_8306,N_2651,N_346);
nor U8307 (N_8307,N_461,N_3788);
nand U8308 (N_8308,N_697,N_4031);
or U8309 (N_8309,N_4896,N_1467);
nand U8310 (N_8310,N_2016,N_887);
and U8311 (N_8311,N_4189,N_3776);
nand U8312 (N_8312,N_3945,N_4904);
xor U8313 (N_8313,N_4468,N_1602);
nand U8314 (N_8314,N_515,N_3694);
or U8315 (N_8315,N_4104,N_3797);
and U8316 (N_8316,N_3447,N_4678);
nand U8317 (N_8317,N_3309,N_4879);
nor U8318 (N_8318,N_874,N_595);
and U8319 (N_8319,N_2419,N_2921);
and U8320 (N_8320,N_2972,N_1519);
and U8321 (N_8321,N_3458,N_3552);
or U8322 (N_8322,N_2941,N_3310);
nor U8323 (N_8323,N_1557,N_2578);
nor U8324 (N_8324,N_213,N_896);
or U8325 (N_8325,N_2878,N_2475);
and U8326 (N_8326,N_1268,N_1897);
and U8327 (N_8327,N_1632,N_610);
nor U8328 (N_8328,N_2163,N_3297);
or U8329 (N_8329,N_468,N_3790);
and U8330 (N_8330,N_1120,N_1441);
or U8331 (N_8331,N_3523,N_4494);
and U8332 (N_8332,N_2725,N_173);
nand U8333 (N_8333,N_3961,N_2059);
nand U8334 (N_8334,N_3863,N_3969);
nor U8335 (N_8335,N_868,N_4069);
nand U8336 (N_8336,N_2059,N_4372);
and U8337 (N_8337,N_3407,N_1393);
and U8338 (N_8338,N_4810,N_3952);
nor U8339 (N_8339,N_246,N_4823);
and U8340 (N_8340,N_592,N_2155);
xor U8341 (N_8341,N_2271,N_2744);
xor U8342 (N_8342,N_147,N_4);
nor U8343 (N_8343,N_3937,N_3644);
or U8344 (N_8344,N_225,N_2502);
nand U8345 (N_8345,N_3704,N_330);
xor U8346 (N_8346,N_626,N_51);
nor U8347 (N_8347,N_2779,N_1209);
and U8348 (N_8348,N_3365,N_662);
nor U8349 (N_8349,N_4680,N_678);
or U8350 (N_8350,N_2467,N_196);
nand U8351 (N_8351,N_626,N_2046);
nand U8352 (N_8352,N_2509,N_2716);
or U8353 (N_8353,N_2784,N_2160);
and U8354 (N_8354,N_480,N_4195);
xnor U8355 (N_8355,N_673,N_4963);
or U8356 (N_8356,N_2076,N_4256);
or U8357 (N_8357,N_1917,N_4663);
and U8358 (N_8358,N_65,N_211);
and U8359 (N_8359,N_938,N_1273);
and U8360 (N_8360,N_2840,N_3114);
nor U8361 (N_8361,N_828,N_754);
xnor U8362 (N_8362,N_4763,N_789);
nor U8363 (N_8363,N_4973,N_2370);
and U8364 (N_8364,N_4699,N_2975);
and U8365 (N_8365,N_1787,N_2152);
nor U8366 (N_8366,N_1297,N_3557);
or U8367 (N_8367,N_3855,N_2346);
xnor U8368 (N_8368,N_318,N_4747);
nand U8369 (N_8369,N_1523,N_4964);
and U8370 (N_8370,N_3965,N_1907);
and U8371 (N_8371,N_3302,N_4618);
and U8372 (N_8372,N_2339,N_2956);
or U8373 (N_8373,N_2082,N_2096);
nand U8374 (N_8374,N_1884,N_4336);
or U8375 (N_8375,N_3191,N_2977);
and U8376 (N_8376,N_2786,N_4533);
and U8377 (N_8377,N_2426,N_2222);
nor U8378 (N_8378,N_4360,N_1106);
nand U8379 (N_8379,N_4126,N_2762);
nand U8380 (N_8380,N_1070,N_3924);
nor U8381 (N_8381,N_2516,N_2572);
nor U8382 (N_8382,N_4693,N_1898);
nor U8383 (N_8383,N_3735,N_794);
and U8384 (N_8384,N_1624,N_346);
and U8385 (N_8385,N_2161,N_4359);
and U8386 (N_8386,N_4641,N_1582);
and U8387 (N_8387,N_3348,N_1400);
nor U8388 (N_8388,N_1348,N_4215);
nor U8389 (N_8389,N_3866,N_1799);
and U8390 (N_8390,N_2864,N_2177);
or U8391 (N_8391,N_4006,N_2239);
nand U8392 (N_8392,N_4975,N_4416);
or U8393 (N_8393,N_278,N_1469);
nand U8394 (N_8394,N_3595,N_928);
or U8395 (N_8395,N_685,N_1021);
nor U8396 (N_8396,N_3196,N_3664);
and U8397 (N_8397,N_2039,N_4384);
or U8398 (N_8398,N_1226,N_1348);
and U8399 (N_8399,N_3937,N_3411);
and U8400 (N_8400,N_1523,N_1979);
and U8401 (N_8401,N_2082,N_2649);
xor U8402 (N_8402,N_264,N_1211);
and U8403 (N_8403,N_1920,N_1150);
and U8404 (N_8404,N_53,N_321);
nand U8405 (N_8405,N_981,N_4607);
nor U8406 (N_8406,N_4843,N_923);
nor U8407 (N_8407,N_3664,N_207);
nand U8408 (N_8408,N_4744,N_1051);
nor U8409 (N_8409,N_4192,N_532);
and U8410 (N_8410,N_714,N_1394);
nor U8411 (N_8411,N_168,N_3163);
or U8412 (N_8412,N_2426,N_4354);
or U8413 (N_8413,N_110,N_1755);
xnor U8414 (N_8414,N_4387,N_4273);
nand U8415 (N_8415,N_2065,N_2472);
or U8416 (N_8416,N_168,N_2668);
or U8417 (N_8417,N_3777,N_3684);
or U8418 (N_8418,N_1862,N_4257);
nand U8419 (N_8419,N_731,N_1630);
xnor U8420 (N_8420,N_4091,N_793);
and U8421 (N_8421,N_2873,N_3122);
or U8422 (N_8422,N_571,N_4517);
and U8423 (N_8423,N_1866,N_4846);
nor U8424 (N_8424,N_1813,N_3758);
nor U8425 (N_8425,N_554,N_969);
or U8426 (N_8426,N_438,N_4630);
and U8427 (N_8427,N_2094,N_359);
nand U8428 (N_8428,N_3821,N_209);
nand U8429 (N_8429,N_44,N_4565);
nand U8430 (N_8430,N_341,N_3967);
or U8431 (N_8431,N_2502,N_2621);
or U8432 (N_8432,N_4820,N_1774);
xor U8433 (N_8433,N_2678,N_1826);
or U8434 (N_8434,N_1717,N_1322);
nand U8435 (N_8435,N_864,N_1159);
and U8436 (N_8436,N_1557,N_3633);
nor U8437 (N_8437,N_4454,N_1890);
or U8438 (N_8438,N_29,N_4542);
nor U8439 (N_8439,N_562,N_1706);
or U8440 (N_8440,N_884,N_2135);
or U8441 (N_8441,N_4643,N_3860);
nor U8442 (N_8442,N_2108,N_1395);
and U8443 (N_8443,N_1132,N_3619);
nand U8444 (N_8444,N_216,N_3833);
nand U8445 (N_8445,N_2568,N_1509);
or U8446 (N_8446,N_1825,N_4625);
nand U8447 (N_8447,N_4283,N_226);
nor U8448 (N_8448,N_1404,N_4938);
nand U8449 (N_8449,N_3513,N_4115);
nand U8450 (N_8450,N_1241,N_1450);
nand U8451 (N_8451,N_3232,N_1285);
nor U8452 (N_8452,N_4631,N_1115);
and U8453 (N_8453,N_4669,N_3792);
and U8454 (N_8454,N_3370,N_2093);
and U8455 (N_8455,N_224,N_4970);
nor U8456 (N_8456,N_3449,N_112);
nor U8457 (N_8457,N_4270,N_1669);
nand U8458 (N_8458,N_3232,N_1978);
or U8459 (N_8459,N_927,N_3425);
nor U8460 (N_8460,N_1570,N_4617);
nor U8461 (N_8461,N_4078,N_4538);
or U8462 (N_8462,N_2734,N_4232);
or U8463 (N_8463,N_2442,N_308);
or U8464 (N_8464,N_3608,N_2097);
and U8465 (N_8465,N_4400,N_4882);
or U8466 (N_8466,N_1808,N_2030);
or U8467 (N_8467,N_3346,N_4482);
nor U8468 (N_8468,N_597,N_109);
xor U8469 (N_8469,N_1323,N_1666);
xnor U8470 (N_8470,N_2700,N_676);
or U8471 (N_8471,N_3122,N_4574);
nor U8472 (N_8472,N_2032,N_4712);
nor U8473 (N_8473,N_3637,N_4118);
xor U8474 (N_8474,N_3401,N_2823);
and U8475 (N_8475,N_1998,N_822);
nor U8476 (N_8476,N_1593,N_3976);
nor U8477 (N_8477,N_1039,N_1978);
xor U8478 (N_8478,N_300,N_18);
nand U8479 (N_8479,N_225,N_3172);
xnor U8480 (N_8480,N_4306,N_1519);
nor U8481 (N_8481,N_181,N_3494);
nor U8482 (N_8482,N_133,N_3951);
nor U8483 (N_8483,N_2738,N_3446);
xor U8484 (N_8484,N_2086,N_485);
or U8485 (N_8485,N_82,N_681);
nor U8486 (N_8486,N_2568,N_1012);
and U8487 (N_8487,N_4178,N_4310);
nand U8488 (N_8488,N_1382,N_3468);
or U8489 (N_8489,N_1213,N_311);
nor U8490 (N_8490,N_140,N_4629);
nor U8491 (N_8491,N_4797,N_343);
nand U8492 (N_8492,N_1058,N_4905);
nor U8493 (N_8493,N_3174,N_3958);
xnor U8494 (N_8494,N_602,N_2370);
or U8495 (N_8495,N_4794,N_2191);
nor U8496 (N_8496,N_1471,N_501);
or U8497 (N_8497,N_515,N_134);
or U8498 (N_8498,N_4455,N_2570);
nand U8499 (N_8499,N_669,N_1592);
nand U8500 (N_8500,N_2891,N_3744);
nand U8501 (N_8501,N_932,N_548);
xor U8502 (N_8502,N_4799,N_2990);
nor U8503 (N_8503,N_588,N_3091);
nand U8504 (N_8504,N_2086,N_107);
or U8505 (N_8505,N_999,N_1149);
nor U8506 (N_8506,N_4366,N_922);
nand U8507 (N_8507,N_3872,N_1819);
and U8508 (N_8508,N_3251,N_4567);
xnor U8509 (N_8509,N_730,N_1042);
nor U8510 (N_8510,N_574,N_4430);
and U8511 (N_8511,N_1022,N_1752);
or U8512 (N_8512,N_2031,N_636);
nand U8513 (N_8513,N_1258,N_1463);
nor U8514 (N_8514,N_1722,N_4315);
nor U8515 (N_8515,N_3534,N_4126);
or U8516 (N_8516,N_3080,N_4461);
and U8517 (N_8517,N_2005,N_3020);
nand U8518 (N_8518,N_883,N_3240);
and U8519 (N_8519,N_4136,N_2156);
and U8520 (N_8520,N_3008,N_120);
and U8521 (N_8521,N_4837,N_2881);
nand U8522 (N_8522,N_1078,N_2188);
or U8523 (N_8523,N_1452,N_3881);
nand U8524 (N_8524,N_1295,N_851);
xor U8525 (N_8525,N_210,N_4755);
nand U8526 (N_8526,N_3419,N_2088);
nor U8527 (N_8527,N_1308,N_220);
or U8528 (N_8528,N_3348,N_3715);
and U8529 (N_8529,N_232,N_3304);
xor U8530 (N_8530,N_4082,N_2685);
nor U8531 (N_8531,N_723,N_3912);
or U8532 (N_8532,N_320,N_580);
nor U8533 (N_8533,N_262,N_4022);
nor U8534 (N_8534,N_1295,N_434);
or U8535 (N_8535,N_4724,N_1447);
nor U8536 (N_8536,N_4899,N_4097);
xor U8537 (N_8537,N_1161,N_1633);
nand U8538 (N_8538,N_221,N_1484);
or U8539 (N_8539,N_682,N_4658);
or U8540 (N_8540,N_3655,N_3861);
xor U8541 (N_8541,N_3896,N_2492);
and U8542 (N_8542,N_4539,N_3542);
and U8543 (N_8543,N_4780,N_186);
xnor U8544 (N_8544,N_3573,N_4448);
nand U8545 (N_8545,N_1924,N_4543);
nand U8546 (N_8546,N_3751,N_2955);
and U8547 (N_8547,N_1485,N_3370);
or U8548 (N_8548,N_2102,N_3253);
and U8549 (N_8549,N_3035,N_923);
nor U8550 (N_8550,N_1867,N_1694);
nor U8551 (N_8551,N_4956,N_4135);
nor U8552 (N_8552,N_2837,N_4831);
or U8553 (N_8553,N_2905,N_4270);
nor U8554 (N_8554,N_2579,N_2974);
nor U8555 (N_8555,N_769,N_4204);
or U8556 (N_8556,N_2729,N_539);
nand U8557 (N_8557,N_3339,N_672);
or U8558 (N_8558,N_2073,N_2572);
and U8559 (N_8559,N_4310,N_2204);
and U8560 (N_8560,N_4812,N_214);
and U8561 (N_8561,N_4752,N_648);
or U8562 (N_8562,N_4840,N_2493);
and U8563 (N_8563,N_1422,N_1818);
and U8564 (N_8564,N_2384,N_3195);
nor U8565 (N_8565,N_2446,N_3552);
and U8566 (N_8566,N_2423,N_82);
or U8567 (N_8567,N_3591,N_520);
nand U8568 (N_8568,N_4853,N_2352);
nor U8569 (N_8569,N_1199,N_2979);
xnor U8570 (N_8570,N_4344,N_4194);
or U8571 (N_8571,N_4389,N_3816);
nand U8572 (N_8572,N_4028,N_2916);
or U8573 (N_8573,N_1179,N_1778);
nor U8574 (N_8574,N_492,N_4783);
or U8575 (N_8575,N_3049,N_2898);
xnor U8576 (N_8576,N_2579,N_1336);
xor U8577 (N_8577,N_2361,N_2230);
and U8578 (N_8578,N_2068,N_2636);
or U8579 (N_8579,N_3862,N_2509);
nand U8580 (N_8580,N_1716,N_1614);
or U8581 (N_8581,N_3018,N_3006);
and U8582 (N_8582,N_4860,N_1849);
nand U8583 (N_8583,N_2594,N_3652);
and U8584 (N_8584,N_4407,N_4033);
or U8585 (N_8585,N_1011,N_888);
xor U8586 (N_8586,N_1764,N_1470);
or U8587 (N_8587,N_2557,N_751);
and U8588 (N_8588,N_3612,N_2526);
and U8589 (N_8589,N_629,N_880);
or U8590 (N_8590,N_4926,N_2353);
and U8591 (N_8591,N_3052,N_2050);
nor U8592 (N_8592,N_2814,N_2384);
and U8593 (N_8593,N_3409,N_4183);
nor U8594 (N_8594,N_1279,N_1354);
or U8595 (N_8595,N_2241,N_3615);
and U8596 (N_8596,N_640,N_970);
xnor U8597 (N_8597,N_1667,N_393);
nor U8598 (N_8598,N_1606,N_456);
or U8599 (N_8599,N_301,N_4373);
or U8600 (N_8600,N_4612,N_4730);
xor U8601 (N_8601,N_2257,N_646);
nand U8602 (N_8602,N_1949,N_1006);
nand U8603 (N_8603,N_2547,N_560);
nand U8604 (N_8604,N_3703,N_1683);
nand U8605 (N_8605,N_4193,N_2346);
xor U8606 (N_8606,N_4805,N_3830);
and U8607 (N_8607,N_72,N_1280);
nor U8608 (N_8608,N_2455,N_1666);
or U8609 (N_8609,N_3191,N_4211);
or U8610 (N_8610,N_2005,N_3620);
or U8611 (N_8611,N_323,N_3469);
nor U8612 (N_8612,N_1781,N_1395);
nor U8613 (N_8613,N_2853,N_322);
nand U8614 (N_8614,N_628,N_3860);
xor U8615 (N_8615,N_1573,N_816);
nor U8616 (N_8616,N_3453,N_867);
nor U8617 (N_8617,N_1629,N_749);
or U8618 (N_8618,N_2865,N_1413);
and U8619 (N_8619,N_3075,N_2872);
nand U8620 (N_8620,N_1086,N_4406);
xnor U8621 (N_8621,N_2958,N_1550);
xnor U8622 (N_8622,N_369,N_1350);
or U8623 (N_8623,N_135,N_3003);
or U8624 (N_8624,N_1888,N_1648);
and U8625 (N_8625,N_1951,N_3632);
and U8626 (N_8626,N_2745,N_3845);
xor U8627 (N_8627,N_820,N_852);
nor U8628 (N_8628,N_3578,N_3011);
nor U8629 (N_8629,N_286,N_2218);
or U8630 (N_8630,N_3322,N_4582);
and U8631 (N_8631,N_1301,N_175);
nand U8632 (N_8632,N_3971,N_3401);
nand U8633 (N_8633,N_4699,N_166);
or U8634 (N_8634,N_4880,N_3374);
or U8635 (N_8635,N_3029,N_1627);
and U8636 (N_8636,N_3673,N_485);
nand U8637 (N_8637,N_1091,N_2633);
nor U8638 (N_8638,N_3330,N_707);
and U8639 (N_8639,N_4757,N_1981);
or U8640 (N_8640,N_2275,N_778);
nor U8641 (N_8641,N_626,N_1522);
or U8642 (N_8642,N_2707,N_1446);
nand U8643 (N_8643,N_3788,N_4052);
and U8644 (N_8644,N_2424,N_4697);
nor U8645 (N_8645,N_4175,N_3162);
and U8646 (N_8646,N_2382,N_4042);
nor U8647 (N_8647,N_3262,N_160);
and U8648 (N_8648,N_2071,N_2304);
or U8649 (N_8649,N_3676,N_2227);
nand U8650 (N_8650,N_4669,N_652);
and U8651 (N_8651,N_2877,N_744);
or U8652 (N_8652,N_4329,N_4608);
nor U8653 (N_8653,N_1236,N_2191);
nor U8654 (N_8654,N_184,N_3280);
nand U8655 (N_8655,N_1022,N_1691);
or U8656 (N_8656,N_24,N_4622);
xnor U8657 (N_8657,N_4677,N_2428);
nor U8658 (N_8658,N_2081,N_4630);
nor U8659 (N_8659,N_919,N_3009);
xor U8660 (N_8660,N_1018,N_642);
and U8661 (N_8661,N_213,N_2040);
nand U8662 (N_8662,N_2969,N_3216);
nand U8663 (N_8663,N_3703,N_4364);
nand U8664 (N_8664,N_2495,N_2993);
nand U8665 (N_8665,N_1255,N_4030);
and U8666 (N_8666,N_2116,N_3219);
nand U8667 (N_8667,N_3552,N_2056);
or U8668 (N_8668,N_3814,N_2833);
and U8669 (N_8669,N_3980,N_1096);
nand U8670 (N_8670,N_4019,N_3801);
nand U8671 (N_8671,N_861,N_4083);
and U8672 (N_8672,N_4949,N_1270);
or U8673 (N_8673,N_3279,N_3311);
nor U8674 (N_8674,N_1875,N_4861);
nand U8675 (N_8675,N_425,N_4172);
xnor U8676 (N_8676,N_1469,N_1134);
or U8677 (N_8677,N_1884,N_983);
nand U8678 (N_8678,N_2401,N_2392);
nand U8679 (N_8679,N_419,N_1839);
nor U8680 (N_8680,N_3369,N_3894);
nand U8681 (N_8681,N_3019,N_3288);
nor U8682 (N_8682,N_4130,N_4943);
nand U8683 (N_8683,N_4946,N_1644);
and U8684 (N_8684,N_1864,N_2127);
nor U8685 (N_8685,N_3817,N_3993);
and U8686 (N_8686,N_1090,N_4505);
and U8687 (N_8687,N_2876,N_3410);
and U8688 (N_8688,N_4062,N_3299);
nand U8689 (N_8689,N_2752,N_2894);
or U8690 (N_8690,N_243,N_2146);
nand U8691 (N_8691,N_2065,N_1102);
nor U8692 (N_8692,N_4921,N_3898);
xnor U8693 (N_8693,N_3761,N_1104);
nand U8694 (N_8694,N_3635,N_2844);
and U8695 (N_8695,N_178,N_4412);
nand U8696 (N_8696,N_4722,N_381);
nand U8697 (N_8697,N_2688,N_2218);
nor U8698 (N_8698,N_4461,N_1403);
nand U8699 (N_8699,N_1091,N_4613);
nor U8700 (N_8700,N_407,N_3736);
or U8701 (N_8701,N_2144,N_4569);
nand U8702 (N_8702,N_169,N_1237);
and U8703 (N_8703,N_864,N_586);
and U8704 (N_8704,N_205,N_3820);
or U8705 (N_8705,N_730,N_1889);
nand U8706 (N_8706,N_4626,N_1970);
nand U8707 (N_8707,N_3848,N_2100);
nand U8708 (N_8708,N_3978,N_2034);
nand U8709 (N_8709,N_3430,N_3621);
and U8710 (N_8710,N_2838,N_628);
and U8711 (N_8711,N_658,N_3769);
nor U8712 (N_8712,N_1270,N_2867);
and U8713 (N_8713,N_2094,N_3204);
and U8714 (N_8714,N_794,N_972);
nand U8715 (N_8715,N_954,N_1047);
and U8716 (N_8716,N_297,N_3165);
xor U8717 (N_8717,N_138,N_2240);
nor U8718 (N_8718,N_3020,N_2823);
and U8719 (N_8719,N_4259,N_3076);
nand U8720 (N_8720,N_2794,N_618);
or U8721 (N_8721,N_3473,N_3342);
nand U8722 (N_8722,N_1834,N_4182);
or U8723 (N_8723,N_2494,N_3705);
and U8724 (N_8724,N_2867,N_4464);
or U8725 (N_8725,N_494,N_3037);
and U8726 (N_8726,N_3255,N_2372);
nor U8727 (N_8727,N_3182,N_3642);
or U8728 (N_8728,N_2694,N_3091);
or U8729 (N_8729,N_1500,N_714);
and U8730 (N_8730,N_2129,N_4034);
and U8731 (N_8731,N_1958,N_164);
and U8732 (N_8732,N_1806,N_4490);
and U8733 (N_8733,N_4818,N_2910);
or U8734 (N_8734,N_2012,N_4464);
nor U8735 (N_8735,N_2473,N_2293);
xor U8736 (N_8736,N_2842,N_3815);
nand U8737 (N_8737,N_1574,N_3521);
and U8738 (N_8738,N_3743,N_2540);
nor U8739 (N_8739,N_1969,N_3526);
nor U8740 (N_8740,N_3843,N_2352);
or U8741 (N_8741,N_4062,N_998);
xnor U8742 (N_8742,N_4012,N_1657);
or U8743 (N_8743,N_4754,N_1459);
nand U8744 (N_8744,N_1666,N_4096);
nand U8745 (N_8745,N_3102,N_1857);
or U8746 (N_8746,N_2243,N_1736);
and U8747 (N_8747,N_1837,N_4069);
nand U8748 (N_8748,N_4281,N_4691);
and U8749 (N_8749,N_3852,N_679);
or U8750 (N_8750,N_2372,N_611);
nand U8751 (N_8751,N_3795,N_710);
or U8752 (N_8752,N_4325,N_4889);
and U8753 (N_8753,N_2926,N_3278);
nor U8754 (N_8754,N_4208,N_3949);
and U8755 (N_8755,N_4558,N_1730);
nand U8756 (N_8756,N_1744,N_1870);
and U8757 (N_8757,N_3371,N_3039);
nor U8758 (N_8758,N_4981,N_4045);
or U8759 (N_8759,N_2733,N_803);
or U8760 (N_8760,N_2163,N_1705);
nand U8761 (N_8761,N_4128,N_1304);
xor U8762 (N_8762,N_2806,N_4713);
xor U8763 (N_8763,N_1074,N_3975);
nor U8764 (N_8764,N_2810,N_4640);
nand U8765 (N_8765,N_834,N_3094);
nor U8766 (N_8766,N_933,N_333);
and U8767 (N_8767,N_78,N_3981);
nand U8768 (N_8768,N_4745,N_683);
nor U8769 (N_8769,N_4706,N_2694);
nand U8770 (N_8770,N_1366,N_688);
nor U8771 (N_8771,N_3416,N_3015);
or U8772 (N_8772,N_4852,N_3622);
or U8773 (N_8773,N_3871,N_1517);
nor U8774 (N_8774,N_4345,N_1089);
nor U8775 (N_8775,N_4877,N_2889);
and U8776 (N_8776,N_636,N_1823);
nor U8777 (N_8777,N_755,N_1962);
nand U8778 (N_8778,N_3467,N_1208);
or U8779 (N_8779,N_805,N_2845);
nor U8780 (N_8780,N_2228,N_1822);
and U8781 (N_8781,N_1949,N_2696);
nor U8782 (N_8782,N_909,N_959);
or U8783 (N_8783,N_890,N_1175);
nand U8784 (N_8784,N_3513,N_963);
nand U8785 (N_8785,N_540,N_4737);
nor U8786 (N_8786,N_3722,N_3841);
nand U8787 (N_8787,N_4126,N_95);
nand U8788 (N_8788,N_1401,N_3173);
nand U8789 (N_8789,N_2863,N_2070);
or U8790 (N_8790,N_1198,N_2870);
nor U8791 (N_8791,N_2223,N_2329);
nor U8792 (N_8792,N_3761,N_1629);
xor U8793 (N_8793,N_679,N_697);
and U8794 (N_8794,N_2730,N_2876);
and U8795 (N_8795,N_3287,N_826);
nor U8796 (N_8796,N_2128,N_1038);
nand U8797 (N_8797,N_3499,N_2440);
xor U8798 (N_8798,N_941,N_3943);
or U8799 (N_8799,N_2463,N_4393);
and U8800 (N_8800,N_2437,N_2155);
nand U8801 (N_8801,N_4732,N_2443);
xnor U8802 (N_8802,N_1901,N_1091);
nand U8803 (N_8803,N_3309,N_4388);
or U8804 (N_8804,N_1100,N_1081);
nor U8805 (N_8805,N_398,N_4667);
nand U8806 (N_8806,N_3808,N_785);
xnor U8807 (N_8807,N_556,N_1519);
nor U8808 (N_8808,N_4089,N_4179);
or U8809 (N_8809,N_2859,N_305);
xor U8810 (N_8810,N_3481,N_4441);
nor U8811 (N_8811,N_4895,N_904);
nor U8812 (N_8812,N_51,N_1081);
nand U8813 (N_8813,N_2061,N_4941);
nand U8814 (N_8814,N_3080,N_1118);
or U8815 (N_8815,N_649,N_4203);
and U8816 (N_8816,N_1638,N_669);
or U8817 (N_8817,N_1803,N_1717);
and U8818 (N_8818,N_1057,N_1869);
and U8819 (N_8819,N_3267,N_1331);
nand U8820 (N_8820,N_1774,N_3752);
nor U8821 (N_8821,N_2654,N_4601);
nor U8822 (N_8822,N_4545,N_2490);
and U8823 (N_8823,N_2209,N_4145);
nor U8824 (N_8824,N_2638,N_847);
nor U8825 (N_8825,N_3057,N_1530);
and U8826 (N_8826,N_3916,N_21);
or U8827 (N_8827,N_1061,N_854);
or U8828 (N_8828,N_4103,N_166);
nand U8829 (N_8829,N_3518,N_2712);
nor U8830 (N_8830,N_1060,N_3529);
nand U8831 (N_8831,N_3462,N_498);
or U8832 (N_8832,N_2474,N_3456);
nand U8833 (N_8833,N_1385,N_1617);
nor U8834 (N_8834,N_2376,N_3221);
nor U8835 (N_8835,N_1480,N_966);
nand U8836 (N_8836,N_3704,N_2380);
nand U8837 (N_8837,N_2070,N_942);
nand U8838 (N_8838,N_3373,N_4576);
xnor U8839 (N_8839,N_1170,N_3845);
nor U8840 (N_8840,N_1184,N_1208);
and U8841 (N_8841,N_1536,N_2123);
nor U8842 (N_8842,N_1782,N_721);
nor U8843 (N_8843,N_901,N_4367);
nor U8844 (N_8844,N_3128,N_637);
or U8845 (N_8845,N_1940,N_314);
nor U8846 (N_8846,N_755,N_594);
nor U8847 (N_8847,N_3969,N_4516);
nand U8848 (N_8848,N_1060,N_507);
and U8849 (N_8849,N_2515,N_3228);
and U8850 (N_8850,N_3273,N_1155);
xnor U8851 (N_8851,N_1291,N_4088);
and U8852 (N_8852,N_4248,N_3820);
nor U8853 (N_8853,N_4757,N_4031);
nor U8854 (N_8854,N_3273,N_3010);
nand U8855 (N_8855,N_3065,N_4433);
nand U8856 (N_8856,N_487,N_1275);
nor U8857 (N_8857,N_1836,N_3088);
xor U8858 (N_8858,N_3714,N_4633);
and U8859 (N_8859,N_4362,N_3453);
xnor U8860 (N_8860,N_1331,N_1537);
xor U8861 (N_8861,N_4445,N_1953);
or U8862 (N_8862,N_2892,N_4551);
and U8863 (N_8863,N_4407,N_463);
nand U8864 (N_8864,N_212,N_3156);
nand U8865 (N_8865,N_4202,N_752);
nor U8866 (N_8866,N_2779,N_4583);
or U8867 (N_8867,N_3192,N_4110);
and U8868 (N_8868,N_2249,N_2442);
xor U8869 (N_8869,N_1008,N_2351);
nor U8870 (N_8870,N_2441,N_595);
nand U8871 (N_8871,N_43,N_2438);
and U8872 (N_8872,N_1313,N_77);
xnor U8873 (N_8873,N_4675,N_1045);
or U8874 (N_8874,N_3178,N_208);
and U8875 (N_8875,N_1328,N_3250);
and U8876 (N_8876,N_2066,N_2919);
nand U8877 (N_8877,N_3971,N_730);
nand U8878 (N_8878,N_376,N_336);
nor U8879 (N_8879,N_3083,N_3063);
nand U8880 (N_8880,N_2332,N_1013);
and U8881 (N_8881,N_4005,N_343);
or U8882 (N_8882,N_1954,N_2765);
and U8883 (N_8883,N_1567,N_98);
and U8884 (N_8884,N_1264,N_182);
nand U8885 (N_8885,N_4357,N_4188);
and U8886 (N_8886,N_4791,N_986);
or U8887 (N_8887,N_2000,N_3274);
and U8888 (N_8888,N_4153,N_613);
nor U8889 (N_8889,N_103,N_2837);
nand U8890 (N_8890,N_2824,N_1123);
nor U8891 (N_8891,N_1553,N_2371);
and U8892 (N_8892,N_1187,N_4166);
and U8893 (N_8893,N_3417,N_2510);
and U8894 (N_8894,N_827,N_4131);
or U8895 (N_8895,N_3509,N_1538);
nor U8896 (N_8896,N_777,N_367);
and U8897 (N_8897,N_375,N_3671);
nor U8898 (N_8898,N_157,N_4530);
nand U8899 (N_8899,N_1548,N_3138);
nor U8900 (N_8900,N_4844,N_3259);
or U8901 (N_8901,N_4840,N_4234);
or U8902 (N_8902,N_2813,N_1357);
and U8903 (N_8903,N_2472,N_4306);
xor U8904 (N_8904,N_1255,N_309);
nor U8905 (N_8905,N_1648,N_662);
or U8906 (N_8906,N_659,N_2232);
nor U8907 (N_8907,N_2948,N_1620);
and U8908 (N_8908,N_4676,N_3758);
nand U8909 (N_8909,N_3792,N_2474);
nor U8910 (N_8910,N_4635,N_4992);
and U8911 (N_8911,N_4849,N_3683);
and U8912 (N_8912,N_3475,N_3885);
xor U8913 (N_8913,N_4179,N_86);
and U8914 (N_8914,N_4953,N_915);
nor U8915 (N_8915,N_154,N_4141);
or U8916 (N_8916,N_1146,N_1170);
and U8917 (N_8917,N_538,N_3069);
and U8918 (N_8918,N_3631,N_4034);
and U8919 (N_8919,N_61,N_2853);
nor U8920 (N_8920,N_1960,N_4406);
and U8921 (N_8921,N_3419,N_915);
xnor U8922 (N_8922,N_403,N_2593);
nand U8923 (N_8923,N_2525,N_4044);
or U8924 (N_8924,N_722,N_4810);
and U8925 (N_8925,N_3942,N_4504);
and U8926 (N_8926,N_530,N_3719);
nand U8927 (N_8927,N_3951,N_4110);
and U8928 (N_8928,N_648,N_4075);
nor U8929 (N_8929,N_659,N_1513);
nand U8930 (N_8930,N_1944,N_1875);
xnor U8931 (N_8931,N_908,N_4292);
or U8932 (N_8932,N_4287,N_2709);
or U8933 (N_8933,N_1532,N_3037);
or U8934 (N_8934,N_2589,N_1023);
and U8935 (N_8935,N_908,N_9);
and U8936 (N_8936,N_3783,N_2795);
nand U8937 (N_8937,N_1872,N_329);
xor U8938 (N_8938,N_2788,N_519);
nor U8939 (N_8939,N_4339,N_2760);
and U8940 (N_8940,N_835,N_4585);
xor U8941 (N_8941,N_3055,N_1714);
nand U8942 (N_8942,N_260,N_967);
xnor U8943 (N_8943,N_395,N_1284);
and U8944 (N_8944,N_342,N_1886);
nand U8945 (N_8945,N_183,N_2017);
and U8946 (N_8946,N_1418,N_2658);
or U8947 (N_8947,N_1938,N_197);
xor U8948 (N_8948,N_4738,N_4845);
and U8949 (N_8949,N_3127,N_1267);
nor U8950 (N_8950,N_892,N_3753);
nor U8951 (N_8951,N_4951,N_3084);
nor U8952 (N_8952,N_1184,N_1916);
nor U8953 (N_8953,N_554,N_3277);
or U8954 (N_8954,N_4198,N_1005);
or U8955 (N_8955,N_1759,N_4068);
nand U8956 (N_8956,N_4555,N_215);
or U8957 (N_8957,N_2584,N_4513);
xnor U8958 (N_8958,N_2380,N_940);
nand U8959 (N_8959,N_530,N_4849);
or U8960 (N_8960,N_2973,N_789);
or U8961 (N_8961,N_3417,N_3973);
or U8962 (N_8962,N_4196,N_3239);
or U8963 (N_8963,N_3748,N_1679);
nor U8964 (N_8964,N_1087,N_4547);
or U8965 (N_8965,N_685,N_4608);
or U8966 (N_8966,N_2165,N_470);
nand U8967 (N_8967,N_3653,N_2483);
nand U8968 (N_8968,N_2818,N_3531);
nand U8969 (N_8969,N_2569,N_4203);
and U8970 (N_8970,N_3129,N_4476);
nand U8971 (N_8971,N_419,N_413);
or U8972 (N_8972,N_1298,N_1809);
nand U8973 (N_8973,N_4282,N_3639);
nand U8974 (N_8974,N_3263,N_1583);
or U8975 (N_8975,N_2647,N_649);
nand U8976 (N_8976,N_3296,N_1440);
nor U8977 (N_8977,N_4909,N_4311);
nand U8978 (N_8978,N_81,N_3859);
xor U8979 (N_8979,N_2533,N_4610);
and U8980 (N_8980,N_2630,N_4021);
or U8981 (N_8981,N_2096,N_2501);
and U8982 (N_8982,N_4502,N_1914);
nand U8983 (N_8983,N_1204,N_4527);
xnor U8984 (N_8984,N_4390,N_4682);
or U8985 (N_8985,N_784,N_2041);
and U8986 (N_8986,N_46,N_1041);
or U8987 (N_8987,N_3460,N_1754);
or U8988 (N_8988,N_1051,N_2899);
and U8989 (N_8989,N_4671,N_2858);
or U8990 (N_8990,N_3351,N_2497);
nand U8991 (N_8991,N_1872,N_2078);
and U8992 (N_8992,N_224,N_4675);
or U8993 (N_8993,N_4186,N_2136);
and U8994 (N_8994,N_2329,N_2877);
nand U8995 (N_8995,N_4388,N_462);
nand U8996 (N_8996,N_4472,N_3114);
nor U8997 (N_8997,N_4133,N_1952);
nor U8998 (N_8998,N_724,N_139);
nor U8999 (N_8999,N_3068,N_2614);
nand U9000 (N_9000,N_694,N_1170);
and U9001 (N_9001,N_961,N_1549);
or U9002 (N_9002,N_565,N_3438);
nor U9003 (N_9003,N_2262,N_2303);
and U9004 (N_9004,N_4154,N_1937);
or U9005 (N_9005,N_2191,N_3455);
and U9006 (N_9006,N_542,N_4111);
and U9007 (N_9007,N_4549,N_3335);
and U9008 (N_9008,N_1828,N_4069);
nand U9009 (N_9009,N_1445,N_3649);
nand U9010 (N_9010,N_2203,N_2131);
xnor U9011 (N_9011,N_3475,N_490);
nor U9012 (N_9012,N_2037,N_439);
xor U9013 (N_9013,N_829,N_1703);
nand U9014 (N_9014,N_1540,N_4409);
nand U9015 (N_9015,N_4911,N_1217);
and U9016 (N_9016,N_3648,N_4922);
nand U9017 (N_9017,N_440,N_2924);
nor U9018 (N_9018,N_2191,N_2111);
nand U9019 (N_9019,N_1766,N_3362);
or U9020 (N_9020,N_3202,N_3770);
or U9021 (N_9021,N_868,N_1881);
nand U9022 (N_9022,N_823,N_202);
nand U9023 (N_9023,N_1822,N_3622);
nor U9024 (N_9024,N_2580,N_2452);
nor U9025 (N_9025,N_2296,N_2461);
or U9026 (N_9026,N_364,N_629);
and U9027 (N_9027,N_2944,N_2795);
and U9028 (N_9028,N_4673,N_3526);
or U9029 (N_9029,N_3611,N_3501);
or U9030 (N_9030,N_2536,N_805);
nand U9031 (N_9031,N_1533,N_275);
or U9032 (N_9032,N_3385,N_4067);
nand U9033 (N_9033,N_4225,N_2782);
nor U9034 (N_9034,N_2860,N_1372);
nor U9035 (N_9035,N_1360,N_3695);
xnor U9036 (N_9036,N_1152,N_296);
nor U9037 (N_9037,N_2367,N_2941);
and U9038 (N_9038,N_3351,N_2034);
and U9039 (N_9039,N_179,N_4123);
or U9040 (N_9040,N_2718,N_3258);
and U9041 (N_9041,N_4384,N_4789);
or U9042 (N_9042,N_533,N_2147);
and U9043 (N_9043,N_3078,N_4943);
or U9044 (N_9044,N_4796,N_4855);
nor U9045 (N_9045,N_479,N_698);
xnor U9046 (N_9046,N_1974,N_2821);
or U9047 (N_9047,N_683,N_3146);
nor U9048 (N_9048,N_853,N_3952);
and U9049 (N_9049,N_4510,N_4029);
xnor U9050 (N_9050,N_4891,N_2229);
nand U9051 (N_9051,N_32,N_2136);
or U9052 (N_9052,N_2313,N_588);
or U9053 (N_9053,N_2102,N_4961);
nand U9054 (N_9054,N_4353,N_483);
and U9055 (N_9055,N_3188,N_3292);
or U9056 (N_9056,N_4514,N_4915);
or U9057 (N_9057,N_710,N_4682);
and U9058 (N_9058,N_2443,N_3163);
and U9059 (N_9059,N_596,N_630);
nor U9060 (N_9060,N_504,N_4501);
nor U9061 (N_9061,N_4973,N_524);
nand U9062 (N_9062,N_1013,N_3500);
nor U9063 (N_9063,N_2550,N_2340);
xor U9064 (N_9064,N_3991,N_259);
xor U9065 (N_9065,N_4524,N_751);
and U9066 (N_9066,N_4197,N_23);
or U9067 (N_9067,N_4307,N_3611);
nand U9068 (N_9068,N_283,N_4102);
and U9069 (N_9069,N_127,N_1997);
nand U9070 (N_9070,N_3719,N_1658);
xnor U9071 (N_9071,N_1098,N_2092);
nor U9072 (N_9072,N_4874,N_305);
nand U9073 (N_9073,N_2592,N_2054);
nor U9074 (N_9074,N_2622,N_4597);
and U9075 (N_9075,N_4199,N_2161);
or U9076 (N_9076,N_4835,N_2386);
and U9077 (N_9077,N_1308,N_3088);
or U9078 (N_9078,N_3004,N_1005);
nand U9079 (N_9079,N_939,N_1526);
nand U9080 (N_9080,N_738,N_1091);
and U9081 (N_9081,N_4285,N_720);
nor U9082 (N_9082,N_4672,N_4478);
nand U9083 (N_9083,N_736,N_2428);
and U9084 (N_9084,N_1400,N_898);
nand U9085 (N_9085,N_2374,N_380);
xnor U9086 (N_9086,N_3412,N_4532);
nand U9087 (N_9087,N_965,N_4293);
nand U9088 (N_9088,N_1034,N_2628);
and U9089 (N_9089,N_1378,N_3436);
nor U9090 (N_9090,N_4435,N_3287);
nand U9091 (N_9091,N_892,N_3217);
nor U9092 (N_9092,N_4900,N_3230);
and U9093 (N_9093,N_1423,N_506);
nor U9094 (N_9094,N_749,N_4689);
nand U9095 (N_9095,N_2589,N_859);
nor U9096 (N_9096,N_688,N_2745);
nor U9097 (N_9097,N_2509,N_4283);
or U9098 (N_9098,N_290,N_4532);
nor U9099 (N_9099,N_47,N_609);
and U9100 (N_9100,N_3405,N_4909);
nand U9101 (N_9101,N_4638,N_1113);
nor U9102 (N_9102,N_4173,N_4461);
nor U9103 (N_9103,N_334,N_3361);
and U9104 (N_9104,N_2629,N_4871);
and U9105 (N_9105,N_4207,N_634);
nand U9106 (N_9106,N_3543,N_3910);
or U9107 (N_9107,N_3706,N_4315);
and U9108 (N_9108,N_4826,N_4488);
nand U9109 (N_9109,N_725,N_1287);
nor U9110 (N_9110,N_3121,N_1375);
nand U9111 (N_9111,N_1280,N_70);
or U9112 (N_9112,N_55,N_1905);
nor U9113 (N_9113,N_1988,N_719);
nor U9114 (N_9114,N_4868,N_1745);
nand U9115 (N_9115,N_2286,N_4637);
nor U9116 (N_9116,N_1151,N_1576);
nor U9117 (N_9117,N_3999,N_3159);
nand U9118 (N_9118,N_621,N_2831);
nand U9119 (N_9119,N_2906,N_3303);
xor U9120 (N_9120,N_335,N_2373);
or U9121 (N_9121,N_1502,N_843);
and U9122 (N_9122,N_3579,N_4198);
nor U9123 (N_9123,N_4171,N_1954);
nand U9124 (N_9124,N_2011,N_1784);
nor U9125 (N_9125,N_3107,N_4569);
nor U9126 (N_9126,N_2808,N_1884);
nand U9127 (N_9127,N_1257,N_4399);
and U9128 (N_9128,N_3713,N_2644);
nand U9129 (N_9129,N_4059,N_2066);
or U9130 (N_9130,N_2531,N_4562);
or U9131 (N_9131,N_1184,N_3170);
nand U9132 (N_9132,N_637,N_4586);
and U9133 (N_9133,N_4836,N_1306);
nor U9134 (N_9134,N_2659,N_3040);
or U9135 (N_9135,N_569,N_1760);
nand U9136 (N_9136,N_737,N_4773);
and U9137 (N_9137,N_44,N_4214);
and U9138 (N_9138,N_1271,N_1630);
nor U9139 (N_9139,N_642,N_3203);
or U9140 (N_9140,N_2444,N_2726);
or U9141 (N_9141,N_2470,N_4714);
nor U9142 (N_9142,N_4794,N_3548);
nor U9143 (N_9143,N_1343,N_4330);
xor U9144 (N_9144,N_150,N_2332);
xor U9145 (N_9145,N_178,N_4842);
nor U9146 (N_9146,N_4298,N_1092);
nor U9147 (N_9147,N_3352,N_3875);
nor U9148 (N_9148,N_4893,N_719);
nand U9149 (N_9149,N_2725,N_4829);
and U9150 (N_9150,N_2131,N_4048);
nor U9151 (N_9151,N_869,N_961);
xnor U9152 (N_9152,N_883,N_2029);
nand U9153 (N_9153,N_320,N_1171);
nor U9154 (N_9154,N_311,N_1097);
and U9155 (N_9155,N_3874,N_3227);
or U9156 (N_9156,N_280,N_560);
nand U9157 (N_9157,N_2038,N_235);
xnor U9158 (N_9158,N_2651,N_2036);
or U9159 (N_9159,N_3192,N_614);
or U9160 (N_9160,N_4476,N_1482);
nand U9161 (N_9161,N_4970,N_3061);
and U9162 (N_9162,N_2515,N_4538);
nor U9163 (N_9163,N_993,N_4655);
nor U9164 (N_9164,N_3314,N_4998);
or U9165 (N_9165,N_3089,N_704);
nor U9166 (N_9166,N_109,N_4193);
nor U9167 (N_9167,N_3033,N_2985);
nand U9168 (N_9168,N_671,N_2662);
and U9169 (N_9169,N_3908,N_1867);
nand U9170 (N_9170,N_4996,N_4830);
and U9171 (N_9171,N_4540,N_865);
and U9172 (N_9172,N_4772,N_2447);
xnor U9173 (N_9173,N_2604,N_3765);
or U9174 (N_9174,N_4814,N_4704);
and U9175 (N_9175,N_44,N_2419);
nor U9176 (N_9176,N_115,N_3941);
nor U9177 (N_9177,N_2694,N_1770);
or U9178 (N_9178,N_2231,N_52);
and U9179 (N_9179,N_2766,N_3790);
nor U9180 (N_9180,N_3238,N_2421);
or U9181 (N_9181,N_2348,N_1527);
or U9182 (N_9182,N_2643,N_4345);
or U9183 (N_9183,N_2299,N_1235);
xor U9184 (N_9184,N_3609,N_1371);
xnor U9185 (N_9185,N_2064,N_4910);
nor U9186 (N_9186,N_1463,N_639);
or U9187 (N_9187,N_3271,N_3645);
or U9188 (N_9188,N_4081,N_4761);
nand U9189 (N_9189,N_3668,N_3291);
nor U9190 (N_9190,N_2327,N_3335);
nand U9191 (N_9191,N_3393,N_3607);
xor U9192 (N_9192,N_4005,N_4602);
xor U9193 (N_9193,N_3439,N_1081);
nand U9194 (N_9194,N_2128,N_1522);
nand U9195 (N_9195,N_3208,N_1983);
xnor U9196 (N_9196,N_138,N_2626);
and U9197 (N_9197,N_4151,N_2559);
nand U9198 (N_9198,N_3910,N_1187);
nand U9199 (N_9199,N_4569,N_3157);
or U9200 (N_9200,N_4758,N_2918);
nor U9201 (N_9201,N_2155,N_3027);
or U9202 (N_9202,N_2679,N_1424);
nor U9203 (N_9203,N_456,N_969);
or U9204 (N_9204,N_310,N_2918);
or U9205 (N_9205,N_537,N_2940);
and U9206 (N_9206,N_4340,N_2192);
nand U9207 (N_9207,N_4769,N_4146);
nor U9208 (N_9208,N_1368,N_2647);
nand U9209 (N_9209,N_665,N_3670);
nor U9210 (N_9210,N_848,N_2841);
and U9211 (N_9211,N_4714,N_1121);
nand U9212 (N_9212,N_3080,N_3774);
or U9213 (N_9213,N_3806,N_432);
or U9214 (N_9214,N_2639,N_1525);
nor U9215 (N_9215,N_3080,N_2620);
nor U9216 (N_9216,N_497,N_2629);
nand U9217 (N_9217,N_1465,N_1421);
and U9218 (N_9218,N_4090,N_3681);
nand U9219 (N_9219,N_3681,N_4140);
nand U9220 (N_9220,N_1491,N_4948);
nor U9221 (N_9221,N_1887,N_1152);
or U9222 (N_9222,N_53,N_2572);
nor U9223 (N_9223,N_1784,N_574);
and U9224 (N_9224,N_102,N_1222);
or U9225 (N_9225,N_1144,N_3380);
nor U9226 (N_9226,N_2849,N_1847);
nand U9227 (N_9227,N_3544,N_2839);
nand U9228 (N_9228,N_2257,N_3691);
or U9229 (N_9229,N_3625,N_3933);
nor U9230 (N_9230,N_1782,N_699);
or U9231 (N_9231,N_4996,N_3141);
or U9232 (N_9232,N_4553,N_2608);
nand U9233 (N_9233,N_4322,N_4291);
or U9234 (N_9234,N_2948,N_162);
nand U9235 (N_9235,N_3941,N_2066);
nor U9236 (N_9236,N_3228,N_2112);
or U9237 (N_9237,N_1232,N_3258);
or U9238 (N_9238,N_147,N_2985);
or U9239 (N_9239,N_1687,N_2768);
or U9240 (N_9240,N_3647,N_2239);
and U9241 (N_9241,N_49,N_3147);
nor U9242 (N_9242,N_904,N_306);
nand U9243 (N_9243,N_4422,N_3573);
or U9244 (N_9244,N_2622,N_2378);
nand U9245 (N_9245,N_3517,N_4886);
and U9246 (N_9246,N_2645,N_293);
nor U9247 (N_9247,N_2741,N_1049);
nor U9248 (N_9248,N_4084,N_3962);
xor U9249 (N_9249,N_668,N_4104);
and U9250 (N_9250,N_112,N_4781);
and U9251 (N_9251,N_2352,N_1476);
or U9252 (N_9252,N_1245,N_1247);
nand U9253 (N_9253,N_1139,N_4541);
and U9254 (N_9254,N_3428,N_567);
xnor U9255 (N_9255,N_2608,N_1113);
xor U9256 (N_9256,N_3709,N_4321);
and U9257 (N_9257,N_4316,N_4750);
nor U9258 (N_9258,N_1106,N_3488);
nand U9259 (N_9259,N_210,N_2562);
xor U9260 (N_9260,N_2151,N_1975);
nand U9261 (N_9261,N_4112,N_406);
or U9262 (N_9262,N_1971,N_4807);
nor U9263 (N_9263,N_4350,N_3523);
and U9264 (N_9264,N_4356,N_1644);
and U9265 (N_9265,N_4106,N_3870);
and U9266 (N_9266,N_1748,N_9);
or U9267 (N_9267,N_4092,N_766);
nand U9268 (N_9268,N_2776,N_2476);
or U9269 (N_9269,N_4025,N_3803);
nor U9270 (N_9270,N_1151,N_2348);
nand U9271 (N_9271,N_1236,N_3218);
nor U9272 (N_9272,N_1730,N_2765);
or U9273 (N_9273,N_2573,N_488);
and U9274 (N_9274,N_3576,N_1345);
nand U9275 (N_9275,N_174,N_4606);
nand U9276 (N_9276,N_1787,N_107);
xor U9277 (N_9277,N_2823,N_4946);
and U9278 (N_9278,N_932,N_2264);
and U9279 (N_9279,N_3795,N_2068);
and U9280 (N_9280,N_2885,N_1990);
and U9281 (N_9281,N_2643,N_2863);
nor U9282 (N_9282,N_741,N_2394);
xor U9283 (N_9283,N_1231,N_1343);
and U9284 (N_9284,N_4911,N_3157);
nor U9285 (N_9285,N_173,N_4052);
nor U9286 (N_9286,N_1280,N_2208);
or U9287 (N_9287,N_2303,N_2097);
and U9288 (N_9288,N_3433,N_4274);
nor U9289 (N_9289,N_4330,N_236);
nor U9290 (N_9290,N_4343,N_1292);
nor U9291 (N_9291,N_4467,N_3082);
nand U9292 (N_9292,N_1751,N_4894);
or U9293 (N_9293,N_1199,N_3289);
xor U9294 (N_9294,N_2736,N_923);
nor U9295 (N_9295,N_3061,N_3994);
nor U9296 (N_9296,N_4159,N_4739);
nand U9297 (N_9297,N_3959,N_1705);
and U9298 (N_9298,N_4034,N_1135);
nor U9299 (N_9299,N_30,N_2978);
or U9300 (N_9300,N_4895,N_3930);
or U9301 (N_9301,N_4980,N_4390);
xnor U9302 (N_9302,N_4503,N_1658);
and U9303 (N_9303,N_2547,N_929);
nor U9304 (N_9304,N_1164,N_413);
nor U9305 (N_9305,N_4669,N_2344);
nor U9306 (N_9306,N_2676,N_920);
nand U9307 (N_9307,N_2069,N_4720);
nand U9308 (N_9308,N_2211,N_88);
and U9309 (N_9309,N_194,N_2057);
nor U9310 (N_9310,N_2453,N_4428);
or U9311 (N_9311,N_1532,N_4239);
or U9312 (N_9312,N_4597,N_694);
nor U9313 (N_9313,N_848,N_783);
or U9314 (N_9314,N_3291,N_2778);
nor U9315 (N_9315,N_144,N_1936);
or U9316 (N_9316,N_2618,N_3536);
or U9317 (N_9317,N_845,N_2495);
nand U9318 (N_9318,N_3630,N_4453);
nor U9319 (N_9319,N_1106,N_1590);
nand U9320 (N_9320,N_3689,N_643);
and U9321 (N_9321,N_2554,N_352);
nor U9322 (N_9322,N_2357,N_3146);
nor U9323 (N_9323,N_1140,N_349);
and U9324 (N_9324,N_1182,N_4801);
nor U9325 (N_9325,N_3177,N_467);
or U9326 (N_9326,N_346,N_3108);
or U9327 (N_9327,N_3534,N_4447);
nand U9328 (N_9328,N_4605,N_4659);
nand U9329 (N_9329,N_4878,N_1290);
nor U9330 (N_9330,N_4188,N_2459);
nor U9331 (N_9331,N_4555,N_3569);
nor U9332 (N_9332,N_2079,N_490);
nor U9333 (N_9333,N_964,N_1077);
nor U9334 (N_9334,N_1802,N_1838);
and U9335 (N_9335,N_3674,N_4368);
or U9336 (N_9336,N_4510,N_4781);
nor U9337 (N_9337,N_4380,N_4460);
and U9338 (N_9338,N_655,N_2699);
and U9339 (N_9339,N_507,N_2508);
nand U9340 (N_9340,N_618,N_3753);
nor U9341 (N_9341,N_1642,N_3830);
or U9342 (N_9342,N_3560,N_1300);
nor U9343 (N_9343,N_1847,N_488);
or U9344 (N_9344,N_4074,N_2507);
nand U9345 (N_9345,N_4699,N_2785);
or U9346 (N_9346,N_1457,N_2559);
or U9347 (N_9347,N_3204,N_991);
or U9348 (N_9348,N_3735,N_4887);
nand U9349 (N_9349,N_4031,N_3162);
nor U9350 (N_9350,N_3130,N_3537);
xnor U9351 (N_9351,N_1873,N_690);
nor U9352 (N_9352,N_2653,N_789);
nor U9353 (N_9353,N_2206,N_3581);
nand U9354 (N_9354,N_4656,N_3061);
nand U9355 (N_9355,N_4869,N_2205);
or U9356 (N_9356,N_1746,N_180);
nor U9357 (N_9357,N_543,N_746);
nand U9358 (N_9358,N_4349,N_982);
or U9359 (N_9359,N_2388,N_3341);
nor U9360 (N_9360,N_1724,N_2996);
xnor U9361 (N_9361,N_828,N_1367);
nor U9362 (N_9362,N_790,N_1286);
nand U9363 (N_9363,N_1957,N_554);
nand U9364 (N_9364,N_1392,N_1269);
and U9365 (N_9365,N_1507,N_3424);
nand U9366 (N_9366,N_4109,N_52);
and U9367 (N_9367,N_3140,N_4848);
xor U9368 (N_9368,N_1142,N_4590);
nand U9369 (N_9369,N_3958,N_3405);
nor U9370 (N_9370,N_965,N_1545);
nor U9371 (N_9371,N_2113,N_3144);
or U9372 (N_9372,N_2033,N_337);
or U9373 (N_9373,N_1673,N_4916);
and U9374 (N_9374,N_3936,N_3298);
or U9375 (N_9375,N_316,N_2066);
nand U9376 (N_9376,N_207,N_1679);
and U9377 (N_9377,N_1039,N_184);
or U9378 (N_9378,N_4883,N_2615);
and U9379 (N_9379,N_2353,N_1838);
nor U9380 (N_9380,N_1074,N_1063);
and U9381 (N_9381,N_175,N_304);
or U9382 (N_9382,N_2018,N_2914);
and U9383 (N_9383,N_388,N_4506);
nor U9384 (N_9384,N_540,N_838);
nor U9385 (N_9385,N_87,N_2770);
and U9386 (N_9386,N_18,N_747);
or U9387 (N_9387,N_752,N_4760);
nand U9388 (N_9388,N_2064,N_1785);
nand U9389 (N_9389,N_1454,N_1080);
or U9390 (N_9390,N_849,N_1067);
nand U9391 (N_9391,N_1903,N_3797);
and U9392 (N_9392,N_4476,N_1391);
nor U9393 (N_9393,N_3039,N_739);
nand U9394 (N_9394,N_3921,N_4616);
and U9395 (N_9395,N_3252,N_616);
nor U9396 (N_9396,N_4988,N_3819);
or U9397 (N_9397,N_836,N_2208);
and U9398 (N_9398,N_746,N_4134);
nor U9399 (N_9399,N_3884,N_2836);
nand U9400 (N_9400,N_2813,N_2826);
or U9401 (N_9401,N_1890,N_4822);
or U9402 (N_9402,N_3310,N_2754);
and U9403 (N_9403,N_2371,N_4497);
nor U9404 (N_9404,N_1243,N_4129);
or U9405 (N_9405,N_357,N_3789);
or U9406 (N_9406,N_2936,N_3421);
and U9407 (N_9407,N_2941,N_2932);
or U9408 (N_9408,N_1451,N_923);
and U9409 (N_9409,N_1343,N_53);
and U9410 (N_9410,N_4205,N_162);
and U9411 (N_9411,N_221,N_2845);
nor U9412 (N_9412,N_311,N_376);
and U9413 (N_9413,N_4856,N_3362);
nor U9414 (N_9414,N_1321,N_4229);
or U9415 (N_9415,N_3049,N_2268);
nand U9416 (N_9416,N_4372,N_1742);
or U9417 (N_9417,N_3968,N_2931);
and U9418 (N_9418,N_279,N_1991);
and U9419 (N_9419,N_3394,N_4414);
or U9420 (N_9420,N_1160,N_1756);
nand U9421 (N_9421,N_1088,N_3850);
and U9422 (N_9422,N_2494,N_2086);
nor U9423 (N_9423,N_666,N_4164);
or U9424 (N_9424,N_4157,N_2030);
and U9425 (N_9425,N_3351,N_2429);
nor U9426 (N_9426,N_808,N_2594);
and U9427 (N_9427,N_2364,N_396);
and U9428 (N_9428,N_4067,N_3465);
nor U9429 (N_9429,N_1094,N_2234);
or U9430 (N_9430,N_1080,N_2488);
or U9431 (N_9431,N_4586,N_4275);
and U9432 (N_9432,N_2707,N_1406);
or U9433 (N_9433,N_4713,N_1158);
or U9434 (N_9434,N_3918,N_2850);
or U9435 (N_9435,N_831,N_2917);
nand U9436 (N_9436,N_3896,N_4951);
nand U9437 (N_9437,N_2989,N_4651);
or U9438 (N_9438,N_1378,N_871);
nor U9439 (N_9439,N_3926,N_2845);
or U9440 (N_9440,N_134,N_1274);
nor U9441 (N_9441,N_3929,N_4007);
or U9442 (N_9442,N_1337,N_4153);
or U9443 (N_9443,N_534,N_1053);
nand U9444 (N_9444,N_1250,N_2579);
and U9445 (N_9445,N_404,N_393);
nor U9446 (N_9446,N_1742,N_4362);
nor U9447 (N_9447,N_384,N_3262);
nand U9448 (N_9448,N_632,N_490);
nor U9449 (N_9449,N_891,N_3774);
nor U9450 (N_9450,N_2525,N_196);
nand U9451 (N_9451,N_4147,N_1370);
or U9452 (N_9452,N_1306,N_1923);
nor U9453 (N_9453,N_4364,N_797);
and U9454 (N_9454,N_2164,N_2917);
nor U9455 (N_9455,N_3,N_717);
or U9456 (N_9456,N_4020,N_1223);
or U9457 (N_9457,N_1228,N_1555);
xor U9458 (N_9458,N_4261,N_3138);
or U9459 (N_9459,N_2172,N_871);
nor U9460 (N_9460,N_2998,N_3064);
nor U9461 (N_9461,N_1613,N_2353);
nor U9462 (N_9462,N_30,N_4731);
or U9463 (N_9463,N_2464,N_988);
and U9464 (N_9464,N_264,N_2090);
or U9465 (N_9465,N_3407,N_874);
nand U9466 (N_9466,N_3424,N_2888);
nand U9467 (N_9467,N_238,N_1164);
and U9468 (N_9468,N_4404,N_607);
nor U9469 (N_9469,N_551,N_3853);
nor U9470 (N_9470,N_1612,N_3968);
nand U9471 (N_9471,N_2575,N_213);
and U9472 (N_9472,N_723,N_1616);
xnor U9473 (N_9473,N_1587,N_1101);
nand U9474 (N_9474,N_3164,N_635);
nor U9475 (N_9475,N_650,N_2366);
and U9476 (N_9476,N_3325,N_3888);
nor U9477 (N_9477,N_4143,N_3316);
nand U9478 (N_9478,N_1831,N_4326);
nor U9479 (N_9479,N_4372,N_4927);
nand U9480 (N_9480,N_1728,N_1965);
or U9481 (N_9481,N_3179,N_556);
and U9482 (N_9482,N_313,N_3935);
nand U9483 (N_9483,N_2051,N_4463);
nand U9484 (N_9484,N_4020,N_1740);
nand U9485 (N_9485,N_921,N_2463);
nor U9486 (N_9486,N_906,N_2248);
nor U9487 (N_9487,N_4360,N_3603);
nand U9488 (N_9488,N_1074,N_2530);
and U9489 (N_9489,N_4181,N_2696);
nand U9490 (N_9490,N_2155,N_4146);
nor U9491 (N_9491,N_3426,N_4444);
or U9492 (N_9492,N_2122,N_1222);
xor U9493 (N_9493,N_189,N_3538);
nand U9494 (N_9494,N_3213,N_901);
nand U9495 (N_9495,N_4993,N_2806);
and U9496 (N_9496,N_985,N_3409);
or U9497 (N_9497,N_3742,N_1795);
or U9498 (N_9498,N_4975,N_2310);
or U9499 (N_9499,N_1552,N_3933);
or U9500 (N_9500,N_3497,N_273);
nor U9501 (N_9501,N_52,N_2429);
xor U9502 (N_9502,N_1706,N_3386);
and U9503 (N_9503,N_2834,N_3053);
and U9504 (N_9504,N_3379,N_4652);
nor U9505 (N_9505,N_4696,N_1675);
or U9506 (N_9506,N_1801,N_175);
nand U9507 (N_9507,N_2464,N_4265);
xor U9508 (N_9508,N_624,N_100);
nand U9509 (N_9509,N_3783,N_1575);
nor U9510 (N_9510,N_1086,N_2826);
and U9511 (N_9511,N_2384,N_2182);
nor U9512 (N_9512,N_3098,N_2083);
and U9513 (N_9513,N_467,N_4588);
nand U9514 (N_9514,N_3217,N_1860);
or U9515 (N_9515,N_2461,N_3533);
or U9516 (N_9516,N_3724,N_3987);
and U9517 (N_9517,N_1742,N_4066);
and U9518 (N_9518,N_3025,N_2023);
and U9519 (N_9519,N_3053,N_2097);
and U9520 (N_9520,N_3502,N_384);
or U9521 (N_9521,N_4915,N_1687);
or U9522 (N_9522,N_321,N_2030);
or U9523 (N_9523,N_1961,N_3817);
nor U9524 (N_9524,N_2270,N_1086);
nand U9525 (N_9525,N_4842,N_401);
xnor U9526 (N_9526,N_4500,N_3086);
and U9527 (N_9527,N_1523,N_1860);
or U9528 (N_9528,N_409,N_4344);
and U9529 (N_9529,N_4826,N_2703);
nor U9530 (N_9530,N_4190,N_1599);
nor U9531 (N_9531,N_4530,N_3483);
and U9532 (N_9532,N_1382,N_1776);
and U9533 (N_9533,N_2858,N_2310);
nor U9534 (N_9534,N_3323,N_488);
nand U9535 (N_9535,N_440,N_411);
or U9536 (N_9536,N_3906,N_14);
nor U9537 (N_9537,N_4342,N_2723);
and U9538 (N_9538,N_1479,N_277);
nor U9539 (N_9539,N_1955,N_78);
or U9540 (N_9540,N_620,N_4097);
or U9541 (N_9541,N_4502,N_981);
or U9542 (N_9542,N_4437,N_4979);
and U9543 (N_9543,N_2321,N_3694);
xor U9544 (N_9544,N_3786,N_1270);
nor U9545 (N_9545,N_3016,N_2240);
and U9546 (N_9546,N_496,N_2021);
nor U9547 (N_9547,N_3859,N_604);
nand U9548 (N_9548,N_2030,N_1064);
nor U9549 (N_9549,N_2009,N_928);
nand U9550 (N_9550,N_2690,N_783);
xor U9551 (N_9551,N_3188,N_2405);
or U9552 (N_9552,N_1343,N_2196);
and U9553 (N_9553,N_4248,N_3725);
nor U9554 (N_9554,N_3079,N_2442);
or U9555 (N_9555,N_3634,N_2603);
nor U9556 (N_9556,N_1380,N_2100);
and U9557 (N_9557,N_2371,N_4529);
or U9558 (N_9558,N_4365,N_3676);
or U9559 (N_9559,N_523,N_22);
nor U9560 (N_9560,N_29,N_3448);
and U9561 (N_9561,N_3550,N_78);
nor U9562 (N_9562,N_3153,N_1716);
nand U9563 (N_9563,N_4743,N_4699);
nor U9564 (N_9564,N_1522,N_686);
nor U9565 (N_9565,N_1979,N_1085);
nor U9566 (N_9566,N_1393,N_4508);
or U9567 (N_9567,N_4944,N_1919);
or U9568 (N_9568,N_2008,N_1999);
or U9569 (N_9569,N_4410,N_498);
nand U9570 (N_9570,N_92,N_3170);
or U9571 (N_9571,N_450,N_172);
or U9572 (N_9572,N_1896,N_2224);
nor U9573 (N_9573,N_897,N_3087);
nand U9574 (N_9574,N_3009,N_1516);
or U9575 (N_9575,N_4479,N_1845);
nor U9576 (N_9576,N_3816,N_1161);
nand U9577 (N_9577,N_365,N_976);
nand U9578 (N_9578,N_4713,N_4411);
nand U9579 (N_9579,N_2453,N_3070);
nor U9580 (N_9580,N_2369,N_3407);
or U9581 (N_9581,N_3664,N_2969);
and U9582 (N_9582,N_453,N_1104);
or U9583 (N_9583,N_3581,N_234);
xor U9584 (N_9584,N_634,N_4377);
and U9585 (N_9585,N_3869,N_1748);
nand U9586 (N_9586,N_2406,N_4029);
or U9587 (N_9587,N_676,N_2840);
nor U9588 (N_9588,N_979,N_2337);
and U9589 (N_9589,N_3164,N_3963);
nand U9590 (N_9590,N_720,N_173);
nor U9591 (N_9591,N_29,N_933);
or U9592 (N_9592,N_2070,N_3660);
nand U9593 (N_9593,N_3820,N_1050);
xnor U9594 (N_9594,N_1632,N_2153);
and U9595 (N_9595,N_1907,N_3918);
and U9596 (N_9596,N_3661,N_4273);
or U9597 (N_9597,N_413,N_450);
and U9598 (N_9598,N_498,N_2564);
and U9599 (N_9599,N_3649,N_696);
xor U9600 (N_9600,N_1012,N_33);
or U9601 (N_9601,N_2378,N_4366);
and U9602 (N_9602,N_4851,N_4911);
and U9603 (N_9603,N_4965,N_4384);
nor U9604 (N_9604,N_3860,N_786);
and U9605 (N_9605,N_2353,N_3096);
and U9606 (N_9606,N_2469,N_3037);
nor U9607 (N_9607,N_1977,N_4366);
and U9608 (N_9608,N_267,N_4018);
nand U9609 (N_9609,N_4979,N_1593);
and U9610 (N_9610,N_2622,N_1236);
or U9611 (N_9611,N_3188,N_1691);
or U9612 (N_9612,N_4942,N_3092);
or U9613 (N_9613,N_4106,N_2229);
nand U9614 (N_9614,N_4,N_4514);
xnor U9615 (N_9615,N_4793,N_2011);
and U9616 (N_9616,N_1204,N_3585);
and U9617 (N_9617,N_3077,N_4737);
and U9618 (N_9618,N_2591,N_4199);
nor U9619 (N_9619,N_4078,N_970);
and U9620 (N_9620,N_4592,N_573);
xor U9621 (N_9621,N_3870,N_4685);
or U9622 (N_9622,N_918,N_688);
nand U9623 (N_9623,N_3914,N_1503);
nand U9624 (N_9624,N_96,N_3837);
nand U9625 (N_9625,N_1920,N_1108);
nand U9626 (N_9626,N_198,N_1971);
and U9627 (N_9627,N_1747,N_1448);
nor U9628 (N_9628,N_4873,N_1848);
or U9629 (N_9629,N_3382,N_3174);
nor U9630 (N_9630,N_3474,N_1388);
nand U9631 (N_9631,N_2643,N_2731);
or U9632 (N_9632,N_3397,N_1973);
and U9633 (N_9633,N_2419,N_921);
and U9634 (N_9634,N_2905,N_3540);
and U9635 (N_9635,N_1788,N_3070);
nand U9636 (N_9636,N_3523,N_3588);
and U9637 (N_9637,N_2568,N_1417);
nor U9638 (N_9638,N_4114,N_3609);
and U9639 (N_9639,N_2218,N_3805);
nand U9640 (N_9640,N_4557,N_2204);
nor U9641 (N_9641,N_2462,N_3805);
and U9642 (N_9642,N_3769,N_2454);
nor U9643 (N_9643,N_4497,N_2035);
xor U9644 (N_9644,N_3061,N_2959);
and U9645 (N_9645,N_4056,N_3656);
nor U9646 (N_9646,N_13,N_841);
nor U9647 (N_9647,N_1042,N_3116);
xor U9648 (N_9648,N_4677,N_2418);
xnor U9649 (N_9649,N_2444,N_248);
or U9650 (N_9650,N_4548,N_1139);
nor U9651 (N_9651,N_1930,N_148);
or U9652 (N_9652,N_1903,N_3583);
nor U9653 (N_9653,N_2933,N_72);
xnor U9654 (N_9654,N_873,N_3673);
and U9655 (N_9655,N_3628,N_1198);
xor U9656 (N_9656,N_2229,N_299);
nor U9657 (N_9657,N_2030,N_4949);
or U9658 (N_9658,N_659,N_2820);
xor U9659 (N_9659,N_745,N_4637);
nor U9660 (N_9660,N_625,N_3660);
nand U9661 (N_9661,N_3699,N_3412);
nor U9662 (N_9662,N_1443,N_4240);
or U9663 (N_9663,N_2188,N_3861);
nor U9664 (N_9664,N_131,N_2302);
nand U9665 (N_9665,N_4539,N_842);
xnor U9666 (N_9666,N_237,N_3138);
nor U9667 (N_9667,N_2403,N_1283);
xor U9668 (N_9668,N_4689,N_2649);
xnor U9669 (N_9669,N_1857,N_2148);
nand U9670 (N_9670,N_1270,N_2035);
and U9671 (N_9671,N_4798,N_2231);
or U9672 (N_9672,N_4624,N_1856);
nand U9673 (N_9673,N_3762,N_4473);
or U9674 (N_9674,N_3840,N_1845);
or U9675 (N_9675,N_1669,N_2323);
nand U9676 (N_9676,N_887,N_3215);
xnor U9677 (N_9677,N_4250,N_579);
xnor U9678 (N_9678,N_749,N_12);
nor U9679 (N_9679,N_1255,N_2820);
or U9680 (N_9680,N_3667,N_3443);
nand U9681 (N_9681,N_3088,N_120);
or U9682 (N_9682,N_1973,N_2662);
and U9683 (N_9683,N_2169,N_2322);
nand U9684 (N_9684,N_933,N_4060);
or U9685 (N_9685,N_1689,N_169);
or U9686 (N_9686,N_2240,N_3744);
nand U9687 (N_9687,N_1896,N_1232);
and U9688 (N_9688,N_591,N_3417);
and U9689 (N_9689,N_4214,N_4344);
nor U9690 (N_9690,N_1834,N_1611);
and U9691 (N_9691,N_85,N_4414);
or U9692 (N_9692,N_2466,N_2905);
or U9693 (N_9693,N_3506,N_4186);
or U9694 (N_9694,N_4682,N_3231);
and U9695 (N_9695,N_2345,N_3180);
nor U9696 (N_9696,N_3857,N_483);
and U9697 (N_9697,N_4609,N_434);
xor U9698 (N_9698,N_2059,N_1851);
nor U9699 (N_9699,N_4405,N_2361);
or U9700 (N_9700,N_3198,N_1001);
nand U9701 (N_9701,N_1207,N_1536);
or U9702 (N_9702,N_2544,N_3461);
nor U9703 (N_9703,N_2846,N_97);
nor U9704 (N_9704,N_4908,N_4826);
nand U9705 (N_9705,N_107,N_1225);
nor U9706 (N_9706,N_1992,N_940);
or U9707 (N_9707,N_882,N_1704);
and U9708 (N_9708,N_1029,N_1167);
nand U9709 (N_9709,N_4025,N_4003);
or U9710 (N_9710,N_3820,N_2682);
xnor U9711 (N_9711,N_1401,N_1913);
or U9712 (N_9712,N_329,N_3255);
and U9713 (N_9713,N_1064,N_4837);
nand U9714 (N_9714,N_2708,N_2894);
nand U9715 (N_9715,N_3880,N_3661);
nand U9716 (N_9716,N_4611,N_608);
and U9717 (N_9717,N_4501,N_2431);
or U9718 (N_9718,N_1418,N_303);
xnor U9719 (N_9719,N_574,N_4297);
or U9720 (N_9720,N_2011,N_3976);
and U9721 (N_9721,N_2571,N_1919);
nor U9722 (N_9722,N_2614,N_4763);
nor U9723 (N_9723,N_1635,N_4480);
nor U9724 (N_9724,N_2271,N_4998);
nand U9725 (N_9725,N_4003,N_4470);
xnor U9726 (N_9726,N_1513,N_3574);
nand U9727 (N_9727,N_4031,N_1206);
nand U9728 (N_9728,N_2463,N_1520);
and U9729 (N_9729,N_2020,N_1836);
nand U9730 (N_9730,N_507,N_2942);
nand U9731 (N_9731,N_2670,N_1180);
nand U9732 (N_9732,N_1924,N_4317);
and U9733 (N_9733,N_2283,N_3450);
and U9734 (N_9734,N_1536,N_1408);
nor U9735 (N_9735,N_1724,N_786);
nor U9736 (N_9736,N_1656,N_3410);
nand U9737 (N_9737,N_1750,N_2071);
and U9738 (N_9738,N_4664,N_891);
and U9739 (N_9739,N_1587,N_4481);
nand U9740 (N_9740,N_3050,N_1522);
xnor U9741 (N_9741,N_4211,N_3954);
or U9742 (N_9742,N_1334,N_1928);
or U9743 (N_9743,N_1445,N_290);
xor U9744 (N_9744,N_3832,N_986);
xnor U9745 (N_9745,N_3520,N_4014);
xnor U9746 (N_9746,N_1660,N_245);
and U9747 (N_9747,N_3176,N_3989);
xor U9748 (N_9748,N_2902,N_4613);
nand U9749 (N_9749,N_983,N_2632);
nand U9750 (N_9750,N_927,N_4396);
or U9751 (N_9751,N_1984,N_3927);
and U9752 (N_9752,N_897,N_3389);
nor U9753 (N_9753,N_104,N_3787);
and U9754 (N_9754,N_1641,N_2094);
or U9755 (N_9755,N_4705,N_1391);
or U9756 (N_9756,N_4119,N_3823);
or U9757 (N_9757,N_3094,N_2104);
nand U9758 (N_9758,N_1793,N_742);
nand U9759 (N_9759,N_876,N_589);
xnor U9760 (N_9760,N_4709,N_2022);
nand U9761 (N_9761,N_3026,N_2987);
or U9762 (N_9762,N_4881,N_378);
nor U9763 (N_9763,N_3019,N_496);
or U9764 (N_9764,N_2640,N_673);
or U9765 (N_9765,N_1065,N_3558);
or U9766 (N_9766,N_2909,N_4835);
xor U9767 (N_9767,N_2071,N_4507);
nor U9768 (N_9768,N_1728,N_2620);
or U9769 (N_9769,N_4379,N_302);
nor U9770 (N_9770,N_1032,N_1274);
nor U9771 (N_9771,N_139,N_3942);
or U9772 (N_9772,N_1627,N_3080);
and U9773 (N_9773,N_4830,N_2310);
or U9774 (N_9774,N_1675,N_3565);
or U9775 (N_9775,N_2087,N_3730);
or U9776 (N_9776,N_2333,N_2294);
nand U9777 (N_9777,N_4911,N_2947);
nor U9778 (N_9778,N_241,N_3011);
or U9779 (N_9779,N_627,N_836);
nand U9780 (N_9780,N_4933,N_4386);
or U9781 (N_9781,N_2183,N_3620);
nand U9782 (N_9782,N_4279,N_3639);
and U9783 (N_9783,N_2705,N_4738);
nand U9784 (N_9784,N_1619,N_4956);
and U9785 (N_9785,N_4335,N_3457);
nand U9786 (N_9786,N_796,N_2064);
and U9787 (N_9787,N_3167,N_2267);
nor U9788 (N_9788,N_3839,N_756);
and U9789 (N_9789,N_2945,N_1557);
and U9790 (N_9790,N_4274,N_260);
or U9791 (N_9791,N_468,N_1319);
and U9792 (N_9792,N_2882,N_1531);
and U9793 (N_9793,N_3744,N_1423);
and U9794 (N_9794,N_4681,N_885);
nor U9795 (N_9795,N_4566,N_2281);
nand U9796 (N_9796,N_953,N_896);
and U9797 (N_9797,N_1664,N_2060);
or U9798 (N_9798,N_0,N_3348);
nor U9799 (N_9799,N_1270,N_3329);
nor U9800 (N_9800,N_921,N_2519);
or U9801 (N_9801,N_4065,N_748);
nand U9802 (N_9802,N_3440,N_2032);
or U9803 (N_9803,N_3130,N_4854);
or U9804 (N_9804,N_1662,N_350);
and U9805 (N_9805,N_858,N_3855);
nor U9806 (N_9806,N_1254,N_3195);
xnor U9807 (N_9807,N_1798,N_1512);
or U9808 (N_9808,N_2288,N_503);
xor U9809 (N_9809,N_3179,N_1957);
and U9810 (N_9810,N_3560,N_3689);
nand U9811 (N_9811,N_1381,N_596);
and U9812 (N_9812,N_3258,N_2736);
and U9813 (N_9813,N_3605,N_2477);
or U9814 (N_9814,N_4349,N_1467);
nor U9815 (N_9815,N_1339,N_2899);
nor U9816 (N_9816,N_1304,N_4138);
or U9817 (N_9817,N_1753,N_3272);
nor U9818 (N_9818,N_2255,N_4418);
nand U9819 (N_9819,N_4902,N_4070);
nand U9820 (N_9820,N_3804,N_1425);
nand U9821 (N_9821,N_3974,N_3386);
xor U9822 (N_9822,N_506,N_4341);
nor U9823 (N_9823,N_856,N_2912);
and U9824 (N_9824,N_1145,N_4095);
nor U9825 (N_9825,N_1200,N_3770);
nand U9826 (N_9826,N_2928,N_4027);
xnor U9827 (N_9827,N_1140,N_4404);
and U9828 (N_9828,N_3174,N_4988);
and U9829 (N_9829,N_2733,N_355);
and U9830 (N_9830,N_1649,N_688);
and U9831 (N_9831,N_290,N_2301);
nand U9832 (N_9832,N_486,N_2403);
and U9833 (N_9833,N_4421,N_2966);
or U9834 (N_9834,N_2421,N_3017);
or U9835 (N_9835,N_1549,N_4065);
xnor U9836 (N_9836,N_3466,N_936);
nor U9837 (N_9837,N_2630,N_3697);
nor U9838 (N_9838,N_2914,N_1685);
nand U9839 (N_9839,N_4853,N_1381);
nor U9840 (N_9840,N_3037,N_408);
xor U9841 (N_9841,N_1543,N_1373);
and U9842 (N_9842,N_3989,N_2580);
and U9843 (N_9843,N_3557,N_485);
and U9844 (N_9844,N_130,N_2724);
nor U9845 (N_9845,N_3861,N_2487);
nand U9846 (N_9846,N_3105,N_4930);
nand U9847 (N_9847,N_1772,N_584);
or U9848 (N_9848,N_43,N_331);
or U9849 (N_9849,N_4048,N_1483);
or U9850 (N_9850,N_4611,N_1546);
nand U9851 (N_9851,N_4951,N_1538);
nand U9852 (N_9852,N_3932,N_4219);
or U9853 (N_9853,N_2900,N_3626);
nand U9854 (N_9854,N_2324,N_3581);
or U9855 (N_9855,N_4400,N_3321);
nand U9856 (N_9856,N_4347,N_3204);
xor U9857 (N_9857,N_2504,N_2053);
nand U9858 (N_9858,N_3822,N_1650);
nand U9859 (N_9859,N_366,N_1772);
and U9860 (N_9860,N_1706,N_4927);
nand U9861 (N_9861,N_1780,N_3538);
nor U9862 (N_9862,N_188,N_1031);
nand U9863 (N_9863,N_2597,N_507);
nor U9864 (N_9864,N_4225,N_2391);
nor U9865 (N_9865,N_3590,N_1895);
or U9866 (N_9866,N_192,N_3609);
nand U9867 (N_9867,N_4540,N_3445);
nand U9868 (N_9868,N_328,N_1312);
nor U9869 (N_9869,N_1849,N_4674);
nor U9870 (N_9870,N_4743,N_970);
or U9871 (N_9871,N_544,N_1678);
nor U9872 (N_9872,N_1785,N_1028);
and U9873 (N_9873,N_1623,N_126);
nand U9874 (N_9874,N_4323,N_2218);
nand U9875 (N_9875,N_4651,N_3944);
or U9876 (N_9876,N_2990,N_787);
and U9877 (N_9877,N_83,N_3650);
and U9878 (N_9878,N_4090,N_1846);
nand U9879 (N_9879,N_3788,N_4369);
nand U9880 (N_9880,N_1063,N_50);
xnor U9881 (N_9881,N_1026,N_2972);
xor U9882 (N_9882,N_326,N_148);
nor U9883 (N_9883,N_4947,N_2207);
or U9884 (N_9884,N_3638,N_2838);
or U9885 (N_9885,N_2561,N_590);
nand U9886 (N_9886,N_3758,N_3293);
xnor U9887 (N_9887,N_3201,N_2332);
nor U9888 (N_9888,N_2788,N_2102);
nor U9889 (N_9889,N_3075,N_576);
and U9890 (N_9890,N_619,N_380);
nor U9891 (N_9891,N_4621,N_1317);
nor U9892 (N_9892,N_3697,N_4258);
and U9893 (N_9893,N_4037,N_4106);
nand U9894 (N_9894,N_4106,N_287);
nor U9895 (N_9895,N_4864,N_353);
xor U9896 (N_9896,N_298,N_1723);
nor U9897 (N_9897,N_3943,N_1678);
and U9898 (N_9898,N_4599,N_1647);
nand U9899 (N_9899,N_3545,N_1136);
nand U9900 (N_9900,N_1220,N_4469);
or U9901 (N_9901,N_4196,N_1394);
nand U9902 (N_9902,N_1746,N_2618);
nor U9903 (N_9903,N_190,N_131);
nor U9904 (N_9904,N_951,N_1022);
nand U9905 (N_9905,N_2653,N_4161);
xor U9906 (N_9906,N_3073,N_35);
nor U9907 (N_9907,N_1165,N_2462);
and U9908 (N_9908,N_1304,N_4133);
nor U9909 (N_9909,N_4776,N_4852);
or U9910 (N_9910,N_2086,N_2138);
and U9911 (N_9911,N_2109,N_1558);
nand U9912 (N_9912,N_2199,N_3878);
or U9913 (N_9913,N_4279,N_2443);
xnor U9914 (N_9914,N_4339,N_2657);
nand U9915 (N_9915,N_3638,N_4732);
or U9916 (N_9916,N_2809,N_3570);
and U9917 (N_9917,N_4498,N_3745);
nor U9918 (N_9918,N_3696,N_4862);
nand U9919 (N_9919,N_1289,N_2636);
nand U9920 (N_9920,N_1131,N_4660);
nand U9921 (N_9921,N_1120,N_1471);
nand U9922 (N_9922,N_2847,N_1447);
or U9923 (N_9923,N_3773,N_1439);
or U9924 (N_9924,N_4346,N_279);
nand U9925 (N_9925,N_4887,N_808);
nand U9926 (N_9926,N_4491,N_4127);
nor U9927 (N_9927,N_2924,N_3782);
and U9928 (N_9928,N_1764,N_4144);
and U9929 (N_9929,N_3626,N_557);
or U9930 (N_9930,N_4627,N_3551);
nor U9931 (N_9931,N_2053,N_631);
nor U9932 (N_9932,N_695,N_2431);
and U9933 (N_9933,N_3379,N_3802);
or U9934 (N_9934,N_202,N_2135);
nor U9935 (N_9935,N_1205,N_3291);
and U9936 (N_9936,N_3503,N_789);
nand U9937 (N_9937,N_1682,N_3123);
xnor U9938 (N_9938,N_4058,N_386);
and U9939 (N_9939,N_2741,N_2738);
nand U9940 (N_9940,N_696,N_455);
or U9941 (N_9941,N_3859,N_4741);
and U9942 (N_9942,N_215,N_1727);
xnor U9943 (N_9943,N_4864,N_2115);
xor U9944 (N_9944,N_3068,N_1990);
nand U9945 (N_9945,N_2177,N_4254);
or U9946 (N_9946,N_4498,N_1829);
xnor U9947 (N_9947,N_4537,N_3956);
nor U9948 (N_9948,N_456,N_1665);
and U9949 (N_9949,N_2999,N_4292);
nor U9950 (N_9950,N_194,N_3933);
xor U9951 (N_9951,N_3226,N_4758);
and U9952 (N_9952,N_1393,N_3073);
and U9953 (N_9953,N_1673,N_1072);
xor U9954 (N_9954,N_3161,N_925);
or U9955 (N_9955,N_3512,N_2295);
nand U9956 (N_9956,N_1267,N_2980);
nand U9957 (N_9957,N_441,N_3582);
and U9958 (N_9958,N_3631,N_4480);
nand U9959 (N_9959,N_716,N_3413);
xnor U9960 (N_9960,N_971,N_3554);
nor U9961 (N_9961,N_3367,N_1507);
or U9962 (N_9962,N_1742,N_563);
or U9963 (N_9963,N_3182,N_4396);
xnor U9964 (N_9964,N_4416,N_4202);
or U9965 (N_9965,N_3372,N_328);
or U9966 (N_9966,N_4364,N_1937);
and U9967 (N_9967,N_2997,N_1246);
and U9968 (N_9968,N_2422,N_1461);
nor U9969 (N_9969,N_4383,N_513);
and U9970 (N_9970,N_4242,N_3632);
nand U9971 (N_9971,N_3816,N_29);
or U9972 (N_9972,N_1355,N_2289);
or U9973 (N_9973,N_3257,N_2238);
nand U9974 (N_9974,N_308,N_1185);
nand U9975 (N_9975,N_3273,N_4621);
and U9976 (N_9976,N_1699,N_3244);
xor U9977 (N_9977,N_4920,N_1789);
and U9978 (N_9978,N_1789,N_4335);
xor U9979 (N_9979,N_635,N_1450);
or U9980 (N_9980,N_3041,N_4252);
and U9981 (N_9981,N_16,N_781);
xnor U9982 (N_9982,N_102,N_1679);
or U9983 (N_9983,N_3963,N_2687);
and U9984 (N_9984,N_428,N_1882);
and U9985 (N_9985,N_2095,N_145);
nand U9986 (N_9986,N_2297,N_1561);
and U9987 (N_9987,N_4872,N_908);
and U9988 (N_9988,N_4492,N_2006);
nand U9989 (N_9989,N_539,N_159);
nor U9990 (N_9990,N_3740,N_98);
nand U9991 (N_9991,N_2257,N_1964);
and U9992 (N_9992,N_4008,N_1861);
nor U9993 (N_9993,N_174,N_2455);
nor U9994 (N_9994,N_3534,N_244);
nor U9995 (N_9995,N_4227,N_3171);
or U9996 (N_9996,N_3275,N_4195);
and U9997 (N_9997,N_4121,N_477);
nor U9998 (N_9998,N_3625,N_77);
nor U9999 (N_9999,N_4060,N_295);
nand U10000 (N_10000,N_5633,N_7609);
nand U10001 (N_10001,N_7547,N_9746);
and U10002 (N_10002,N_6596,N_9900);
nor U10003 (N_10003,N_5636,N_6945);
nand U10004 (N_10004,N_6850,N_8247);
nand U10005 (N_10005,N_7523,N_7568);
nand U10006 (N_10006,N_8824,N_7915);
nand U10007 (N_10007,N_9224,N_9338);
or U10008 (N_10008,N_7938,N_9182);
nand U10009 (N_10009,N_5419,N_7322);
nor U10010 (N_10010,N_5192,N_8384);
or U10011 (N_10011,N_9892,N_6910);
nand U10012 (N_10012,N_8147,N_7425);
or U10013 (N_10013,N_6592,N_7186);
nand U10014 (N_10014,N_9492,N_7646);
and U10015 (N_10015,N_7517,N_7197);
nand U10016 (N_10016,N_5058,N_9260);
and U10017 (N_10017,N_5473,N_6389);
and U10018 (N_10018,N_8726,N_5816);
and U10019 (N_10019,N_6434,N_5513);
and U10020 (N_10020,N_7670,N_9793);
and U10021 (N_10021,N_5977,N_9572);
and U10022 (N_10022,N_9763,N_9841);
xor U10023 (N_10023,N_6301,N_7126);
and U10024 (N_10024,N_6009,N_8815);
or U10025 (N_10025,N_9490,N_6161);
and U10026 (N_10026,N_9945,N_6673);
nor U10027 (N_10027,N_7434,N_8919);
or U10028 (N_10028,N_8684,N_9227);
or U10029 (N_10029,N_5908,N_8124);
and U10030 (N_10030,N_5549,N_6285);
nand U10031 (N_10031,N_8568,N_8050);
nand U10032 (N_10032,N_8282,N_7628);
nand U10033 (N_10033,N_6004,N_9919);
nor U10034 (N_10034,N_9167,N_6267);
and U10035 (N_10035,N_8425,N_7157);
xor U10036 (N_10036,N_8757,N_6474);
and U10037 (N_10037,N_5729,N_6560);
or U10038 (N_10038,N_7129,N_5857);
nor U10039 (N_10039,N_9136,N_6635);
nor U10040 (N_10040,N_9020,N_6441);
nor U10041 (N_10041,N_5066,N_7992);
or U10042 (N_10042,N_8764,N_6737);
and U10043 (N_10043,N_6594,N_7785);
nor U10044 (N_10044,N_7716,N_5631);
or U10045 (N_10045,N_9935,N_9842);
nand U10046 (N_10046,N_6143,N_7767);
nand U10047 (N_10047,N_9201,N_6032);
or U10048 (N_10048,N_5936,N_9160);
and U10049 (N_10049,N_8920,N_8604);
nor U10050 (N_10050,N_8819,N_9152);
nor U10051 (N_10051,N_6805,N_9869);
xor U10052 (N_10052,N_5585,N_6196);
xnor U10053 (N_10053,N_7748,N_7557);
or U10054 (N_10054,N_5276,N_6528);
or U10055 (N_10055,N_8867,N_7514);
nor U10056 (N_10056,N_7274,N_5503);
or U10057 (N_10057,N_9520,N_8771);
or U10058 (N_10058,N_7688,N_6972);
nor U10059 (N_10059,N_6199,N_8118);
xor U10060 (N_10060,N_9239,N_6062);
or U10061 (N_10061,N_9649,N_7311);
nor U10062 (N_10062,N_9506,N_8523);
nor U10063 (N_10063,N_5806,N_6706);
nand U10064 (N_10064,N_5042,N_8422);
xnor U10065 (N_10065,N_6549,N_8679);
nor U10066 (N_10066,N_6626,N_6776);
xor U10067 (N_10067,N_9665,N_7980);
nand U10068 (N_10068,N_5368,N_6869);
nand U10069 (N_10069,N_6558,N_9786);
or U10070 (N_10070,N_9782,N_7765);
and U10071 (N_10071,N_7860,N_7820);
nand U10072 (N_10072,N_6812,N_8090);
nand U10073 (N_10073,N_5254,N_7367);
and U10074 (N_10074,N_9186,N_9871);
xnor U10075 (N_10075,N_5367,N_6977);
nand U10076 (N_10076,N_7313,N_8791);
and U10077 (N_10077,N_6343,N_5040);
nor U10078 (N_10078,N_6992,N_5380);
nor U10079 (N_10079,N_8650,N_5583);
or U10080 (N_10080,N_9736,N_8811);
or U10081 (N_10081,N_8250,N_8715);
nor U10082 (N_10082,N_9192,N_8735);
nor U10083 (N_10083,N_7028,N_8538);
nor U10084 (N_10084,N_5502,N_5379);
xnor U10085 (N_10085,N_6183,N_9659);
and U10086 (N_10086,N_6382,N_6197);
and U10087 (N_10087,N_8439,N_8777);
and U10088 (N_10088,N_7083,N_6215);
nor U10089 (N_10089,N_9911,N_5768);
nor U10090 (N_10090,N_9585,N_6356);
or U10091 (N_10091,N_9255,N_8915);
nand U10092 (N_10092,N_8412,N_6732);
or U10093 (N_10093,N_9840,N_8891);
or U10094 (N_10094,N_8693,N_9593);
nor U10095 (N_10095,N_7303,N_7435);
nand U10096 (N_10096,N_5798,N_7344);
xor U10097 (N_10097,N_7436,N_8946);
and U10098 (N_10098,N_6958,N_7082);
nand U10099 (N_10099,N_6281,N_9323);
nor U10100 (N_10100,N_7396,N_9683);
and U10101 (N_10101,N_5797,N_5378);
or U10102 (N_10102,N_5021,N_5597);
nor U10103 (N_10103,N_8302,N_9985);
nor U10104 (N_10104,N_8228,N_7105);
and U10105 (N_10105,N_7775,N_5870);
nand U10106 (N_10106,N_9744,N_8647);
or U10107 (N_10107,N_5125,N_5226);
and U10108 (N_10108,N_9729,N_7706);
nand U10109 (N_10109,N_8851,N_9609);
or U10110 (N_10110,N_5693,N_5669);
xor U10111 (N_10111,N_8541,N_7232);
nand U10112 (N_10112,N_6785,N_5846);
and U10113 (N_10113,N_9624,N_7960);
or U10114 (N_10114,N_5655,N_5975);
nor U10115 (N_10115,N_7247,N_5123);
nor U10116 (N_10116,N_5582,N_7546);
xnor U10117 (N_10117,N_5707,N_9371);
or U10118 (N_10118,N_7725,N_9463);
or U10119 (N_10119,N_5682,N_8685);
and U10120 (N_10120,N_9602,N_9413);
xor U10121 (N_10121,N_5619,N_8185);
nand U10122 (N_10122,N_7442,N_8544);
and U10123 (N_10123,N_8455,N_8584);
and U10124 (N_10124,N_9159,N_6472);
nand U10125 (N_10125,N_6276,N_5894);
xnor U10126 (N_10126,N_8033,N_9843);
xnor U10127 (N_10127,N_5350,N_9686);
or U10128 (N_10128,N_6676,N_7164);
nor U10129 (N_10129,N_6541,N_6533);
nand U10130 (N_10130,N_5081,N_8136);
xnor U10131 (N_10131,N_8183,N_8786);
or U10132 (N_10132,N_6550,N_9180);
and U10133 (N_10133,N_7168,N_5759);
nand U10134 (N_10134,N_5364,N_6035);
nand U10135 (N_10135,N_8769,N_7993);
nand U10136 (N_10136,N_7520,N_5712);
or U10137 (N_10137,N_7804,N_7294);
and U10138 (N_10138,N_9590,N_9105);
nand U10139 (N_10139,N_5777,N_9493);
and U10140 (N_10140,N_5931,N_5644);
nand U10141 (N_10141,N_7707,N_6045);
or U10142 (N_10142,N_7862,N_8535);
xnor U10143 (N_10143,N_7299,N_8525);
nand U10144 (N_10144,N_9670,N_6361);
or U10145 (N_10145,N_7064,N_8901);
and U10146 (N_10146,N_7250,N_7985);
nand U10147 (N_10147,N_6930,N_9329);
nor U10148 (N_10148,N_6054,N_9417);
or U10149 (N_10149,N_8407,N_8960);
nand U10150 (N_10150,N_9934,N_5043);
nand U10151 (N_10151,N_6693,N_7917);
and U10152 (N_10152,N_5608,N_5264);
nand U10153 (N_10153,N_5457,N_6109);
nand U10154 (N_10154,N_6037,N_7438);
and U10155 (N_10155,N_7167,N_6688);
and U10156 (N_10156,N_9115,N_7477);
nor U10157 (N_10157,N_8334,N_7638);
xor U10158 (N_10158,N_8035,N_8415);
xor U10159 (N_10159,N_8609,N_8507);
and U10160 (N_10160,N_8103,N_6520);
nor U10161 (N_10161,N_8567,N_6671);
or U10162 (N_10162,N_6367,N_5389);
nor U10163 (N_10163,N_6999,N_5903);
and U10164 (N_10164,N_8619,N_5735);
nor U10165 (N_10165,N_5382,N_7682);
nor U10166 (N_10166,N_9570,N_5191);
xor U10167 (N_10167,N_7280,N_6717);
or U10168 (N_10168,N_5520,N_9545);
and U10169 (N_10169,N_7615,N_6911);
xnor U10170 (N_10170,N_5454,N_8238);
nor U10171 (N_10171,N_7097,N_6544);
and U10172 (N_10172,N_9563,N_5667);
nor U10173 (N_10173,N_5885,N_9281);
nor U10174 (N_10174,N_6595,N_7658);
nand U10175 (N_10175,N_7850,N_7673);
xnor U10176 (N_10176,N_6213,N_9719);
or U10177 (N_10177,N_9519,N_6255);
and U10178 (N_10178,N_9090,N_7573);
nor U10179 (N_10179,N_8040,N_5994);
nand U10180 (N_10180,N_8747,N_8374);
and U10181 (N_10181,N_8266,N_6324);
or U10182 (N_10182,N_8338,N_7950);
nand U10183 (N_10183,N_5688,N_8408);
nor U10184 (N_10184,N_9203,N_6208);
and U10185 (N_10185,N_9794,N_5565);
and U10186 (N_10186,N_8830,N_7269);
xnor U10187 (N_10187,N_8220,N_6535);
nor U10188 (N_10188,N_8027,N_8128);
nand U10189 (N_10189,N_9132,N_6269);
or U10190 (N_10190,N_9808,N_5322);
and U10191 (N_10191,N_8972,N_8102);
nor U10192 (N_10192,N_7637,N_5055);
xnor U10193 (N_10193,N_7249,N_5801);
nand U10194 (N_10194,N_8270,N_7233);
or U10195 (N_10195,N_7404,N_9314);
nand U10196 (N_10196,N_7761,N_7360);
nand U10197 (N_10197,N_9299,N_7034);
or U10198 (N_10198,N_5696,N_7086);
nor U10199 (N_10199,N_8037,N_7101);
and U10200 (N_10200,N_7751,N_6099);
nand U10201 (N_10201,N_9393,N_9799);
and U10202 (N_10202,N_5165,N_9282);
and U10203 (N_10203,N_6942,N_8914);
nor U10204 (N_10204,N_7224,N_5620);
nor U10205 (N_10205,N_6968,N_6657);
and U10206 (N_10206,N_9163,N_9824);
and U10207 (N_10207,N_5629,N_9515);
or U10208 (N_10208,N_8468,N_9213);
nor U10209 (N_10209,N_5711,N_9185);
and U10210 (N_10210,N_9967,N_7752);
nor U10211 (N_10211,N_8341,N_5321);
nand U10212 (N_10212,N_8293,N_8717);
or U10213 (N_10213,N_7834,N_8746);
xor U10214 (N_10214,N_6725,N_9994);
or U10215 (N_10215,N_7887,N_8838);
nor U10216 (N_10216,N_8962,N_9327);
and U10217 (N_10217,N_5157,N_5762);
and U10218 (N_10218,N_8004,N_7339);
and U10219 (N_10219,N_6493,N_9081);
xnor U10220 (N_10220,N_8913,N_8518);
xnor U10221 (N_10221,N_6959,N_5240);
or U10222 (N_10222,N_6397,N_6905);
nor U10223 (N_10223,N_6616,N_9689);
or U10224 (N_10224,N_5106,N_9938);
nor U10225 (N_10225,N_7465,N_9025);
nand U10226 (N_10226,N_5437,N_7629);
nor U10227 (N_10227,N_7192,N_8804);
nor U10228 (N_10228,N_7553,N_9846);
and U10229 (N_10229,N_9425,N_8024);
or U10230 (N_10230,N_5463,N_8194);
nor U10231 (N_10231,N_6814,N_7512);
xnor U10232 (N_10232,N_7920,N_6902);
xnor U10233 (N_10233,N_6753,N_5934);
nand U10234 (N_10234,N_5329,N_5199);
nand U10235 (N_10235,N_9755,N_7596);
nor U10236 (N_10236,N_9031,N_5630);
nor U10237 (N_10237,N_9370,N_6490);
and U10238 (N_10238,N_6606,N_9447);
nand U10239 (N_10239,N_6678,N_7945);
nor U10240 (N_10240,N_9284,N_9028);
or U10241 (N_10241,N_9923,N_9962);
nor U10242 (N_10242,N_6920,N_8506);
and U10243 (N_10243,N_5691,N_7409);
and U10244 (N_10244,N_5131,N_5887);
nand U10245 (N_10245,N_8259,N_5578);
nor U10246 (N_10246,N_9863,N_5646);
and U10247 (N_10247,N_6100,N_8780);
nor U10248 (N_10248,N_6387,N_8706);
xnor U10249 (N_10249,N_8158,N_6980);
nand U10250 (N_10250,N_5536,N_6284);
nand U10251 (N_10251,N_7014,N_8431);
and U10252 (N_10252,N_8470,N_8770);
xnor U10253 (N_10253,N_9331,N_7015);
nand U10254 (N_10254,N_8104,N_9470);
xor U10255 (N_10255,N_5219,N_6427);
nand U10256 (N_10256,N_9150,N_7555);
nor U10257 (N_10257,N_8042,N_9672);
nor U10258 (N_10258,N_7237,N_6921);
or U10259 (N_10259,N_7933,N_5738);
nor U10260 (N_10260,N_6426,N_6574);
or U10261 (N_10261,N_8774,N_5283);
nand U10262 (N_10262,N_8078,N_5054);
xnor U10263 (N_10263,N_5401,N_9802);
nand U10264 (N_10264,N_7412,N_8475);
xor U10265 (N_10265,N_7229,N_5640);
nand U10266 (N_10266,N_9956,N_5727);
and U10267 (N_10267,N_5788,N_9355);
nand U10268 (N_10268,N_7213,N_9748);
and U10269 (N_10269,N_5957,N_8421);
or U10270 (N_10270,N_7439,N_8833);
nand U10271 (N_10271,N_7782,N_8643);
or U10272 (N_10272,N_9170,N_6797);
and U10273 (N_10273,N_5493,N_9086);
and U10274 (N_10274,N_7732,N_5360);
and U10275 (N_10275,N_6642,N_6615);
or U10276 (N_10276,N_6080,N_7784);
and U10277 (N_10277,N_7591,N_6176);
and U10278 (N_10278,N_9715,N_9523);
and U10279 (N_10279,N_7709,N_6365);
and U10280 (N_10280,N_9703,N_7899);
xor U10281 (N_10281,N_7429,N_5399);
and U10282 (N_10282,N_5002,N_7398);
and U10283 (N_10283,N_5197,N_8054);
nor U10284 (N_10284,N_8386,N_7332);
or U10285 (N_10285,N_9998,N_7444);
or U10286 (N_10286,N_7925,N_6844);
or U10287 (N_10287,N_5900,N_9975);
nand U10288 (N_10288,N_9830,N_5819);
nand U10289 (N_10289,N_9676,N_6128);
nand U10290 (N_10290,N_9701,N_9884);
nand U10291 (N_10291,N_6150,N_7558);
and U10292 (N_10292,N_5815,N_8285);
and U10293 (N_10293,N_6271,N_8836);
nor U10294 (N_10294,N_5796,N_6572);
nand U10295 (N_10295,N_5188,N_6491);
or U10296 (N_10296,N_5449,N_5769);
nand U10297 (N_10297,N_5476,N_9087);
nor U10298 (N_10298,N_5882,N_7457);
or U10299 (N_10299,N_5821,N_6492);
nand U10300 (N_10300,N_9639,N_5172);
and U10301 (N_10301,N_9601,N_5892);
xnor U10302 (N_10302,N_6457,N_7330);
and U10303 (N_10303,N_5731,N_5627);
nand U10304 (N_10304,N_8283,N_9548);
nand U10305 (N_10305,N_8566,N_5778);
nor U10306 (N_10306,N_7946,N_7541);
nand U10307 (N_10307,N_8474,N_7117);
nor U10308 (N_10308,N_7759,N_6392);
xnor U10309 (N_10309,N_9635,N_5460);
nor U10310 (N_10310,N_8986,N_6107);
and U10311 (N_10311,N_7348,N_7453);
xor U10312 (N_10312,N_6681,N_6901);
and U10313 (N_10313,N_5924,N_7421);
nand U10314 (N_10314,N_8980,N_9457);
nor U10315 (N_10315,N_6826,N_9142);
and U10316 (N_10316,N_9288,N_5345);
nand U10317 (N_10317,N_5490,N_9754);
nor U10318 (N_10318,N_5407,N_9677);
xnor U10319 (N_10319,N_6880,N_6458);
nand U10320 (N_10320,N_6257,N_8835);
xnor U10321 (N_10321,N_7800,N_6647);
nor U10322 (N_10322,N_9172,N_9146);
and U10323 (N_10323,N_9606,N_7238);
nand U10324 (N_10324,N_8448,N_8072);
or U10325 (N_10325,N_5875,N_7495);
and U10326 (N_10326,N_9997,N_9818);
nand U10327 (N_10327,N_6971,N_8443);
nand U10328 (N_10328,N_8359,N_6345);
nand U10329 (N_10329,N_9075,N_7900);
nor U10330 (N_10330,N_7809,N_7908);
and U10331 (N_10331,N_5461,N_7802);
nand U10332 (N_10332,N_9138,N_8089);
or U10333 (N_10333,N_9711,N_5852);
xor U10334 (N_10334,N_6141,N_7559);
nand U10335 (N_10335,N_6652,N_8973);
and U10336 (N_10336,N_9610,N_6848);
nor U10337 (N_10337,N_6772,N_6148);
and U10338 (N_10338,N_7494,N_9249);
nand U10339 (N_10339,N_7108,N_9247);
xor U10340 (N_10340,N_9315,N_8383);
or U10341 (N_10341,N_8932,N_7058);
and U10342 (N_10342,N_9758,N_8736);
and U10343 (N_10343,N_8827,N_7585);
and U10344 (N_10344,N_8893,N_6242);
and U10345 (N_10345,N_8536,N_9381);
xor U10346 (N_10346,N_5466,N_5413);
xor U10347 (N_10347,N_6154,N_9801);
or U10348 (N_10348,N_8364,N_5039);
nand U10349 (N_10349,N_5668,N_6130);
or U10350 (N_10350,N_7216,N_9021);
and U10351 (N_10351,N_8257,N_9403);
nand U10352 (N_10352,N_7198,N_6299);
and U10353 (N_10353,N_5073,N_9243);
and U10354 (N_10354,N_8694,N_5530);
nor U10355 (N_10355,N_7866,N_9819);
nor U10356 (N_10356,N_7605,N_6125);
or U10357 (N_10357,N_5726,N_6542);
or U10358 (N_10358,N_9716,N_6579);
or U10359 (N_10359,N_7895,N_9456);
xnor U10360 (N_10360,N_6039,N_5860);
nand U10361 (N_10361,N_9891,N_5167);
nand U10362 (N_10362,N_5372,N_5077);
nor U10363 (N_10363,N_5293,N_8180);
nor U10364 (N_10364,N_5514,N_8157);
and U10365 (N_10365,N_9278,N_7867);
nor U10366 (N_10366,N_8292,N_6714);
nand U10367 (N_10367,N_6879,N_8320);
nand U10368 (N_10368,N_6769,N_6863);
and U10369 (N_10369,N_8298,N_7273);
or U10370 (N_10370,N_5333,N_6584);
nand U10371 (N_10371,N_5772,N_6747);
and U10372 (N_10372,N_9580,N_7050);
nand U10373 (N_10373,N_8351,N_7600);
nor U10374 (N_10374,N_5375,N_6620);
nor U10375 (N_10375,N_7454,N_6842);
and U10376 (N_10376,N_5132,N_7369);
nor U10377 (N_10377,N_7272,N_8435);
or U10378 (N_10378,N_7528,N_6318);
xor U10379 (N_10379,N_9931,N_6118);
xnor U10380 (N_10380,N_7057,N_6656);
xnor U10381 (N_10381,N_5112,N_7692);
nor U10382 (N_10382,N_6177,N_8006);
nor U10383 (N_10383,N_7031,N_6899);
or U10384 (N_10384,N_8930,N_9272);
xnor U10385 (N_10385,N_9310,N_7290);
nor U10386 (N_10386,N_6277,N_9294);
nor U10387 (N_10387,N_8713,N_6494);
and U10388 (N_10388,N_8343,N_9140);
nor U10389 (N_10389,N_8989,N_6881);
and U10390 (N_10390,N_8303,N_8308);
or U10391 (N_10391,N_8918,N_9981);
or U10392 (N_10392,N_7019,N_7723);
nand U10393 (N_10393,N_8816,N_9398);
or U10394 (N_10394,N_9768,N_5196);
and U10395 (N_10395,N_8012,N_6425);
and U10396 (N_10396,N_8842,N_7305);
and U10397 (N_10397,N_7407,N_8545);
or U10398 (N_10398,N_8553,N_9194);
nor U10399 (N_10399,N_5573,N_9268);
and U10400 (N_10400,N_6133,N_7210);
and U10401 (N_10401,N_5932,N_8317);
xnor U10402 (N_10402,N_7262,N_7861);
nor U10403 (N_10403,N_9231,N_7947);
nand U10404 (N_10404,N_5678,N_9321);
or U10405 (N_10405,N_6888,N_7169);
nand U10406 (N_10406,N_6697,N_6847);
or U10407 (N_10407,N_9207,N_8683);
or U10408 (N_10408,N_5153,N_9861);
xor U10409 (N_10409,N_5517,N_5044);
or U10410 (N_10410,N_8822,N_6226);
and U10411 (N_10411,N_5059,N_8192);
or U10412 (N_10412,N_8911,N_8190);
nand U10413 (N_10413,N_7118,N_5786);
or U10414 (N_10414,N_7479,N_6687);
xnor U10415 (N_10415,N_6212,N_5940);
and U10416 (N_10416,N_5773,N_7486);
or U10417 (N_10417,N_8592,N_6916);
and U10418 (N_10418,N_8875,N_5397);
nand U10419 (N_10419,N_9277,N_5862);
and U10420 (N_10420,N_9353,N_5969);
nand U10421 (N_10421,N_7973,N_5465);
nand U10422 (N_10422,N_8406,N_8401);
nand U10423 (N_10423,N_5866,N_6023);
or U10424 (N_10424,N_5858,N_8275);
or U10425 (N_10425,N_8597,N_5434);
and U10426 (N_10426,N_6084,N_7854);
and U10427 (N_10427,N_5947,N_5259);
nand U10428 (N_10428,N_9502,N_6286);
xor U10429 (N_10429,N_5019,N_8971);
nand U10430 (N_10430,N_8278,N_9219);
or U10431 (N_10431,N_8079,N_6346);
nor U10432 (N_10432,N_9798,N_8928);
and U10433 (N_10433,N_6588,N_9559);
or U10434 (N_10434,N_9054,N_5291);
xnor U10435 (N_10435,N_7987,N_9472);
and U10436 (N_10436,N_9106,N_9034);
nor U10437 (N_10437,N_5448,N_6781);
nand U10438 (N_10438,N_7951,N_6857);
and U10439 (N_10439,N_6347,N_8397);
nor U10440 (N_10440,N_8887,N_8982);
nor U10441 (N_10441,N_7134,N_6895);
or U10442 (N_10442,N_8227,N_8909);
xor U10443 (N_10443,N_6946,N_9474);
or U10444 (N_10444,N_6344,N_8339);
and U10445 (N_10445,N_5151,N_8086);
nor U10446 (N_10446,N_8755,N_6264);
nor U10447 (N_10447,N_7368,N_9805);
nor U10448 (N_10448,N_8613,N_6378);
nand U10449 (N_10449,N_9209,N_9103);
and U10450 (N_10450,N_6309,N_6931);
or U10451 (N_10451,N_5552,N_8896);
xor U10452 (N_10452,N_9354,N_6654);
and U10453 (N_10453,N_8625,N_6385);
and U10454 (N_10454,N_9694,N_7515);
nand U10455 (N_10455,N_8127,N_6225);
and U10456 (N_10456,N_7092,N_8105);
or U10457 (N_10457,N_8016,N_9762);
or U10458 (N_10458,N_8554,N_6423);
nor U10459 (N_10459,N_6679,N_6178);
or U10460 (N_10460,N_6698,N_5704);
or U10461 (N_10461,N_9365,N_5498);
and U10462 (N_10462,N_8612,N_6906);
nor U10463 (N_10463,N_7848,N_5596);
xor U10464 (N_10464,N_7783,N_7584);
nor U10465 (N_10465,N_8623,N_5046);
nor U10466 (N_10466,N_7631,N_9014);
xor U10467 (N_10467,N_8288,N_9814);
or U10468 (N_10468,N_5232,N_6582);
nor U10469 (N_10469,N_5544,N_8603);
nor U10470 (N_10470,N_8454,N_7753);
nor U10471 (N_10471,N_7024,N_7141);
xnor U10472 (N_10472,N_9179,N_9048);
nand U10473 (N_10473,N_8274,N_6867);
nor U10474 (N_10474,N_6988,N_5236);
nor U10475 (N_10475,N_6686,N_9684);
nor U10476 (N_10476,N_9778,N_9378);
nor U10477 (N_10477,N_8219,N_5351);
nor U10478 (N_10478,N_7567,N_9018);
nor U10479 (N_10479,N_8120,N_8528);
or U10480 (N_10480,N_8514,N_6082);
or U10481 (N_10481,N_9541,N_9107);
and U10482 (N_10482,N_9796,N_5220);
nand U10483 (N_10483,N_9850,N_6973);
and U10484 (N_10484,N_7155,N_7450);
or U10485 (N_10485,N_6648,N_8916);
or U10486 (N_10486,N_5826,N_9072);
nand U10487 (N_10487,N_8659,N_6862);
or U10488 (N_10488,N_7284,N_6187);
nor U10489 (N_10489,N_7524,N_9154);
or U10490 (N_10490,N_6764,N_5231);
or U10491 (N_10491,N_5625,N_7380);
nor U10492 (N_10492,N_8141,N_6085);
or U10493 (N_10493,N_8179,N_6012);
nor U10494 (N_10494,N_8993,N_7162);
xor U10495 (N_10495,N_5805,N_8286);
nand U10496 (N_10496,N_7844,N_5657);
nor U10497 (N_10497,N_6914,N_7415);
nand U10498 (N_10498,N_7679,N_7279);
or U10499 (N_10499,N_7869,N_6578);
and U10500 (N_10500,N_9921,N_8908);
nor U10501 (N_10501,N_5812,N_6131);
nor U10502 (N_10502,N_5586,N_5005);
or U10503 (N_10503,N_7045,N_6522);
and U10504 (N_10504,N_9943,N_5981);
and U10505 (N_10505,N_5302,N_5859);
or U10506 (N_10506,N_9301,N_9550);
or U10507 (N_10507,N_6031,N_7929);
xnor U10508 (N_10508,N_7622,N_9628);
xor U10509 (N_10509,N_6892,N_9236);
and U10510 (N_10510,N_6724,N_7794);
xnor U10511 (N_10511,N_5546,N_6719);
nor U10512 (N_10512,N_6248,N_5921);
xor U10513 (N_10513,N_6750,N_7466);
nand U10514 (N_10514,N_7483,N_7347);
nand U10515 (N_10515,N_7599,N_6223);
xor U10516 (N_10516,N_9908,N_9347);
and U10517 (N_10517,N_8322,N_7109);
nand U10518 (N_10518,N_9330,N_7686);
nand U10519 (N_10519,N_7840,N_8043);
nand U10520 (N_10520,N_9554,N_7264);
or U10521 (N_10521,N_8926,N_5270);
nor U10522 (N_10522,N_8246,N_7768);
and U10523 (N_10523,N_8823,N_7107);
nor U10524 (N_10524,N_5110,N_9747);
or U10525 (N_10525,N_7543,N_6254);
and U10526 (N_10526,N_9894,N_6617);
and U10527 (N_10527,N_7026,N_8013);
nand U10528 (N_10528,N_7661,N_8752);
or U10529 (N_10529,N_5609,N_6481);
or U10530 (N_10530,N_5150,N_6399);
nor U10531 (N_10531,N_7029,N_6803);
or U10532 (N_10532,N_6241,N_6138);
and U10533 (N_10533,N_8297,N_6782);
nand U10534 (N_10534,N_6630,N_5521);
nor U10535 (N_10535,N_8843,N_6184);
or U10536 (N_10536,N_6855,N_8030);
and U10537 (N_10537,N_8229,N_5484);
or U10538 (N_10538,N_5576,N_9913);
nand U10539 (N_10539,N_9560,N_7063);
nand U10540 (N_10540,N_9101,N_6153);
nor U10541 (N_10541,N_9661,N_9085);
and U10542 (N_10542,N_6500,N_7674);
or U10543 (N_10543,N_9721,N_6022);
nand U10544 (N_10544,N_5366,N_9316);
xnor U10545 (N_10545,N_6110,N_5650);
nor U10546 (N_10546,N_7762,N_5622);
or U10547 (N_10547,N_8108,N_5140);
nand U10548 (N_10548,N_6108,N_6722);
and U10549 (N_10549,N_7132,N_6440);
and U10550 (N_10550,N_6735,N_8071);
and U10551 (N_10551,N_7357,N_9372);
and U10552 (N_10552,N_6758,N_6214);
nor U10553 (N_10553,N_9383,N_6552);
or U10554 (N_10554,N_7597,N_5218);
nand U10555 (N_10555,N_8565,N_7750);
nand U10556 (N_10556,N_5730,N_7545);
and U10557 (N_10557,N_6624,N_5984);
and U10558 (N_10558,N_6876,N_7373);
nand U10559 (N_10559,N_7563,N_9924);
nor U10560 (N_10560,N_6919,N_5888);
and U10561 (N_10561,N_9787,N_7292);
or U10562 (N_10562,N_8754,N_5825);
or U10563 (N_10563,N_9242,N_8376);
nand U10564 (N_10564,N_6231,N_6875);
or U10565 (N_10565,N_8018,N_9109);
nand U10566 (N_10566,N_6447,N_8877);
nand U10567 (N_10567,N_9379,N_7475);
nand U10568 (N_10568,N_5637,N_7352);
or U10569 (N_10569,N_8145,N_6989);
nand U10570 (N_10570,N_8204,N_9060);
nor U10571 (N_10571,N_8702,N_6433);
nor U10572 (N_10572,N_5170,N_9037);
and U10573 (N_10573,N_8903,N_7540);
nand U10574 (N_10574,N_7140,N_9654);
or U10575 (N_10575,N_7041,N_7691);
nor U10576 (N_10576,N_6290,N_8205);
or U10577 (N_10577,N_9435,N_7610);
nor U10578 (N_10578,N_9681,N_5120);
or U10579 (N_10579,N_6236,N_6889);
or U10580 (N_10580,N_9141,N_5238);
or U10581 (N_10581,N_9223,N_5227);
and U10582 (N_10582,N_7392,N_7417);
or U10583 (N_10583,N_7703,N_6868);
and U10584 (N_10584,N_9749,N_7401);
and U10585 (N_10585,N_6088,N_6244);
nand U10586 (N_10586,N_5724,N_6870);
and U10587 (N_10587,N_5803,N_7955);
nand U10588 (N_10588,N_6097,N_7910);
and U10589 (N_10589,N_8447,N_7544);
nor U10590 (N_10590,N_9134,N_7002);
and U10591 (N_10591,N_7342,N_7714);
nand U10592 (N_10592,N_9445,N_7764);
xor U10593 (N_10593,N_8074,N_9764);
and U10594 (N_10594,N_5925,N_5049);
and U10595 (N_10595,N_8954,N_7548);
nor U10596 (N_10596,N_7626,N_5307);
nor U10597 (N_10597,N_8064,N_9627);
and U10598 (N_10598,N_7037,N_9196);
and U10599 (N_10599,N_9961,N_8997);
or U10600 (N_10600,N_9704,N_6794);
or U10601 (N_10601,N_5251,N_8299);
or U10602 (N_10602,N_7075,N_6338);
xor U10603 (N_10603,N_5510,N_7183);
nand U10604 (N_10604,N_8898,N_6741);
nor U10605 (N_10605,N_8426,N_7253);
and U10606 (N_10606,N_7267,N_8311);
or U10607 (N_10607,N_6279,N_5013);
or U10608 (N_10608,N_6027,N_6415);
nand U10609 (N_10609,N_6562,N_7940);
nor U10610 (N_10610,N_7754,N_6538);
and U10611 (N_10611,N_9633,N_6024);
or U10612 (N_10612,N_6330,N_7013);
or U10613 (N_10613,N_7770,N_7989);
xor U10614 (N_10614,N_9306,N_5325);
or U10615 (N_10615,N_6300,N_8052);
and U10616 (N_10616,N_6135,N_9455);
nor U10617 (N_10617,N_6120,N_5838);
nand U10618 (N_10618,N_6775,N_9468);
or U10619 (N_10619,N_9139,N_7766);
nor U10620 (N_10620,N_7131,N_5158);
nor U10621 (N_10621,N_6288,N_8549);
xor U10622 (N_10622,N_9737,N_8495);
nand U10623 (N_10623,N_5080,N_7418);
nand U10624 (N_10624,N_7289,N_7983);
or U10625 (N_10625,N_5898,N_6104);
and U10626 (N_10626,N_8629,N_6707);
nand U10627 (N_10627,N_5808,N_9759);
nand U10628 (N_10628,N_5960,N_8917);
or U10629 (N_10629,N_7846,N_6638);
and U10630 (N_10630,N_7113,N_5734);
nand U10631 (N_10631,N_6777,N_9057);
and U10632 (N_10632,N_9770,N_9734);
nand U10633 (N_10633,N_7093,N_5943);
nand U10634 (N_10634,N_5317,N_6936);
xor U10635 (N_10635,N_5779,N_5694);
nand U10636 (N_10636,N_7506,N_5928);
and U10637 (N_10637,N_5015,N_5168);
and U10638 (N_10638,N_6155,N_7067);
or U10639 (N_10639,N_7776,N_6795);
nor U10640 (N_10640,N_5766,N_5405);
nor U10641 (N_10641,N_9581,N_5478);
and U10642 (N_10642,N_8487,N_6185);
nor U10643 (N_10643,N_7868,N_7316);
and U10644 (N_10644,N_6092,N_9982);
and U10645 (N_10645,N_5353,N_7667);
and U10646 (N_10646,N_8853,N_6071);
nand U10647 (N_10647,N_7128,N_6190);
and U10648 (N_10648,N_5385,N_7678);
nand U10649 (N_10649,N_9708,N_5215);
or U10650 (N_10650,N_6026,N_9643);
xnor U10651 (N_10651,N_6165,N_9983);
and U10652 (N_10652,N_6090,N_6163);
xnor U10653 (N_10653,N_9887,N_6180);
nor U10654 (N_10654,N_5332,N_6543);
or U10655 (N_10655,N_8848,N_5346);
or U10656 (N_10656,N_6349,N_8451);
nor U10657 (N_10657,N_5971,N_6953);
or U10658 (N_10658,N_7496,N_6829);
nor U10659 (N_10659,N_7207,N_5050);
or U10660 (N_10660,N_9458,N_6576);
xnor U10661 (N_10661,N_6537,N_6967);
or U10662 (N_10662,N_5343,N_5872);
nand U10663 (N_10663,N_9812,N_6705);
nor U10664 (N_10664,N_6061,N_9091);
and U10665 (N_10665,N_7923,N_6536);
nand U10666 (N_10666,N_9384,N_5717);
and U10667 (N_10667,N_8888,N_8633);
and U10668 (N_10668,N_7577,N_5338);
and U10669 (N_10669,N_6838,N_9577);
and U10670 (N_10670,N_6547,N_8420);
nor U10671 (N_10671,N_7046,N_9880);
nand U10672 (N_10672,N_6728,N_5086);
nor U10673 (N_10673,N_5745,N_8358);
nand U10674 (N_10674,N_8000,N_8516);
and U10675 (N_10675,N_6115,N_7906);
nand U10676 (N_10676,N_5893,N_8213);
nand U10677 (N_10677,N_5844,N_8345);
nand U10678 (N_10678,N_5889,N_7381);
nor U10679 (N_10679,N_7158,N_9495);
nand U10680 (N_10680,N_9939,N_7801);
or U10681 (N_10681,N_5304,N_7885);
or U10682 (N_10682,N_9195,N_9866);
and U10683 (N_10683,N_5459,N_9626);
nand U10684 (N_10684,N_7098,N_6329);
nand U10685 (N_10685,N_5728,N_6602);
and U10686 (N_10686,N_6052,N_7255);
and U10687 (N_10687,N_7423,N_6274);
and U10688 (N_10688,N_8244,N_9565);
or U10689 (N_10689,N_5946,N_6368);
or U10690 (N_10690,N_5000,N_7571);
nor U10691 (N_10691,N_9752,N_6820);
nor U10692 (N_10692,N_8277,N_5676);
nor U10693 (N_10693,N_5301,N_7831);
xor U10694 (N_10694,N_9827,N_8944);
or U10695 (N_10695,N_6674,N_5403);
xor U10696 (N_10696,N_9757,N_5250);
nor U10697 (N_10697,N_9271,N_8890);
nand U10698 (N_10698,N_8477,N_6036);
or U10699 (N_10699,N_8862,N_7217);
and U10700 (N_10700,N_6997,N_7135);
and U10701 (N_10701,N_5482,N_5263);
xor U10702 (N_10702,N_9868,N_5245);
nand U10703 (N_10703,N_7077,N_6508);
and U10704 (N_10704,N_8437,N_6792);
xnor U10705 (N_10705,N_5268,N_7124);
nand U10706 (N_10706,N_6256,N_8645);
xnor U10707 (N_10707,N_5365,N_7227);
and U10708 (N_10708,N_8931,N_7254);
and U10709 (N_10709,N_5376,N_8646);
nand U10710 (N_10710,N_6406,N_8366);
and U10711 (N_10711,N_7651,N_7073);
and U10712 (N_10712,N_9144,N_9546);
nand U10713 (N_10713,N_9251,N_7345);
xnor U10714 (N_10714,N_5791,N_8607);
nor U10715 (N_10715,N_8142,N_9623);
nand U10716 (N_10716,N_7588,N_6677);
or U10717 (N_10717,N_5292,N_7729);
nand U10718 (N_10718,N_7011,N_5643);
nor U10719 (N_10719,N_7713,N_9250);
or U10720 (N_10720,N_5371,N_8876);
and U10721 (N_10721,N_7395,N_8109);
and U10722 (N_10722,N_5286,N_9854);
xor U10723 (N_10723,N_8864,N_7919);
nor U10724 (N_10724,N_7318,N_5904);
and U10725 (N_10725,N_6418,N_8059);
nand U10726 (N_10726,N_7656,N_9464);
nand U10727 (N_10727,N_6828,N_9629);
nor U10728 (N_10728,N_9412,N_9888);
and U10729 (N_10729,N_7319,N_6072);
or U10730 (N_10730,N_5051,N_5319);
nand U10731 (N_10731,N_7248,N_7358);
nand U10732 (N_10732,N_9148,N_9188);
or U10733 (N_10733,N_5700,N_5659);
nor U10734 (N_10734,N_7047,N_6825);
nor U10735 (N_10735,N_8846,N_8153);
nand U10736 (N_10736,N_7156,N_9467);
and U10737 (N_10737,N_5228,N_7315);
and U10738 (N_10738,N_5820,N_9149);
nand U10739 (N_10739,N_6710,N_7565);
or U10740 (N_10740,N_8527,N_6789);
nor U10741 (N_10741,N_9387,N_5979);
nor U10742 (N_10742,N_7076,N_8240);
xnor U10743 (N_10743,N_7810,N_6651);
nor U10744 (N_10744,N_6394,N_8135);
and U10745 (N_10745,N_5010,N_7587);
nor U10746 (N_10746,N_7564,N_7972);
or U10747 (N_10747,N_9774,N_8765);
and U10748 (N_10748,N_6599,N_7633);
nand U10749 (N_10749,N_6532,N_5628);
and U10750 (N_10750,N_6370,N_9904);
nand U10751 (N_10751,N_5527,N_9110);
and U10752 (N_10752,N_8718,N_6809);
nand U10753 (N_10753,N_6655,N_8201);
xor U10754 (N_10754,N_5752,N_8709);
xor U10755 (N_10755,N_6704,N_7455);
nand U10756 (N_10756,N_5097,N_6323);
and U10757 (N_10757,N_6122,N_8854);
or U10758 (N_10758,N_6608,N_5408);
or U10759 (N_10759,N_6164,N_7693);
and U10760 (N_10760,N_5913,N_6234);
nor U10761 (N_10761,N_7355,N_7190);
xnor U10762 (N_10762,N_9636,N_7163);
xnor U10763 (N_10763,N_5524,N_7089);
nor U10764 (N_10764,N_6939,N_9705);
or U10765 (N_10765,N_6604,N_7185);
and U10766 (N_10766,N_9421,N_8557);
nor U10767 (N_10767,N_9655,N_6293);
nand U10768 (N_10768,N_5634,N_5126);
nor U10769 (N_10769,N_9183,N_7538);
xor U10770 (N_10770,N_9886,N_6216);
xnor U10771 (N_10771,N_7136,N_8344);
nor U10772 (N_10772,N_8253,N_9356);
nand U10773 (N_10773,N_9816,N_5809);
nor U10774 (N_10774,N_6049,N_9269);
nand U10775 (N_10775,N_7575,N_6307);
nand U10776 (N_10776,N_7205,N_7350);
and U10777 (N_10777,N_8844,N_6436);
xnor U10778 (N_10778,N_9679,N_6593);
or U10779 (N_10779,N_9429,N_7662);
nand U10780 (N_10780,N_9077,N_6044);
and U10781 (N_10781,N_6912,N_8014);
nor U10782 (N_10782,N_7956,N_8522);
or U10783 (N_10783,N_9855,N_5613);
nand U10784 (N_10784,N_9088,N_9930);
or U10785 (N_10785,N_7952,N_8137);
nand U10786 (N_10786,N_8241,N_9158);
nand U10787 (N_10787,N_7283,N_7874);
or U10788 (N_10788,N_8939,N_7888);
nor U10789 (N_10789,N_6695,N_8391);
xnor U10790 (N_10790,N_5431,N_8007);
or U10791 (N_10791,N_6477,N_8464);
nand U10792 (N_10792,N_5201,N_9702);
or U10793 (N_10793,N_5193,N_6915);
and U10794 (N_10794,N_6075,N_8690);
or U10795 (N_10795,N_8382,N_6832);
nor U10796 (N_10796,N_7968,N_5985);
xnor U10797 (N_10797,N_9199,N_5337);
xnor U10798 (N_10798,N_7364,N_5243);
and U10799 (N_10799,N_9588,N_9475);
nor U10800 (N_10800,N_5817,N_5062);
and U10801 (N_10801,N_8589,N_9168);
or U10802 (N_10802,N_7642,N_6952);
and U10803 (N_10803,N_5014,N_8865);
nand U10804 (N_10804,N_7664,N_7779);
and U10805 (N_10805,N_9454,N_7592);
nand U10806 (N_10806,N_9517,N_6454);
and U10807 (N_10807,N_6317,N_8342);
xnor U10808 (N_10808,N_8417,N_5308);
nor U10809 (N_10809,N_7499,N_9465);
nor U10810 (N_10810,N_6060,N_9415);
nand U10811 (N_10811,N_5835,N_5804);
nand U10812 (N_10812,N_5632,N_6209);
or U10813 (N_10813,N_5171,N_6557);
nand U10814 (N_10814,N_8624,N_8121);
nor U10815 (N_10815,N_9273,N_5452);
and U10816 (N_10816,N_6974,N_9392);
nand U10817 (N_10817,N_7103,N_6103);
or U10818 (N_10818,N_8818,N_6424);
and U10819 (N_10819,N_6002,N_7880);
and U10820 (N_10820,N_9418,N_9295);
and U10821 (N_10821,N_8635,N_8850);
nor U10822 (N_10822,N_5756,N_5910);
xnor U10823 (N_10823,N_7671,N_6924);
nor U10824 (N_10824,N_5446,N_8268);
and U10825 (N_10825,N_5901,N_7737);
xnor U10826 (N_10826,N_6796,N_8360);
nand U10827 (N_10827,N_9232,N_9728);
nand U10828 (N_10828,N_9399,N_8362);
or U10829 (N_10829,N_6941,N_9241);
nor U10830 (N_10830,N_8430,N_5677);
nor U10831 (N_10831,N_6121,N_8594);
nand U10832 (N_10832,N_9489,N_6393);
xnor U10833 (N_10833,N_7876,N_9369);
xor U10834 (N_10834,N_7617,N_5675);
or U10835 (N_10835,N_7230,N_9831);
or U10836 (N_10836,N_5539,N_7321);
nand U10837 (N_10837,N_9527,N_8682);
and U10838 (N_10838,N_9096,N_5899);
nand U10839 (N_10839,N_7665,N_5743);
and U10840 (N_10840,N_8775,N_6833);
and U10841 (N_10841,N_9668,N_5162);
and U10842 (N_10842,N_9389,N_7606);
and U10843 (N_10843,N_6456,N_7463);
nand U10844 (N_10844,N_7180,N_9311);
nor U10845 (N_10845,N_5288,N_6355);
xnor U10846 (N_10846,N_9187,N_8262);
nor U10847 (N_10847,N_9882,N_5849);
nor U10848 (N_10848,N_5200,N_8252);
nor U10849 (N_10849,N_7341,N_6230);
or U10850 (N_10850,N_9837,N_9806);
nand U10851 (N_10851,N_8001,N_5349);
or U10852 (N_10852,N_8305,N_7121);
nand U10853 (N_10853,N_5877,N_8154);
or U10854 (N_10854,N_5248,N_8895);
nand U10855 (N_10855,N_8019,N_5753);
or U10856 (N_10856,N_7389,N_5203);
and U10857 (N_10857,N_6237,N_7569);
or U10858 (N_10858,N_9124,N_7531);
or U10859 (N_10859,N_7824,N_5600);
or U10860 (N_10860,N_8562,N_9325);
nor U10861 (N_10861,N_9448,N_5982);
nor U10862 (N_10862,N_7090,N_7441);
and U10863 (N_10863,N_6247,N_9875);
or U10864 (N_10864,N_8729,N_9303);
nor U10865 (N_10865,N_5374,N_7427);
or U10866 (N_10866,N_5426,N_6824);
and U10867 (N_10867,N_7151,N_8585);
nor U10868 (N_10868,N_5177,N_8073);
nor U10869 (N_10869,N_5922,N_5159);
and U10870 (N_10870,N_8794,N_6756);
and U10871 (N_10871,N_8587,N_7979);
and U10872 (N_10872,N_5592,N_5068);
xor U10873 (N_10873,N_5685,N_9350);
nand U10874 (N_10874,N_7997,N_5289);
and U10875 (N_10875,N_9647,N_6667);
nand U10876 (N_10876,N_6067,N_9127);
or U10877 (N_10877,N_5135,N_7268);
nand U10878 (N_10878,N_5435,N_5535);
or U10879 (N_10879,N_8129,N_6860);
and U10880 (N_10880,N_7096,N_7604);
nor U10881 (N_10881,N_7489,N_8996);
or U10882 (N_10882,N_8689,N_5869);
nand U10883 (N_10883,N_8463,N_9712);
and U10884 (N_10884,N_7849,N_7668);
or U10885 (N_10885,N_8296,N_9300);
or U10886 (N_10886,N_7309,N_6251);
or U10887 (N_10887,N_9486,N_7030);
nor U10888 (N_10888,N_5684,N_8999);
nand U10889 (N_10889,N_9976,N_5941);
nand U10890 (N_10890,N_9488,N_8611);
xor U10891 (N_10891,N_5939,N_6981);
nand U10892 (N_10892,N_7701,N_8497);
nor U10893 (N_10893,N_9505,N_8498);
and U10894 (N_10894,N_6504,N_7161);
and U10895 (N_10895,N_6463,N_6745);
and U10896 (N_10896,N_9484,N_6413);
nor U10897 (N_10897,N_6438,N_6801);
xnor U10898 (N_10898,N_8602,N_7102);
nor U10899 (N_10899,N_8392,N_9446);
nand U10900 (N_10900,N_7595,N_9530);
and U10901 (N_10901,N_8365,N_8148);
nand U10902 (N_10902,N_9411,N_9373);
nand U10903 (N_10903,N_8003,N_5886);
or U10904 (N_10904,N_6448,N_8748);
and U10905 (N_10905,N_5130,N_9817);
or U10906 (N_10906,N_7513,N_9656);
nand U10907 (N_10907,N_8077,N_5952);
and U10908 (N_10908,N_6711,N_5381);
and U10909 (N_10909,N_8287,N_8882);
or U10910 (N_10910,N_7149,N_9596);
or U10911 (N_10911,N_7902,N_8967);
and U10912 (N_10912,N_6034,N_5793);
nand U10913 (N_10913,N_7209,N_8953);
and U10914 (N_10914,N_9427,N_8314);
nor U10915 (N_10915,N_6662,N_8656);
and U10916 (N_10916,N_7659,N_7239);
or U10917 (N_10917,N_7695,N_9500);
xor U10918 (N_10918,N_9952,N_8663);
and U10919 (N_10919,N_9925,N_7053);
or U10920 (N_10920,N_6613,N_5179);
nand U10921 (N_10921,N_7091,N_9761);
and U10922 (N_10922,N_9780,N_9262);
nor U10923 (N_10923,N_9735,N_7650);
or U10924 (N_10924,N_5210,N_7975);
or U10925 (N_10925,N_5807,N_6933);
nand U10926 (N_10926,N_7133,N_5763);
nand U10927 (N_10927,N_6835,N_5025);
or U10928 (N_10928,N_7903,N_9348);
xor U10929 (N_10929,N_9181,N_9293);
nand U10930 (N_10930,N_9929,N_5755);
and U10931 (N_10931,N_9026,N_5450);
or U10932 (N_10932,N_8797,N_9002);
or U10933 (N_10933,N_7377,N_7172);
or U10934 (N_10934,N_9996,N_9946);
nand U10935 (N_10935,N_7791,N_9166);
nand U10936 (N_10936,N_8781,N_7334);
nor U10937 (N_10937,N_7510,N_8760);
or U10938 (N_10938,N_7122,N_9029);
nor U10939 (N_10939,N_9408,N_8768);
nand U10940 (N_10940,N_9699,N_7242);
and U10941 (N_10941,N_5523,N_8977);
or U10942 (N_10942,N_6569,N_8106);
and U10943 (N_10943,N_7422,N_6013);
xnor U10944 (N_10944,N_8773,N_7586);
nor U10945 (N_10945,N_9424,N_7769);
nor U10946 (N_10946,N_8419,N_8318);
or U10947 (N_10947,N_9420,N_5285);
nand U10948 (N_10948,N_8446,N_6011);
and U10949 (N_10949,N_6885,N_6970);
or U10950 (N_10950,N_5129,N_6404);
nand U10951 (N_10951,N_5702,N_9491);
or U10952 (N_10952,N_5344,N_6482);
or U10953 (N_10953,N_6051,N_5775);
and U10954 (N_10954,N_5318,N_8793);
nor U10955 (N_10955,N_8955,N_9302);
xor U10956 (N_10956,N_9619,N_6147);
xor U10957 (N_10957,N_6375,N_5421);
and U10958 (N_10958,N_8332,N_9394);
xor U10959 (N_10959,N_5560,N_8581);
nor U10960 (N_10960,N_9351,N_6419);
nor U10961 (N_10961,N_6112,N_8779);
nor U10962 (N_10962,N_5221,N_5362);
or U10963 (N_10963,N_5519,N_8295);
or U10964 (N_10964,N_9177,N_6331);
nor U10965 (N_10965,N_8216,N_7504);
and U10966 (N_10966,N_6830,N_6431);
or U10967 (N_10967,N_9480,N_8301);
nand U10968 (N_10968,N_9339,N_5567);
nand U10969 (N_10969,N_8191,N_8456);
nand U10970 (N_10970,N_9745,N_9972);
and U10971 (N_10971,N_8859,N_6040);
or U10972 (N_10972,N_9532,N_5716);
nor U10973 (N_10973,N_8138,N_5313);
nor U10974 (N_10974,N_7006,N_6843);
or U10975 (N_10975,N_6157,N_9312);
or U10976 (N_10976,N_5761,N_9033);
nor U10977 (N_10977,N_5944,N_6771);
or U10978 (N_10978,N_5926,N_9191);
nor U10979 (N_10979,N_5674,N_6918);
nor U10980 (N_10980,N_6259,N_9918);
or U10981 (N_10981,N_8476,N_5718);
and U10982 (N_10982,N_5223,N_8563);
nor U10983 (N_10983,N_5906,N_8494);
or U10984 (N_10984,N_6696,N_5602);
or U10985 (N_10985,N_7301,N_8837);
or U10986 (N_10986,N_8692,N_7746);
nor U10987 (N_10987,N_8524,N_5271);
or U10988 (N_10988,N_9773,N_6252);
nand U10989 (N_10989,N_7154,N_6407);
and U10990 (N_10990,N_6087,N_7744);
or U10991 (N_10991,N_6139,N_7386);
or U10992 (N_10992,N_9332,N_9717);
and U10993 (N_10993,N_6621,N_7556);
nand U10994 (N_10994,N_9008,N_5570);
or U10995 (N_10995,N_8036,N_6291);
and U10996 (N_10996,N_6282,N_8375);
xnor U10997 (N_10997,N_7928,N_5056);
or U10998 (N_10998,N_5525,N_6612);
and U10999 (N_10999,N_9438,N_7864);
and U11000 (N_11000,N_5469,N_7445);
and U11001 (N_11001,N_8405,N_8598);
and U11002 (N_11002,N_6752,N_9874);
or U11003 (N_11003,N_6336,N_9986);
and U11004 (N_11004,N_6788,N_9386);
and U11005 (N_11005,N_8025,N_5453);
nor U11006 (N_11006,N_5938,N_9594);
and U11007 (N_11007,N_8665,N_5485);
or U11008 (N_11008,N_5146,N_5591);
nand U11009 (N_11009,N_5087,N_6193);
nand U11010 (N_11010,N_9147,N_7731);
nand U11011 (N_11011,N_6462,N_5714);
or U11012 (N_11012,N_7865,N_6762);
or U11013 (N_11013,N_8502,N_6377);
or U11014 (N_11014,N_7000,N_6038);
nand U11015 (N_11015,N_7836,N_5672);
xnor U11016 (N_11016,N_8675,N_5395);
or U11017 (N_11017,N_9336,N_8616);
nor U11018 (N_11018,N_8547,N_8789);
and U11019 (N_11019,N_5189,N_8175);
or U11020 (N_11020,N_6495,N_5137);
nand U11021 (N_11021,N_7562,N_9902);
or U11022 (N_11022,N_6682,N_6770);
or U11023 (N_11023,N_6079,N_5933);
nor U11024 (N_11024,N_7153,N_6219);
nor U11025 (N_11025,N_7623,N_9557);
nor U11026 (N_11026,N_9889,N_5004);
and U11027 (N_11027,N_6995,N_7413);
or U11028 (N_11028,N_9221,N_5182);
xor U11029 (N_11029,N_5265,N_5736);
nor U11030 (N_11030,N_8796,N_6089);
nand U11031 (N_11031,N_7270,N_5008);
or U11032 (N_11032,N_9978,N_5275);
and U11033 (N_11033,N_5986,N_7580);
or U11034 (N_11034,N_7666,N_5456);
or U11035 (N_11035,N_9042,N_8719);
xnor U11036 (N_11036,N_8723,N_5679);
nand U11037 (N_11037,N_9112,N_5853);
and U11038 (N_11038,N_6567,N_7612);
and U11039 (N_11039,N_8762,N_9313);
or U11040 (N_11040,N_8482,N_8369);
or U11041 (N_11041,N_6817,N_5951);
xnor U11042 (N_11042,N_9222,N_5999);
and U11043 (N_11043,N_8324,N_5373);
or U11044 (N_11044,N_6744,N_9750);
nor U11045 (N_11045,N_9155,N_6691);
xor U11046 (N_11046,N_5785,N_7464);
nor U11047 (N_11047,N_8115,N_5710);
nand U11048 (N_11048,N_7627,N_5038);
nor U11049 (N_11049,N_5508,N_8208);
nand U11050 (N_11050,N_8427,N_6467);
or U11051 (N_11051,N_6700,N_8648);
and U11052 (N_11052,N_7618,N_8251);
nor U11053 (N_11053,N_7116,N_8438);
and U11054 (N_11054,N_6390,N_8680);
and U11055 (N_11055,N_5723,N_6813);
nor U11056 (N_11056,N_7038,N_8133);
nand U11057 (N_11057,N_9176,N_6731);
or U11058 (N_11058,N_9437,N_8393);
xor U11059 (N_11059,N_8491,N_9973);
or U11060 (N_11060,N_8840,N_8708);
or U11061 (N_11061,N_8965,N_9977);
and U11062 (N_11062,N_7325,N_9586);
and U11063 (N_11063,N_9598,N_9259);
or U11064 (N_11064,N_7297,N_9274);
nand U11065 (N_11065,N_5064,N_9131);
nand U11066 (N_11066,N_5532,N_6018);
or U11067 (N_11067,N_7889,N_6173);
nor U11068 (N_11068,N_7040,N_5660);
nand U11069 (N_11069,N_6239,N_5911);
and U11070 (N_11070,N_5229,N_7677);
or U11071 (N_11071,N_5022,N_7852);
nor U11072 (N_11072,N_5443,N_5742);
nand U11073 (N_11073,N_7410,N_7958);
and U11074 (N_11074,N_9864,N_6748);
or U11075 (N_11075,N_7170,N_8044);
and U11076 (N_11076,N_9164,N_9582);
and U11077 (N_11077,N_8783,N_6886);
or U11078 (N_11078,N_5173,N_8564);
and U11079 (N_11079,N_6858,N_7856);
and U11080 (N_11080,N_6929,N_6000);
nor U11081 (N_11081,N_6306,N_5198);
or U11082 (N_11082,N_9993,N_6333);
or U11083 (N_11083,N_7799,N_8889);
nand U11084 (N_11084,N_8957,N_6006);
xor U11085 (N_11085,N_5031,N_6546);
or U11086 (N_11086,N_9725,N_7921);
nand U11087 (N_11087,N_8574,N_5222);
nor U11088 (N_11088,N_5085,N_9605);
nor U11089 (N_11089,N_7023,N_5776);
and U11090 (N_11090,N_6132,N_7937);
and U11091 (N_11091,N_8057,N_6149);
nor U11092 (N_11092,N_6073,N_6320);
xor U11093 (N_11093,N_7472,N_6527);
nor U11094 (N_11094,N_7579,N_6831);
nand U11095 (N_11095,N_7397,N_5758);
or U11096 (N_11096,N_6391,N_5260);
xor U11097 (N_11097,N_6408,N_8478);
nand U11098 (N_11098,N_5708,N_8022);
or U11099 (N_11099,N_9094,N_6708);
and U11100 (N_11100,N_5314,N_5690);
and U11101 (N_11101,N_9245,N_5656);
nand U11102 (N_11102,N_5309,N_8276);
xnor U11103 (N_11103,N_5715,N_7704);
and U11104 (N_11104,N_7833,N_7705);
nor U11105 (N_11105,N_6897,N_7226);
and U11106 (N_11106,N_8348,N_5929);
nand U11107 (N_11107,N_5436,N_6316);
or U11108 (N_11108,N_7007,N_8258);
nand U11109 (N_11109,N_9592,N_8099);
nand U11110 (N_11110,N_7437,N_9341);
nand U11111 (N_11111,N_9476,N_8481);
nor U11112 (N_11112,N_7244,N_5564);
xor U11113 (N_11113,N_6873,N_8668);
nand U11114 (N_11114,N_8513,N_5494);
nor U11115 (N_11115,N_8490,N_6718);
and U11116 (N_11116,N_9416,N_6437);
nor U11117 (N_11117,N_8666,N_9775);
or U11118 (N_11118,N_8860,N_6096);
or U11119 (N_11119,N_5635,N_7473);
and U11120 (N_11120,N_7460,N_8732);
xor U11121 (N_11121,N_7663,N_8187);
and U11122 (N_11122,N_8380,N_9622);
nor U11123 (N_11123,N_8271,N_7907);
nand U11124 (N_11124,N_8812,N_5424);
or U11125 (N_11125,N_5078,N_6432);
nand U11126 (N_11126,N_5538,N_8622);
or U11127 (N_11127,N_9214,N_7106);
and U11128 (N_11128,N_6488,N_7331);
nor U11129 (N_11129,N_5787,N_5865);
nor U11130 (N_11130,N_5433,N_6505);
nor U11131 (N_11131,N_5516,N_7886);
nand U11132 (N_11132,N_8123,N_7470);
or U11133 (N_11133,N_8505,N_6793);
or U11134 (N_11134,N_9766,N_8534);
or U11135 (N_11135,N_7419,N_5749);
and U11136 (N_11136,N_9825,N_6742);
or U11137 (N_11137,N_6258,N_9265);
or U11138 (N_11138,N_5581,N_8669);
nand U11139 (N_11139,N_5280,N_7481);
nor U11140 (N_11140,N_5638,N_5406);
and U11141 (N_11141,N_6715,N_8899);
nand U11142 (N_11142,N_9257,N_8211);
nand U11143 (N_11143,N_5483,N_7502);
nor U11144 (N_11144,N_9129,N_9807);
and U11145 (N_11145,N_8510,N_8125);
nor U11146 (N_11146,N_7788,N_9410);
and U11147 (N_11147,N_8792,N_5230);
and U11148 (N_11148,N_5504,N_9567);
nand U11149 (N_11149,N_8330,N_5083);
or U11150 (N_11150,N_5737,N_7376);
nand U11151 (N_11151,N_8432,N_8508);
xor U11152 (N_11152,N_5065,N_7372);
and U11153 (N_11153,N_8224,N_8152);
nor U11154 (N_11154,N_8981,N_9584);
or U11155 (N_11155,N_9079,N_5225);
nand U11156 (N_11156,N_5363,N_6954);
xor U11157 (N_11157,N_6669,N_7145);
or U11158 (N_11158,N_5282,N_8202);
or U11159 (N_11159,N_6763,N_9208);
xor U11160 (N_11160,N_7740,N_7416);
or U11161 (N_11161,N_5722,N_5001);
or U11162 (N_11162,N_6619,N_8966);
nand U11163 (N_11163,N_5195,N_7786);
nor U11164 (N_11164,N_6818,N_8107);
xnor U11165 (N_11165,N_5836,N_9125);
xor U11166 (N_11166,N_5439,N_5027);
and U11167 (N_11167,N_8740,N_6152);
nand U11168 (N_11168,N_6222,N_9267);
and U11169 (N_11169,N_5964,N_7446);
nand U11170 (N_11170,N_7080,N_7391);
nand U11171 (N_11171,N_6001,N_6702);
or U11172 (N_11172,N_8480,N_6416);
nand U11173 (N_11173,N_6106,N_9111);
and U11174 (N_11174,N_6503,N_5134);
or U11175 (N_11175,N_5937,N_7821);
and U11176 (N_11176,N_7079,N_7700);
or U11177 (N_11177,N_6311,N_8834);
or U11178 (N_11178,N_7771,N_9220);
nor U11179 (N_11179,N_8323,N_6294);
or U11180 (N_11180,N_7246,N_7503);
nand U11181 (N_11181,N_5063,N_6221);
and U11182 (N_11182,N_7110,N_7259);
or U11183 (N_11183,N_8701,N_5501);
nand U11184 (N_11184,N_6428,N_7147);
nor U11185 (N_11185,N_7060,N_5830);
or U11186 (N_11186,N_6784,N_8239);
nor U11187 (N_11187,N_8807,N_8658);
and U11188 (N_11188,N_9212,N_5183);
nand U11189 (N_11189,N_7378,N_7807);
or U11190 (N_11190,N_5542,N_9409);
or U11191 (N_11191,N_9873,N_8559);
xnor U11192 (N_11192,N_6371,N_6791);
nand U11193 (N_11193,N_7984,N_8539);
and U11194 (N_11194,N_5361,N_5326);
xnor U11195 (N_11195,N_6709,N_8852);
nand U11196 (N_11196,N_5425,N_5868);
nor U11197 (N_11197,N_8467,N_5967);
nand U11198 (N_11198,N_8600,N_7211);
nand U11199 (N_11199,N_6273,N_6268);
and U11200 (N_11200,N_7721,N_9660);
nand U11201 (N_11201,N_8378,N_8168);
and U11202 (N_11202,N_7815,N_6422);
nand U11203 (N_11203,N_9650,N_8550);
and U11204 (N_11204,N_8924,N_8093);
nand U11205 (N_11205,N_7490,N_5915);
or U11206 (N_11206,N_7986,N_6479);
xnor U11207 (N_11207,N_8182,N_9906);
nand U11208 (N_11208,N_5814,N_7349);
and U11209 (N_11209,N_7672,N_5699);
nand U11210 (N_11210,N_7461,N_9452);
nor U11211 (N_11211,N_5036,N_9504);
nand U11212 (N_11212,N_6633,N_9074);
or U11213 (N_11213,N_8657,N_9360);
nor U11214 (N_11214,N_9388,N_8642);
nand U11215 (N_11215,N_5124,N_9693);
nor U11216 (N_11216,N_9781,N_6443);
and U11217 (N_11217,N_5789,N_5607);
nand U11218 (N_11218,N_6475,N_9375);
xor U11219 (N_11219,N_8200,N_6810);
or U11220 (N_11220,N_6322,N_7970);
or U11221 (N_11221,N_8785,N_7314);
nor U11222 (N_11222,N_7813,N_9834);
and U11223 (N_11223,N_8697,N_9095);
nor U11224 (N_11224,N_7578,N_9440);
nand U11225 (N_11225,N_7293,N_5330);
or U11226 (N_11226,N_8943,N_6932);
nor U11227 (N_11227,N_5765,N_9200);
xor U11228 (N_11228,N_5178,N_5506);
xnor U11229 (N_11229,N_8452,N_5571);
and U11230 (N_11230,N_6746,N_9400);
and U11231 (N_11231,N_8444,N_8031);
nand U11232 (N_11232,N_6123,N_7991);
xor U11233 (N_11233,N_6799,N_9507);
nor U11234 (N_11234,N_5441,N_7018);
nand U11235 (N_11235,N_5388,N_8745);
nor U11236 (N_11236,N_5095,N_6341);
or U11237 (N_11237,N_9358,N_8558);
or U11238 (N_11238,N_9815,N_8161);
or U11239 (N_11239,N_9190,N_8849);
and U11240 (N_11240,N_6598,N_8654);
nor U11241 (N_11241,N_7003,N_8114);
nor U11242 (N_11242,N_9732,N_9434);
and U11243 (N_11243,N_6162,N_9653);
and U11244 (N_11244,N_9756,N_6083);
and U11245 (N_11245,N_8520,N_7074);
and U11246 (N_11246,N_7056,N_5878);
xor U11247 (N_11247,N_6739,N_6585);
or U11248 (N_11248,N_7061,N_8313);
or U11249 (N_11249,N_9835,N_6802);
and U11250 (N_11250,N_8217,N_5617);
and U11251 (N_11251,N_9320,N_9171);
and U11252 (N_11252,N_8703,N_5295);
and U11253 (N_11253,N_6804,N_7104);
xnor U11254 (N_11254,N_6235,N_9328);
nand U11255 (N_11255,N_9036,N_7052);
nor U11256 (N_11256,N_5347,N_9664);
nor U11257 (N_11257,N_8349,N_7468);
and U11258 (N_11258,N_5611,N_7222);
and U11259 (N_11259,N_9616,N_7932);
and U11260 (N_11260,N_6189,N_9992);
nor U11261 (N_11261,N_8503,N_7957);
nand U11262 (N_11262,N_8336,N_6086);
or U11263 (N_11263,N_7125,N_6566);
or U11264 (N_11264,N_9405,N_8041);
nor U11265 (N_11265,N_6156,N_7051);
nand U11266 (N_11266,N_6926,N_8800);
xnor U11267 (N_11267,N_7790,N_7724);
and U11268 (N_11268,N_5061,N_7998);
or U11269 (N_11269,N_5320,N_5016);
or U11270 (N_11270,N_8950,N_5695);
nand U11271 (N_11271,N_5445,N_5300);
or U11272 (N_11272,N_6765,N_6689);
nor U11273 (N_11273,N_9175,N_6653);
or U11274 (N_11274,N_9286,N_5194);
and U11275 (N_11275,N_5108,N_5883);
nand U11276 (N_11276,N_8871,N_7394);
nor U11277 (N_11277,N_5090,N_9524);
nand U11278 (N_11278,N_6761,N_9538);
and U11279 (N_11279,N_6837,N_9509);
nor U11280 (N_11280,N_9552,N_6821);
nor U11281 (N_11281,N_5781,N_5795);
xor U11282 (N_11282,N_7291,N_9540);
and U11283 (N_11283,N_6064,N_8577);
and U11284 (N_11284,N_8593,N_6405);
and U11285 (N_11285,N_8742,N_5400);
xor U11286 (N_11286,N_7756,N_8912);
and U11287 (N_11287,N_5606,N_7184);
nand U11288 (N_11288,N_5687,N_6116);
xnor U11289 (N_11289,N_6174,N_8699);
nand U11290 (N_11290,N_7070,N_9914);
nor U11291 (N_11291,N_8803,N_7639);
nand U11292 (N_11292,N_7276,N_8450);
xnor U11293 (N_11293,N_6129,N_8218);
nor U11294 (N_11294,N_7221,N_7402);
nand U11295 (N_11295,N_6021,N_5615);
or U11296 (N_11296,N_7215,N_8601);
nor U11297 (N_11297,N_8473,N_8938);
nor U11298 (N_11298,N_7780,N_8309);
xnor U11299 (N_11299,N_7505,N_5980);
nor U11300 (N_11300,N_9867,N_9279);
nand U11301 (N_11301,N_7049,N_6339);
xnor U11302 (N_11302,N_5955,N_9829);
or U11303 (N_11303,N_7822,N_9045);
and U11304 (N_11304,N_7462,N_8767);
nor U11305 (N_11305,N_8355,N_5874);
nor U11306 (N_11306,N_9791,N_6632);
nor U11307 (N_11307,N_9954,N_7072);
xor U11308 (N_11308,N_6400,N_9634);
and U11309 (N_11309,N_7570,N_6854);
or U11310 (N_11310,N_6043,N_9518);
nor U11311 (N_11311,N_6618,N_6721);
nor U11312 (N_11312,N_5105,N_5927);
nand U11313 (N_11313,N_6699,N_5587);
or U11314 (N_11314,N_9963,N_6468);
or U11315 (N_11315,N_7669,N_7777);
and U11316 (N_11316,N_9206,N_9121);
nor U11317 (N_11317,N_5500,N_8483);
and U11318 (N_11318,N_5873,N_7882);
nor U11319 (N_11319,N_7036,N_7977);
nor U11320 (N_11320,N_5420,N_8881);
or U11321 (N_11321,N_5212,N_8029);
nor U11322 (N_11322,N_9697,N_5907);
xnor U11323 (N_11323,N_9357,N_8795);
xnor U11324 (N_11324,N_5335,N_7493);
nor U11325 (N_11325,N_6773,N_7476);
nor U11326 (N_11326,N_6521,N_8988);
nand U11327 (N_11327,N_6314,N_9174);
xnor U11328 (N_11328,N_6364,N_8618);
nand U11329 (N_11329,N_8925,N_6511);
and U11330 (N_11330,N_9675,N_6589);
nor U11331 (N_11331,N_8787,N_9631);
or U11332 (N_11332,N_9630,N_5471);
and U11333 (N_11333,N_9511,N_7491);
nand U11334 (N_11334,N_6372,N_6228);
nor U11335 (N_11335,N_8661,N_9444);
and U11336 (N_11336,N_9007,N_8974);
or U11337 (N_11337,N_5580,N_6767);
or U11338 (N_11338,N_7371,N_9771);
or U11339 (N_11339,N_6469,N_9723);
and U11340 (N_11340,N_5834,N_5475);
nor U11341 (N_11341,N_6729,N_6925);
xor U11342 (N_11342,N_9915,N_9010);
nand U11343 (N_11343,N_6249,N_7304);
xnor U11344 (N_11344,N_8810,N_6913);
and U11345 (N_11345,N_8061,N_7008);
xnor U11346 (N_11346,N_9450,N_6078);
or U11347 (N_11347,N_7728,N_8552);
and U11348 (N_11348,N_5298,N_9926);
nand U11349 (N_11349,N_8172,N_8458);
and U11350 (N_11350,N_8733,N_5096);
nor U11351 (N_11351,N_7803,N_7062);
nor U11352 (N_11352,N_9528,N_7393);
nand U11353 (N_11353,N_9100,N_8504);
nand U11354 (N_11354,N_7877,N_6145);
nand U11355 (N_11355,N_7308,N_8377);
nand U11356 (N_11356,N_6168,N_9253);
or U11357 (N_11357,N_8724,N_7400);
nand U11358 (N_11358,N_6640,N_9513);
xnor U11359 (N_11359,N_7208,N_8416);
or U11360 (N_11360,N_8281,N_7387);
nor U11361 (N_11361,N_5733,N_6683);
nand U11362 (N_11362,N_5048,N_7696);
or U11363 (N_11363,N_9760,N_5562);
and U11364 (N_11364,N_9788,N_9551);
nand U11365 (N_11365,N_5185,N_6900);
xor U11366 (N_11366,N_6287,N_7760);
and U11367 (N_11367,N_6098,N_7223);
or U11368 (N_11368,N_5554,N_8166);
or U11369 (N_11369,N_9319,N_5721);
nor U11370 (N_11370,N_5247,N_8676);
nand U11371 (N_11371,N_9189,N_7351);
xnor U11372 (N_11372,N_7534,N_7530);
nand U11373 (N_11373,N_8493,N_8941);
or U11374 (N_11374,N_9642,N_6478);
or U11375 (N_11375,N_9005,N_9508);
and U11376 (N_11376,N_5954,N_5012);
nand U11377 (N_11377,N_6246,N_8969);
nor U11378 (N_11378,N_7296,N_9828);
xor U11379 (N_11379,N_9032,N_5447);
or U11380 (N_11380,N_8171,N_8652);
nand U11381 (N_11381,N_7271,N_5839);
nor U11382 (N_11382,N_7959,N_9625);
nand U11383 (N_11383,N_9948,N_7916);
nor U11384 (N_11384,N_7027,N_7883);
or U11385 (N_11385,N_7819,N_6465);
xnor U11386 (N_11386,N_7326,N_6877);
xnor U11387 (N_11387,N_9322,N_9632);
nor U11388 (N_11388,N_8537,N_9682);
nand U11389 (N_11389,N_7924,N_8813);
and U11390 (N_11390,N_7990,N_8381);
and U11391 (N_11391,N_6526,N_8151);
or U11392 (N_11392,N_6580,N_5680);
and U11393 (N_11393,N_8131,N_6170);
nor U11394 (N_11394,N_8005,N_6751);
and U11395 (N_11395,N_7922,N_7825);
nor U11396 (N_11396,N_9334,N_8847);
or U11397 (N_11397,N_8714,N_9813);
nand U11398 (N_11398,N_7111,N_8110);
xnor U11399 (N_11399,N_6302,N_8511);
and U11400 (N_11400,N_9226,N_6029);
xor U11401 (N_11401,N_7632,N_6556);
xnor U11402 (N_11402,N_8905,N_6417);
or U11403 (N_11403,N_9852,N_7699);
nor U11404 (N_11404,N_8639,N_8738);
nor U11405 (N_11405,N_5697,N_9061);
and U11406 (N_11406,N_5410,N_9385);
and U11407 (N_11407,N_5681,N_6922);
and U11408 (N_11408,N_7507,N_9430);
xnor U11409 (N_11409,N_6059,N_9145);
nor U11410 (N_11410,N_6986,N_7225);
nand U11411 (N_11411,N_9960,N_6142);
and U11412 (N_11412,N_9423,N_6518);
and U11413 (N_11413,N_6319,N_8101);
or U11414 (N_11414,N_6993,N_8372);
or U11415 (N_11415,N_7655,N_9726);
nand U11416 (N_11416,N_5296,N_5102);
nand U11417 (N_11417,N_7519,N_9404);
and U11418 (N_11418,N_9851,N_6401);
nor U11419 (N_11419,N_7941,N_6816);
nor U11420 (N_11420,N_9307,N_7551);
and U11421 (N_11421,N_5800,N_9860);
and U11422 (N_11422,N_8011,N_5966);
nand U11423 (N_11423,N_8653,N_8671);
nor U11424 (N_11424,N_5464,N_8790);
and U11425 (N_11425,N_5122,N_6348);
and U11426 (N_11426,N_6449,N_9700);
or U11427 (N_11427,N_5430,N_9951);
xor U11428 (N_11428,N_8698,N_8578);
or U11429 (N_11429,N_5144,N_6649);
and U11430 (N_11430,N_9979,N_6716);
or U11431 (N_11431,N_7048,N_6819);
or U11432 (N_11432,N_6194,N_5920);
and U11433 (N_11433,N_7069,N_8599);
or U11434 (N_11434,N_8469,N_6065);
and U11435 (N_11435,N_7787,N_6030);
and U11436 (N_11436,N_5774,N_8975);
or U11437 (N_11437,N_5496,N_8140);
or U11438 (N_11438,N_5047,N_8892);
and U11439 (N_11439,N_8531,N_7194);
and U11440 (N_11440,N_6664,N_7747);
xor U11441 (N_11441,N_9308,N_7608);
or U11442 (N_11442,N_6025,N_6383);
or U11443 (N_11443,N_6966,N_7022);
nand U11444 (N_11444,N_5472,N_8866);
nor U11445 (N_11445,N_9055,N_5327);
and U11446 (N_11446,N_6851,N_6253);
nor U11447 (N_11447,N_6937,N_8126);
or U11448 (N_11448,N_6159,N_9966);
and U11449 (N_11449,N_8453,N_7328);
nand U11450 (N_11450,N_8651,N_8096);
or U11451 (N_11451,N_5855,N_7757);
or U11452 (N_11452,N_6811,N_7763);
nand U11453 (N_11453,N_9858,N_7583);
nor U11454 (N_11454,N_7177,N_8160);
nor U11455 (N_11455,N_7365,N_9289);
nor U11456 (N_11456,N_9657,N_9959);
or U11457 (N_11457,N_6265,N_5840);
nor U11458 (N_11458,N_9116,N_9442);
and U11459 (N_11459,N_9165,N_6233);
nor U11460 (N_11460,N_7282,N_5412);
nor U11461 (N_11461,N_5750,N_9753);
nand U11462 (N_11462,N_8711,N_6430);
or U11463 (N_11463,N_6046,N_7428);
and U11464 (N_11464,N_7838,N_8605);
xnor U11465 (N_11465,N_8829,N_5850);
nor U11466 (N_11466,N_5396,N_8053);
nor U11467 (N_11467,N_9741,N_9363);
and U11468 (N_11468,N_8828,N_8315);
nor U11469 (N_11469,N_8499,N_7182);
or U11470 (N_11470,N_8879,N_9376);
nor U11471 (N_11471,N_6295,N_8434);
or U11472 (N_11472,N_6464,N_9258);
or U11473 (N_11473,N_9169,N_7181);
or U11474 (N_11474,N_6591,N_5563);
xor U11475 (N_11475,N_7878,N_8267);
or U11476 (N_11476,N_8307,N_5923);
or U11477 (N_11477,N_6484,N_6201);
nand U11478 (N_11478,N_8571,N_6663);
nand U11479 (N_11479,N_6539,N_7277);
and U11480 (N_11480,N_9248,N_8923);
xnor U11481 (N_11481,N_9256,N_7745);
nand U11482 (N_11482,N_7200,N_9246);
or U11483 (N_11483,N_6471,N_7948);
nand U11484 (N_11484,N_8831,N_6094);
or U11485 (N_11485,N_9391,N_6325);
and U11486 (N_11486,N_6446,N_7204);
or U11487 (N_11487,N_8026,N_8051);
or U11488 (N_11488,N_7212,N_6238);
nand U11489 (N_11489,N_9512,N_8484);
nand U11490 (N_11490,N_5831,N_6105);
nor U11491 (N_11491,N_5507,N_7456);
or U11492 (N_11492,N_6486,N_7403);
nor U11493 (N_11493,N_6102,N_5257);
or U11494 (N_11494,N_6192,N_8399);
and U11495 (N_11495,N_5109,N_5848);
or U11496 (N_11496,N_8060,N_8164);
nor U11497 (N_11497,N_8198,N_5792);
or U11498 (N_11498,N_6531,N_7335);
or U11499 (N_11499,N_6362,N_6866);
nor U11500 (N_11500,N_7452,N_9291);
nand U11501 (N_11501,N_8116,N_5007);
nand U11502 (N_11502,N_8111,N_6614);
or U11503 (N_11503,N_6003,N_5497);
nand U11504 (N_11504,N_9352,N_6342);
and U11505 (N_11505,N_5829,N_8636);
xnor U11506 (N_11506,N_5462,N_6641);
and U11507 (N_11507,N_8722,N_5930);
and U11508 (N_11508,N_8614,N_9970);
or U11509 (N_11509,N_5748,N_9568);
or U11510 (N_11510,N_9162,N_6220);
nor U11511 (N_11511,N_6665,N_6581);
or U11512 (N_11512,N_6296,N_7730);
nor U11513 (N_11513,N_5206,N_5216);
and U11514 (N_11514,N_9608,N_6310);
or U11515 (N_11515,N_8390,N_7964);
and U11516 (N_11516,N_6601,N_5026);
nand U11517 (N_11517,N_8034,N_7601);
and U11518 (N_11518,N_8555,N_8496);
and U11519 (N_11519,N_8310,N_7220);
and U11520 (N_11520,N_6461,N_9362);
nand U11521 (N_11521,N_5052,N_8529);
and U11522 (N_11522,N_5402,N_6646);
nand U11523 (N_11523,N_5970,N_5336);
or U11524 (N_11524,N_7443,N_9396);
nor U11525 (N_11525,N_7518,N_9263);
nand U11526 (N_11526,N_9795,N_7324);
nor U11527 (N_11527,N_8580,N_9666);
or U11528 (N_11528,N_6987,N_5269);
nand U11529 (N_11529,N_5306,N_7982);
and U11530 (N_11530,N_8626,N_9275);
nor U11531 (N_11531,N_9767,N_8112);
and U11532 (N_11532,N_8328,N_7988);
and U11533 (N_11533,N_9685,N_5818);
nor U11534 (N_11534,N_6957,N_5202);
and U11535 (N_11535,N_7384,N_6357);
nor U11536 (N_11536,N_6017,N_8233);
nand U11537 (N_11537,N_5354,N_7333);
or U11538 (N_11538,N_8961,N_8731);
nand U11539 (N_11539,N_5780,N_6376);
nand U11540 (N_11540,N_5998,N_9638);
nor U11541 (N_11541,N_6452,N_5088);
nand U11542 (N_11542,N_7675,N_6275);
and U11543 (N_11543,N_7798,N_9870);
nand U11544 (N_11544,N_6028,N_8627);
and U11545 (N_11545,N_8207,N_9989);
or U11546 (N_11546,N_5316,N_6016);
xor U11547 (N_11547,N_9453,N_8084);
nand U11548 (N_11548,N_9958,N_7337);
nand U11549 (N_11549,N_9514,N_8479);
nand U11550 (N_11550,N_6056,N_5213);
xor U11551 (N_11551,N_9944,N_7607);
and U11552 (N_11552,N_8284,N_5355);
xnor U11553 (N_11553,N_7323,N_5118);
or U11554 (N_11554,N_6514,N_6948);
and U11555 (N_11555,N_8049,N_7356);
and U11556 (N_11556,N_7179,N_6668);
and U11557 (N_11557,N_8424,N_6884);
nand U11558 (N_11558,N_8968,N_5281);
and U11559 (N_11559,N_5658,N_8519);
xor U11560 (N_11560,N_9905,N_5942);
and U11561 (N_11561,N_6529,N_9335);
nor U11562 (N_11562,N_8196,N_7044);
and U11563 (N_11563,N_6498,N_8163);
or U11564 (N_11564,N_7201,N_7375);
or U11565 (N_11565,N_5357,N_9620);
xor U11566 (N_11566,N_8225,N_8910);
xor U11567 (N_11567,N_9709,N_5654);
or U11568 (N_11568,N_6701,N_9407);
or U11569 (N_11569,N_9536,N_8462);
and U11570 (N_11570,N_6218,N_5444);
or U11571 (N_11571,N_9496,N_6409);
nand U11572 (N_11572,N_8674,N_6007);
nor U11573 (N_11573,N_8756,N_7936);
and U11574 (N_11574,N_6923,N_7366);
or U11575 (N_11575,N_9607,N_7855);
or U11576 (N_11576,N_7758,N_9252);
or U11577 (N_11577,N_6091,N_5919);
or U11578 (N_11578,N_5673,N_8744);
nand U11579 (N_11579,N_5612,N_6499);
or U11580 (N_11580,N_8047,N_5989);
and U11581 (N_11581,N_6827,N_7020);
or U11582 (N_11582,N_5029,N_7853);
or U11583 (N_11583,N_8515,N_6421);
and U11584 (N_11584,N_5662,N_7370);
or U11585 (N_11585,N_5028,N_7363);
nand U11586 (N_11586,N_7742,N_6380);
and U11587 (N_11587,N_9876,N_8091);
or U11588 (N_11588,N_5492,N_6442);
or U11589 (N_11589,N_9126,N_9287);
or U11590 (N_11590,N_9235,N_5489);
and U11591 (N_11591,N_5891,N_5861);
and U11592 (N_11592,N_5557,N_8501);
xnor U11593 (N_11593,N_9879,N_5890);
and U11594 (N_11594,N_9783,N_5166);
xor U11595 (N_11595,N_5235,N_8353);
or U11596 (N_11596,N_8806,N_9899);
or U11597 (N_11597,N_9575,N_9023);
nor U11598 (N_11598,N_8367,N_7285);
and U11599 (N_11599,N_7789,N_5988);
nand U11600 (N_11600,N_5671,N_8326);
and U11601 (N_11601,N_6790,N_9083);
nor U11602 (N_11602,N_7405,N_7755);
nand U11603 (N_11603,N_5837,N_7736);
nand U11604 (N_11604,N_6587,N_6849);
nand U11605 (N_11605,N_5548,N_5155);
nor U11606 (N_11606,N_7837,N_8132);
and U11607 (N_11607,N_6126,N_7590);
or U11608 (N_11608,N_5739,N_8532);
xnor U11609 (N_11609,N_7965,N_6555);
or U11610 (N_11610,N_6048,N_5871);
or U11611 (N_11611,N_9836,N_9390);
and U11612 (N_11612,N_6907,N_5032);
nand U11613 (N_11613,N_8460,N_6351);
nand U11614 (N_11614,N_9035,N_7645);
nor U11615 (N_11615,N_9123,N_5468);
and U11616 (N_11616,N_9669,N_5556);
or U11617 (N_11617,N_7894,N_7652);
nor U11618 (N_11618,N_5383,N_5972);
nor U11619 (N_11619,N_7884,N_9696);
nand U11620 (N_11620,N_6243,N_8411);
nand U11621 (N_11621,N_5589,N_9482);
nand U11622 (N_11622,N_9928,N_5474);
or U11623 (N_11623,N_5686,N_8081);
or U11624 (N_11624,N_5370,N_7066);
and U11625 (N_11625,N_6069,N_9068);
or U11626 (N_11626,N_7176,N_7458);
nand U11627 (N_11627,N_8691,N_6672);
and U11628 (N_11628,N_6846,N_8687);
nor U11629 (N_11629,N_7278,N_7516);
xnor U11630 (N_11630,N_6603,N_7812);
or U11631 (N_11631,N_8186,N_7624);
and U11632 (N_11632,N_8874,N_6720);
and U11633 (N_11633,N_7025,N_5616);
nand U11634 (N_11634,N_9809,N_8155);
nor U11635 (N_11635,N_7252,N_7613);
nor U11636 (N_11636,N_9254,N_8788);
nor U11637 (N_11637,N_7594,N_6502);
nand U11638 (N_11638,N_9922,N_8226);
and U11639 (N_11639,N_5312,N_9473);
nor U11640 (N_11640,N_6350,N_7214);
nor U11641 (N_11641,N_5561,N_7265);
nor U11642 (N_11642,N_7875,N_5701);
nor U11643 (N_11643,N_8543,N_6563);
nor U11644 (N_11644,N_6515,N_5117);
or U11645 (N_11645,N_9687,N_6874);
xnor U11646 (N_11646,N_8134,N_8028);
and U11647 (N_11647,N_7839,N_8256);
nor U11648 (N_11648,N_6496,N_7488);
xnor U11649 (N_11649,N_8725,N_8398);
or U11650 (N_11650,N_8070,N_5740);
and U11651 (N_11651,N_7143,N_8264);
and U11652 (N_11652,N_6272,N_9920);
nand U11653 (N_11653,N_7733,N_7266);
nor U11654 (N_11654,N_6841,N_7690);
nand U11655 (N_11655,N_9883,N_8548);
nand U11656 (N_11656,N_7702,N_6005);
xnor U11657 (N_11657,N_7166,N_7054);
nor U11658 (N_11658,N_7005,N_9720);
and U11659 (N_11659,N_6070,N_8436);
or U11660 (N_11660,N_6836,N_8994);
nand U11661 (N_11661,N_8280,N_9204);
xor U11662 (N_11662,N_5467,N_5041);
xor U11663 (N_11663,N_6117,N_8144);
and U11664 (N_11664,N_8023,N_9893);
or U11665 (N_11665,N_9050,N_7017);
nand U11666 (N_11666,N_9080,N_6840);
xor U11667 (N_11667,N_5487,N_9326);
and U11668 (N_11668,N_9535,N_6470);
or U11669 (N_11669,N_5023,N_9422);
nor U11670 (N_11670,N_5845,N_9361);
nor U11671 (N_11671,N_7817,N_9133);
and U11672 (N_11672,N_6260,N_9678);
or U11673 (N_11673,N_9234,N_7635);
and U11674 (N_11674,N_6134,N_9599);
or U11675 (N_11675,N_6366,N_7432);
nand U11676 (N_11676,N_8082,N_7826);
or U11677 (N_11677,N_6917,N_8236);
nand U11678 (N_11678,N_5057,N_5997);
and U11679 (N_11679,N_5550,N_9402);
nor U11680 (N_11680,N_8579,N_5030);
nand U11681 (N_11681,N_8243,N_7814);
nand U11682 (N_11682,N_5584,N_6340);
nand U11683 (N_11683,N_9478,N_9093);
and U11684 (N_11684,N_5342,N_6053);
nor U11685 (N_11685,N_7694,N_9707);
and U11686 (N_11686,N_9995,N_7636);
or U11687 (N_11687,N_8471,N_6151);
and U11688 (N_11688,N_5393,N_9459);
nor U11689 (N_11689,N_5568,N_9161);
or U11690 (N_11690,N_7712,N_9058);
nor U11691 (N_11691,N_6712,N_7897);
or U11692 (N_11692,N_7362,N_9614);
and U11693 (N_11693,N_8949,N_9290);
xor U11694 (N_11694,N_9397,N_8235);
xnor U11695 (N_11695,N_9521,N_6206);
and U11696 (N_11696,N_9853,N_9822);
nor U11697 (N_11697,N_7698,N_9848);
nand U11698 (N_11698,N_8087,N_9556);
and U11699 (N_11699,N_7726,N_5211);
or U11700 (N_11700,N_6292,N_8203);
nor U11701 (N_11701,N_5479,N_5842);
xor U11702 (N_11702,N_9999,N_9012);
nand U11703 (N_11703,N_6650,N_6757);
or U11704 (N_11704,N_9730,N_6066);
and U11705 (N_11705,N_5034,N_5648);
xor U11706 (N_11706,N_7630,N_7537);
nor U11707 (N_11707,N_6144,N_5601);
or U11708 (N_11708,N_7653,N_5488);
and U11709 (N_11709,N_9215,N_8948);
nor U11710 (N_11710,N_5790,N_5075);
nor U11711 (N_11711,N_6113,N_5481);
or U11712 (N_11712,N_8272,N_6636);
xnor U11713 (N_11713,N_8173,N_5902);
and U11714 (N_11714,N_7346,N_5237);
or U11715 (N_11715,N_6554,N_6859);
nor U11716 (N_11716,N_6545,N_7872);
or U11717 (N_11717,N_8075,N_7408);
or U11718 (N_11718,N_8832,N_7433);
nand U11719 (N_11719,N_9862,N_5529);
or U11720 (N_11720,N_9414,N_9076);
or U11721 (N_11721,N_9932,N_8825);
or U11722 (N_11722,N_6127,N_5833);
or U11723 (N_11723,N_9600,N_5595);
nand U11724 (N_11724,N_7084,N_7722);
nor U11725 (N_11725,N_6570,N_6358);
and U11726 (N_11726,N_8630,N_5092);
and U11727 (N_11727,N_7178,N_7302);
or U11728 (N_11728,N_8400,N_5094);
nand U11729 (N_11729,N_8015,N_5757);
xnor U11730 (N_11730,N_9349,N_8809);
nand U11731 (N_11731,N_6779,N_9229);
xor U11732 (N_11732,N_6182,N_9483);
nand U11733 (N_11733,N_7863,N_7286);
or U11734 (N_11734,N_7522,N_9595);
nand U11735 (N_11735,N_9084,N_6864);
or U11736 (N_11736,N_8357,N_6985);
nand U11737 (N_11737,N_7281,N_9637);
nor U11738 (N_11738,N_8641,N_7035);
and U11739 (N_11739,N_9120,N_7485);
or U11740 (N_11740,N_8352,N_8820);
and U11741 (N_11741,N_7288,N_8863);
and U11742 (N_11742,N_6321,N_8232);
nand U11743 (N_11743,N_8978,N_7430);
and U11744 (N_11744,N_6670,N_9564);
nand U11745 (N_11745,N_9401,N_9013);
xor U11746 (N_11746,N_9940,N_9082);
nand U11747 (N_11747,N_7718,N_7912);
nor U11748 (N_11748,N_6690,N_9789);
nand U11749 (N_11749,N_8092,N_5261);
nor U11750 (N_11750,N_7203,N_7088);
nand U11751 (N_11751,N_9739,N_6459);
nor U11752 (N_11752,N_9942,N_6308);
nor U11753 (N_11753,N_5440,N_9612);
or U11754 (N_11754,N_6949,N_9872);
nand U11755 (N_11755,N_6312,N_6229);
and U11756 (N_11756,N_6507,N_5341);
nor U11757 (N_11757,N_5369,N_9971);
and U11758 (N_11758,N_7240,N_6660);
or U11759 (N_11759,N_5574,N_5719);
and U11760 (N_11760,N_5121,N_7603);
nand U11761 (N_11761,N_6853,N_7406);
or U11762 (N_11762,N_9439,N_7188);
nor U11763 (N_11763,N_6074,N_5076);
nand U11764 (N_11764,N_7087,N_7100);
nand U11765 (N_11765,N_8576,N_6548);
and U11766 (N_11766,N_7379,N_5963);
and U11767 (N_11767,N_7778,N_9718);
and U11768 (N_11768,N_6610,N_8181);
xor U11769 (N_11769,N_9553,N_8215);
or U11770 (N_11770,N_7497,N_9157);
and U11771 (N_11771,N_6675,N_9907);
nor U11772 (N_11772,N_8710,N_9344);
xnor U11773 (N_11773,N_5751,N_7719);
and U11774 (N_11774,N_6093,N_8237);
nand U11775 (N_11775,N_9173,N_5053);
nand U11776 (N_11776,N_7500,N_5991);
and U11777 (N_11777,N_9547,N_5356);
and U11778 (N_11778,N_8143,N_9885);
nand U11779 (N_11779,N_9043,N_6188);
nand U11780 (N_11780,N_8583,N_5398);
or U11781 (N_11781,N_7943,N_7343);
or U11782 (N_11782,N_9337,N_8234);
and U11783 (N_11783,N_9003,N_8193);
and U11784 (N_11784,N_9738,N_8707);
and U11785 (N_11785,N_6278,N_8039);
and U11786 (N_11786,N_8249,N_6402);
xor U11787 (N_11787,N_9617,N_5810);
or U11788 (N_11788,N_6713,N_9305);
nand U11789 (N_11789,N_8984,N_8934);
nor U11790 (N_11790,N_5480,N_5961);
or U11791 (N_11791,N_9537,N_6335);
or U11792 (N_11792,N_8206,N_6658);
nor U11793 (N_11793,N_8410,N_9821);
nand U11794 (N_11794,N_6172,N_7978);
and U11795 (N_11795,N_5091,N_5072);
nand U11796 (N_11796,N_8396,N_8637);
nand U11797 (N_11797,N_8970,N_6534);
nor U11798 (N_11798,N_9503,N_6685);
xnor U11799 (N_11799,N_5239,N_7043);
nor U11800 (N_11800,N_7969,N_8610);
or U11801 (N_11801,N_5411,N_6564);
nand U11802 (N_11802,N_6297,N_9297);
nor U11803 (N_11803,N_7420,N_7808);
and U11804 (N_11804,N_5905,N_7243);
nor U11805 (N_11805,N_7927,N_5604);
nand U11806 (N_11806,N_6181,N_8582);
or U11807 (N_11807,N_8337,N_9671);
or U11808 (N_11808,N_6639,N_8122);
nor U11809 (N_11809,N_7256,N_9276);
nand U11810 (N_11810,N_6774,N_7961);
or U11811 (N_11811,N_9047,N_5642);
nand U11812 (N_11812,N_7526,N_5884);
nor U11813 (N_11813,N_8990,N_5340);
nand U11814 (N_11814,N_6360,N_9784);
and U11815 (N_11815,N_6994,N_7942);
xor U11816 (N_11816,N_9713,N_8721);
or U11817 (N_11817,N_7459,N_9779);
and U11818 (N_11818,N_5978,N_7542);
nor U11819 (N_11819,N_9296,N_9479);
nor U11820 (N_11820,N_6961,N_8492);
xnor U11821 (N_11821,N_5880,N_5992);
nand U11822 (N_11822,N_6487,N_8660);
nor U11823 (N_11823,N_9533,N_9611);
or U11824 (N_11824,N_8869,N_7159);
and U11825 (N_11825,N_7236,N_5555);
nor U11826 (N_11826,N_9449,N_5113);
and U11827 (N_11827,N_7382,N_5645);
or U11828 (N_11828,N_8170,N_5284);
nor U11829 (N_11829,N_6298,N_8667);
or U11830 (N_11830,N_6694,N_7228);
and U11831 (N_11831,N_5169,N_7081);
or U11832 (N_11832,N_5017,N_5242);
xnor U11833 (N_11833,N_7114,N_5610);
nor U11834 (N_11834,N_9016,N_7039);
or U11835 (N_11835,N_8664,N_7085);
xor U11836 (N_11836,N_9156,N_5863);
and U11837 (N_11837,N_5451,N_9980);
nor U11838 (N_11838,N_8094,N_6996);
nand U11839 (N_11839,N_7967,N_7994);
and U11840 (N_11840,N_6114,N_6403);
nor U11841 (N_11841,N_6111,N_5754);
or U11842 (N_11842,N_9804,N_5732);
nand U11843 (N_11843,N_5116,N_7963);
nor U11844 (N_11844,N_9731,N_7647);
nand U11845 (N_11845,N_5069,N_9304);
and U11846 (N_11846,N_5175,N_6943);
and U11847 (N_11847,N_5827,N_5190);
nand U11848 (N_11848,N_5664,N_7845);
nor U11849 (N_11849,N_8595,N_6388);
nand U11850 (N_11850,N_9558,N_7320);
and U11851 (N_11851,N_8379,N_8009);
or U11852 (N_11852,N_6733,N_7042);
nor U11853 (N_11853,N_5771,N_5119);
and U11854 (N_11854,N_8394,N_8291);
nand U11855 (N_11855,N_8387,N_6047);
nor U11856 (N_11856,N_8561,N_5764);
and U11857 (N_11857,N_8929,N_6191);
nand U11858 (N_11858,N_9471,N_9820);
or U11859 (N_11859,N_8068,N_9104);
or U11860 (N_11860,N_6058,N_8165);
xnor U11861 (N_11861,N_5843,N_5391);
xnor U11862 (N_11862,N_6186,N_7139);
nor U11863 (N_11863,N_6590,N_8935);
nor U11864 (N_11864,N_5099,N_6179);
or U11865 (N_11865,N_8870,N_6894);
nor U11866 (N_11866,N_9451,N_5246);
and U11867 (N_11867,N_5647,N_8750);
nor U11868 (N_11868,N_5623,N_8020);
nor U11869 (N_11869,N_8254,N_5149);
and U11870 (N_11870,N_8963,N_8737);
or U11871 (N_11871,N_6483,N_6684);
nor U11872 (N_11872,N_9833,N_5377);
and U11873 (N_11873,N_8279,N_8696);
nor U11874 (N_11874,N_7689,N_7842);
nand U11875 (N_11875,N_8799,N_5128);
and U11876 (N_11876,N_6798,N_5160);
or U11877 (N_11877,N_8440,N_8441);
nand U11878 (N_11878,N_5127,N_9947);
nor U11879 (N_11879,N_8255,N_9856);
and U11880 (N_11880,N_7995,N_7619);
nand U11881 (N_11881,N_7566,N_8167);
nor U11882 (N_11882,N_5071,N_5164);
nand U11883 (N_11883,N_6960,N_8776);
nor U11884 (N_11884,N_6978,N_6352);
and U11885 (N_11885,N_5767,N_7914);
and U11886 (N_11886,N_5491,N_8590);
and U11887 (N_11887,N_7654,N_9135);
or U11888 (N_11888,N_9663,N_7687);
nor U11889 (N_11889,N_5020,N_9597);
and U11890 (N_11890,N_5744,N_5741);
nand U11891 (N_11891,N_9217,N_6891);
and U11892 (N_11892,N_7773,N_6395);
or U11893 (N_11893,N_9690,N_5945);
xor U11894 (N_11894,N_6871,N_5626);
or U11895 (N_11895,N_7996,N_5303);
and U11896 (N_11896,N_9205,N_5217);
and U11897 (N_11897,N_8347,N_9652);
nor U11898 (N_11898,N_6755,N_7684);
nand U11899 (N_11899,N_9066,N_6506);
and U11900 (N_11900,N_6740,N_7482);
nor U11901 (N_11901,N_6410,N_9137);
and U11902 (N_11902,N_5138,N_5176);
nor U11903 (N_11903,N_9964,N_5515);
and U11904 (N_11904,N_6063,N_5142);
xor U11905 (N_11905,N_7572,N_8983);
nor U11906 (N_11906,N_7552,N_9832);
and U11907 (N_11907,N_7511,N_6379);
or U11908 (N_11908,N_9847,N_8640);
and U11909 (N_11909,N_8489,N_9618);
or U11910 (N_11910,N_5187,N_7918);
nor U11911 (N_11911,N_7593,N_9615);
and U11912 (N_11912,N_5896,N_8517);
nor U11913 (N_11913,N_5990,N_8902);
nor U11914 (N_11914,N_6480,N_5147);
nand U11915 (N_11915,N_9143,N_8414);
nor U11916 (N_11916,N_9481,N_9432);
or U11917 (N_11917,N_7195,N_9542);
or U11918 (N_11918,N_5414,N_8959);
and U11919 (N_11919,N_6963,N_7625);
nand U11920 (N_11920,N_7338,N_8395);
nor U11921 (N_11921,N_7898,N_8556);
nor U11922 (N_11922,N_6878,N_6577);
and U11923 (N_11923,N_8294,N_5528);
xnor U11924 (N_11924,N_5698,N_7710);
xnor U11925 (N_11925,N_6766,N_7251);
xnor U11926 (N_11926,N_9644,N_7554);
nand U11927 (N_11927,N_5152,N_5649);
or U11928 (N_11928,N_9377,N_9070);
or U11929 (N_11929,N_6645,N_7399);
nor U11930 (N_11930,N_9497,N_5115);
or U11931 (N_11931,N_5418,N_6489);
and U11932 (N_11932,N_9015,N_8772);
and U11933 (N_11933,N_5244,N_5856);
xnor U11934 (N_11934,N_8904,N_8316);
nand U11935 (N_11935,N_6898,N_6327);
xnor U11936 (N_11936,N_7680,N_6510);
or U11937 (N_11937,N_6955,N_9062);
and U11938 (N_11938,N_7202,N_7469);
and U11939 (N_11939,N_6786,N_5477);
nand U11940 (N_11940,N_6396,N_8540);
nor U11941 (N_11941,N_9990,N_6661);
or U11942 (N_11942,N_8269,N_6727);
or U11943 (N_11943,N_7574,N_9969);
and U11944 (N_11944,N_8223,N_6856);
and U11945 (N_11945,N_8759,N_8841);
nand U11946 (N_11946,N_5841,N_5802);
nor U11947 (N_11947,N_8319,N_6998);
nor U11948 (N_11948,N_5725,N_8886);
or U11949 (N_11949,N_5390,N_6553);
or U11950 (N_11950,N_7648,N_7772);
nand U11951 (N_11951,N_6207,N_8221);
xnor U11952 (N_11952,N_8560,N_9613);
nand U11953 (N_11953,N_7911,N_7385);
and U11954 (N_11954,N_8766,N_9443);
xnor U11955 (N_11955,N_8802,N_8038);
xor U11956 (N_11956,N_6808,N_9065);
or U11957 (N_11957,N_7300,N_7191);
nand U11958 (N_11958,N_9130,N_9797);
or U11959 (N_11959,N_7539,N_5423);
nor U11960 (N_11960,N_5747,N_7896);
or U11961 (N_11961,N_5917,N_6976);
nand U11962 (N_11962,N_8856,N_5234);
or U11963 (N_11963,N_9878,N_6010);
and U11964 (N_11964,N_7307,N_8329);
and U11965 (N_11965,N_6666,N_6734);
nand U11966 (N_11966,N_8312,N_7173);
nor U11967 (N_11967,N_8956,N_5438);
and U11968 (N_11968,N_6014,N_9069);
nor U11969 (N_11969,N_6951,N_9714);
nor U11970 (N_11970,N_7146,N_7123);
nor U11971 (N_11971,N_5241,N_7535);
nand U11972 (N_11972,N_5599,N_9674);
and U11973 (N_11973,N_9844,N_5746);
and U11974 (N_11974,N_6204,N_9589);
or U11975 (N_11975,N_6439,N_9431);
nor U11976 (N_11976,N_8150,N_5641);
or U11977 (N_11977,N_8389,N_8265);
nand U11978 (N_11978,N_6210,N_9122);
and U11979 (N_11979,N_7095,N_9574);
nand U11980 (N_11980,N_9692,N_6451);
nand U11981 (N_11981,N_7231,N_8008);
nand U11982 (N_11982,N_7099,N_6627);
nand U11983 (N_11983,N_5359,N_5070);
and U11984 (N_11984,N_7550,N_7697);
nor U11985 (N_11985,N_5653,N_5522);
or U11986 (N_11986,N_8058,N_8985);
nor U11987 (N_11987,N_6476,N_8176);
nand U11988 (N_11988,N_9426,N_6865);
and U11989 (N_11989,N_6326,N_7683);
nor U11990 (N_11990,N_7589,N_8174);
or U11991 (N_11991,N_5114,N_5569);
or U11992 (N_11992,N_5956,N_7717);
nor U11993 (N_11993,N_7999,N_8100);
nand U11994 (N_11994,N_9792,N_9193);
or U11995 (N_11995,N_8734,N_8521);
nor U11996 (N_11996,N_5832,N_5278);
nand U11997 (N_11997,N_5918,N_6303);
and U11998 (N_11998,N_7904,N_7676);
and U11999 (N_11999,N_8325,N_8046);
nor U12000 (N_12000,N_9909,N_6787);
nor U12001 (N_12001,N_5074,N_8940);
nor U12002 (N_12002,N_5541,N_9092);
nor U12003 (N_12003,N_8632,N_8686);
nand U12004 (N_12004,N_8321,N_9790);
and U12005 (N_12005,N_5881,N_5093);
and U12006 (N_12006,N_8991,N_6068);
or U12007 (N_12007,N_7263,N_7749);
and U12008 (N_12008,N_8512,N_8987);
nor U12009 (N_12009,N_7234,N_7306);
nand U12010 (N_12010,N_5323,N_7174);
nor U12011 (N_12011,N_9742,N_9710);
nor U12012 (N_12012,N_6703,N_9046);
and U12013 (N_12013,N_9071,N_8509);
nand U12014 (N_12014,N_5593,N_9803);
and U12015 (N_12015,N_8551,N_9098);
or U12016 (N_12016,N_8861,N_8370);
nand U12017 (N_12017,N_8080,N_8197);
and U12018 (N_12018,N_6969,N_7858);
nand U12019 (N_12019,N_7774,N_6845);
nor U12020 (N_12020,N_7576,N_6778);
xnor U12021 (N_12021,N_9544,N_5851);
nor U12022 (N_12022,N_5794,N_5352);
nor U12023 (N_12023,N_8937,N_5060);
and U12024 (N_12024,N_5387,N_7805);
or U12025 (N_12025,N_8010,N_8677);
nor U12026 (N_12026,N_5255,N_5588);
and U12027 (N_12027,N_9346,N_9317);
nor U12028 (N_12028,N_9695,N_7828);
nor U12029 (N_12029,N_9522,N_8958);
nor U12030 (N_12030,N_6975,N_9113);
nand U12031 (N_12031,N_7901,N_5214);
and U12032 (N_12032,N_8488,N_8655);
or U12033 (N_12033,N_6381,N_6077);
xnor U12034 (N_12034,N_7870,N_7792);
and U12035 (N_12035,N_9237,N_5621);
and U12036 (N_12036,N_7340,N_8608);
nor U12037 (N_12037,N_9382,N_6313);
xor U12038 (N_12038,N_9743,N_6019);
xor U12039 (N_12039,N_9499,N_9838);
nand U12040 (N_12040,N_8992,N_8678);
and U12041 (N_12041,N_6140,N_7245);
nor U12042 (N_12042,N_8533,N_6927);
and U12043 (N_12043,N_6903,N_6008);
nand U12044 (N_12044,N_9881,N_7130);
nand U12045 (N_12045,N_8210,N_6956);
nand U12046 (N_12046,N_8634,N_8936);
nand U12047 (N_12047,N_8883,N_6373);
and U12048 (N_12048,N_6896,N_9004);
nand U12049 (N_12049,N_7796,N_8067);
and U12050 (N_12050,N_6101,N_6807);
or U12051 (N_12051,N_9724,N_7260);
nand U12052 (N_12052,N_9051,N_5358);
and U12053 (N_12053,N_8720,N_5339);
and U12054 (N_12054,N_5854,N_8821);
nor U12055 (N_12055,N_6749,N_6815);
xor U12056 (N_12056,N_7218,N_8098);
nor U12057 (N_12057,N_8751,N_9901);
nor U12058 (N_12058,N_5262,N_5499);
nor U12059 (N_12059,N_7484,N_9555);
or U12060 (N_12060,N_9529,N_8606);
nor U12061 (N_12061,N_9461,N_5163);
nor U12062 (N_12062,N_5267,N_7144);
and U12063 (N_12063,N_6328,N_7944);
or U12064 (N_12064,N_7374,N_9984);
and U12065 (N_12065,N_5348,N_8596);
nor U12066 (N_12066,N_7641,N_7426);
xnor U12067 (N_12067,N_5709,N_8433);
or U12068 (N_12068,N_9561,N_5666);
xor U12069 (N_12069,N_7353,N_6374);
or U12070 (N_12070,N_5579,N_9950);
nor U12071 (N_12071,N_9800,N_9573);
and U12072 (N_12072,N_5311,N_7981);
or U12073 (N_12073,N_7424,N_5689);
or U12074 (N_12074,N_5545,N_7962);
nand U12075 (N_12075,N_7611,N_9769);
nor U12076 (N_12076,N_9501,N_6909);
nor U12077 (N_12077,N_9477,N_7501);
nor U12078 (N_12078,N_8189,N_8873);
nand U12079 (N_12079,N_7640,N_9228);
or U12080 (N_12080,N_7295,N_9064);
and U12081 (N_12081,N_9865,N_5277);
and U12082 (N_12082,N_6634,N_8906);
and U12083 (N_12083,N_9526,N_8459);
or U12084 (N_12084,N_8261,N_9722);
and U12085 (N_12085,N_6565,N_6597);
xnor U12086 (N_12086,N_5518,N_7685);
nor U12087 (N_12087,N_6460,N_7949);
and U12088 (N_12088,N_8021,N_9826);
and U12089 (N_12089,N_8995,N_8485);
or U12090 (N_12090,N_6780,N_9044);
and U12091 (N_12091,N_6453,N_8872);
and U12092 (N_12092,N_5024,N_9364);
nor U12093 (N_12093,N_9428,N_9988);
and U12094 (N_12094,N_6659,N_7189);
nor U12095 (N_12095,N_8361,N_9244);
nor U12096 (N_12096,N_9270,N_6414);
or U12097 (N_12097,N_6205,N_7873);
nor U12098 (N_12098,N_7827,N_6730);
and U12099 (N_12099,N_8214,N_7449);
nand U12100 (N_12100,N_9114,N_9197);
and U12101 (N_12101,N_7001,N_6166);
and U12102 (N_12102,N_7931,N_5067);
and U12103 (N_12103,N_8245,N_8672);
and U12104 (N_12104,N_7841,N_8808);
nand U12105 (N_12105,N_9343,N_8798);
nand U12106 (N_12106,N_6146,N_5205);
xnor U12107 (N_12107,N_6171,N_7954);
nor U12108 (N_12108,N_8922,N_7811);
or U12109 (N_12109,N_5422,N_7905);
nand U12110 (N_12110,N_9576,N_6450);
and U12111 (N_12111,N_8002,N_6262);
nor U12112 (N_12112,N_9839,N_8673);
nand U12113 (N_12113,N_7913,N_6754);
xor U12114 (N_12114,N_8429,N_5107);
and U12115 (N_12115,N_7287,N_6305);
and U12116 (N_12116,N_7930,N_8817);
or U12117 (N_12117,N_8248,N_5156);
nand U12118 (N_12118,N_7440,N_9280);
or U12119 (N_12119,N_8273,N_8617);
and U12120 (N_12120,N_8045,N_6224);
nand U12121 (N_12121,N_6445,N_5590);
or U12122 (N_12122,N_8076,N_9587);
nor U12123 (N_12123,N_5639,N_8927);
nor U12124 (N_12124,N_9462,N_9680);
nor U12125 (N_12125,N_6743,N_5427);
or U12126 (N_12126,N_5101,N_5442);
nor U12127 (N_12127,N_7536,N_5098);
and U12128 (N_12128,N_6600,N_5409);
nand U12129 (N_12129,N_6517,N_6261);
xor U12130 (N_12130,N_8304,N_7743);
nor U12131 (N_12131,N_6928,N_7193);
or U12132 (N_12132,N_6607,N_8878);
and U12133 (N_12133,N_8199,N_8184);
nand U12134 (N_12134,N_9011,N_5045);
nand U12135 (N_12135,N_9571,N_9225);
nand U12136 (N_12136,N_5505,N_8230);
nand U12137 (N_12137,N_6573,N_6203);
or U12138 (N_12138,N_6568,N_9108);
nor U12139 (N_12139,N_6020,N_7739);
xor U12140 (N_12140,N_6444,N_6270);
and U12141 (N_12141,N_7859,N_5823);
and U12142 (N_12142,N_8327,N_9073);
or U12143 (N_12143,N_8704,N_9099);
nand U12144 (N_12144,N_7492,N_5294);
nand U12145 (N_12145,N_9367,N_5897);
nor U12146 (N_12146,N_7383,N_8388);
or U12147 (N_12147,N_9292,N_6455);
or U12148 (N_12148,N_8363,N_7532);
nor U12149 (N_12149,N_7467,N_8300);
xnor U12150 (N_12150,N_5224,N_7738);
and U12151 (N_12151,N_9531,N_6289);
nand U12152 (N_12152,N_6195,N_5876);
nor U12153 (N_12153,N_6908,N_5540);
nor U12154 (N_12154,N_5652,N_9936);
and U12155 (N_12155,N_5154,N_5603);
nand U12156 (N_12156,N_7016,N_9897);
nand U12157 (N_12157,N_8442,N_5959);
nand U12158 (N_12158,N_8356,N_5537);
and U12159 (N_12159,N_8569,N_5968);
and U12160 (N_12160,N_9151,N_7582);
and U12161 (N_12161,N_7206,N_5614);
or U12162 (N_12162,N_8964,N_9903);
or U12163 (N_12163,N_6015,N_5799);
or U12164 (N_12164,N_8289,N_8331);
or U12165 (N_12165,N_6334,N_9543);
and U12166 (N_12166,N_9469,N_9751);
nor U12167 (N_12167,N_5533,N_9968);
and U12168 (N_12168,N_6991,N_7317);
nor U12169 (N_12169,N_9000,N_9368);
nand U12170 (N_12170,N_6523,N_5895);
nor U12171 (N_12171,N_8778,N_7830);
and U12172 (N_12172,N_9498,N_6760);
nand U12173 (N_12173,N_8615,N_8212);
nor U12174 (N_12174,N_9765,N_6736);
nand U12175 (N_12175,N_5386,N_6337);
xor U12176 (N_12176,N_8065,N_7298);
nor U12177 (N_12177,N_7561,N_7021);
nor U12178 (N_12178,N_7359,N_9645);
or U12179 (N_12179,N_7857,N_7823);
and U12180 (N_12180,N_7451,N_9579);
or U12181 (N_12181,N_5315,N_9941);
nor U12182 (N_12182,N_6473,N_9441);
nand U12183 (N_12183,N_6680,N_9562);
nand U12184 (N_12184,N_9153,N_8169);
nor U12185 (N_12185,N_6304,N_8700);
and U12186 (N_12186,N_5103,N_9240);
nor U12187 (N_12187,N_5033,N_6525);
nand U12188 (N_12188,N_8681,N_7649);
nor U12189 (N_12189,N_6983,N_6095);
nand U12190 (N_12190,N_5253,N_9953);
nand U12191 (N_12191,N_9896,N_7012);
xor U12192 (N_12192,N_7529,N_7004);
nand U12193 (N_12193,N_8945,N_6055);
and U12194 (N_12194,N_8088,N_9017);
nand U12195 (N_12195,N_5551,N_5864);
nor U12196 (N_12196,N_9052,N_8743);
xor U12197 (N_12197,N_8095,N_9019);
xor U12198 (N_12198,N_9022,N_9333);
xnor U12199 (N_12199,N_9059,N_8649);
and U12200 (N_12200,N_7414,N_8575);
xnor U12201 (N_12201,N_8097,N_6882);
xnor U12202 (N_12202,N_8900,N_5953);
xnor U12203 (N_12203,N_5995,N_5100);
or U12204 (N_12204,N_7327,N_8894);
nor U12205 (N_12205,N_5912,N_7832);
or U12206 (N_12206,N_7708,N_7581);
or U12207 (N_12207,N_5828,N_5432);
and U12208 (N_12208,N_7893,N_9102);
nor U12209 (N_12209,N_7119,N_8346);
nand U12210 (N_12210,N_8763,N_6609);
or U12211 (N_12211,N_5782,N_6137);
nor U12212 (N_12212,N_5575,N_8620);
nand U12213 (N_12213,N_6119,N_8350);
nand U12214 (N_12214,N_7148,N_7614);
and U12215 (N_12215,N_7795,N_8784);
nand U12216 (N_12216,N_7974,N_6033);
nand U12217 (N_12217,N_7478,N_9283);
nor U12218 (N_12218,N_9001,N_5558);
and U12219 (N_12219,N_7935,N_9823);
nor U12220 (N_12220,N_6984,N_6738);
nor U12221 (N_12221,N_5470,N_9485);
nor U12222 (N_12222,N_9673,N_9727);
and U12223 (N_12223,N_9117,N_8546);
and U12224 (N_12224,N_8149,N_5692);
and U12225 (N_12225,N_6622,N_5328);
or U12226 (N_12226,N_6947,N_6883);
nand U12227 (N_12227,N_8423,N_8177);
and U12228 (N_12228,N_6198,N_7120);
nor U12229 (N_12229,N_6783,N_7055);
nor U12230 (N_12230,N_7137,N_8195);
nand U12231 (N_12231,N_9877,N_5266);
nor U12232 (N_12232,N_7966,N_5181);
xor U12233 (N_12233,N_5813,N_8716);
or U12234 (N_12234,N_5208,N_6412);
xnor U12235 (N_12235,N_5139,N_8570);
nor U12236 (N_12236,N_5618,N_9395);
or U12237 (N_12237,N_6834,N_6839);
nand U12238 (N_12238,N_6962,N_7851);
or U12239 (N_12239,N_8670,N_5079);
nor U12240 (N_12240,N_9030,N_8413);
nand U12241 (N_12241,N_8465,N_5916);
nor U12242 (N_12242,N_9987,N_9646);
nand U12243 (N_12243,N_9890,N_6890);
nor U12244 (N_12244,N_5543,N_8500);
nand U12245 (N_12245,N_9927,N_5287);
nand U12246 (N_12246,N_5104,N_6398);
and U12247 (N_12247,N_5811,N_9603);
or U12248 (N_12248,N_8354,N_9949);
xor U12249 (N_12249,N_9785,N_5824);
xnor U12250 (N_12250,N_5962,N_9419);
nor U12251 (N_12251,N_6057,N_5394);
and U12252 (N_12252,N_6631,N_9698);
xnor U12253 (N_12253,N_9974,N_9917);
or U12254 (N_12254,N_5384,N_9937);
or U12255 (N_12255,N_5324,N_5996);
or U12256 (N_12256,N_5566,N_8638);
and U12257 (N_12257,N_8868,N_5909);
nor U12258 (N_12258,N_5665,N_9039);
or U12259 (N_12259,N_7431,N_5331);
nand U12260 (N_12260,N_8063,N_9049);
nor U12261 (N_12261,N_6354,N_9009);
nand U12262 (N_12262,N_8263,N_9078);
and U12263 (N_12263,N_8855,N_9772);
nor U12264 (N_12264,N_6893,N_7616);
and U12265 (N_12265,N_7071,N_9776);
or U12266 (N_12266,N_7261,N_8542);
nand U12267 (N_12267,N_9525,N_6530);
nor U12268 (N_12268,N_6250,N_8428);
nand U12269 (N_12269,N_8695,N_9264);
nor U12270 (N_12270,N_8880,N_8761);
nand U12271 (N_12271,N_6167,N_8727);
nor U12272 (N_12272,N_5965,N_9366);
and U12273 (N_12273,N_9604,N_9211);
and U12274 (N_12274,N_8048,N_9266);
or U12275 (N_12275,N_6332,N_8188);
or U12276 (N_12276,N_5706,N_5273);
nor U12277 (N_12277,N_7199,N_6623);
xor U12278 (N_12278,N_9910,N_5760);
or U12279 (N_12279,N_7498,N_6217);
xor U12280 (N_12280,N_9965,N_8845);
or U12281 (N_12281,N_5184,N_6965);
nand U12282 (N_12282,N_5784,N_8139);
and U12283 (N_12283,N_9053,N_5145);
and U12284 (N_12284,N_8741,N_9298);
nand U12285 (N_12285,N_9380,N_9216);
nand U12286 (N_12286,N_5089,N_5973);
xnor U12287 (N_12287,N_6571,N_5299);
nor U12288 (N_12288,N_8976,N_8178);
nor U12289 (N_12289,N_9309,N_5428);
nand U12290 (N_12290,N_5703,N_7160);
or U12291 (N_12291,N_7634,N_7175);
nor U12292 (N_12292,N_7235,N_7727);
nor U12293 (N_12293,N_8385,N_5204);
and U12294 (N_12294,N_8826,N_7818);
nand U12295 (N_12295,N_9859,N_9097);
xnor U12296 (N_12296,N_7275,N_7681);
nand U12297 (N_12297,N_9569,N_8119);
nor U12298 (N_12298,N_5847,N_8409);
and U12299 (N_12299,N_8586,N_5148);
nand U12300 (N_12300,N_7847,N_7059);
and U12301 (N_12301,N_6551,N_8402);
nor U12302 (N_12302,N_6501,N_8368);
nor U12303 (N_12303,N_9566,N_9359);
and U12304 (N_12304,N_8814,N_5958);
and U12305 (N_12305,N_8418,N_5495);
nor U12306 (N_12306,N_8373,N_9340);
nand U12307 (N_12307,N_6637,N_8146);
nor U12308 (N_12308,N_9583,N_8662);
or U12309 (N_12309,N_8290,N_9433);
and U12310 (N_12310,N_8728,N_9027);
nor U12311 (N_12311,N_6583,N_5180);
or U12312 (N_12312,N_6887,N_6516);
or U12313 (N_12313,N_7474,N_8588);
and U12314 (N_12314,N_9957,N_9916);
nand U12315 (N_12315,N_6124,N_7127);
or U12316 (N_12316,N_7471,N_7621);
and U12317 (N_12317,N_9991,N_5006);
and U12318 (N_12318,N_5252,N_6861);
or U12319 (N_12319,N_5392,N_7711);
nand U12320 (N_12320,N_7509,N_6940);
nor U12321 (N_12321,N_7142,N_7829);
or U12322 (N_12322,N_5272,N_5526);
nand U12323 (N_12323,N_9184,N_9233);
or U12324 (N_12324,N_6158,N_7715);
nor U12325 (N_12325,N_7835,N_8631);
and U12326 (N_12326,N_7843,N_7448);
or U12327 (N_12327,N_8472,N_7734);
nor U12328 (N_12328,N_9740,N_9128);
xnor U12329 (N_12329,N_8942,N_9578);
nand U12330 (N_12330,N_6202,N_5974);
or U12331 (N_12331,N_8162,N_8839);
nor U12332 (N_12332,N_6586,N_9912);
nor U12333 (N_12333,N_8222,N_6386);
or U12334 (N_12334,N_8159,N_5084);
nand U12335 (N_12335,N_6076,N_9119);
nand U12336 (N_12336,N_9202,N_7891);
xor U12337 (N_12337,N_7094,N_9285);
xor U12338 (N_12338,N_9549,N_8340);
nor U12339 (N_12339,N_9041,N_8130);
or U12340 (N_12340,N_5082,N_8335);
or U12341 (N_12341,N_7138,N_5233);
nor U12342 (N_12342,N_5458,N_8885);
nor U12343 (N_12343,N_9849,N_6211);
nand U12344 (N_12344,N_5136,N_6042);
nor U12345 (N_12345,N_5511,N_7939);
xnor U12346 (N_12346,N_6852,N_5256);
nor U12347 (N_12347,N_6485,N_8371);
and U12348 (N_12348,N_6041,N_6934);
xnor U12349 (N_12349,N_7033,N_7602);
nor U12350 (N_12350,N_6823,N_5018);
or U12351 (N_12351,N_9516,N_6232);
and U12352 (N_12352,N_8801,N_7816);
xnor U12353 (N_12353,N_6605,N_5547);
nor U12354 (N_12354,N_6363,N_5509);
or U12355 (N_12355,N_7644,N_6429);
and U12356 (N_12356,N_8907,N_8526);
nor U12357 (N_12357,N_5161,N_8056);
xor U12358 (N_12358,N_8753,N_9777);
nand U12359 (N_12359,N_6806,N_8688);
nand U12360 (N_12360,N_9640,N_8897);
or U12361 (N_12361,N_6519,N_7797);
nor U12362 (N_12362,N_9811,N_7508);
nor U12363 (N_12363,N_8998,N_6611);
nor U12364 (N_12364,N_8457,N_6359);
xor U12365 (N_12365,N_6050,N_7521);
or U12366 (N_12366,N_6315,N_5011);
and U12367 (N_12367,N_5174,N_7065);
or U12368 (N_12368,N_6982,N_6692);
nand U12369 (N_12369,N_5670,N_7549);
nand U12370 (N_12370,N_7892,N_8628);
or U12371 (N_12371,N_9857,N_8805);
or U12372 (N_12372,N_5683,N_6200);
or U12373 (N_12373,N_5950,N_8644);
nand U12374 (N_12374,N_8712,N_5783);
xnor U12375 (N_12375,N_6950,N_6509);
nand U12376 (N_12376,N_6559,N_9345);
and U12377 (N_12377,N_7390,N_7533);
nand U12378 (N_12378,N_9460,N_8621);
xnor U12379 (N_12379,N_8032,N_6160);
nand U12380 (N_12380,N_5713,N_6822);
nor U12381 (N_12381,N_8445,N_7312);
xor U12382 (N_12382,N_5720,N_9006);
nand U12383 (N_12383,N_9318,N_7976);
nor U12384 (N_12384,N_5605,N_7793);
or U12385 (N_12385,N_6497,N_7953);
nor U12386 (N_12386,N_6575,N_6435);
nor U12387 (N_12387,N_9510,N_5249);
nand U12388 (N_12388,N_6872,N_5290);
nor U12389 (N_12389,N_7010,N_9955);
nor U12390 (N_12390,N_5572,N_8782);
xor U12391 (N_12391,N_7171,N_9056);
or U12392 (N_12392,N_9641,N_5867);
nor U12393 (N_12393,N_6411,N_7009);
or U12394 (N_12394,N_6227,N_8758);
nor U12395 (N_12395,N_5661,N_7487);
or U12396 (N_12396,N_7926,N_6944);
nor U12397 (N_12397,N_5651,N_6136);
and U12398 (N_12398,N_9178,N_8858);
and U12399 (N_12399,N_9845,N_7643);
nor U12400 (N_12400,N_7310,N_9210);
xor U12401 (N_12401,N_6245,N_9067);
or U12402 (N_12402,N_7660,N_9810);
nand U12403 (N_12403,N_9621,N_9534);
nand U12404 (N_12404,N_8933,N_5983);
nand U12405 (N_12405,N_5822,N_9933);
xor U12406 (N_12406,N_5976,N_6768);
nor U12407 (N_12407,N_5534,N_7258);
and U12408 (N_12408,N_6513,N_7078);
nand U12409 (N_12409,N_6512,N_9063);
nand U12410 (N_12410,N_9089,N_6629);
and U12411 (N_12411,N_9406,N_6240);
xor U12412 (N_12412,N_9591,N_7806);
nand U12413 (N_12413,N_7741,N_6280);
nand U12414 (N_12414,N_6759,N_9688);
nand U12415 (N_12415,N_7620,N_7598);
and U12416 (N_12416,N_8117,N_5553);
xor U12417 (N_12417,N_9706,N_7150);
nor U12418 (N_12418,N_6628,N_7241);
or U12419 (N_12419,N_7735,N_8705);
nor U12420 (N_12420,N_8242,N_7890);
or U12421 (N_12421,N_9691,N_8156);
xor U12422 (N_12422,N_7361,N_9218);
nand U12423 (N_12423,N_7068,N_6169);
nand U12424 (N_12424,N_8572,N_5948);
nand U12425 (N_12425,N_5009,N_7781);
or U12426 (N_12426,N_8979,N_8403);
xnor U12427 (N_12427,N_9487,N_7329);
or U12428 (N_12428,N_5624,N_8591);
xnor U12429 (N_12429,N_8530,N_9342);
or U12430 (N_12430,N_8113,N_7971);
or U12431 (N_12431,N_5209,N_6369);
or U12432 (N_12432,N_5663,N_8466);
nor U12433 (N_12433,N_8066,N_8884);
nand U12434 (N_12434,N_6266,N_6904);
nor U12435 (N_12435,N_5559,N_5455);
and U12436 (N_12436,N_8951,N_6263);
nand U12437 (N_12437,N_7527,N_9230);
and U12438 (N_12438,N_8055,N_9324);
and U12439 (N_12439,N_6524,N_5037);
xnor U12440 (N_12440,N_5949,N_9539);
nand U12441 (N_12441,N_7165,N_9198);
or U12442 (N_12442,N_7187,N_8085);
nand U12443 (N_12443,N_8083,N_5003);
nor U12444 (N_12444,N_8333,N_5415);
nor U12445 (N_12445,N_7196,N_7560);
nor U12446 (N_12446,N_7871,N_6420);
nand U12447 (N_12447,N_7879,N_5531);
nor U12448 (N_12448,N_5987,N_8062);
or U12449 (N_12449,N_7480,N_8449);
and U12450 (N_12450,N_8573,N_5577);
xor U12451 (N_12451,N_9040,N_9038);
nor U12452 (N_12452,N_9648,N_8306);
or U12453 (N_12453,N_5305,N_8947);
or U12454 (N_12454,N_9733,N_9651);
nand U12455 (N_12455,N_9238,N_7354);
xnor U12456 (N_12456,N_6643,N_5417);
or U12457 (N_12457,N_6625,N_5404);
nor U12458 (N_12458,N_9895,N_8069);
nand U12459 (N_12459,N_5310,N_8461);
or U12460 (N_12460,N_9118,N_6990);
and U12461 (N_12461,N_6540,N_5879);
xnor U12462 (N_12462,N_7881,N_8404);
and U12463 (N_12463,N_8739,N_5035);
nor U12464 (N_12464,N_5416,N_5186);
or U12465 (N_12465,N_9436,N_7657);
nand U12466 (N_12466,N_5279,N_8017);
or U12467 (N_12467,N_6979,N_6466);
nand U12468 (N_12468,N_8952,N_5993);
nand U12469 (N_12469,N_7112,N_7257);
nor U12470 (N_12470,N_5598,N_6561);
nor U12471 (N_12471,N_9662,N_8857);
nor U12472 (N_12472,N_7388,N_5297);
xor U12473 (N_12473,N_6935,N_7720);
or U12474 (N_12474,N_9667,N_7411);
nand U12475 (N_12475,N_6800,N_8486);
nor U12476 (N_12476,N_8260,N_6726);
nor U12477 (N_12477,N_7934,N_7219);
nor U12478 (N_12478,N_5705,N_5207);
and U12479 (N_12479,N_7336,N_8730);
or U12480 (N_12480,N_9261,N_6964);
or U12481 (N_12481,N_9658,N_5935);
nor U12482 (N_12482,N_7447,N_7032);
or U12483 (N_12483,N_5486,N_5770);
nand U12484 (N_12484,N_5133,N_6081);
nor U12485 (N_12485,N_5111,N_5274);
nand U12486 (N_12486,N_6353,N_6175);
or U12487 (N_12487,N_5914,N_9024);
xnor U12488 (N_12488,N_6938,N_6283);
nor U12489 (N_12489,N_9374,N_5141);
xnor U12490 (N_12490,N_6384,N_5512);
or U12491 (N_12491,N_7115,N_9494);
nor U12492 (N_12492,N_8921,N_8749);
and U12493 (N_12493,N_7152,N_7909);
nor U12494 (N_12494,N_8209,N_9466);
or U12495 (N_12495,N_5143,N_6723);
nand U12496 (N_12496,N_5429,N_6644);
or U12497 (N_12497,N_5258,N_5594);
and U12498 (N_12498,N_9898,N_7525);
or U12499 (N_12499,N_8231,N_5334);
or U12500 (N_12500,N_9456,N_6619);
xor U12501 (N_12501,N_7259,N_9171);
or U12502 (N_12502,N_6808,N_8250);
and U12503 (N_12503,N_7123,N_8177);
or U12504 (N_12504,N_8280,N_7558);
nand U12505 (N_12505,N_6813,N_5320);
or U12506 (N_12506,N_8590,N_5855);
nand U12507 (N_12507,N_8171,N_9851);
and U12508 (N_12508,N_5531,N_8416);
or U12509 (N_12509,N_5542,N_9056);
or U12510 (N_12510,N_5360,N_8593);
xor U12511 (N_12511,N_7972,N_7360);
or U12512 (N_12512,N_9411,N_7648);
and U12513 (N_12513,N_6159,N_5738);
xor U12514 (N_12514,N_7597,N_7128);
nor U12515 (N_12515,N_6468,N_8766);
nand U12516 (N_12516,N_6204,N_9287);
nor U12517 (N_12517,N_5557,N_8593);
and U12518 (N_12518,N_9521,N_7072);
and U12519 (N_12519,N_9626,N_9360);
nand U12520 (N_12520,N_7704,N_8149);
or U12521 (N_12521,N_9934,N_5148);
or U12522 (N_12522,N_8022,N_7455);
and U12523 (N_12523,N_8065,N_5091);
and U12524 (N_12524,N_5255,N_5307);
and U12525 (N_12525,N_9889,N_7735);
nor U12526 (N_12526,N_8018,N_8661);
nand U12527 (N_12527,N_6625,N_5921);
nand U12528 (N_12528,N_7174,N_6366);
and U12529 (N_12529,N_6486,N_8219);
and U12530 (N_12530,N_5127,N_9834);
and U12531 (N_12531,N_8214,N_5432);
nand U12532 (N_12532,N_8537,N_5342);
and U12533 (N_12533,N_6779,N_7253);
nand U12534 (N_12534,N_5508,N_9475);
or U12535 (N_12535,N_5557,N_6821);
nand U12536 (N_12536,N_7858,N_6411);
nor U12537 (N_12537,N_8722,N_8602);
xor U12538 (N_12538,N_9607,N_9940);
xor U12539 (N_12539,N_9000,N_6980);
nand U12540 (N_12540,N_5679,N_6491);
nor U12541 (N_12541,N_9278,N_8378);
and U12542 (N_12542,N_9975,N_6307);
nand U12543 (N_12543,N_8561,N_5159);
nand U12544 (N_12544,N_6666,N_6058);
xor U12545 (N_12545,N_8667,N_5155);
nand U12546 (N_12546,N_5883,N_6584);
nand U12547 (N_12547,N_6683,N_6544);
nand U12548 (N_12548,N_9510,N_8851);
or U12549 (N_12549,N_8893,N_9265);
nand U12550 (N_12550,N_5306,N_8259);
nor U12551 (N_12551,N_6184,N_9622);
nor U12552 (N_12552,N_6731,N_7047);
xnor U12553 (N_12553,N_6748,N_9429);
nor U12554 (N_12554,N_8985,N_5820);
and U12555 (N_12555,N_8770,N_7390);
nor U12556 (N_12556,N_7387,N_9456);
or U12557 (N_12557,N_5819,N_7346);
or U12558 (N_12558,N_9769,N_8982);
and U12559 (N_12559,N_6966,N_9202);
or U12560 (N_12560,N_8237,N_6580);
xnor U12561 (N_12561,N_8094,N_6801);
nor U12562 (N_12562,N_5951,N_8196);
xnor U12563 (N_12563,N_8697,N_5298);
or U12564 (N_12564,N_5061,N_7347);
and U12565 (N_12565,N_7952,N_8602);
or U12566 (N_12566,N_5703,N_6304);
nor U12567 (N_12567,N_7680,N_8946);
or U12568 (N_12568,N_5186,N_8939);
or U12569 (N_12569,N_9013,N_5748);
and U12570 (N_12570,N_6338,N_9425);
and U12571 (N_12571,N_8753,N_6489);
nand U12572 (N_12572,N_8640,N_8998);
or U12573 (N_12573,N_9108,N_9324);
nand U12574 (N_12574,N_8303,N_5402);
and U12575 (N_12575,N_6193,N_7041);
or U12576 (N_12576,N_9587,N_6896);
xnor U12577 (N_12577,N_5445,N_5372);
or U12578 (N_12578,N_9430,N_7529);
nand U12579 (N_12579,N_6298,N_9901);
nand U12580 (N_12580,N_6194,N_5391);
nor U12581 (N_12581,N_7208,N_8103);
and U12582 (N_12582,N_5226,N_7793);
nand U12583 (N_12583,N_5992,N_5284);
or U12584 (N_12584,N_8893,N_6126);
nand U12585 (N_12585,N_8801,N_5578);
and U12586 (N_12586,N_7383,N_7376);
or U12587 (N_12587,N_8236,N_7019);
and U12588 (N_12588,N_8990,N_6116);
nand U12589 (N_12589,N_7998,N_6239);
and U12590 (N_12590,N_7498,N_7130);
nor U12591 (N_12591,N_8623,N_8049);
nor U12592 (N_12592,N_5836,N_6325);
and U12593 (N_12593,N_8753,N_8708);
nand U12594 (N_12594,N_5246,N_8817);
nand U12595 (N_12595,N_8970,N_8683);
nand U12596 (N_12596,N_6463,N_5429);
or U12597 (N_12597,N_8026,N_9447);
nand U12598 (N_12598,N_9485,N_7695);
and U12599 (N_12599,N_6028,N_6451);
and U12600 (N_12600,N_6646,N_8542);
nor U12601 (N_12601,N_6458,N_9522);
nor U12602 (N_12602,N_9789,N_8692);
and U12603 (N_12603,N_8107,N_6942);
and U12604 (N_12604,N_5541,N_5202);
nor U12605 (N_12605,N_9781,N_6919);
nand U12606 (N_12606,N_7535,N_6951);
or U12607 (N_12607,N_5495,N_8070);
nor U12608 (N_12608,N_5953,N_8560);
nor U12609 (N_12609,N_5650,N_6339);
nand U12610 (N_12610,N_8906,N_5773);
and U12611 (N_12611,N_8295,N_7803);
and U12612 (N_12612,N_8968,N_8380);
or U12613 (N_12613,N_8961,N_6454);
and U12614 (N_12614,N_7216,N_7068);
and U12615 (N_12615,N_5202,N_8280);
nand U12616 (N_12616,N_8179,N_6523);
or U12617 (N_12617,N_6945,N_9182);
nor U12618 (N_12618,N_8581,N_9397);
and U12619 (N_12619,N_5644,N_9144);
and U12620 (N_12620,N_6330,N_6541);
nand U12621 (N_12621,N_7530,N_5981);
xnor U12622 (N_12622,N_5224,N_9862);
or U12623 (N_12623,N_6362,N_9672);
xor U12624 (N_12624,N_8627,N_8373);
and U12625 (N_12625,N_7958,N_6607);
or U12626 (N_12626,N_6161,N_5525);
or U12627 (N_12627,N_7554,N_6912);
or U12628 (N_12628,N_8113,N_6461);
and U12629 (N_12629,N_8955,N_5079);
and U12630 (N_12630,N_9585,N_6931);
or U12631 (N_12631,N_7141,N_9984);
nor U12632 (N_12632,N_5872,N_5217);
nor U12633 (N_12633,N_6682,N_9253);
nand U12634 (N_12634,N_8275,N_9639);
nand U12635 (N_12635,N_6227,N_7348);
xor U12636 (N_12636,N_7796,N_9464);
and U12637 (N_12637,N_9575,N_6336);
nand U12638 (N_12638,N_7683,N_6328);
nor U12639 (N_12639,N_5561,N_5752);
nor U12640 (N_12640,N_5428,N_8955);
nand U12641 (N_12641,N_6600,N_8430);
nor U12642 (N_12642,N_9086,N_5443);
and U12643 (N_12643,N_9636,N_5495);
xor U12644 (N_12644,N_5925,N_7113);
and U12645 (N_12645,N_7798,N_5375);
or U12646 (N_12646,N_8548,N_6936);
nor U12647 (N_12647,N_6864,N_8730);
and U12648 (N_12648,N_5797,N_5241);
nand U12649 (N_12649,N_9241,N_9571);
nand U12650 (N_12650,N_9883,N_8269);
nand U12651 (N_12651,N_5445,N_7236);
or U12652 (N_12652,N_9579,N_8523);
xor U12653 (N_12653,N_5893,N_6840);
and U12654 (N_12654,N_6446,N_5530);
nand U12655 (N_12655,N_6219,N_8418);
xor U12656 (N_12656,N_9562,N_6122);
xor U12657 (N_12657,N_7787,N_8874);
nor U12658 (N_12658,N_5970,N_7862);
nor U12659 (N_12659,N_9696,N_8907);
nand U12660 (N_12660,N_9958,N_7984);
and U12661 (N_12661,N_7222,N_5978);
or U12662 (N_12662,N_8324,N_6326);
xor U12663 (N_12663,N_7972,N_5386);
or U12664 (N_12664,N_8376,N_9221);
nor U12665 (N_12665,N_7755,N_9205);
or U12666 (N_12666,N_9342,N_7563);
and U12667 (N_12667,N_8437,N_7533);
and U12668 (N_12668,N_9302,N_8843);
nand U12669 (N_12669,N_5266,N_7222);
nor U12670 (N_12670,N_8344,N_9837);
or U12671 (N_12671,N_6474,N_6409);
nand U12672 (N_12672,N_9629,N_7093);
nand U12673 (N_12673,N_5065,N_9270);
or U12674 (N_12674,N_6843,N_5278);
and U12675 (N_12675,N_9268,N_8519);
and U12676 (N_12676,N_7540,N_6612);
or U12677 (N_12677,N_8248,N_6469);
xnor U12678 (N_12678,N_8008,N_9917);
or U12679 (N_12679,N_6341,N_9219);
nor U12680 (N_12680,N_6738,N_9716);
and U12681 (N_12681,N_6787,N_7262);
or U12682 (N_12682,N_5555,N_7785);
nand U12683 (N_12683,N_8762,N_8781);
and U12684 (N_12684,N_8924,N_5330);
and U12685 (N_12685,N_8508,N_8217);
or U12686 (N_12686,N_7667,N_8979);
and U12687 (N_12687,N_7431,N_5662);
nor U12688 (N_12688,N_8026,N_9871);
xnor U12689 (N_12689,N_7603,N_8412);
and U12690 (N_12690,N_6403,N_8434);
or U12691 (N_12691,N_9983,N_5101);
xnor U12692 (N_12692,N_6001,N_8927);
and U12693 (N_12693,N_5441,N_8137);
and U12694 (N_12694,N_5645,N_7109);
nand U12695 (N_12695,N_6616,N_5354);
xor U12696 (N_12696,N_7956,N_9429);
nand U12697 (N_12697,N_6203,N_8762);
nor U12698 (N_12698,N_6060,N_5337);
nor U12699 (N_12699,N_7097,N_9895);
and U12700 (N_12700,N_5402,N_7511);
nor U12701 (N_12701,N_8846,N_5531);
and U12702 (N_12702,N_9072,N_7175);
or U12703 (N_12703,N_6638,N_5371);
and U12704 (N_12704,N_5593,N_6093);
nor U12705 (N_12705,N_9042,N_6229);
or U12706 (N_12706,N_6592,N_6471);
and U12707 (N_12707,N_6379,N_7309);
and U12708 (N_12708,N_9038,N_7616);
nand U12709 (N_12709,N_8402,N_6908);
nor U12710 (N_12710,N_5656,N_7356);
nor U12711 (N_12711,N_5309,N_8581);
nor U12712 (N_12712,N_5737,N_7611);
xor U12713 (N_12713,N_7218,N_9967);
nand U12714 (N_12714,N_9275,N_6827);
nand U12715 (N_12715,N_6448,N_9737);
nor U12716 (N_12716,N_5409,N_7452);
nor U12717 (N_12717,N_6493,N_5718);
or U12718 (N_12718,N_9251,N_7243);
nand U12719 (N_12719,N_8250,N_8422);
xnor U12720 (N_12720,N_9783,N_5880);
and U12721 (N_12721,N_5924,N_7348);
nand U12722 (N_12722,N_6256,N_5715);
nor U12723 (N_12723,N_7412,N_9861);
or U12724 (N_12724,N_5038,N_5411);
nor U12725 (N_12725,N_8638,N_8741);
nand U12726 (N_12726,N_5362,N_5410);
and U12727 (N_12727,N_7945,N_5421);
xor U12728 (N_12728,N_6298,N_5881);
nand U12729 (N_12729,N_6080,N_5498);
nand U12730 (N_12730,N_9397,N_9366);
and U12731 (N_12731,N_6630,N_8027);
nor U12732 (N_12732,N_6515,N_6175);
nor U12733 (N_12733,N_5985,N_9737);
xor U12734 (N_12734,N_6176,N_6528);
nor U12735 (N_12735,N_8028,N_6907);
and U12736 (N_12736,N_6438,N_9669);
or U12737 (N_12737,N_8408,N_9365);
nor U12738 (N_12738,N_8098,N_5341);
nand U12739 (N_12739,N_5601,N_8715);
or U12740 (N_12740,N_7601,N_8077);
xnor U12741 (N_12741,N_7196,N_9420);
and U12742 (N_12742,N_6342,N_7202);
and U12743 (N_12743,N_8249,N_9964);
xnor U12744 (N_12744,N_6197,N_8909);
xnor U12745 (N_12745,N_9163,N_9028);
nand U12746 (N_12746,N_6663,N_6906);
or U12747 (N_12747,N_8825,N_5920);
or U12748 (N_12748,N_6911,N_8979);
or U12749 (N_12749,N_7392,N_6857);
xnor U12750 (N_12750,N_5396,N_7039);
nand U12751 (N_12751,N_8020,N_6738);
or U12752 (N_12752,N_6360,N_9559);
nor U12753 (N_12753,N_8009,N_6365);
xor U12754 (N_12754,N_6593,N_7213);
nand U12755 (N_12755,N_7404,N_5726);
or U12756 (N_12756,N_9034,N_8542);
nor U12757 (N_12757,N_8449,N_8169);
or U12758 (N_12758,N_8588,N_7049);
and U12759 (N_12759,N_8224,N_9892);
nor U12760 (N_12760,N_5119,N_9679);
nor U12761 (N_12761,N_5505,N_9959);
nor U12762 (N_12762,N_7894,N_7827);
and U12763 (N_12763,N_8952,N_6873);
nor U12764 (N_12764,N_5261,N_9432);
and U12765 (N_12765,N_6024,N_5649);
or U12766 (N_12766,N_9659,N_6164);
or U12767 (N_12767,N_5415,N_7867);
nor U12768 (N_12768,N_7846,N_6206);
nor U12769 (N_12769,N_7595,N_6457);
nand U12770 (N_12770,N_5986,N_7833);
nor U12771 (N_12771,N_8372,N_6711);
and U12772 (N_12772,N_5526,N_9407);
or U12773 (N_12773,N_8264,N_7576);
and U12774 (N_12774,N_5531,N_5353);
and U12775 (N_12775,N_5104,N_8853);
or U12776 (N_12776,N_9405,N_9053);
nor U12777 (N_12777,N_8537,N_7959);
nor U12778 (N_12778,N_5296,N_7898);
nor U12779 (N_12779,N_5373,N_6723);
or U12780 (N_12780,N_8365,N_5286);
nor U12781 (N_12781,N_6763,N_6933);
or U12782 (N_12782,N_6666,N_9678);
nor U12783 (N_12783,N_5769,N_6503);
and U12784 (N_12784,N_9712,N_6636);
or U12785 (N_12785,N_5572,N_8624);
and U12786 (N_12786,N_9688,N_7006);
nand U12787 (N_12787,N_7489,N_7852);
nand U12788 (N_12788,N_9913,N_7846);
nand U12789 (N_12789,N_7832,N_7847);
or U12790 (N_12790,N_7701,N_9297);
nor U12791 (N_12791,N_6656,N_5223);
and U12792 (N_12792,N_8105,N_8326);
nor U12793 (N_12793,N_8128,N_8322);
nand U12794 (N_12794,N_7461,N_5529);
and U12795 (N_12795,N_9430,N_6455);
xnor U12796 (N_12796,N_7371,N_5853);
and U12797 (N_12797,N_9590,N_5493);
nor U12798 (N_12798,N_8537,N_5272);
xnor U12799 (N_12799,N_7059,N_7383);
or U12800 (N_12800,N_6987,N_8462);
nor U12801 (N_12801,N_6665,N_8641);
and U12802 (N_12802,N_8568,N_8904);
nand U12803 (N_12803,N_8663,N_5323);
xor U12804 (N_12804,N_6495,N_5087);
nor U12805 (N_12805,N_8430,N_5801);
nand U12806 (N_12806,N_9302,N_9534);
xor U12807 (N_12807,N_8104,N_7898);
and U12808 (N_12808,N_6263,N_7736);
nand U12809 (N_12809,N_7677,N_8204);
nor U12810 (N_12810,N_8556,N_7625);
xnor U12811 (N_12811,N_9607,N_8412);
and U12812 (N_12812,N_7809,N_7212);
nand U12813 (N_12813,N_5818,N_6218);
nand U12814 (N_12814,N_8995,N_8564);
or U12815 (N_12815,N_5913,N_5145);
nor U12816 (N_12816,N_7493,N_8528);
or U12817 (N_12817,N_8808,N_7081);
and U12818 (N_12818,N_8250,N_8404);
nand U12819 (N_12819,N_9901,N_6107);
and U12820 (N_12820,N_5825,N_6778);
and U12821 (N_12821,N_9545,N_8690);
and U12822 (N_12822,N_9631,N_5248);
nand U12823 (N_12823,N_7850,N_8054);
and U12824 (N_12824,N_9343,N_8256);
xor U12825 (N_12825,N_8091,N_5600);
nor U12826 (N_12826,N_5664,N_5881);
or U12827 (N_12827,N_7065,N_7593);
or U12828 (N_12828,N_7675,N_5726);
nand U12829 (N_12829,N_8456,N_9547);
and U12830 (N_12830,N_7834,N_7938);
or U12831 (N_12831,N_7908,N_6698);
or U12832 (N_12832,N_8155,N_5242);
xor U12833 (N_12833,N_5600,N_9923);
and U12834 (N_12834,N_7080,N_5705);
nand U12835 (N_12835,N_5674,N_8168);
and U12836 (N_12836,N_5258,N_7207);
nor U12837 (N_12837,N_6330,N_7851);
nor U12838 (N_12838,N_5273,N_9284);
and U12839 (N_12839,N_8243,N_6040);
nor U12840 (N_12840,N_6714,N_6638);
or U12841 (N_12841,N_5907,N_6366);
xnor U12842 (N_12842,N_5840,N_6272);
and U12843 (N_12843,N_5449,N_9863);
nor U12844 (N_12844,N_7014,N_9167);
and U12845 (N_12845,N_9564,N_8794);
nor U12846 (N_12846,N_6254,N_6595);
xnor U12847 (N_12847,N_8076,N_8648);
or U12848 (N_12848,N_7028,N_5100);
nor U12849 (N_12849,N_9191,N_8948);
and U12850 (N_12850,N_9443,N_5653);
nor U12851 (N_12851,N_8641,N_9845);
nand U12852 (N_12852,N_6400,N_8989);
and U12853 (N_12853,N_5254,N_9304);
nor U12854 (N_12854,N_9769,N_5329);
xor U12855 (N_12855,N_6639,N_6170);
nor U12856 (N_12856,N_8961,N_6254);
nand U12857 (N_12857,N_9103,N_5181);
xnor U12858 (N_12858,N_7199,N_9342);
nand U12859 (N_12859,N_7823,N_8692);
nand U12860 (N_12860,N_7628,N_8136);
or U12861 (N_12861,N_9830,N_5409);
nor U12862 (N_12862,N_6209,N_8515);
nand U12863 (N_12863,N_9472,N_9547);
nand U12864 (N_12864,N_8489,N_9454);
and U12865 (N_12865,N_7829,N_5275);
nand U12866 (N_12866,N_8651,N_9106);
nand U12867 (N_12867,N_7254,N_8140);
and U12868 (N_12868,N_8230,N_5015);
nor U12869 (N_12869,N_7292,N_5021);
and U12870 (N_12870,N_8206,N_8506);
nor U12871 (N_12871,N_8274,N_5611);
nor U12872 (N_12872,N_7437,N_9474);
nand U12873 (N_12873,N_6448,N_5267);
and U12874 (N_12874,N_8212,N_9343);
or U12875 (N_12875,N_8748,N_5239);
and U12876 (N_12876,N_8914,N_9763);
nand U12877 (N_12877,N_7005,N_7959);
and U12878 (N_12878,N_6386,N_7078);
xor U12879 (N_12879,N_6756,N_9549);
nor U12880 (N_12880,N_8928,N_8855);
and U12881 (N_12881,N_7055,N_8988);
or U12882 (N_12882,N_9345,N_8016);
nor U12883 (N_12883,N_7417,N_5089);
or U12884 (N_12884,N_8676,N_8389);
nor U12885 (N_12885,N_6953,N_6469);
and U12886 (N_12886,N_6716,N_6038);
and U12887 (N_12887,N_7846,N_9396);
or U12888 (N_12888,N_7140,N_6216);
or U12889 (N_12889,N_8721,N_9717);
or U12890 (N_12890,N_6054,N_5289);
or U12891 (N_12891,N_8778,N_7921);
or U12892 (N_12892,N_7053,N_9069);
nand U12893 (N_12893,N_9220,N_8512);
xor U12894 (N_12894,N_8313,N_6827);
nand U12895 (N_12895,N_6786,N_5091);
or U12896 (N_12896,N_7384,N_5051);
nor U12897 (N_12897,N_8060,N_9508);
nand U12898 (N_12898,N_8532,N_7758);
or U12899 (N_12899,N_8185,N_9463);
or U12900 (N_12900,N_9131,N_8216);
and U12901 (N_12901,N_7718,N_6981);
or U12902 (N_12902,N_8543,N_5171);
and U12903 (N_12903,N_9374,N_7690);
nor U12904 (N_12904,N_5466,N_7119);
xor U12905 (N_12905,N_6860,N_5470);
and U12906 (N_12906,N_8244,N_9156);
or U12907 (N_12907,N_6823,N_6066);
nand U12908 (N_12908,N_9242,N_9115);
nand U12909 (N_12909,N_5325,N_8732);
nand U12910 (N_12910,N_9659,N_5318);
and U12911 (N_12911,N_8515,N_8263);
nand U12912 (N_12912,N_5128,N_9541);
xor U12913 (N_12913,N_7016,N_5159);
nand U12914 (N_12914,N_8163,N_8171);
nor U12915 (N_12915,N_8600,N_9520);
or U12916 (N_12916,N_7300,N_9513);
nor U12917 (N_12917,N_7651,N_8563);
or U12918 (N_12918,N_7675,N_9176);
nor U12919 (N_12919,N_6433,N_6774);
nor U12920 (N_12920,N_6185,N_7810);
xor U12921 (N_12921,N_8572,N_8134);
nor U12922 (N_12922,N_7198,N_7129);
xor U12923 (N_12923,N_7526,N_5828);
and U12924 (N_12924,N_8722,N_9426);
or U12925 (N_12925,N_5929,N_8997);
nand U12926 (N_12926,N_8120,N_7348);
nand U12927 (N_12927,N_9352,N_5975);
nor U12928 (N_12928,N_5027,N_8843);
nand U12929 (N_12929,N_5491,N_9473);
or U12930 (N_12930,N_9897,N_7318);
and U12931 (N_12931,N_6842,N_7077);
or U12932 (N_12932,N_7958,N_9576);
nor U12933 (N_12933,N_5254,N_5583);
nor U12934 (N_12934,N_5046,N_9024);
and U12935 (N_12935,N_6987,N_8134);
xor U12936 (N_12936,N_7601,N_5686);
and U12937 (N_12937,N_5678,N_9934);
xnor U12938 (N_12938,N_9459,N_8979);
nor U12939 (N_12939,N_7025,N_5179);
or U12940 (N_12940,N_6138,N_7118);
and U12941 (N_12941,N_7954,N_5608);
and U12942 (N_12942,N_5256,N_6200);
or U12943 (N_12943,N_9723,N_9361);
nor U12944 (N_12944,N_8597,N_5821);
and U12945 (N_12945,N_7960,N_7887);
nor U12946 (N_12946,N_7200,N_8230);
or U12947 (N_12947,N_6501,N_7572);
or U12948 (N_12948,N_6691,N_8916);
nand U12949 (N_12949,N_7754,N_9514);
or U12950 (N_12950,N_8969,N_5113);
xnor U12951 (N_12951,N_8934,N_5480);
xnor U12952 (N_12952,N_6538,N_8175);
nand U12953 (N_12953,N_5303,N_5135);
and U12954 (N_12954,N_6674,N_8508);
nand U12955 (N_12955,N_7041,N_9911);
xnor U12956 (N_12956,N_9611,N_5839);
nor U12957 (N_12957,N_9958,N_5963);
nor U12958 (N_12958,N_7869,N_8747);
or U12959 (N_12959,N_8813,N_5966);
nand U12960 (N_12960,N_8736,N_7071);
or U12961 (N_12961,N_6229,N_6973);
nor U12962 (N_12962,N_6893,N_8273);
and U12963 (N_12963,N_8233,N_6451);
nand U12964 (N_12964,N_8862,N_8198);
nor U12965 (N_12965,N_8346,N_7751);
or U12966 (N_12966,N_9112,N_7812);
nand U12967 (N_12967,N_6734,N_9125);
nand U12968 (N_12968,N_8641,N_8741);
nor U12969 (N_12969,N_9176,N_6770);
and U12970 (N_12970,N_6994,N_7393);
nor U12971 (N_12971,N_8402,N_8768);
nand U12972 (N_12972,N_7977,N_6186);
nand U12973 (N_12973,N_5010,N_9439);
nand U12974 (N_12974,N_9715,N_6295);
nand U12975 (N_12975,N_5450,N_8392);
nor U12976 (N_12976,N_8540,N_8166);
xnor U12977 (N_12977,N_6559,N_8014);
or U12978 (N_12978,N_6708,N_7606);
and U12979 (N_12979,N_8204,N_6580);
xor U12980 (N_12980,N_5224,N_8126);
and U12981 (N_12981,N_6224,N_9388);
or U12982 (N_12982,N_6669,N_5173);
and U12983 (N_12983,N_9400,N_7351);
or U12984 (N_12984,N_8278,N_9747);
xor U12985 (N_12985,N_5594,N_9278);
or U12986 (N_12986,N_6288,N_7013);
and U12987 (N_12987,N_9142,N_6083);
and U12988 (N_12988,N_9508,N_6943);
xor U12989 (N_12989,N_5693,N_8955);
and U12990 (N_12990,N_5906,N_8659);
nor U12991 (N_12991,N_6519,N_9866);
nor U12992 (N_12992,N_7496,N_9107);
or U12993 (N_12993,N_9852,N_8865);
nor U12994 (N_12994,N_6356,N_7811);
xor U12995 (N_12995,N_7404,N_6328);
and U12996 (N_12996,N_5968,N_6098);
nand U12997 (N_12997,N_7026,N_6446);
or U12998 (N_12998,N_8413,N_9233);
or U12999 (N_12999,N_7499,N_5953);
nor U13000 (N_13000,N_9954,N_9527);
and U13001 (N_13001,N_6789,N_8245);
nand U13002 (N_13002,N_6278,N_7391);
xnor U13003 (N_13003,N_8226,N_7411);
or U13004 (N_13004,N_9854,N_7528);
xor U13005 (N_13005,N_5112,N_7663);
nor U13006 (N_13006,N_9933,N_5120);
or U13007 (N_13007,N_8458,N_9954);
nand U13008 (N_13008,N_6573,N_8793);
nand U13009 (N_13009,N_7993,N_8606);
nor U13010 (N_13010,N_6441,N_8439);
or U13011 (N_13011,N_5760,N_8507);
or U13012 (N_13012,N_8174,N_9088);
nor U13013 (N_13013,N_9463,N_7500);
and U13014 (N_13014,N_8583,N_7160);
and U13015 (N_13015,N_8362,N_5297);
or U13016 (N_13016,N_5667,N_6430);
and U13017 (N_13017,N_7057,N_9365);
nor U13018 (N_13018,N_7927,N_7784);
or U13019 (N_13019,N_6642,N_6043);
or U13020 (N_13020,N_5035,N_7058);
nor U13021 (N_13021,N_8245,N_9949);
and U13022 (N_13022,N_6835,N_5533);
or U13023 (N_13023,N_9411,N_6870);
nand U13024 (N_13024,N_7035,N_7810);
and U13025 (N_13025,N_7758,N_8338);
or U13026 (N_13026,N_6787,N_7387);
nor U13027 (N_13027,N_6890,N_7148);
or U13028 (N_13028,N_5377,N_8819);
xor U13029 (N_13029,N_6146,N_9036);
nand U13030 (N_13030,N_7952,N_8530);
or U13031 (N_13031,N_8579,N_5254);
or U13032 (N_13032,N_8347,N_7205);
nor U13033 (N_13033,N_9277,N_9771);
nor U13034 (N_13034,N_6762,N_5896);
nand U13035 (N_13035,N_6195,N_6766);
xor U13036 (N_13036,N_8614,N_5361);
nor U13037 (N_13037,N_9527,N_7753);
nand U13038 (N_13038,N_6594,N_5061);
and U13039 (N_13039,N_9333,N_6780);
nor U13040 (N_13040,N_5447,N_8144);
xnor U13041 (N_13041,N_9828,N_9515);
nor U13042 (N_13042,N_8371,N_9619);
nor U13043 (N_13043,N_7291,N_8989);
nand U13044 (N_13044,N_8920,N_6839);
xnor U13045 (N_13045,N_5163,N_5882);
or U13046 (N_13046,N_5908,N_6545);
or U13047 (N_13047,N_6735,N_6419);
nor U13048 (N_13048,N_6671,N_5761);
and U13049 (N_13049,N_9327,N_5768);
and U13050 (N_13050,N_9119,N_9639);
and U13051 (N_13051,N_6389,N_7826);
nand U13052 (N_13052,N_7676,N_6284);
xor U13053 (N_13053,N_9520,N_6312);
nor U13054 (N_13054,N_6546,N_6101);
and U13055 (N_13055,N_5949,N_7166);
nor U13056 (N_13056,N_8128,N_8849);
nand U13057 (N_13057,N_8318,N_6773);
nor U13058 (N_13058,N_7655,N_7827);
and U13059 (N_13059,N_8612,N_9098);
and U13060 (N_13060,N_6084,N_5182);
or U13061 (N_13061,N_7013,N_5018);
or U13062 (N_13062,N_8584,N_7900);
xnor U13063 (N_13063,N_8651,N_7414);
and U13064 (N_13064,N_5093,N_7000);
xor U13065 (N_13065,N_7251,N_9503);
and U13066 (N_13066,N_5759,N_7040);
nor U13067 (N_13067,N_9599,N_5051);
nand U13068 (N_13068,N_8525,N_8510);
and U13069 (N_13069,N_5281,N_8801);
and U13070 (N_13070,N_9188,N_5420);
nor U13071 (N_13071,N_9535,N_9984);
xnor U13072 (N_13072,N_6969,N_9701);
and U13073 (N_13073,N_9731,N_8401);
nand U13074 (N_13074,N_5729,N_9073);
nand U13075 (N_13075,N_7143,N_9050);
nand U13076 (N_13076,N_7505,N_6986);
and U13077 (N_13077,N_5709,N_5481);
xor U13078 (N_13078,N_9412,N_9414);
or U13079 (N_13079,N_5770,N_8826);
or U13080 (N_13080,N_7076,N_6084);
nor U13081 (N_13081,N_8265,N_7999);
or U13082 (N_13082,N_6245,N_6065);
xnor U13083 (N_13083,N_6199,N_6480);
nor U13084 (N_13084,N_7023,N_7809);
or U13085 (N_13085,N_6523,N_8755);
or U13086 (N_13086,N_9711,N_7460);
xor U13087 (N_13087,N_6166,N_5107);
nand U13088 (N_13088,N_7142,N_5030);
nand U13089 (N_13089,N_9361,N_8565);
and U13090 (N_13090,N_5166,N_7818);
nand U13091 (N_13091,N_5996,N_5367);
nand U13092 (N_13092,N_8062,N_6387);
nand U13093 (N_13093,N_9373,N_9281);
nor U13094 (N_13094,N_6837,N_8322);
or U13095 (N_13095,N_8985,N_8678);
nor U13096 (N_13096,N_8201,N_5294);
nand U13097 (N_13097,N_9657,N_8421);
nand U13098 (N_13098,N_6601,N_5385);
nand U13099 (N_13099,N_7124,N_9402);
nand U13100 (N_13100,N_6947,N_8364);
xnor U13101 (N_13101,N_8151,N_5510);
xnor U13102 (N_13102,N_9897,N_8462);
and U13103 (N_13103,N_9304,N_8091);
xnor U13104 (N_13104,N_9171,N_6608);
nor U13105 (N_13105,N_8924,N_7668);
and U13106 (N_13106,N_5137,N_6635);
or U13107 (N_13107,N_5128,N_6605);
nor U13108 (N_13108,N_7435,N_9573);
nor U13109 (N_13109,N_9663,N_8462);
or U13110 (N_13110,N_6102,N_8788);
or U13111 (N_13111,N_5873,N_8700);
nand U13112 (N_13112,N_8642,N_7113);
nor U13113 (N_13113,N_8840,N_5801);
and U13114 (N_13114,N_5114,N_8815);
or U13115 (N_13115,N_8017,N_6709);
nor U13116 (N_13116,N_5912,N_6957);
xor U13117 (N_13117,N_9316,N_8912);
xnor U13118 (N_13118,N_9904,N_7809);
and U13119 (N_13119,N_8943,N_9999);
nand U13120 (N_13120,N_5315,N_9895);
or U13121 (N_13121,N_8149,N_8288);
or U13122 (N_13122,N_9403,N_9309);
or U13123 (N_13123,N_7158,N_8485);
xnor U13124 (N_13124,N_7915,N_7243);
nand U13125 (N_13125,N_8741,N_9739);
xnor U13126 (N_13126,N_5950,N_5569);
xnor U13127 (N_13127,N_7719,N_7724);
nor U13128 (N_13128,N_8944,N_6787);
xor U13129 (N_13129,N_7766,N_7284);
nand U13130 (N_13130,N_7712,N_9966);
or U13131 (N_13131,N_8712,N_8390);
or U13132 (N_13132,N_5926,N_8437);
or U13133 (N_13133,N_5741,N_9220);
or U13134 (N_13134,N_8924,N_7341);
nand U13135 (N_13135,N_7931,N_5418);
and U13136 (N_13136,N_7759,N_7203);
xor U13137 (N_13137,N_6340,N_5040);
nand U13138 (N_13138,N_9499,N_9520);
nand U13139 (N_13139,N_7611,N_6650);
and U13140 (N_13140,N_8296,N_6199);
nand U13141 (N_13141,N_6308,N_5348);
nor U13142 (N_13142,N_8813,N_7716);
or U13143 (N_13143,N_9342,N_9191);
and U13144 (N_13144,N_6939,N_8347);
nand U13145 (N_13145,N_7639,N_8951);
and U13146 (N_13146,N_6658,N_6680);
or U13147 (N_13147,N_5348,N_8137);
nand U13148 (N_13148,N_6743,N_9281);
nor U13149 (N_13149,N_9032,N_6748);
nand U13150 (N_13150,N_5122,N_9710);
nor U13151 (N_13151,N_9738,N_6650);
or U13152 (N_13152,N_6026,N_7492);
xnor U13153 (N_13153,N_5883,N_8094);
nand U13154 (N_13154,N_7183,N_8134);
and U13155 (N_13155,N_8882,N_8495);
nand U13156 (N_13156,N_6741,N_9649);
nand U13157 (N_13157,N_7483,N_9967);
nor U13158 (N_13158,N_9100,N_9073);
or U13159 (N_13159,N_6804,N_6507);
and U13160 (N_13160,N_8743,N_9623);
nor U13161 (N_13161,N_6414,N_9265);
nor U13162 (N_13162,N_5848,N_9212);
and U13163 (N_13163,N_5231,N_5952);
nand U13164 (N_13164,N_5072,N_6341);
nor U13165 (N_13165,N_8072,N_9192);
and U13166 (N_13166,N_9424,N_6189);
nor U13167 (N_13167,N_6442,N_7248);
nand U13168 (N_13168,N_6797,N_9333);
nand U13169 (N_13169,N_9310,N_9226);
nand U13170 (N_13170,N_5810,N_7810);
xor U13171 (N_13171,N_9247,N_7948);
nor U13172 (N_13172,N_7649,N_7902);
or U13173 (N_13173,N_5261,N_6922);
nor U13174 (N_13174,N_7453,N_5774);
nand U13175 (N_13175,N_6680,N_9998);
and U13176 (N_13176,N_8072,N_7428);
nand U13177 (N_13177,N_8991,N_7657);
nor U13178 (N_13178,N_5270,N_7346);
nor U13179 (N_13179,N_7852,N_6630);
or U13180 (N_13180,N_7866,N_5177);
and U13181 (N_13181,N_6398,N_6347);
nand U13182 (N_13182,N_6679,N_6306);
or U13183 (N_13183,N_9891,N_7149);
nor U13184 (N_13184,N_9914,N_5587);
nand U13185 (N_13185,N_6837,N_7954);
and U13186 (N_13186,N_5033,N_9574);
and U13187 (N_13187,N_7077,N_7302);
nand U13188 (N_13188,N_5815,N_8795);
or U13189 (N_13189,N_7536,N_7906);
or U13190 (N_13190,N_6012,N_9113);
and U13191 (N_13191,N_5243,N_5173);
nand U13192 (N_13192,N_7261,N_5627);
and U13193 (N_13193,N_6515,N_9569);
and U13194 (N_13194,N_7312,N_8343);
and U13195 (N_13195,N_9443,N_8806);
or U13196 (N_13196,N_8224,N_7279);
xor U13197 (N_13197,N_6693,N_9486);
and U13198 (N_13198,N_9473,N_7977);
nand U13199 (N_13199,N_7705,N_6351);
nor U13200 (N_13200,N_7039,N_9735);
xnor U13201 (N_13201,N_5163,N_6505);
nand U13202 (N_13202,N_8213,N_6791);
nor U13203 (N_13203,N_6874,N_7544);
or U13204 (N_13204,N_8075,N_5550);
nor U13205 (N_13205,N_7036,N_6675);
and U13206 (N_13206,N_6258,N_7402);
or U13207 (N_13207,N_6946,N_5599);
nor U13208 (N_13208,N_8139,N_6130);
and U13209 (N_13209,N_6276,N_7944);
nor U13210 (N_13210,N_6511,N_6472);
nor U13211 (N_13211,N_9376,N_5938);
nor U13212 (N_13212,N_9286,N_9808);
or U13213 (N_13213,N_9238,N_8124);
nand U13214 (N_13214,N_7543,N_9098);
and U13215 (N_13215,N_8699,N_9809);
and U13216 (N_13216,N_8841,N_9570);
nand U13217 (N_13217,N_9591,N_7114);
and U13218 (N_13218,N_7008,N_9941);
and U13219 (N_13219,N_9589,N_6119);
xor U13220 (N_13220,N_8859,N_9908);
nand U13221 (N_13221,N_5984,N_5627);
nand U13222 (N_13222,N_5901,N_9754);
nand U13223 (N_13223,N_8375,N_6866);
or U13224 (N_13224,N_7523,N_9708);
xnor U13225 (N_13225,N_7868,N_5094);
xor U13226 (N_13226,N_8606,N_9727);
nor U13227 (N_13227,N_6001,N_9187);
nor U13228 (N_13228,N_7248,N_6260);
nand U13229 (N_13229,N_8856,N_8453);
nor U13230 (N_13230,N_6118,N_8397);
or U13231 (N_13231,N_8904,N_6517);
and U13232 (N_13232,N_5127,N_6650);
and U13233 (N_13233,N_5780,N_7664);
or U13234 (N_13234,N_8872,N_5266);
nand U13235 (N_13235,N_8009,N_8448);
nor U13236 (N_13236,N_9543,N_9779);
nand U13237 (N_13237,N_5309,N_5069);
or U13238 (N_13238,N_8373,N_5369);
nand U13239 (N_13239,N_8376,N_5273);
nor U13240 (N_13240,N_5174,N_5934);
or U13241 (N_13241,N_9954,N_7036);
nand U13242 (N_13242,N_5529,N_9145);
nor U13243 (N_13243,N_6158,N_5224);
nand U13244 (N_13244,N_9228,N_6072);
nand U13245 (N_13245,N_5334,N_6214);
nand U13246 (N_13246,N_6707,N_9800);
nand U13247 (N_13247,N_7124,N_9799);
nor U13248 (N_13248,N_9227,N_6670);
nand U13249 (N_13249,N_6688,N_7388);
and U13250 (N_13250,N_9351,N_5085);
and U13251 (N_13251,N_7361,N_8832);
and U13252 (N_13252,N_8298,N_7277);
or U13253 (N_13253,N_6632,N_9258);
nor U13254 (N_13254,N_8953,N_9952);
or U13255 (N_13255,N_7574,N_7153);
or U13256 (N_13256,N_8182,N_9485);
nor U13257 (N_13257,N_6312,N_5012);
or U13258 (N_13258,N_8658,N_9325);
nand U13259 (N_13259,N_5510,N_9236);
nor U13260 (N_13260,N_6114,N_8748);
or U13261 (N_13261,N_6278,N_8376);
or U13262 (N_13262,N_9245,N_8376);
and U13263 (N_13263,N_7878,N_7435);
or U13264 (N_13264,N_5681,N_5264);
nand U13265 (N_13265,N_7648,N_8162);
or U13266 (N_13266,N_9675,N_9950);
and U13267 (N_13267,N_5971,N_8457);
nand U13268 (N_13268,N_9550,N_8708);
xor U13269 (N_13269,N_9140,N_7535);
or U13270 (N_13270,N_6464,N_7650);
and U13271 (N_13271,N_9462,N_8617);
and U13272 (N_13272,N_5410,N_5949);
and U13273 (N_13273,N_7984,N_7027);
or U13274 (N_13274,N_5200,N_9635);
xnor U13275 (N_13275,N_9083,N_5451);
nor U13276 (N_13276,N_8490,N_5693);
nand U13277 (N_13277,N_8496,N_7286);
nor U13278 (N_13278,N_6717,N_5941);
nor U13279 (N_13279,N_5182,N_9735);
or U13280 (N_13280,N_8668,N_8407);
nor U13281 (N_13281,N_6167,N_6990);
nor U13282 (N_13282,N_6441,N_9448);
nor U13283 (N_13283,N_5571,N_5237);
or U13284 (N_13284,N_9035,N_9864);
xnor U13285 (N_13285,N_7911,N_8556);
nand U13286 (N_13286,N_5569,N_7031);
nor U13287 (N_13287,N_7108,N_7607);
xor U13288 (N_13288,N_9597,N_6446);
or U13289 (N_13289,N_6842,N_7649);
nand U13290 (N_13290,N_8434,N_6650);
xnor U13291 (N_13291,N_9774,N_7920);
and U13292 (N_13292,N_6602,N_5803);
nor U13293 (N_13293,N_9662,N_7308);
and U13294 (N_13294,N_9232,N_9700);
xor U13295 (N_13295,N_9918,N_7794);
xnor U13296 (N_13296,N_9554,N_5189);
nor U13297 (N_13297,N_5359,N_7680);
xnor U13298 (N_13298,N_8199,N_7704);
and U13299 (N_13299,N_9050,N_8954);
nand U13300 (N_13300,N_7223,N_5647);
nor U13301 (N_13301,N_9683,N_7248);
nor U13302 (N_13302,N_6520,N_5301);
nor U13303 (N_13303,N_9328,N_6410);
nor U13304 (N_13304,N_9883,N_7955);
nor U13305 (N_13305,N_9456,N_6079);
xnor U13306 (N_13306,N_6822,N_7279);
or U13307 (N_13307,N_9559,N_7231);
nand U13308 (N_13308,N_9993,N_5133);
nor U13309 (N_13309,N_7029,N_6336);
nand U13310 (N_13310,N_9899,N_8622);
and U13311 (N_13311,N_9199,N_8927);
or U13312 (N_13312,N_9737,N_7717);
or U13313 (N_13313,N_9399,N_5058);
and U13314 (N_13314,N_9625,N_6407);
nor U13315 (N_13315,N_7725,N_7343);
nand U13316 (N_13316,N_6988,N_5528);
nor U13317 (N_13317,N_5366,N_7451);
and U13318 (N_13318,N_6972,N_8371);
nor U13319 (N_13319,N_9518,N_9621);
nor U13320 (N_13320,N_5901,N_9719);
or U13321 (N_13321,N_9175,N_8879);
or U13322 (N_13322,N_5056,N_8174);
nand U13323 (N_13323,N_5844,N_6084);
and U13324 (N_13324,N_6179,N_9860);
nand U13325 (N_13325,N_5139,N_5680);
nand U13326 (N_13326,N_6284,N_6752);
nor U13327 (N_13327,N_6987,N_5750);
or U13328 (N_13328,N_7046,N_6655);
nand U13329 (N_13329,N_9047,N_9590);
and U13330 (N_13330,N_5448,N_9327);
nand U13331 (N_13331,N_5704,N_6713);
or U13332 (N_13332,N_5013,N_5982);
nand U13333 (N_13333,N_9181,N_9833);
nand U13334 (N_13334,N_6834,N_6751);
or U13335 (N_13335,N_9330,N_7807);
or U13336 (N_13336,N_6101,N_9212);
nor U13337 (N_13337,N_8566,N_8038);
nand U13338 (N_13338,N_8143,N_8327);
nor U13339 (N_13339,N_7977,N_8315);
or U13340 (N_13340,N_8993,N_9548);
nor U13341 (N_13341,N_9424,N_9044);
or U13342 (N_13342,N_6686,N_9925);
nor U13343 (N_13343,N_8895,N_9362);
nor U13344 (N_13344,N_7247,N_6830);
nand U13345 (N_13345,N_6147,N_8794);
nor U13346 (N_13346,N_7348,N_6001);
nor U13347 (N_13347,N_8544,N_6426);
and U13348 (N_13348,N_9670,N_9688);
nand U13349 (N_13349,N_7519,N_8183);
and U13350 (N_13350,N_9207,N_6943);
or U13351 (N_13351,N_6816,N_7644);
xnor U13352 (N_13352,N_8684,N_5122);
nor U13353 (N_13353,N_5517,N_8784);
nand U13354 (N_13354,N_7642,N_9761);
xnor U13355 (N_13355,N_8265,N_7997);
nand U13356 (N_13356,N_6421,N_6062);
or U13357 (N_13357,N_6265,N_9880);
xor U13358 (N_13358,N_5671,N_8725);
nand U13359 (N_13359,N_7478,N_6619);
or U13360 (N_13360,N_9171,N_5678);
nor U13361 (N_13361,N_6318,N_7225);
or U13362 (N_13362,N_7039,N_7203);
nor U13363 (N_13363,N_9655,N_8270);
and U13364 (N_13364,N_7775,N_8632);
or U13365 (N_13365,N_7381,N_6985);
and U13366 (N_13366,N_7893,N_9242);
nor U13367 (N_13367,N_8605,N_8898);
nand U13368 (N_13368,N_8573,N_5172);
and U13369 (N_13369,N_5394,N_9566);
xnor U13370 (N_13370,N_7047,N_6594);
or U13371 (N_13371,N_6515,N_9018);
nor U13372 (N_13372,N_8499,N_5747);
nor U13373 (N_13373,N_7430,N_7449);
nor U13374 (N_13374,N_5711,N_8443);
nand U13375 (N_13375,N_5358,N_6403);
nand U13376 (N_13376,N_5653,N_9240);
xor U13377 (N_13377,N_9496,N_6691);
or U13378 (N_13378,N_5437,N_5163);
or U13379 (N_13379,N_8981,N_5074);
nand U13380 (N_13380,N_8369,N_7331);
nand U13381 (N_13381,N_9942,N_8803);
nand U13382 (N_13382,N_7458,N_7247);
and U13383 (N_13383,N_7423,N_5743);
xnor U13384 (N_13384,N_7283,N_8075);
nor U13385 (N_13385,N_7945,N_9538);
and U13386 (N_13386,N_6624,N_8894);
and U13387 (N_13387,N_9468,N_5606);
xor U13388 (N_13388,N_8713,N_6938);
and U13389 (N_13389,N_9860,N_7763);
nor U13390 (N_13390,N_9686,N_8062);
and U13391 (N_13391,N_7575,N_6130);
or U13392 (N_13392,N_6249,N_7773);
nor U13393 (N_13393,N_9501,N_9243);
and U13394 (N_13394,N_9534,N_9799);
or U13395 (N_13395,N_5282,N_7792);
or U13396 (N_13396,N_5672,N_7846);
nor U13397 (N_13397,N_5794,N_6384);
nor U13398 (N_13398,N_8571,N_6750);
nand U13399 (N_13399,N_7490,N_9340);
nand U13400 (N_13400,N_9946,N_7399);
and U13401 (N_13401,N_6397,N_6274);
nor U13402 (N_13402,N_7699,N_8939);
nor U13403 (N_13403,N_8823,N_5379);
nor U13404 (N_13404,N_8207,N_6421);
and U13405 (N_13405,N_6430,N_8471);
or U13406 (N_13406,N_7065,N_8269);
nand U13407 (N_13407,N_9527,N_8788);
and U13408 (N_13408,N_5039,N_7659);
nand U13409 (N_13409,N_5336,N_6790);
nor U13410 (N_13410,N_8700,N_8648);
or U13411 (N_13411,N_6268,N_8532);
xor U13412 (N_13412,N_6162,N_8087);
nand U13413 (N_13413,N_9407,N_8622);
xor U13414 (N_13414,N_7502,N_5626);
and U13415 (N_13415,N_7414,N_7930);
nand U13416 (N_13416,N_6485,N_9966);
xnor U13417 (N_13417,N_8220,N_7504);
nand U13418 (N_13418,N_7912,N_7940);
or U13419 (N_13419,N_7239,N_6140);
and U13420 (N_13420,N_6992,N_5163);
nor U13421 (N_13421,N_6440,N_5982);
and U13422 (N_13422,N_7325,N_9893);
nand U13423 (N_13423,N_7218,N_5608);
and U13424 (N_13424,N_5319,N_9143);
and U13425 (N_13425,N_8320,N_8204);
and U13426 (N_13426,N_9413,N_7551);
xnor U13427 (N_13427,N_8834,N_5623);
xnor U13428 (N_13428,N_6135,N_7053);
or U13429 (N_13429,N_9597,N_6813);
nor U13430 (N_13430,N_6175,N_7190);
xor U13431 (N_13431,N_5045,N_9177);
nor U13432 (N_13432,N_9764,N_6375);
or U13433 (N_13433,N_5394,N_8229);
and U13434 (N_13434,N_5849,N_9053);
xnor U13435 (N_13435,N_6538,N_7883);
or U13436 (N_13436,N_7905,N_7516);
xor U13437 (N_13437,N_9560,N_9490);
nand U13438 (N_13438,N_7114,N_9992);
and U13439 (N_13439,N_7297,N_9533);
or U13440 (N_13440,N_5450,N_8230);
and U13441 (N_13441,N_7693,N_6926);
and U13442 (N_13442,N_7471,N_5832);
nand U13443 (N_13443,N_8304,N_8370);
nand U13444 (N_13444,N_6331,N_9731);
nand U13445 (N_13445,N_7773,N_6109);
and U13446 (N_13446,N_8196,N_8839);
nand U13447 (N_13447,N_7129,N_5575);
nand U13448 (N_13448,N_8610,N_6511);
nor U13449 (N_13449,N_5393,N_8075);
or U13450 (N_13450,N_5480,N_7240);
and U13451 (N_13451,N_6072,N_5665);
nor U13452 (N_13452,N_7391,N_8565);
nor U13453 (N_13453,N_7117,N_6540);
or U13454 (N_13454,N_7044,N_7042);
nor U13455 (N_13455,N_6616,N_6352);
and U13456 (N_13456,N_9843,N_9527);
xor U13457 (N_13457,N_8681,N_9591);
or U13458 (N_13458,N_8469,N_9921);
and U13459 (N_13459,N_6465,N_8038);
nand U13460 (N_13460,N_9671,N_6059);
nand U13461 (N_13461,N_5695,N_7187);
nor U13462 (N_13462,N_6676,N_9995);
xnor U13463 (N_13463,N_9491,N_7642);
or U13464 (N_13464,N_5775,N_7545);
xor U13465 (N_13465,N_8077,N_8794);
nor U13466 (N_13466,N_6167,N_6332);
nor U13467 (N_13467,N_9828,N_7764);
nand U13468 (N_13468,N_5448,N_9460);
nand U13469 (N_13469,N_6623,N_6385);
or U13470 (N_13470,N_7012,N_8309);
or U13471 (N_13471,N_9331,N_8364);
nor U13472 (N_13472,N_8851,N_6584);
and U13473 (N_13473,N_6761,N_9763);
or U13474 (N_13474,N_5011,N_9613);
nor U13475 (N_13475,N_8664,N_6581);
nor U13476 (N_13476,N_6853,N_5306);
or U13477 (N_13477,N_9764,N_6309);
and U13478 (N_13478,N_6359,N_8074);
nand U13479 (N_13479,N_5409,N_8769);
nor U13480 (N_13480,N_8751,N_8709);
nand U13481 (N_13481,N_9078,N_6299);
or U13482 (N_13482,N_9131,N_8790);
nor U13483 (N_13483,N_8477,N_6727);
nor U13484 (N_13484,N_8363,N_5158);
and U13485 (N_13485,N_5576,N_8104);
or U13486 (N_13486,N_9938,N_7506);
nor U13487 (N_13487,N_7624,N_7173);
or U13488 (N_13488,N_9745,N_8682);
and U13489 (N_13489,N_7236,N_9169);
xnor U13490 (N_13490,N_8118,N_7988);
or U13491 (N_13491,N_8488,N_5139);
or U13492 (N_13492,N_9254,N_8223);
xnor U13493 (N_13493,N_8631,N_6942);
or U13494 (N_13494,N_8278,N_9488);
nor U13495 (N_13495,N_7141,N_5017);
nor U13496 (N_13496,N_8365,N_9295);
nor U13497 (N_13497,N_5636,N_7834);
nor U13498 (N_13498,N_7821,N_5318);
nand U13499 (N_13499,N_6943,N_6750);
nor U13500 (N_13500,N_8230,N_6498);
nor U13501 (N_13501,N_5391,N_8289);
or U13502 (N_13502,N_7523,N_6805);
or U13503 (N_13503,N_8630,N_9595);
and U13504 (N_13504,N_9768,N_9069);
nand U13505 (N_13505,N_7956,N_6656);
nand U13506 (N_13506,N_8907,N_7442);
and U13507 (N_13507,N_8008,N_7300);
nor U13508 (N_13508,N_7897,N_8369);
nand U13509 (N_13509,N_9898,N_7223);
xor U13510 (N_13510,N_6910,N_5085);
nand U13511 (N_13511,N_6556,N_5829);
and U13512 (N_13512,N_6006,N_7684);
or U13513 (N_13513,N_6689,N_9158);
and U13514 (N_13514,N_6408,N_7454);
and U13515 (N_13515,N_7557,N_5957);
xnor U13516 (N_13516,N_9017,N_9843);
or U13517 (N_13517,N_7024,N_6536);
nand U13518 (N_13518,N_5706,N_8672);
or U13519 (N_13519,N_9162,N_9053);
nand U13520 (N_13520,N_5368,N_8430);
xnor U13521 (N_13521,N_8306,N_9872);
or U13522 (N_13522,N_5650,N_5509);
nor U13523 (N_13523,N_6055,N_6151);
and U13524 (N_13524,N_7632,N_5373);
nor U13525 (N_13525,N_9039,N_9643);
nand U13526 (N_13526,N_8122,N_8087);
nand U13527 (N_13527,N_7223,N_9536);
nor U13528 (N_13528,N_5578,N_5567);
nand U13529 (N_13529,N_9075,N_9427);
or U13530 (N_13530,N_9753,N_5266);
nor U13531 (N_13531,N_6097,N_6083);
nand U13532 (N_13532,N_7286,N_9973);
nand U13533 (N_13533,N_5831,N_8900);
or U13534 (N_13534,N_6398,N_9275);
nor U13535 (N_13535,N_8395,N_6777);
or U13536 (N_13536,N_8394,N_6428);
or U13537 (N_13537,N_9541,N_9084);
nor U13538 (N_13538,N_8638,N_8991);
nand U13539 (N_13539,N_8738,N_6742);
nor U13540 (N_13540,N_8353,N_8435);
and U13541 (N_13541,N_8995,N_6060);
and U13542 (N_13542,N_9611,N_9031);
nand U13543 (N_13543,N_8770,N_5743);
nor U13544 (N_13544,N_9448,N_7538);
nor U13545 (N_13545,N_5529,N_6185);
and U13546 (N_13546,N_6714,N_6850);
nor U13547 (N_13547,N_7427,N_8156);
xor U13548 (N_13548,N_5666,N_8260);
or U13549 (N_13549,N_6714,N_9433);
or U13550 (N_13550,N_6571,N_8135);
nand U13551 (N_13551,N_5826,N_7322);
or U13552 (N_13552,N_5049,N_8072);
nand U13553 (N_13553,N_5314,N_7740);
xnor U13554 (N_13554,N_6628,N_5354);
nor U13555 (N_13555,N_9430,N_5726);
and U13556 (N_13556,N_9027,N_6021);
xnor U13557 (N_13557,N_8818,N_7928);
and U13558 (N_13558,N_5314,N_9325);
or U13559 (N_13559,N_5890,N_6811);
xnor U13560 (N_13560,N_5091,N_8161);
or U13561 (N_13561,N_8743,N_6825);
or U13562 (N_13562,N_5096,N_5805);
nor U13563 (N_13563,N_8589,N_5857);
or U13564 (N_13564,N_5485,N_9032);
nand U13565 (N_13565,N_8126,N_8045);
nor U13566 (N_13566,N_7257,N_7441);
and U13567 (N_13567,N_8969,N_8966);
nand U13568 (N_13568,N_8401,N_6248);
nand U13569 (N_13569,N_5733,N_8629);
or U13570 (N_13570,N_5730,N_5594);
and U13571 (N_13571,N_5112,N_7914);
nor U13572 (N_13572,N_7817,N_8247);
nor U13573 (N_13573,N_6219,N_6153);
xor U13574 (N_13574,N_8525,N_6373);
nand U13575 (N_13575,N_9656,N_8634);
nand U13576 (N_13576,N_5378,N_9641);
or U13577 (N_13577,N_6332,N_9992);
and U13578 (N_13578,N_5438,N_8374);
nor U13579 (N_13579,N_8960,N_9057);
or U13580 (N_13580,N_7202,N_7638);
and U13581 (N_13581,N_8718,N_9106);
xor U13582 (N_13582,N_5383,N_5170);
or U13583 (N_13583,N_6401,N_7295);
or U13584 (N_13584,N_6848,N_6458);
and U13585 (N_13585,N_5755,N_9666);
or U13586 (N_13586,N_6494,N_7835);
and U13587 (N_13587,N_5652,N_7852);
nand U13588 (N_13588,N_8588,N_8453);
nand U13589 (N_13589,N_9339,N_7206);
nor U13590 (N_13590,N_7584,N_5141);
xor U13591 (N_13591,N_8624,N_9771);
and U13592 (N_13592,N_5430,N_5774);
or U13593 (N_13593,N_6642,N_7529);
nand U13594 (N_13594,N_9353,N_7526);
or U13595 (N_13595,N_5924,N_9221);
nor U13596 (N_13596,N_5551,N_8318);
or U13597 (N_13597,N_6342,N_6638);
nor U13598 (N_13598,N_6612,N_9862);
nand U13599 (N_13599,N_8660,N_9587);
and U13600 (N_13600,N_7650,N_9552);
nor U13601 (N_13601,N_7639,N_9160);
nand U13602 (N_13602,N_5489,N_8761);
and U13603 (N_13603,N_5933,N_5508);
nor U13604 (N_13604,N_8034,N_6854);
nor U13605 (N_13605,N_6202,N_9483);
or U13606 (N_13606,N_9771,N_9351);
nor U13607 (N_13607,N_5786,N_5560);
and U13608 (N_13608,N_7030,N_8418);
and U13609 (N_13609,N_9775,N_9046);
xnor U13610 (N_13610,N_9807,N_8844);
xor U13611 (N_13611,N_5304,N_5246);
xor U13612 (N_13612,N_8616,N_7211);
or U13613 (N_13613,N_9857,N_8757);
nor U13614 (N_13614,N_8205,N_8730);
nand U13615 (N_13615,N_5270,N_9266);
nor U13616 (N_13616,N_8201,N_9435);
or U13617 (N_13617,N_8700,N_7903);
nand U13618 (N_13618,N_7455,N_7872);
nor U13619 (N_13619,N_8366,N_7901);
or U13620 (N_13620,N_9524,N_5332);
and U13621 (N_13621,N_8356,N_5723);
nand U13622 (N_13622,N_9902,N_7264);
nor U13623 (N_13623,N_9379,N_6738);
and U13624 (N_13624,N_9498,N_9637);
nor U13625 (N_13625,N_6801,N_6170);
nand U13626 (N_13626,N_8492,N_9022);
nor U13627 (N_13627,N_5291,N_8630);
xor U13628 (N_13628,N_5440,N_6086);
or U13629 (N_13629,N_7749,N_9875);
nor U13630 (N_13630,N_6714,N_7798);
nand U13631 (N_13631,N_8235,N_7242);
nand U13632 (N_13632,N_6695,N_6168);
and U13633 (N_13633,N_9934,N_8049);
and U13634 (N_13634,N_5976,N_8392);
nand U13635 (N_13635,N_8665,N_9490);
and U13636 (N_13636,N_7203,N_7685);
nand U13637 (N_13637,N_7102,N_5167);
nor U13638 (N_13638,N_9731,N_6221);
or U13639 (N_13639,N_5483,N_6438);
and U13640 (N_13640,N_5626,N_8190);
or U13641 (N_13641,N_5496,N_6503);
nand U13642 (N_13642,N_6348,N_6764);
or U13643 (N_13643,N_8737,N_6410);
nor U13644 (N_13644,N_6946,N_9175);
and U13645 (N_13645,N_8487,N_8177);
nand U13646 (N_13646,N_7185,N_7547);
or U13647 (N_13647,N_6773,N_8441);
nor U13648 (N_13648,N_9570,N_5474);
and U13649 (N_13649,N_8156,N_8594);
nand U13650 (N_13650,N_7024,N_6138);
or U13651 (N_13651,N_8111,N_7237);
or U13652 (N_13652,N_9016,N_9969);
nand U13653 (N_13653,N_8334,N_6711);
or U13654 (N_13654,N_7588,N_8762);
nand U13655 (N_13655,N_7985,N_6179);
nand U13656 (N_13656,N_9527,N_9294);
and U13657 (N_13657,N_9659,N_9447);
and U13658 (N_13658,N_8850,N_8719);
nand U13659 (N_13659,N_8433,N_9300);
nand U13660 (N_13660,N_7645,N_9616);
nor U13661 (N_13661,N_5420,N_5886);
and U13662 (N_13662,N_8155,N_6356);
nand U13663 (N_13663,N_7686,N_5722);
nand U13664 (N_13664,N_6030,N_6244);
and U13665 (N_13665,N_7285,N_6321);
or U13666 (N_13666,N_9885,N_5231);
nand U13667 (N_13667,N_7207,N_5718);
nor U13668 (N_13668,N_7785,N_7766);
and U13669 (N_13669,N_6336,N_8113);
nand U13670 (N_13670,N_7232,N_8188);
or U13671 (N_13671,N_5917,N_9777);
nand U13672 (N_13672,N_9433,N_8344);
nand U13673 (N_13673,N_9034,N_9012);
or U13674 (N_13674,N_7823,N_9625);
nand U13675 (N_13675,N_5813,N_6229);
xor U13676 (N_13676,N_6340,N_9521);
and U13677 (N_13677,N_8302,N_7725);
and U13678 (N_13678,N_8053,N_7384);
or U13679 (N_13679,N_5393,N_8493);
nor U13680 (N_13680,N_8148,N_8473);
nor U13681 (N_13681,N_7439,N_8819);
nor U13682 (N_13682,N_7462,N_6859);
or U13683 (N_13683,N_5267,N_9200);
xnor U13684 (N_13684,N_7749,N_7484);
xnor U13685 (N_13685,N_6454,N_6082);
xor U13686 (N_13686,N_6859,N_8470);
nor U13687 (N_13687,N_7399,N_6762);
or U13688 (N_13688,N_8289,N_7627);
and U13689 (N_13689,N_5924,N_5409);
nand U13690 (N_13690,N_9349,N_8498);
nor U13691 (N_13691,N_8271,N_8291);
xnor U13692 (N_13692,N_8489,N_5098);
nand U13693 (N_13693,N_9007,N_6210);
nor U13694 (N_13694,N_6484,N_7915);
or U13695 (N_13695,N_7886,N_8741);
nand U13696 (N_13696,N_8915,N_9451);
or U13697 (N_13697,N_5247,N_6683);
nor U13698 (N_13698,N_5801,N_7887);
nand U13699 (N_13699,N_7126,N_7680);
nor U13700 (N_13700,N_7691,N_5201);
and U13701 (N_13701,N_7809,N_8749);
nor U13702 (N_13702,N_7344,N_9669);
and U13703 (N_13703,N_9388,N_7061);
nand U13704 (N_13704,N_7332,N_9503);
nor U13705 (N_13705,N_9693,N_8598);
nand U13706 (N_13706,N_7919,N_7771);
or U13707 (N_13707,N_5873,N_8709);
nor U13708 (N_13708,N_7188,N_6243);
nor U13709 (N_13709,N_6547,N_9864);
xnor U13710 (N_13710,N_6928,N_8973);
nand U13711 (N_13711,N_6939,N_9936);
and U13712 (N_13712,N_9958,N_5651);
or U13713 (N_13713,N_8233,N_6025);
or U13714 (N_13714,N_7307,N_8320);
and U13715 (N_13715,N_7072,N_8963);
nand U13716 (N_13716,N_9699,N_5631);
or U13717 (N_13717,N_5628,N_5832);
nand U13718 (N_13718,N_5069,N_6174);
and U13719 (N_13719,N_5807,N_8977);
or U13720 (N_13720,N_6337,N_7887);
and U13721 (N_13721,N_6048,N_8358);
nand U13722 (N_13722,N_7140,N_5349);
nand U13723 (N_13723,N_8684,N_5921);
and U13724 (N_13724,N_5660,N_5690);
xnor U13725 (N_13725,N_5173,N_9941);
or U13726 (N_13726,N_6252,N_7003);
and U13727 (N_13727,N_6124,N_9242);
and U13728 (N_13728,N_8245,N_6030);
and U13729 (N_13729,N_8749,N_5165);
and U13730 (N_13730,N_9953,N_8490);
and U13731 (N_13731,N_6405,N_9213);
and U13732 (N_13732,N_9911,N_8218);
nor U13733 (N_13733,N_9050,N_8118);
or U13734 (N_13734,N_6194,N_7882);
or U13735 (N_13735,N_9259,N_6976);
and U13736 (N_13736,N_5923,N_7762);
nor U13737 (N_13737,N_8672,N_9669);
and U13738 (N_13738,N_7903,N_5740);
nand U13739 (N_13739,N_7547,N_9521);
nand U13740 (N_13740,N_7973,N_5536);
nand U13741 (N_13741,N_9328,N_9758);
xnor U13742 (N_13742,N_8663,N_7126);
and U13743 (N_13743,N_5486,N_6143);
nor U13744 (N_13744,N_5495,N_5034);
or U13745 (N_13745,N_6684,N_7955);
nor U13746 (N_13746,N_8690,N_8734);
or U13747 (N_13747,N_8394,N_9548);
or U13748 (N_13748,N_7139,N_6992);
and U13749 (N_13749,N_7538,N_6469);
nor U13750 (N_13750,N_8286,N_6434);
or U13751 (N_13751,N_7139,N_6941);
or U13752 (N_13752,N_5334,N_6754);
nor U13753 (N_13753,N_7691,N_7145);
xnor U13754 (N_13754,N_5213,N_6133);
nand U13755 (N_13755,N_9575,N_8779);
xor U13756 (N_13756,N_6339,N_8855);
and U13757 (N_13757,N_6773,N_8928);
xnor U13758 (N_13758,N_8259,N_8832);
and U13759 (N_13759,N_7757,N_6871);
or U13760 (N_13760,N_5337,N_5479);
and U13761 (N_13761,N_6532,N_8074);
and U13762 (N_13762,N_8223,N_9782);
or U13763 (N_13763,N_8290,N_5953);
or U13764 (N_13764,N_5408,N_5221);
xor U13765 (N_13765,N_9158,N_5774);
nand U13766 (N_13766,N_9602,N_6272);
and U13767 (N_13767,N_7570,N_8729);
nand U13768 (N_13768,N_5925,N_6586);
or U13769 (N_13769,N_8990,N_6539);
or U13770 (N_13770,N_8940,N_6905);
or U13771 (N_13771,N_5421,N_8590);
or U13772 (N_13772,N_9493,N_8969);
or U13773 (N_13773,N_9987,N_9235);
nand U13774 (N_13774,N_8366,N_9532);
or U13775 (N_13775,N_7566,N_7516);
or U13776 (N_13776,N_6113,N_5061);
or U13777 (N_13777,N_6215,N_5980);
and U13778 (N_13778,N_6549,N_8333);
nor U13779 (N_13779,N_8109,N_6668);
nor U13780 (N_13780,N_5355,N_9397);
nor U13781 (N_13781,N_8511,N_6367);
nor U13782 (N_13782,N_7364,N_8806);
nor U13783 (N_13783,N_6031,N_5244);
and U13784 (N_13784,N_6114,N_5307);
nor U13785 (N_13785,N_8898,N_5180);
and U13786 (N_13786,N_5227,N_6820);
nor U13787 (N_13787,N_6274,N_7530);
and U13788 (N_13788,N_5585,N_8321);
nand U13789 (N_13789,N_7822,N_7387);
nor U13790 (N_13790,N_7063,N_5351);
or U13791 (N_13791,N_5822,N_7758);
xnor U13792 (N_13792,N_5135,N_8204);
nor U13793 (N_13793,N_8835,N_6568);
and U13794 (N_13794,N_9399,N_5088);
or U13795 (N_13795,N_8660,N_5052);
nand U13796 (N_13796,N_8620,N_5822);
nor U13797 (N_13797,N_6521,N_7430);
nor U13798 (N_13798,N_8435,N_9975);
and U13799 (N_13799,N_8136,N_8246);
or U13800 (N_13800,N_7621,N_8364);
nor U13801 (N_13801,N_7931,N_6904);
nand U13802 (N_13802,N_8912,N_9811);
and U13803 (N_13803,N_9216,N_7277);
nand U13804 (N_13804,N_9925,N_6856);
nand U13805 (N_13805,N_6069,N_7580);
nand U13806 (N_13806,N_8879,N_6430);
nor U13807 (N_13807,N_8507,N_6940);
or U13808 (N_13808,N_9351,N_7141);
nor U13809 (N_13809,N_6588,N_9921);
nand U13810 (N_13810,N_8774,N_8903);
and U13811 (N_13811,N_9757,N_7813);
nor U13812 (N_13812,N_6888,N_7597);
nand U13813 (N_13813,N_7083,N_8197);
or U13814 (N_13814,N_8108,N_5564);
nor U13815 (N_13815,N_7366,N_6830);
nor U13816 (N_13816,N_7649,N_7563);
xor U13817 (N_13817,N_7644,N_9370);
and U13818 (N_13818,N_7654,N_8845);
xor U13819 (N_13819,N_6375,N_9896);
and U13820 (N_13820,N_7777,N_7194);
nand U13821 (N_13821,N_9869,N_7281);
nand U13822 (N_13822,N_8943,N_7384);
or U13823 (N_13823,N_8227,N_6472);
xor U13824 (N_13824,N_5926,N_9234);
or U13825 (N_13825,N_9183,N_6733);
or U13826 (N_13826,N_7883,N_6268);
nor U13827 (N_13827,N_7894,N_5511);
and U13828 (N_13828,N_5140,N_5641);
or U13829 (N_13829,N_7691,N_8858);
xnor U13830 (N_13830,N_9451,N_6807);
xnor U13831 (N_13831,N_6719,N_9361);
and U13832 (N_13832,N_9752,N_5516);
nor U13833 (N_13833,N_5056,N_9153);
and U13834 (N_13834,N_5764,N_8479);
nand U13835 (N_13835,N_7884,N_9955);
or U13836 (N_13836,N_8944,N_7381);
nand U13837 (N_13837,N_5194,N_6080);
nand U13838 (N_13838,N_5704,N_7873);
nor U13839 (N_13839,N_5959,N_6033);
nor U13840 (N_13840,N_8275,N_5512);
nor U13841 (N_13841,N_8573,N_8220);
or U13842 (N_13842,N_9595,N_6989);
and U13843 (N_13843,N_6758,N_6149);
xor U13844 (N_13844,N_7920,N_8322);
or U13845 (N_13845,N_6986,N_9467);
nor U13846 (N_13846,N_9214,N_8977);
or U13847 (N_13847,N_6668,N_6143);
xor U13848 (N_13848,N_8857,N_7908);
and U13849 (N_13849,N_7582,N_5464);
nand U13850 (N_13850,N_8540,N_6672);
or U13851 (N_13851,N_7866,N_6280);
and U13852 (N_13852,N_5424,N_9307);
nor U13853 (N_13853,N_9447,N_9888);
xnor U13854 (N_13854,N_8755,N_8761);
or U13855 (N_13855,N_7412,N_8667);
and U13856 (N_13856,N_9947,N_9100);
nor U13857 (N_13857,N_7896,N_9002);
and U13858 (N_13858,N_8934,N_8396);
or U13859 (N_13859,N_6348,N_8480);
nand U13860 (N_13860,N_6725,N_6216);
or U13861 (N_13861,N_7766,N_7591);
or U13862 (N_13862,N_9935,N_8128);
nand U13863 (N_13863,N_7132,N_9048);
or U13864 (N_13864,N_6697,N_9238);
nand U13865 (N_13865,N_9177,N_9520);
and U13866 (N_13866,N_9148,N_5576);
or U13867 (N_13867,N_9253,N_9429);
xnor U13868 (N_13868,N_7283,N_7400);
nand U13869 (N_13869,N_6347,N_7818);
nand U13870 (N_13870,N_8314,N_5891);
or U13871 (N_13871,N_8955,N_6246);
nor U13872 (N_13872,N_9752,N_8272);
xnor U13873 (N_13873,N_5117,N_7731);
or U13874 (N_13874,N_6887,N_9699);
and U13875 (N_13875,N_6844,N_9364);
and U13876 (N_13876,N_5020,N_7752);
or U13877 (N_13877,N_5114,N_9348);
or U13878 (N_13878,N_8177,N_7579);
xor U13879 (N_13879,N_6200,N_8269);
xnor U13880 (N_13880,N_8991,N_5310);
or U13881 (N_13881,N_5297,N_7751);
nand U13882 (N_13882,N_9658,N_8014);
nor U13883 (N_13883,N_7713,N_9467);
or U13884 (N_13884,N_6642,N_5371);
or U13885 (N_13885,N_5368,N_5920);
or U13886 (N_13886,N_9507,N_7160);
or U13887 (N_13887,N_9348,N_6041);
nand U13888 (N_13888,N_6038,N_8095);
or U13889 (N_13889,N_6064,N_6798);
nor U13890 (N_13890,N_6703,N_8009);
nand U13891 (N_13891,N_9228,N_6116);
nand U13892 (N_13892,N_8089,N_8398);
nor U13893 (N_13893,N_8578,N_5781);
and U13894 (N_13894,N_5216,N_9535);
nor U13895 (N_13895,N_7878,N_9676);
nand U13896 (N_13896,N_8889,N_8696);
nand U13897 (N_13897,N_5446,N_6267);
nand U13898 (N_13898,N_5512,N_9147);
or U13899 (N_13899,N_5080,N_5320);
nor U13900 (N_13900,N_5864,N_8550);
xor U13901 (N_13901,N_6905,N_6936);
or U13902 (N_13902,N_8100,N_8384);
nand U13903 (N_13903,N_9358,N_9990);
or U13904 (N_13904,N_9875,N_6944);
xor U13905 (N_13905,N_7468,N_6451);
nand U13906 (N_13906,N_8297,N_5118);
nand U13907 (N_13907,N_9868,N_8298);
and U13908 (N_13908,N_8643,N_8809);
nor U13909 (N_13909,N_7555,N_5701);
and U13910 (N_13910,N_8783,N_8424);
nor U13911 (N_13911,N_5931,N_9844);
nand U13912 (N_13912,N_5768,N_8780);
or U13913 (N_13913,N_5886,N_9780);
nand U13914 (N_13914,N_8210,N_8562);
nand U13915 (N_13915,N_8047,N_5292);
nand U13916 (N_13916,N_7712,N_7822);
or U13917 (N_13917,N_5744,N_5141);
or U13918 (N_13918,N_6918,N_5770);
or U13919 (N_13919,N_8088,N_5996);
nand U13920 (N_13920,N_7898,N_5012);
xor U13921 (N_13921,N_7363,N_6889);
nor U13922 (N_13922,N_7917,N_7159);
and U13923 (N_13923,N_9468,N_9541);
or U13924 (N_13924,N_6940,N_7660);
nor U13925 (N_13925,N_8589,N_5328);
xor U13926 (N_13926,N_6574,N_5218);
and U13927 (N_13927,N_8456,N_7221);
nor U13928 (N_13928,N_5322,N_8184);
nand U13929 (N_13929,N_6484,N_8520);
nor U13930 (N_13930,N_8749,N_9736);
nor U13931 (N_13931,N_6533,N_5077);
or U13932 (N_13932,N_5527,N_9046);
nand U13933 (N_13933,N_8194,N_9594);
nor U13934 (N_13934,N_5125,N_5105);
and U13935 (N_13935,N_5241,N_6951);
and U13936 (N_13936,N_6010,N_7811);
and U13937 (N_13937,N_9682,N_7515);
and U13938 (N_13938,N_9744,N_9800);
nand U13939 (N_13939,N_8365,N_8221);
nor U13940 (N_13940,N_6439,N_5671);
nor U13941 (N_13941,N_6368,N_8021);
and U13942 (N_13942,N_8139,N_9457);
and U13943 (N_13943,N_5205,N_9611);
or U13944 (N_13944,N_8202,N_6336);
nand U13945 (N_13945,N_9598,N_8814);
or U13946 (N_13946,N_6606,N_8286);
and U13947 (N_13947,N_6207,N_9887);
nand U13948 (N_13948,N_5000,N_8392);
and U13949 (N_13949,N_7547,N_9844);
nand U13950 (N_13950,N_8272,N_8532);
or U13951 (N_13951,N_9903,N_7374);
and U13952 (N_13952,N_9597,N_6003);
and U13953 (N_13953,N_9642,N_9019);
or U13954 (N_13954,N_5400,N_5771);
and U13955 (N_13955,N_5106,N_8867);
nand U13956 (N_13956,N_8246,N_9839);
nor U13957 (N_13957,N_8107,N_7020);
xor U13958 (N_13958,N_8750,N_5689);
nand U13959 (N_13959,N_5244,N_8298);
and U13960 (N_13960,N_9401,N_7491);
xor U13961 (N_13961,N_9365,N_8546);
nor U13962 (N_13962,N_5541,N_5004);
and U13963 (N_13963,N_5379,N_9545);
or U13964 (N_13964,N_7364,N_7653);
nand U13965 (N_13965,N_5372,N_6293);
or U13966 (N_13966,N_6151,N_5331);
nor U13967 (N_13967,N_7194,N_5402);
or U13968 (N_13968,N_9952,N_5385);
or U13969 (N_13969,N_6835,N_9142);
nand U13970 (N_13970,N_5350,N_8136);
or U13971 (N_13971,N_5958,N_6367);
nand U13972 (N_13972,N_7276,N_8923);
xnor U13973 (N_13973,N_9225,N_9188);
and U13974 (N_13974,N_8635,N_8628);
nand U13975 (N_13975,N_5760,N_8191);
nor U13976 (N_13976,N_9995,N_7857);
nor U13977 (N_13977,N_5171,N_5324);
nor U13978 (N_13978,N_8957,N_6824);
and U13979 (N_13979,N_8362,N_7731);
nand U13980 (N_13980,N_6519,N_5690);
xnor U13981 (N_13981,N_8032,N_6131);
and U13982 (N_13982,N_6745,N_9895);
or U13983 (N_13983,N_8535,N_6615);
nor U13984 (N_13984,N_7793,N_5924);
nand U13985 (N_13985,N_8651,N_6355);
nand U13986 (N_13986,N_6896,N_5542);
and U13987 (N_13987,N_7470,N_9311);
nor U13988 (N_13988,N_7852,N_6231);
and U13989 (N_13989,N_6200,N_5737);
or U13990 (N_13990,N_6663,N_8510);
nor U13991 (N_13991,N_8676,N_7208);
xor U13992 (N_13992,N_9933,N_8496);
nand U13993 (N_13993,N_7736,N_5607);
and U13994 (N_13994,N_7671,N_8589);
or U13995 (N_13995,N_9095,N_5975);
xnor U13996 (N_13996,N_9837,N_8929);
nand U13997 (N_13997,N_7050,N_8963);
and U13998 (N_13998,N_6891,N_5043);
xnor U13999 (N_13999,N_9105,N_8687);
and U14000 (N_14000,N_7513,N_9569);
or U14001 (N_14001,N_9953,N_6762);
and U14002 (N_14002,N_6693,N_7068);
nand U14003 (N_14003,N_5948,N_7804);
and U14004 (N_14004,N_7283,N_6746);
nand U14005 (N_14005,N_7697,N_5234);
or U14006 (N_14006,N_7452,N_6497);
nand U14007 (N_14007,N_7335,N_5921);
or U14008 (N_14008,N_7368,N_9161);
nor U14009 (N_14009,N_9699,N_5195);
and U14010 (N_14010,N_6020,N_8999);
nand U14011 (N_14011,N_8714,N_5056);
or U14012 (N_14012,N_5784,N_9743);
nand U14013 (N_14013,N_8318,N_8060);
nand U14014 (N_14014,N_7945,N_8922);
and U14015 (N_14015,N_7744,N_6492);
nand U14016 (N_14016,N_8002,N_5555);
or U14017 (N_14017,N_5140,N_6751);
or U14018 (N_14018,N_9294,N_8908);
and U14019 (N_14019,N_8829,N_6172);
and U14020 (N_14020,N_7920,N_5542);
and U14021 (N_14021,N_7015,N_5454);
nor U14022 (N_14022,N_8964,N_9250);
nor U14023 (N_14023,N_9656,N_6832);
xnor U14024 (N_14024,N_8478,N_8528);
or U14025 (N_14025,N_9640,N_8248);
or U14026 (N_14026,N_9085,N_8162);
or U14027 (N_14027,N_6093,N_8072);
or U14028 (N_14028,N_9869,N_8506);
or U14029 (N_14029,N_6814,N_7955);
or U14030 (N_14030,N_7790,N_6571);
nand U14031 (N_14031,N_5062,N_6846);
and U14032 (N_14032,N_8411,N_9483);
nor U14033 (N_14033,N_9789,N_8771);
or U14034 (N_14034,N_6589,N_6231);
nand U14035 (N_14035,N_5893,N_5703);
nand U14036 (N_14036,N_6447,N_6425);
or U14037 (N_14037,N_8519,N_5481);
nor U14038 (N_14038,N_6504,N_7609);
or U14039 (N_14039,N_8312,N_6908);
or U14040 (N_14040,N_7745,N_7885);
nand U14041 (N_14041,N_5064,N_7821);
and U14042 (N_14042,N_7070,N_5706);
and U14043 (N_14043,N_9757,N_5205);
nor U14044 (N_14044,N_8981,N_9081);
or U14045 (N_14045,N_8982,N_9668);
nand U14046 (N_14046,N_5636,N_7571);
or U14047 (N_14047,N_9692,N_8108);
nor U14048 (N_14048,N_5168,N_8035);
and U14049 (N_14049,N_8635,N_8505);
and U14050 (N_14050,N_7790,N_7449);
xor U14051 (N_14051,N_7598,N_7736);
or U14052 (N_14052,N_8217,N_8436);
xnor U14053 (N_14053,N_8903,N_6053);
and U14054 (N_14054,N_8609,N_6436);
or U14055 (N_14055,N_6819,N_8560);
nor U14056 (N_14056,N_8563,N_9297);
or U14057 (N_14057,N_6377,N_6461);
nand U14058 (N_14058,N_8759,N_5534);
or U14059 (N_14059,N_7971,N_9841);
nor U14060 (N_14060,N_8995,N_6456);
and U14061 (N_14061,N_7475,N_6323);
and U14062 (N_14062,N_7292,N_5153);
and U14063 (N_14063,N_7169,N_7906);
or U14064 (N_14064,N_8545,N_6817);
nand U14065 (N_14065,N_9505,N_9626);
nor U14066 (N_14066,N_6133,N_5077);
nor U14067 (N_14067,N_6313,N_5332);
nand U14068 (N_14068,N_9064,N_7432);
nor U14069 (N_14069,N_6959,N_7767);
nor U14070 (N_14070,N_5822,N_6271);
xnor U14071 (N_14071,N_6529,N_7822);
or U14072 (N_14072,N_9405,N_5322);
nor U14073 (N_14073,N_8396,N_5748);
nor U14074 (N_14074,N_7221,N_8116);
or U14075 (N_14075,N_5572,N_9904);
nand U14076 (N_14076,N_8350,N_9011);
nor U14077 (N_14077,N_8267,N_6712);
and U14078 (N_14078,N_8635,N_7840);
nor U14079 (N_14079,N_5202,N_8797);
or U14080 (N_14080,N_7139,N_7434);
nor U14081 (N_14081,N_7434,N_7015);
nor U14082 (N_14082,N_9083,N_9505);
nor U14083 (N_14083,N_5231,N_6470);
and U14084 (N_14084,N_8866,N_8051);
and U14085 (N_14085,N_6567,N_7136);
nand U14086 (N_14086,N_5663,N_8472);
and U14087 (N_14087,N_8042,N_9537);
nand U14088 (N_14088,N_5910,N_8909);
and U14089 (N_14089,N_9599,N_7122);
or U14090 (N_14090,N_7540,N_7041);
and U14091 (N_14091,N_9457,N_6125);
nand U14092 (N_14092,N_7704,N_5893);
nor U14093 (N_14093,N_5037,N_6239);
or U14094 (N_14094,N_7380,N_5954);
and U14095 (N_14095,N_6246,N_8212);
and U14096 (N_14096,N_6942,N_9603);
nor U14097 (N_14097,N_7525,N_9515);
nor U14098 (N_14098,N_8466,N_7915);
xnor U14099 (N_14099,N_8799,N_5365);
and U14100 (N_14100,N_8297,N_8066);
nor U14101 (N_14101,N_5128,N_7678);
nor U14102 (N_14102,N_9902,N_7418);
or U14103 (N_14103,N_7691,N_6195);
and U14104 (N_14104,N_8869,N_5042);
or U14105 (N_14105,N_6520,N_8340);
xnor U14106 (N_14106,N_8231,N_7683);
or U14107 (N_14107,N_5299,N_7792);
nor U14108 (N_14108,N_7833,N_9348);
nand U14109 (N_14109,N_8990,N_8678);
and U14110 (N_14110,N_8180,N_8328);
nor U14111 (N_14111,N_7349,N_6829);
and U14112 (N_14112,N_6558,N_9590);
or U14113 (N_14113,N_9793,N_5343);
and U14114 (N_14114,N_5778,N_7682);
or U14115 (N_14115,N_7715,N_7464);
nor U14116 (N_14116,N_6763,N_5255);
nand U14117 (N_14117,N_7525,N_5306);
or U14118 (N_14118,N_6098,N_7511);
or U14119 (N_14119,N_7140,N_9317);
and U14120 (N_14120,N_8533,N_9335);
nor U14121 (N_14121,N_5217,N_6123);
and U14122 (N_14122,N_5904,N_7362);
nand U14123 (N_14123,N_6017,N_7964);
nand U14124 (N_14124,N_5544,N_6823);
xnor U14125 (N_14125,N_7301,N_8778);
nor U14126 (N_14126,N_7614,N_6183);
or U14127 (N_14127,N_6478,N_5646);
and U14128 (N_14128,N_9795,N_8220);
nand U14129 (N_14129,N_6386,N_7815);
xnor U14130 (N_14130,N_6021,N_9015);
xnor U14131 (N_14131,N_6188,N_8195);
and U14132 (N_14132,N_5860,N_6891);
and U14133 (N_14133,N_6434,N_6084);
nand U14134 (N_14134,N_8041,N_8153);
xor U14135 (N_14135,N_8132,N_8768);
nor U14136 (N_14136,N_9993,N_8992);
and U14137 (N_14137,N_7608,N_6925);
or U14138 (N_14138,N_8133,N_8205);
xor U14139 (N_14139,N_9117,N_6563);
and U14140 (N_14140,N_8768,N_9379);
nand U14141 (N_14141,N_7653,N_7067);
nor U14142 (N_14142,N_9306,N_7766);
or U14143 (N_14143,N_5789,N_8944);
or U14144 (N_14144,N_8438,N_6783);
and U14145 (N_14145,N_5472,N_6377);
or U14146 (N_14146,N_9398,N_6280);
and U14147 (N_14147,N_7054,N_5936);
and U14148 (N_14148,N_9721,N_9400);
or U14149 (N_14149,N_8923,N_9060);
nand U14150 (N_14150,N_6365,N_7104);
xnor U14151 (N_14151,N_5587,N_8727);
or U14152 (N_14152,N_6465,N_7839);
xor U14153 (N_14153,N_6728,N_9865);
or U14154 (N_14154,N_6879,N_5480);
or U14155 (N_14155,N_7630,N_7875);
and U14156 (N_14156,N_7602,N_5632);
and U14157 (N_14157,N_8051,N_7303);
or U14158 (N_14158,N_9683,N_9738);
or U14159 (N_14159,N_8702,N_8790);
and U14160 (N_14160,N_7665,N_5681);
or U14161 (N_14161,N_5016,N_5453);
nand U14162 (N_14162,N_9115,N_6669);
or U14163 (N_14163,N_6123,N_8258);
xnor U14164 (N_14164,N_5045,N_8227);
nand U14165 (N_14165,N_7986,N_6982);
or U14166 (N_14166,N_7755,N_8753);
nand U14167 (N_14167,N_7138,N_8137);
or U14168 (N_14168,N_9525,N_5281);
nor U14169 (N_14169,N_7199,N_5072);
nand U14170 (N_14170,N_7898,N_8969);
nand U14171 (N_14171,N_5295,N_7857);
nand U14172 (N_14172,N_5261,N_6293);
nor U14173 (N_14173,N_6738,N_9211);
nor U14174 (N_14174,N_5308,N_7831);
xnor U14175 (N_14175,N_5384,N_5561);
and U14176 (N_14176,N_9659,N_5368);
or U14177 (N_14177,N_6908,N_5774);
and U14178 (N_14178,N_6169,N_7793);
or U14179 (N_14179,N_7059,N_6246);
or U14180 (N_14180,N_8358,N_5578);
xor U14181 (N_14181,N_8439,N_6494);
nor U14182 (N_14182,N_9693,N_8073);
or U14183 (N_14183,N_9098,N_7293);
nor U14184 (N_14184,N_9116,N_6917);
nor U14185 (N_14185,N_8570,N_9950);
or U14186 (N_14186,N_5074,N_6938);
xnor U14187 (N_14187,N_9279,N_7626);
and U14188 (N_14188,N_5638,N_9661);
and U14189 (N_14189,N_5849,N_7423);
nand U14190 (N_14190,N_8987,N_6114);
and U14191 (N_14191,N_7578,N_8067);
nor U14192 (N_14192,N_6349,N_9175);
and U14193 (N_14193,N_9003,N_8440);
and U14194 (N_14194,N_6896,N_5560);
nor U14195 (N_14195,N_7236,N_7337);
nor U14196 (N_14196,N_6680,N_7386);
or U14197 (N_14197,N_8644,N_5443);
or U14198 (N_14198,N_6731,N_8797);
and U14199 (N_14199,N_8994,N_9919);
nand U14200 (N_14200,N_9153,N_8238);
or U14201 (N_14201,N_7428,N_9283);
or U14202 (N_14202,N_9417,N_8844);
or U14203 (N_14203,N_5447,N_8912);
nand U14204 (N_14204,N_7296,N_7119);
and U14205 (N_14205,N_6142,N_8221);
or U14206 (N_14206,N_8375,N_5873);
or U14207 (N_14207,N_8148,N_7466);
and U14208 (N_14208,N_9349,N_7641);
xor U14209 (N_14209,N_9028,N_7451);
and U14210 (N_14210,N_9803,N_5060);
or U14211 (N_14211,N_9811,N_8992);
nor U14212 (N_14212,N_8093,N_9533);
and U14213 (N_14213,N_9776,N_7331);
or U14214 (N_14214,N_8147,N_9576);
nand U14215 (N_14215,N_7087,N_9380);
or U14216 (N_14216,N_6495,N_7028);
and U14217 (N_14217,N_5292,N_5077);
and U14218 (N_14218,N_8828,N_7749);
nand U14219 (N_14219,N_5120,N_8717);
and U14220 (N_14220,N_9368,N_7589);
and U14221 (N_14221,N_5913,N_5340);
or U14222 (N_14222,N_8006,N_8829);
or U14223 (N_14223,N_9694,N_8789);
or U14224 (N_14224,N_5166,N_7013);
nor U14225 (N_14225,N_8303,N_5717);
nor U14226 (N_14226,N_7459,N_7537);
and U14227 (N_14227,N_5069,N_8941);
or U14228 (N_14228,N_7586,N_8859);
xnor U14229 (N_14229,N_6783,N_5251);
nand U14230 (N_14230,N_5469,N_9807);
and U14231 (N_14231,N_7426,N_5819);
or U14232 (N_14232,N_8972,N_9011);
and U14233 (N_14233,N_6154,N_9264);
or U14234 (N_14234,N_6143,N_8055);
nand U14235 (N_14235,N_5467,N_8421);
and U14236 (N_14236,N_9270,N_5330);
nand U14237 (N_14237,N_6268,N_6743);
nor U14238 (N_14238,N_5426,N_5391);
xnor U14239 (N_14239,N_6247,N_8207);
or U14240 (N_14240,N_6317,N_9533);
nor U14241 (N_14241,N_5273,N_6826);
nand U14242 (N_14242,N_6122,N_8399);
nor U14243 (N_14243,N_9626,N_6577);
nand U14244 (N_14244,N_7481,N_6286);
and U14245 (N_14245,N_5225,N_8312);
or U14246 (N_14246,N_6036,N_5289);
and U14247 (N_14247,N_7860,N_7033);
nand U14248 (N_14248,N_5695,N_6211);
and U14249 (N_14249,N_7487,N_5581);
nor U14250 (N_14250,N_8774,N_9978);
xnor U14251 (N_14251,N_5824,N_5454);
nand U14252 (N_14252,N_8052,N_9348);
xnor U14253 (N_14253,N_6683,N_9589);
or U14254 (N_14254,N_6922,N_8250);
nand U14255 (N_14255,N_5350,N_9233);
xnor U14256 (N_14256,N_8565,N_9933);
and U14257 (N_14257,N_7391,N_5092);
and U14258 (N_14258,N_8399,N_6547);
nor U14259 (N_14259,N_6116,N_5023);
xor U14260 (N_14260,N_7704,N_5959);
nor U14261 (N_14261,N_9581,N_6716);
nor U14262 (N_14262,N_9784,N_5820);
nor U14263 (N_14263,N_5158,N_7651);
nor U14264 (N_14264,N_9512,N_7380);
xnor U14265 (N_14265,N_5546,N_5638);
or U14266 (N_14266,N_8737,N_5384);
nand U14267 (N_14267,N_8855,N_8235);
nor U14268 (N_14268,N_8524,N_7423);
nand U14269 (N_14269,N_6441,N_8077);
or U14270 (N_14270,N_7882,N_8390);
nand U14271 (N_14271,N_7047,N_7179);
and U14272 (N_14272,N_8395,N_9625);
nand U14273 (N_14273,N_5506,N_5656);
nor U14274 (N_14274,N_6725,N_5876);
nor U14275 (N_14275,N_7945,N_6355);
or U14276 (N_14276,N_6293,N_8968);
and U14277 (N_14277,N_5424,N_7580);
or U14278 (N_14278,N_6012,N_6358);
and U14279 (N_14279,N_9497,N_5901);
nor U14280 (N_14280,N_6220,N_6928);
nand U14281 (N_14281,N_5477,N_8895);
and U14282 (N_14282,N_6944,N_8597);
and U14283 (N_14283,N_5789,N_7323);
nor U14284 (N_14284,N_6859,N_8139);
or U14285 (N_14285,N_6672,N_8848);
nor U14286 (N_14286,N_7064,N_8819);
nor U14287 (N_14287,N_6549,N_9631);
and U14288 (N_14288,N_5888,N_5569);
and U14289 (N_14289,N_8506,N_5298);
and U14290 (N_14290,N_5266,N_7360);
and U14291 (N_14291,N_7942,N_6553);
and U14292 (N_14292,N_8587,N_9512);
xor U14293 (N_14293,N_8243,N_9822);
nand U14294 (N_14294,N_7446,N_5358);
and U14295 (N_14295,N_9191,N_7231);
nor U14296 (N_14296,N_7946,N_7820);
nand U14297 (N_14297,N_8681,N_7004);
xor U14298 (N_14298,N_9143,N_8618);
or U14299 (N_14299,N_9729,N_7644);
xnor U14300 (N_14300,N_8752,N_8364);
nand U14301 (N_14301,N_7662,N_5555);
nor U14302 (N_14302,N_8998,N_6332);
xor U14303 (N_14303,N_7757,N_5739);
and U14304 (N_14304,N_6079,N_9426);
and U14305 (N_14305,N_7771,N_5604);
or U14306 (N_14306,N_5345,N_7327);
or U14307 (N_14307,N_9064,N_6756);
xor U14308 (N_14308,N_7558,N_9903);
or U14309 (N_14309,N_6758,N_5239);
nand U14310 (N_14310,N_5782,N_8720);
or U14311 (N_14311,N_8898,N_5436);
nand U14312 (N_14312,N_5003,N_5928);
and U14313 (N_14313,N_8454,N_8993);
nand U14314 (N_14314,N_8564,N_6206);
nand U14315 (N_14315,N_5848,N_6099);
nand U14316 (N_14316,N_5266,N_7833);
nand U14317 (N_14317,N_5538,N_6908);
nand U14318 (N_14318,N_9506,N_7976);
or U14319 (N_14319,N_6115,N_5617);
nand U14320 (N_14320,N_6525,N_7886);
or U14321 (N_14321,N_9173,N_7808);
nand U14322 (N_14322,N_5579,N_6408);
and U14323 (N_14323,N_9617,N_6263);
nand U14324 (N_14324,N_8417,N_8398);
and U14325 (N_14325,N_8760,N_9997);
or U14326 (N_14326,N_8994,N_9394);
or U14327 (N_14327,N_7849,N_7561);
nor U14328 (N_14328,N_7602,N_9342);
nand U14329 (N_14329,N_7324,N_6291);
xnor U14330 (N_14330,N_9937,N_5531);
and U14331 (N_14331,N_8741,N_8014);
xor U14332 (N_14332,N_6130,N_9144);
nor U14333 (N_14333,N_5742,N_9920);
nand U14334 (N_14334,N_8031,N_8279);
nand U14335 (N_14335,N_7486,N_6491);
or U14336 (N_14336,N_8001,N_7142);
nor U14337 (N_14337,N_7490,N_6295);
or U14338 (N_14338,N_7064,N_6251);
and U14339 (N_14339,N_9728,N_8606);
nor U14340 (N_14340,N_7690,N_7272);
and U14341 (N_14341,N_5080,N_8380);
xor U14342 (N_14342,N_7935,N_7024);
or U14343 (N_14343,N_5544,N_9841);
nand U14344 (N_14344,N_7343,N_6545);
nand U14345 (N_14345,N_6645,N_8286);
and U14346 (N_14346,N_7593,N_9193);
nor U14347 (N_14347,N_8536,N_7376);
xor U14348 (N_14348,N_7942,N_5746);
and U14349 (N_14349,N_7423,N_6268);
nand U14350 (N_14350,N_6512,N_9001);
nand U14351 (N_14351,N_6098,N_6528);
nor U14352 (N_14352,N_9343,N_8691);
and U14353 (N_14353,N_8239,N_6860);
xor U14354 (N_14354,N_8841,N_8570);
and U14355 (N_14355,N_6913,N_5703);
nor U14356 (N_14356,N_5314,N_5932);
and U14357 (N_14357,N_9566,N_9275);
xor U14358 (N_14358,N_7326,N_8574);
or U14359 (N_14359,N_5018,N_7051);
or U14360 (N_14360,N_7973,N_5802);
and U14361 (N_14361,N_5937,N_9632);
nor U14362 (N_14362,N_7943,N_7619);
nand U14363 (N_14363,N_9818,N_5230);
and U14364 (N_14364,N_8714,N_5553);
nand U14365 (N_14365,N_6617,N_9217);
and U14366 (N_14366,N_8021,N_5854);
and U14367 (N_14367,N_7821,N_9086);
or U14368 (N_14368,N_8191,N_6707);
or U14369 (N_14369,N_9976,N_8984);
or U14370 (N_14370,N_6592,N_5115);
nor U14371 (N_14371,N_9145,N_9216);
or U14372 (N_14372,N_5219,N_6540);
nor U14373 (N_14373,N_9134,N_5694);
xnor U14374 (N_14374,N_6771,N_7651);
or U14375 (N_14375,N_7485,N_9128);
xnor U14376 (N_14376,N_6689,N_5087);
nand U14377 (N_14377,N_5800,N_8853);
nor U14378 (N_14378,N_6949,N_5098);
nand U14379 (N_14379,N_5099,N_5277);
or U14380 (N_14380,N_7648,N_9836);
nor U14381 (N_14381,N_6655,N_5716);
nand U14382 (N_14382,N_7782,N_9690);
nand U14383 (N_14383,N_7982,N_6515);
and U14384 (N_14384,N_9901,N_8654);
xnor U14385 (N_14385,N_8018,N_5251);
nand U14386 (N_14386,N_8661,N_7827);
or U14387 (N_14387,N_5869,N_6699);
nand U14388 (N_14388,N_6283,N_7316);
nor U14389 (N_14389,N_6793,N_5294);
or U14390 (N_14390,N_9193,N_6101);
nand U14391 (N_14391,N_5994,N_7503);
or U14392 (N_14392,N_6668,N_7737);
and U14393 (N_14393,N_7695,N_6887);
nor U14394 (N_14394,N_9172,N_9485);
or U14395 (N_14395,N_5008,N_9328);
and U14396 (N_14396,N_9419,N_9293);
nand U14397 (N_14397,N_9354,N_9771);
nand U14398 (N_14398,N_7824,N_8408);
and U14399 (N_14399,N_9113,N_9905);
nor U14400 (N_14400,N_9328,N_6502);
and U14401 (N_14401,N_8670,N_5581);
and U14402 (N_14402,N_5871,N_8251);
or U14403 (N_14403,N_5015,N_7037);
and U14404 (N_14404,N_7082,N_9337);
nor U14405 (N_14405,N_7268,N_8648);
nor U14406 (N_14406,N_6524,N_7401);
nor U14407 (N_14407,N_8052,N_5075);
and U14408 (N_14408,N_6205,N_5734);
nand U14409 (N_14409,N_9484,N_6740);
or U14410 (N_14410,N_9845,N_8401);
or U14411 (N_14411,N_9056,N_9928);
nor U14412 (N_14412,N_6400,N_8292);
nor U14413 (N_14413,N_8240,N_9248);
or U14414 (N_14414,N_9359,N_5213);
and U14415 (N_14415,N_6715,N_9448);
or U14416 (N_14416,N_5573,N_8680);
nor U14417 (N_14417,N_9004,N_6246);
nor U14418 (N_14418,N_7281,N_6307);
nand U14419 (N_14419,N_6967,N_8973);
or U14420 (N_14420,N_9252,N_7850);
nand U14421 (N_14421,N_8118,N_9259);
or U14422 (N_14422,N_7263,N_8600);
or U14423 (N_14423,N_9413,N_8536);
and U14424 (N_14424,N_7439,N_6808);
nor U14425 (N_14425,N_8311,N_8668);
nand U14426 (N_14426,N_8017,N_8513);
nor U14427 (N_14427,N_9243,N_9336);
nand U14428 (N_14428,N_8118,N_5789);
nor U14429 (N_14429,N_6746,N_6237);
nand U14430 (N_14430,N_8626,N_6186);
and U14431 (N_14431,N_7296,N_6453);
xor U14432 (N_14432,N_5089,N_5755);
nor U14433 (N_14433,N_7619,N_7639);
nor U14434 (N_14434,N_5453,N_8311);
and U14435 (N_14435,N_9157,N_7287);
or U14436 (N_14436,N_8560,N_5519);
or U14437 (N_14437,N_9525,N_7040);
or U14438 (N_14438,N_9541,N_8830);
nand U14439 (N_14439,N_5864,N_9075);
or U14440 (N_14440,N_7736,N_7642);
nor U14441 (N_14441,N_6511,N_9412);
or U14442 (N_14442,N_9596,N_6465);
nand U14443 (N_14443,N_7218,N_7179);
nor U14444 (N_14444,N_8967,N_8707);
or U14445 (N_14445,N_5436,N_8778);
or U14446 (N_14446,N_6540,N_7255);
nor U14447 (N_14447,N_5272,N_9745);
xor U14448 (N_14448,N_8552,N_8029);
nand U14449 (N_14449,N_8172,N_5365);
and U14450 (N_14450,N_8431,N_8539);
and U14451 (N_14451,N_8376,N_6562);
and U14452 (N_14452,N_9649,N_8879);
nand U14453 (N_14453,N_5187,N_7463);
or U14454 (N_14454,N_8428,N_9822);
nand U14455 (N_14455,N_8230,N_6829);
and U14456 (N_14456,N_9822,N_8096);
or U14457 (N_14457,N_9722,N_7300);
nand U14458 (N_14458,N_7398,N_8971);
and U14459 (N_14459,N_9674,N_6042);
nor U14460 (N_14460,N_6142,N_9711);
and U14461 (N_14461,N_6839,N_6902);
and U14462 (N_14462,N_9690,N_5836);
nor U14463 (N_14463,N_7590,N_5792);
nand U14464 (N_14464,N_6743,N_6423);
nand U14465 (N_14465,N_6038,N_6538);
or U14466 (N_14466,N_6010,N_9932);
or U14467 (N_14467,N_6267,N_9683);
and U14468 (N_14468,N_7813,N_5623);
xnor U14469 (N_14469,N_9801,N_8976);
nand U14470 (N_14470,N_8284,N_6491);
nand U14471 (N_14471,N_8044,N_8212);
or U14472 (N_14472,N_7577,N_5017);
xor U14473 (N_14473,N_8060,N_5931);
nand U14474 (N_14474,N_5632,N_9421);
and U14475 (N_14475,N_8172,N_5363);
nand U14476 (N_14476,N_5192,N_8133);
nand U14477 (N_14477,N_7280,N_9814);
nand U14478 (N_14478,N_5349,N_9594);
nand U14479 (N_14479,N_8461,N_8138);
nor U14480 (N_14480,N_7930,N_5066);
or U14481 (N_14481,N_6942,N_6304);
nor U14482 (N_14482,N_8275,N_5446);
nand U14483 (N_14483,N_6421,N_7215);
or U14484 (N_14484,N_6260,N_7559);
or U14485 (N_14485,N_9146,N_9055);
or U14486 (N_14486,N_9298,N_7071);
or U14487 (N_14487,N_5375,N_5835);
nor U14488 (N_14488,N_5841,N_7529);
nand U14489 (N_14489,N_6303,N_9854);
nand U14490 (N_14490,N_7306,N_6101);
and U14491 (N_14491,N_5640,N_9958);
nor U14492 (N_14492,N_8194,N_5472);
nand U14493 (N_14493,N_6946,N_8343);
nand U14494 (N_14494,N_6140,N_5812);
and U14495 (N_14495,N_7374,N_9841);
xnor U14496 (N_14496,N_6071,N_8135);
nand U14497 (N_14497,N_9483,N_9428);
nand U14498 (N_14498,N_8108,N_9033);
or U14499 (N_14499,N_5186,N_6359);
or U14500 (N_14500,N_9423,N_5754);
and U14501 (N_14501,N_5647,N_8099);
and U14502 (N_14502,N_9328,N_6583);
nand U14503 (N_14503,N_9725,N_6755);
and U14504 (N_14504,N_8220,N_8085);
nor U14505 (N_14505,N_7209,N_9054);
xnor U14506 (N_14506,N_5178,N_8524);
or U14507 (N_14507,N_5503,N_7877);
nand U14508 (N_14508,N_6245,N_8612);
and U14509 (N_14509,N_6052,N_5473);
and U14510 (N_14510,N_6593,N_5587);
or U14511 (N_14511,N_6810,N_9785);
or U14512 (N_14512,N_7345,N_5635);
or U14513 (N_14513,N_6155,N_9675);
nand U14514 (N_14514,N_9821,N_8435);
and U14515 (N_14515,N_8712,N_6212);
and U14516 (N_14516,N_6990,N_8010);
nor U14517 (N_14517,N_7924,N_7312);
xor U14518 (N_14518,N_7488,N_9442);
or U14519 (N_14519,N_8491,N_9019);
nor U14520 (N_14520,N_7045,N_5881);
or U14521 (N_14521,N_7980,N_9840);
or U14522 (N_14522,N_6868,N_9077);
and U14523 (N_14523,N_9054,N_7990);
or U14524 (N_14524,N_6185,N_6336);
or U14525 (N_14525,N_6342,N_8515);
nor U14526 (N_14526,N_8171,N_7648);
and U14527 (N_14527,N_6970,N_8053);
or U14528 (N_14528,N_8957,N_6165);
xor U14529 (N_14529,N_5071,N_6448);
nor U14530 (N_14530,N_6509,N_7866);
and U14531 (N_14531,N_5188,N_6519);
or U14532 (N_14532,N_5955,N_6070);
or U14533 (N_14533,N_6591,N_8511);
nor U14534 (N_14534,N_6615,N_8034);
or U14535 (N_14535,N_9018,N_7763);
nor U14536 (N_14536,N_6913,N_9775);
nor U14537 (N_14537,N_8391,N_7006);
nand U14538 (N_14538,N_5224,N_9755);
and U14539 (N_14539,N_5932,N_8148);
and U14540 (N_14540,N_5605,N_8284);
nand U14541 (N_14541,N_7461,N_5650);
xnor U14542 (N_14542,N_6144,N_8186);
nand U14543 (N_14543,N_9084,N_5976);
or U14544 (N_14544,N_8033,N_7135);
nor U14545 (N_14545,N_5387,N_6844);
nand U14546 (N_14546,N_7885,N_7536);
nand U14547 (N_14547,N_8222,N_7747);
nor U14548 (N_14548,N_5531,N_7173);
nand U14549 (N_14549,N_9759,N_5490);
and U14550 (N_14550,N_7106,N_6539);
nor U14551 (N_14551,N_5084,N_7533);
and U14552 (N_14552,N_5493,N_5748);
xor U14553 (N_14553,N_7546,N_6636);
or U14554 (N_14554,N_5281,N_5591);
and U14555 (N_14555,N_8472,N_6368);
nor U14556 (N_14556,N_8771,N_7899);
nor U14557 (N_14557,N_6216,N_6124);
and U14558 (N_14558,N_8779,N_6398);
nand U14559 (N_14559,N_9228,N_6719);
nor U14560 (N_14560,N_6606,N_9860);
or U14561 (N_14561,N_5701,N_5243);
nand U14562 (N_14562,N_7293,N_8631);
or U14563 (N_14563,N_7388,N_6339);
and U14564 (N_14564,N_6029,N_8416);
and U14565 (N_14565,N_8166,N_6888);
and U14566 (N_14566,N_5029,N_5543);
and U14567 (N_14567,N_8136,N_6547);
nor U14568 (N_14568,N_5298,N_8146);
or U14569 (N_14569,N_6578,N_6548);
or U14570 (N_14570,N_9870,N_7788);
and U14571 (N_14571,N_9338,N_9744);
and U14572 (N_14572,N_6094,N_5486);
or U14573 (N_14573,N_7957,N_8335);
and U14574 (N_14574,N_7571,N_8931);
or U14575 (N_14575,N_7496,N_6037);
and U14576 (N_14576,N_8062,N_8125);
or U14577 (N_14577,N_7885,N_6963);
or U14578 (N_14578,N_7536,N_5590);
or U14579 (N_14579,N_5590,N_8940);
and U14580 (N_14580,N_8412,N_6159);
and U14581 (N_14581,N_7092,N_7016);
nand U14582 (N_14582,N_9795,N_9153);
nand U14583 (N_14583,N_9873,N_9724);
xor U14584 (N_14584,N_8454,N_7796);
and U14585 (N_14585,N_6362,N_5227);
and U14586 (N_14586,N_6020,N_7071);
xor U14587 (N_14587,N_5528,N_5836);
or U14588 (N_14588,N_6782,N_5851);
nand U14589 (N_14589,N_5322,N_6359);
xor U14590 (N_14590,N_7253,N_9543);
nor U14591 (N_14591,N_6298,N_6248);
or U14592 (N_14592,N_6433,N_7729);
nand U14593 (N_14593,N_6821,N_8345);
xnor U14594 (N_14594,N_8301,N_5752);
nor U14595 (N_14595,N_8906,N_9730);
nand U14596 (N_14596,N_5950,N_7913);
and U14597 (N_14597,N_7834,N_8883);
nor U14598 (N_14598,N_6956,N_8922);
nand U14599 (N_14599,N_5540,N_5278);
nor U14600 (N_14600,N_7124,N_5895);
nor U14601 (N_14601,N_7928,N_8314);
or U14602 (N_14602,N_7379,N_6760);
nor U14603 (N_14603,N_8039,N_8213);
and U14604 (N_14604,N_7756,N_6388);
or U14605 (N_14605,N_7545,N_6588);
nor U14606 (N_14606,N_5802,N_5541);
and U14607 (N_14607,N_6540,N_5378);
or U14608 (N_14608,N_7629,N_5395);
xor U14609 (N_14609,N_5444,N_6647);
or U14610 (N_14610,N_8077,N_9652);
and U14611 (N_14611,N_5269,N_5897);
or U14612 (N_14612,N_5207,N_5805);
and U14613 (N_14613,N_8849,N_5780);
and U14614 (N_14614,N_7601,N_6166);
nand U14615 (N_14615,N_8595,N_6347);
nor U14616 (N_14616,N_5663,N_9151);
or U14617 (N_14617,N_5280,N_7407);
nor U14618 (N_14618,N_9083,N_5237);
nand U14619 (N_14619,N_9214,N_5598);
nor U14620 (N_14620,N_6771,N_9621);
and U14621 (N_14621,N_5279,N_7239);
nand U14622 (N_14622,N_9694,N_5589);
nor U14623 (N_14623,N_5662,N_7705);
and U14624 (N_14624,N_6787,N_5549);
nor U14625 (N_14625,N_6740,N_8676);
nor U14626 (N_14626,N_6460,N_6573);
and U14627 (N_14627,N_7896,N_8857);
nand U14628 (N_14628,N_5981,N_8583);
and U14629 (N_14629,N_8217,N_6918);
or U14630 (N_14630,N_7767,N_9129);
nand U14631 (N_14631,N_8587,N_7909);
nor U14632 (N_14632,N_8601,N_5790);
or U14633 (N_14633,N_5877,N_8954);
nor U14634 (N_14634,N_6517,N_8475);
or U14635 (N_14635,N_9163,N_6958);
nand U14636 (N_14636,N_8658,N_6161);
or U14637 (N_14637,N_9612,N_7532);
or U14638 (N_14638,N_7498,N_6603);
or U14639 (N_14639,N_9603,N_9058);
xor U14640 (N_14640,N_9944,N_6159);
nor U14641 (N_14641,N_6943,N_8927);
nand U14642 (N_14642,N_5145,N_5591);
nor U14643 (N_14643,N_9813,N_5330);
nand U14644 (N_14644,N_9777,N_8341);
and U14645 (N_14645,N_7709,N_6721);
nand U14646 (N_14646,N_7525,N_6004);
and U14647 (N_14647,N_7503,N_5657);
nand U14648 (N_14648,N_8355,N_7410);
and U14649 (N_14649,N_8397,N_8595);
xor U14650 (N_14650,N_9577,N_9385);
nand U14651 (N_14651,N_7882,N_8361);
or U14652 (N_14652,N_6852,N_9884);
or U14653 (N_14653,N_5652,N_9885);
nor U14654 (N_14654,N_8119,N_8768);
xor U14655 (N_14655,N_9412,N_9231);
or U14656 (N_14656,N_6365,N_6637);
or U14657 (N_14657,N_5768,N_5953);
nor U14658 (N_14658,N_9914,N_7234);
or U14659 (N_14659,N_8999,N_6441);
or U14660 (N_14660,N_8235,N_7041);
nor U14661 (N_14661,N_7860,N_6195);
nand U14662 (N_14662,N_7480,N_7303);
xor U14663 (N_14663,N_7375,N_6023);
or U14664 (N_14664,N_8836,N_7345);
and U14665 (N_14665,N_8207,N_5230);
and U14666 (N_14666,N_6787,N_9040);
and U14667 (N_14667,N_6044,N_5128);
or U14668 (N_14668,N_8651,N_8608);
or U14669 (N_14669,N_5481,N_7723);
or U14670 (N_14670,N_8424,N_9072);
nor U14671 (N_14671,N_6996,N_8635);
nand U14672 (N_14672,N_5987,N_5183);
or U14673 (N_14673,N_7579,N_6653);
nand U14674 (N_14674,N_5151,N_8429);
nor U14675 (N_14675,N_5582,N_5392);
nand U14676 (N_14676,N_9266,N_8515);
xor U14677 (N_14677,N_5995,N_8071);
and U14678 (N_14678,N_6892,N_6689);
nand U14679 (N_14679,N_6538,N_6827);
nand U14680 (N_14680,N_5054,N_7147);
nor U14681 (N_14681,N_8910,N_8396);
nand U14682 (N_14682,N_7764,N_6656);
nor U14683 (N_14683,N_9542,N_6442);
nand U14684 (N_14684,N_6216,N_7229);
nor U14685 (N_14685,N_8943,N_7929);
xnor U14686 (N_14686,N_7878,N_5848);
nor U14687 (N_14687,N_9479,N_9291);
and U14688 (N_14688,N_7075,N_9523);
nor U14689 (N_14689,N_7027,N_7047);
or U14690 (N_14690,N_8816,N_5823);
and U14691 (N_14691,N_6510,N_8872);
nor U14692 (N_14692,N_6689,N_9615);
nor U14693 (N_14693,N_5010,N_5012);
nand U14694 (N_14694,N_8046,N_8964);
xnor U14695 (N_14695,N_9903,N_6730);
and U14696 (N_14696,N_7666,N_9007);
nand U14697 (N_14697,N_6110,N_8111);
nor U14698 (N_14698,N_9801,N_7860);
nor U14699 (N_14699,N_8309,N_6578);
nor U14700 (N_14700,N_8753,N_9667);
or U14701 (N_14701,N_9178,N_9044);
or U14702 (N_14702,N_5310,N_8900);
nand U14703 (N_14703,N_8862,N_9615);
or U14704 (N_14704,N_6154,N_7872);
and U14705 (N_14705,N_6993,N_9921);
nor U14706 (N_14706,N_7640,N_8265);
or U14707 (N_14707,N_6275,N_5405);
and U14708 (N_14708,N_8287,N_9132);
or U14709 (N_14709,N_6641,N_7369);
nor U14710 (N_14710,N_9213,N_5442);
nor U14711 (N_14711,N_6723,N_5064);
nor U14712 (N_14712,N_6951,N_9732);
xnor U14713 (N_14713,N_6700,N_9405);
or U14714 (N_14714,N_7575,N_9826);
nor U14715 (N_14715,N_8287,N_7469);
nand U14716 (N_14716,N_9311,N_9852);
nor U14717 (N_14717,N_9467,N_5539);
nand U14718 (N_14718,N_6241,N_6679);
xnor U14719 (N_14719,N_9367,N_7181);
nand U14720 (N_14720,N_5171,N_7076);
xor U14721 (N_14721,N_9796,N_5743);
nor U14722 (N_14722,N_5431,N_6411);
or U14723 (N_14723,N_8447,N_7262);
nand U14724 (N_14724,N_8306,N_6185);
nand U14725 (N_14725,N_5135,N_6466);
or U14726 (N_14726,N_6461,N_6579);
and U14727 (N_14727,N_8985,N_6923);
nand U14728 (N_14728,N_9691,N_8426);
and U14729 (N_14729,N_8416,N_9633);
or U14730 (N_14730,N_8808,N_9175);
xnor U14731 (N_14731,N_5593,N_6959);
nor U14732 (N_14732,N_6561,N_7044);
or U14733 (N_14733,N_9622,N_7921);
or U14734 (N_14734,N_8024,N_7210);
or U14735 (N_14735,N_7635,N_5018);
or U14736 (N_14736,N_5827,N_5992);
nor U14737 (N_14737,N_9342,N_8263);
or U14738 (N_14738,N_7416,N_9099);
nor U14739 (N_14739,N_8781,N_5252);
nand U14740 (N_14740,N_5140,N_5083);
nor U14741 (N_14741,N_7508,N_7078);
and U14742 (N_14742,N_9942,N_7626);
nor U14743 (N_14743,N_6281,N_9541);
or U14744 (N_14744,N_6368,N_6704);
nand U14745 (N_14745,N_6402,N_8640);
nand U14746 (N_14746,N_7410,N_8726);
nor U14747 (N_14747,N_8478,N_6329);
and U14748 (N_14748,N_7811,N_7631);
or U14749 (N_14749,N_8328,N_7374);
xnor U14750 (N_14750,N_5950,N_6193);
and U14751 (N_14751,N_6205,N_6991);
nand U14752 (N_14752,N_8662,N_6539);
nor U14753 (N_14753,N_9095,N_7187);
or U14754 (N_14754,N_7897,N_7570);
and U14755 (N_14755,N_5990,N_8420);
and U14756 (N_14756,N_5125,N_8040);
or U14757 (N_14757,N_5718,N_5644);
and U14758 (N_14758,N_6787,N_6501);
xor U14759 (N_14759,N_7809,N_7541);
nor U14760 (N_14760,N_7384,N_6758);
or U14761 (N_14761,N_7070,N_6392);
or U14762 (N_14762,N_8444,N_8057);
nand U14763 (N_14763,N_8749,N_8394);
or U14764 (N_14764,N_5296,N_9045);
or U14765 (N_14765,N_5749,N_7934);
nand U14766 (N_14766,N_8113,N_6458);
and U14767 (N_14767,N_7280,N_8783);
nor U14768 (N_14768,N_7946,N_7281);
nand U14769 (N_14769,N_8649,N_7803);
nor U14770 (N_14770,N_5050,N_8794);
and U14771 (N_14771,N_8809,N_5702);
and U14772 (N_14772,N_8608,N_7803);
or U14773 (N_14773,N_9475,N_9372);
or U14774 (N_14774,N_6895,N_5821);
nand U14775 (N_14775,N_5707,N_8103);
nand U14776 (N_14776,N_5325,N_6509);
nand U14777 (N_14777,N_6016,N_5829);
or U14778 (N_14778,N_5978,N_9300);
nor U14779 (N_14779,N_6927,N_7807);
nand U14780 (N_14780,N_7523,N_7020);
or U14781 (N_14781,N_8006,N_5377);
xnor U14782 (N_14782,N_5665,N_8918);
nor U14783 (N_14783,N_7821,N_6440);
xnor U14784 (N_14784,N_6487,N_9055);
nor U14785 (N_14785,N_8911,N_7902);
nor U14786 (N_14786,N_9342,N_5638);
nand U14787 (N_14787,N_6387,N_8099);
and U14788 (N_14788,N_6131,N_7385);
and U14789 (N_14789,N_9865,N_6060);
and U14790 (N_14790,N_5032,N_6434);
nand U14791 (N_14791,N_9682,N_7446);
or U14792 (N_14792,N_8849,N_7891);
or U14793 (N_14793,N_5515,N_8960);
nand U14794 (N_14794,N_7145,N_6660);
or U14795 (N_14795,N_6577,N_8546);
and U14796 (N_14796,N_6572,N_8433);
xnor U14797 (N_14797,N_7288,N_8421);
and U14798 (N_14798,N_8347,N_6478);
and U14799 (N_14799,N_5902,N_6641);
and U14800 (N_14800,N_6547,N_7198);
nor U14801 (N_14801,N_8441,N_5287);
xor U14802 (N_14802,N_5630,N_8686);
nor U14803 (N_14803,N_5842,N_8768);
nor U14804 (N_14804,N_8238,N_7786);
nand U14805 (N_14805,N_7198,N_9211);
and U14806 (N_14806,N_5946,N_8455);
nand U14807 (N_14807,N_8076,N_9582);
xor U14808 (N_14808,N_5434,N_9680);
nand U14809 (N_14809,N_8407,N_5266);
or U14810 (N_14810,N_7953,N_5854);
nand U14811 (N_14811,N_5932,N_7258);
or U14812 (N_14812,N_6158,N_7905);
nor U14813 (N_14813,N_5387,N_8769);
and U14814 (N_14814,N_5497,N_5690);
nor U14815 (N_14815,N_9835,N_8789);
and U14816 (N_14816,N_8096,N_9891);
nor U14817 (N_14817,N_6996,N_6586);
nor U14818 (N_14818,N_5947,N_7153);
or U14819 (N_14819,N_9366,N_8110);
nand U14820 (N_14820,N_9059,N_5774);
nand U14821 (N_14821,N_5957,N_6127);
nor U14822 (N_14822,N_5634,N_6282);
or U14823 (N_14823,N_7963,N_8912);
and U14824 (N_14824,N_7855,N_9772);
nor U14825 (N_14825,N_5709,N_8221);
and U14826 (N_14826,N_7926,N_9279);
nor U14827 (N_14827,N_9636,N_5506);
nand U14828 (N_14828,N_6226,N_7540);
nor U14829 (N_14829,N_6363,N_7806);
or U14830 (N_14830,N_9971,N_8479);
xor U14831 (N_14831,N_7224,N_8226);
nand U14832 (N_14832,N_8786,N_6109);
and U14833 (N_14833,N_8210,N_9173);
xor U14834 (N_14834,N_9870,N_8956);
or U14835 (N_14835,N_7237,N_8937);
or U14836 (N_14836,N_6485,N_5088);
or U14837 (N_14837,N_6178,N_7682);
nand U14838 (N_14838,N_9691,N_5536);
nor U14839 (N_14839,N_7430,N_8155);
or U14840 (N_14840,N_6114,N_8505);
nor U14841 (N_14841,N_8930,N_7516);
and U14842 (N_14842,N_7109,N_9540);
nor U14843 (N_14843,N_5470,N_7917);
xnor U14844 (N_14844,N_7511,N_9462);
and U14845 (N_14845,N_9877,N_7909);
nor U14846 (N_14846,N_8033,N_7887);
xnor U14847 (N_14847,N_8003,N_5467);
and U14848 (N_14848,N_8248,N_9010);
nor U14849 (N_14849,N_6622,N_7302);
and U14850 (N_14850,N_7982,N_5368);
or U14851 (N_14851,N_8300,N_9594);
nor U14852 (N_14852,N_6856,N_7622);
nor U14853 (N_14853,N_7292,N_7975);
or U14854 (N_14854,N_8294,N_5510);
nor U14855 (N_14855,N_9399,N_5344);
nand U14856 (N_14856,N_7467,N_7543);
nor U14857 (N_14857,N_9792,N_9886);
and U14858 (N_14858,N_5797,N_9318);
and U14859 (N_14859,N_9859,N_8101);
nand U14860 (N_14860,N_9763,N_5154);
and U14861 (N_14861,N_8848,N_7382);
nand U14862 (N_14862,N_5175,N_6426);
nor U14863 (N_14863,N_9344,N_9134);
nand U14864 (N_14864,N_7274,N_5618);
nor U14865 (N_14865,N_8163,N_8660);
or U14866 (N_14866,N_8777,N_7616);
and U14867 (N_14867,N_8984,N_5768);
nor U14868 (N_14868,N_9735,N_5473);
and U14869 (N_14869,N_7348,N_8397);
nand U14870 (N_14870,N_6388,N_9476);
nand U14871 (N_14871,N_9609,N_8590);
and U14872 (N_14872,N_6938,N_5421);
nor U14873 (N_14873,N_7167,N_8706);
nor U14874 (N_14874,N_7967,N_8501);
or U14875 (N_14875,N_8402,N_6504);
nor U14876 (N_14876,N_7160,N_8648);
or U14877 (N_14877,N_8937,N_7615);
or U14878 (N_14878,N_5489,N_8705);
nand U14879 (N_14879,N_9389,N_9014);
or U14880 (N_14880,N_6442,N_9090);
and U14881 (N_14881,N_7098,N_9647);
nor U14882 (N_14882,N_5862,N_9320);
or U14883 (N_14883,N_6694,N_5413);
and U14884 (N_14884,N_7891,N_9649);
or U14885 (N_14885,N_7391,N_8908);
nand U14886 (N_14886,N_9260,N_9389);
and U14887 (N_14887,N_7911,N_6640);
nand U14888 (N_14888,N_8001,N_7398);
and U14889 (N_14889,N_5088,N_9162);
nand U14890 (N_14890,N_8982,N_9139);
and U14891 (N_14891,N_6186,N_8676);
nand U14892 (N_14892,N_7536,N_9861);
and U14893 (N_14893,N_7431,N_8397);
or U14894 (N_14894,N_9829,N_7089);
and U14895 (N_14895,N_5408,N_9770);
or U14896 (N_14896,N_7698,N_6164);
and U14897 (N_14897,N_8476,N_9555);
or U14898 (N_14898,N_9350,N_9981);
nand U14899 (N_14899,N_6052,N_8553);
and U14900 (N_14900,N_9564,N_5706);
nor U14901 (N_14901,N_5589,N_9097);
xnor U14902 (N_14902,N_5194,N_7804);
or U14903 (N_14903,N_7567,N_5536);
xor U14904 (N_14904,N_5529,N_7915);
nor U14905 (N_14905,N_8470,N_7135);
or U14906 (N_14906,N_6872,N_5161);
or U14907 (N_14907,N_6907,N_7331);
xor U14908 (N_14908,N_9119,N_5832);
nor U14909 (N_14909,N_9014,N_5644);
nor U14910 (N_14910,N_9871,N_9049);
and U14911 (N_14911,N_6452,N_7972);
xnor U14912 (N_14912,N_9519,N_7382);
nor U14913 (N_14913,N_8219,N_8576);
and U14914 (N_14914,N_9830,N_9956);
nand U14915 (N_14915,N_9304,N_8608);
and U14916 (N_14916,N_8890,N_8623);
nor U14917 (N_14917,N_5925,N_6253);
and U14918 (N_14918,N_5145,N_8430);
nor U14919 (N_14919,N_8255,N_9465);
or U14920 (N_14920,N_6753,N_9815);
nand U14921 (N_14921,N_5898,N_8320);
nor U14922 (N_14922,N_7524,N_8152);
and U14923 (N_14923,N_6447,N_8590);
nor U14924 (N_14924,N_5780,N_7546);
nor U14925 (N_14925,N_8708,N_9702);
or U14926 (N_14926,N_5753,N_7785);
nand U14927 (N_14927,N_7716,N_8689);
nand U14928 (N_14928,N_5350,N_8747);
and U14929 (N_14929,N_9476,N_7241);
nor U14930 (N_14930,N_9476,N_7749);
nand U14931 (N_14931,N_5915,N_8997);
nand U14932 (N_14932,N_9740,N_9132);
nand U14933 (N_14933,N_8448,N_8980);
or U14934 (N_14934,N_8806,N_9779);
or U14935 (N_14935,N_7675,N_8631);
and U14936 (N_14936,N_8149,N_6766);
and U14937 (N_14937,N_7423,N_7133);
nor U14938 (N_14938,N_9855,N_6620);
and U14939 (N_14939,N_7370,N_5561);
nand U14940 (N_14940,N_6640,N_6281);
nand U14941 (N_14941,N_7946,N_6271);
nand U14942 (N_14942,N_6280,N_9732);
and U14943 (N_14943,N_5272,N_9225);
xor U14944 (N_14944,N_6557,N_9882);
nand U14945 (N_14945,N_8783,N_5464);
xor U14946 (N_14946,N_5401,N_9974);
or U14947 (N_14947,N_5312,N_9408);
xnor U14948 (N_14948,N_5477,N_5953);
xnor U14949 (N_14949,N_7647,N_5147);
and U14950 (N_14950,N_9680,N_6906);
or U14951 (N_14951,N_5846,N_9466);
or U14952 (N_14952,N_9376,N_7795);
nand U14953 (N_14953,N_6443,N_7160);
or U14954 (N_14954,N_8144,N_8863);
or U14955 (N_14955,N_6817,N_9089);
or U14956 (N_14956,N_5261,N_6720);
xnor U14957 (N_14957,N_7434,N_5589);
xor U14958 (N_14958,N_5010,N_9943);
nor U14959 (N_14959,N_5329,N_9828);
nand U14960 (N_14960,N_5327,N_6449);
or U14961 (N_14961,N_7714,N_8351);
nand U14962 (N_14962,N_7109,N_8323);
or U14963 (N_14963,N_8692,N_6345);
or U14964 (N_14964,N_9659,N_5569);
nand U14965 (N_14965,N_8684,N_5666);
or U14966 (N_14966,N_8105,N_9979);
nor U14967 (N_14967,N_6919,N_8141);
or U14968 (N_14968,N_7339,N_5813);
nand U14969 (N_14969,N_9219,N_6391);
nor U14970 (N_14970,N_5120,N_7213);
and U14971 (N_14971,N_9394,N_6118);
or U14972 (N_14972,N_5104,N_9040);
or U14973 (N_14973,N_5071,N_8020);
nand U14974 (N_14974,N_8273,N_9373);
nor U14975 (N_14975,N_9043,N_7760);
and U14976 (N_14976,N_7079,N_8200);
and U14977 (N_14977,N_7345,N_7166);
xnor U14978 (N_14978,N_8602,N_5826);
or U14979 (N_14979,N_5017,N_8953);
and U14980 (N_14980,N_7056,N_7785);
and U14981 (N_14981,N_8397,N_5302);
nand U14982 (N_14982,N_6537,N_8025);
or U14983 (N_14983,N_9122,N_7654);
nor U14984 (N_14984,N_5327,N_5358);
nor U14985 (N_14985,N_8091,N_6093);
or U14986 (N_14986,N_8785,N_8535);
and U14987 (N_14987,N_8428,N_8998);
and U14988 (N_14988,N_6445,N_7516);
nand U14989 (N_14989,N_9853,N_8371);
and U14990 (N_14990,N_6758,N_8887);
xnor U14991 (N_14991,N_7470,N_6434);
and U14992 (N_14992,N_5844,N_6553);
nor U14993 (N_14993,N_8040,N_9901);
nand U14994 (N_14994,N_5674,N_9493);
nand U14995 (N_14995,N_7558,N_6223);
or U14996 (N_14996,N_5288,N_8036);
and U14997 (N_14997,N_9509,N_6817);
nor U14998 (N_14998,N_5999,N_7946);
and U14999 (N_14999,N_5418,N_8840);
and U15000 (N_15000,N_14514,N_12248);
and U15001 (N_15001,N_11885,N_10036);
nand U15002 (N_15002,N_10852,N_12849);
or U15003 (N_15003,N_11968,N_13915);
nand U15004 (N_15004,N_11772,N_11823);
and U15005 (N_15005,N_14670,N_13632);
and U15006 (N_15006,N_11285,N_14205);
or U15007 (N_15007,N_13939,N_10921);
and U15008 (N_15008,N_12208,N_14575);
and U15009 (N_15009,N_11641,N_11690);
nand U15010 (N_15010,N_14481,N_13207);
nor U15011 (N_15011,N_13869,N_12409);
nand U15012 (N_15012,N_12413,N_14053);
or U15013 (N_15013,N_14144,N_10992);
or U15014 (N_15014,N_10671,N_13304);
nor U15015 (N_15015,N_12156,N_13950);
nand U15016 (N_15016,N_14200,N_11134);
and U15017 (N_15017,N_14213,N_14199);
nand U15018 (N_15018,N_11190,N_10670);
xnor U15019 (N_15019,N_11278,N_13903);
and U15020 (N_15020,N_13369,N_11943);
or U15021 (N_15021,N_10327,N_14339);
and U15022 (N_15022,N_13417,N_10660);
or U15023 (N_15023,N_13587,N_13162);
nand U15024 (N_15024,N_10209,N_11999);
or U15025 (N_15025,N_14028,N_10908);
and U15026 (N_15026,N_11554,N_13171);
or U15027 (N_15027,N_14762,N_10974);
xnor U15028 (N_15028,N_11372,N_14369);
nand U15029 (N_15029,N_13696,N_10196);
or U15030 (N_15030,N_13172,N_13484);
and U15031 (N_15031,N_10693,N_11655);
or U15032 (N_15032,N_11274,N_10580);
nor U15033 (N_15033,N_11514,N_10749);
nor U15034 (N_15034,N_12900,N_11167);
and U15035 (N_15035,N_14054,N_11357);
or U15036 (N_15036,N_13197,N_14447);
nand U15037 (N_15037,N_11337,N_13280);
nor U15038 (N_15038,N_10681,N_13255);
and U15039 (N_15039,N_10453,N_13866);
nand U15040 (N_15040,N_11464,N_11188);
xor U15041 (N_15041,N_14741,N_11938);
nand U15042 (N_15042,N_11391,N_13060);
nor U15043 (N_15043,N_12512,N_14103);
or U15044 (N_15044,N_11273,N_10924);
nand U15045 (N_15045,N_14478,N_12971);
or U15046 (N_15046,N_11863,N_11333);
xor U15047 (N_15047,N_13493,N_12055);
and U15048 (N_15048,N_10228,N_11246);
and U15049 (N_15049,N_14527,N_14999);
nand U15050 (N_15050,N_12330,N_10236);
nand U15051 (N_15051,N_12419,N_10210);
nand U15052 (N_15052,N_13238,N_11922);
nor U15053 (N_15053,N_12963,N_14065);
nor U15054 (N_15054,N_12108,N_14778);
nor U15055 (N_15055,N_12764,N_13966);
nor U15056 (N_15056,N_12891,N_12803);
xnor U15057 (N_15057,N_11792,N_13298);
xnor U15058 (N_15058,N_10790,N_11280);
and U15059 (N_15059,N_12111,N_10116);
nor U15060 (N_15060,N_14457,N_14171);
xnor U15061 (N_15061,N_11515,N_11084);
nor U15062 (N_15062,N_10844,N_14212);
nor U15063 (N_15063,N_10122,N_11635);
and U15064 (N_15064,N_13997,N_12050);
xor U15065 (N_15065,N_12756,N_11776);
nand U15066 (N_15066,N_12358,N_10829);
and U15067 (N_15067,N_11581,N_14105);
and U15068 (N_15068,N_10610,N_10097);
and U15069 (N_15069,N_12661,N_11680);
or U15070 (N_15070,N_10557,N_10630);
nand U15071 (N_15071,N_14554,N_14497);
nand U15072 (N_15072,N_13846,N_10001);
nor U15073 (N_15073,N_14376,N_10450);
nand U15074 (N_15074,N_10898,N_10213);
or U15075 (N_15075,N_12465,N_12493);
xnor U15076 (N_15076,N_12716,N_13196);
xnor U15077 (N_15077,N_11123,N_10917);
nand U15078 (N_15078,N_10423,N_10558);
or U15079 (N_15079,N_10896,N_10202);
or U15080 (N_15080,N_11489,N_12653);
and U15081 (N_15081,N_11936,N_12066);
and U15082 (N_15082,N_13557,N_12595);
nand U15083 (N_15083,N_12198,N_14990);
nand U15084 (N_15084,N_11490,N_12503);
nand U15085 (N_15085,N_14201,N_11013);
nor U15086 (N_15086,N_13621,N_10753);
nor U15087 (N_15087,N_11047,N_13202);
or U15088 (N_15088,N_13935,N_10306);
or U15089 (N_15089,N_10381,N_13439);
or U15090 (N_15090,N_14752,N_14529);
xnor U15091 (N_15091,N_11616,N_14240);
and U15092 (N_15092,N_14971,N_14320);
or U15093 (N_15093,N_11562,N_10851);
nand U15094 (N_15094,N_11801,N_14725);
or U15095 (N_15095,N_11934,N_14433);
and U15096 (N_15096,N_14651,N_13898);
or U15097 (N_15097,N_11098,N_11072);
or U15098 (N_15098,N_12471,N_14794);
and U15099 (N_15099,N_11779,N_11051);
and U15100 (N_15100,N_13148,N_14408);
and U15101 (N_15101,N_10570,N_10076);
and U15102 (N_15102,N_13037,N_13778);
nor U15103 (N_15103,N_10940,N_12860);
nor U15104 (N_15104,N_11668,N_11611);
nand U15105 (N_15105,N_14468,N_14800);
nor U15106 (N_15106,N_11862,N_10165);
or U15107 (N_15107,N_12240,N_11346);
and U15108 (N_15108,N_14170,N_14585);
nand U15109 (N_15109,N_10168,N_11797);
nor U15110 (N_15110,N_14414,N_14252);
nand U15111 (N_15111,N_11079,N_11433);
nor U15112 (N_15112,N_10397,N_14060);
xor U15113 (N_15113,N_13629,N_14063);
or U15114 (N_15114,N_13018,N_13340);
nand U15115 (N_15115,N_12277,N_11971);
nand U15116 (N_15116,N_13194,N_11647);
nand U15117 (N_15117,N_12695,N_10263);
nand U15118 (N_15118,N_11403,N_14963);
or U15119 (N_15119,N_13055,N_14475);
or U15120 (N_15120,N_12366,N_13353);
nand U15121 (N_15121,N_12201,N_11381);
and U15122 (N_15122,N_12027,N_11845);
nand U15123 (N_15123,N_14328,N_11688);
nand U15124 (N_15124,N_10111,N_10089);
nor U15125 (N_15125,N_13333,N_13682);
nand U15126 (N_15126,N_14976,N_12463);
xor U15127 (N_15127,N_12270,N_10041);
and U15128 (N_15128,N_10167,N_14410);
nand U15129 (N_15129,N_13857,N_12416);
and U15130 (N_15130,N_10411,N_12016);
nand U15131 (N_15131,N_12319,N_10909);
xor U15132 (N_15132,N_11130,N_12254);
and U15133 (N_15133,N_12206,N_14982);
and U15134 (N_15134,N_10481,N_10109);
nand U15135 (N_15135,N_13844,N_12130);
nand U15136 (N_15136,N_10374,N_14656);
nor U15137 (N_15137,N_12567,N_10846);
xor U15138 (N_15138,N_11535,N_14018);
nor U15139 (N_15139,N_14790,N_13941);
and U15140 (N_15140,N_14248,N_10810);
and U15141 (N_15141,N_11578,N_13120);
or U15142 (N_15142,N_12781,N_13303);
and U15143 (N_15143,N_10741,N_11457);
and U15144 (N_15144,N_14541,N_14579);
nor U15145 (N_15145,N_12536,N_11220);
or U15146 (N_15146,N_12539,N_13378);
nand U15147 (N_15147,N_10348,N_14469);
or U15148 (N_15148,N_14394,N_10633);
nor U15149 (N_15149,N_13902,N_13998);
nand U15150 (N_15150,N_13085,N_10271);
and U15151 (N_15151,N_10792,N_12407);
and U15152 (N_15152,N_14735,N_11694);
nor U15153 (N_15153,N_13169,N_14487);
and U15154 (N_15154,N_10527,N_10399);
nand U15155 (N_15155,N_11543,N_12826);
or U15156 (N_15156,N_11427,N_10025);
nor U15157 (N_15157,N_11209,N_10010);
or U15158 (N_15158,N_12836,N_14088);
or U15159 (N_15159,N_13039,N_11675);
or U15160 (N_15160,N_14476,N_13927);
or U15161 (N_15161,N_12871,N_11705);
nor U15162 (N_15162,N_14340,N_12968);
nand U15163 (N_15163,N_14090,N_11994);
nor U15164 (N_15164,N_12680,N_13005);
or U15165 (N_15165,N_14025,N_11353);
xnor U15166 (N_15166,N_12025,N_14837);
nand U15167 (N_15167,N_11193,N_10245);
or U15168 (N_15168,N_14445,N_14594);
nand U15169 (N_15169,N_14503,N_13600);
nand U15170 (N_15170,N_13296,N_14626);
and U15171 (N_15171,N_13167,N_11347);
xor U15172 (N_15172,N_11957,N_12932);
xnor U15173 (N_15173,N_13042,N_13359);
nor U15174 (N_15174,N_10538,N_13468);
nor U15175 (N_15175,N_12357,N_10776);
or U15176 (N_15176,N_13134,N_10095);
or U15177 (N_15177,N_14887,N_10482);
or U15178 (N_15178,N_13404,N_14935);
nor U15179 (N_15179,N_10417,N_10048);
nand U15180 (N_15180,N_12802,N_13667);
or U15181 (N_15181,N_13074,N_11715);
and U15182 (N_15182,N_12384,N_10012);
nand U15183 (N_15183,N_10569,N_11410);
or U15184 (N_15184,N_13920,N_13499);
and U15185 (N_15185,N_14006,N_14907);
and U15186 (N_15186,N_10891,N_13412);
and U15187 (N_15187,N_12796,N_10096);
or U15188 (N_15188,N_11361,N_13859);
xnor U15189 (N_15189,N_13899,N_12641);
nor U15190 (N_15190,N_13544,N_13354);
xor U15191 (N_15191,N_13115,N_14304);
nor U15192 (N_15192,N_12943,N_11571);
nand U15193 (N_15193,N_10211,N_12132);
nand U15194 (N_15194,N_11196,N_12866);
or U15195 (N_15195,N_13348,N_10872);
nand U15196 (N_15196,N_10566,N_13580);
or U15197 (N_15197,N_10276,N_12747);
or U15198 (N_15198,N_11055,N_10022);
or U15199 (N_15199,N_12477,N_13441);
and U15200 (N_15200,N_12275,N_10414);
xnor U15201 (N_15201,N_13572,N_11902);
and U15202 (N_15202,N_10328,N_12334);
and U15203 (N_15203,N_14493,N_11370);
and U15204 (N_15204,N_13146,N_11748);
and U15205 (N_15205,N_12785,N_11599);
or U15206 (N_15206,N_14138,N_13765);
xnor U15207 (N_15207,N_10249,N_10581);
nand U15208 (N_15208,N_10579,N_10666);
and U15209 (N_15209,N_14909,N_10442);
nor U15210 (N_15210,N_13474,N_11603);
nor U15211 (N_15211,N_11766,N_13086);
nand U15212 (N_15212,N_13307,N_12501);
nand U15213 (N_15213,N_14062,N_14225);
nand U15214 (N_15214,N_13555,N_13111);
nand U15215 (N_15215,N_10027,N_14513);
nor U15216 (N_15216,N_11470,N_10060);
nor U15217 (N_15217,N_12829,N_14356);
nor U15218 (N_15218,N_10156,N_12320);
nand U15219 (N_15219,N_14986,N_14327);
and U15220 (N_15220,N_11582,N_12189);
nor U15221 (N_15221,N_11369,N_10128);
or U15222 (N_15222,N_11476,N_13106);
and U15223 (N_15223,N_13612,N_13357);
nand U15224 (N_15224,N_13605,N_10293);
or U15225 (N_15225,N_12474,N_12917);
nor U15226 (N_15226,N_12281,N_14037);
nand U15227 (N_15227,N_10448,N_10408);
nand U15228 (N_15228,N_13906,N_11408);
and U15229 (N_15229,N_12942,N_14864);
xor U15230 (N_15230,N_12196,N_13829);
nor U15231 (N_15231,N_14072,N_12739);
nand U15232 (N_15232,N_12318,N_10542);
nor U15233 (N_15233,N_11959,N_11261);
nor U15234 (N_15234,N_10874,N_12522);
xor U15235 (N_15235,N_14903,N_12611);
and U15236 (N_15236,N_10084,N_10410);
or U15237 (N_15237,N_14720,N_12141);
nand U15238 (N_15238,N_13618,N_10008);
nor U15239 (N_15239,N_12734,N_11431);
nor U15240 (N_15240,N_14217,N_14869);
nand U15241 (N_15241,N_12393,N_11471);
or U15242 (N_15242,N_10967,N_12858);
or U15243 (N_15243,N_11711,N_10473);
nand U15244 (N_15244,N_11122,N_10231);
or U15245 (N_15245,N_14486,N_14166);
xnor U15246 (N_15246,N_11678,N_11396);
nor U15247 (N_15247,N_13320,N_10155);
nand U15248 (N_15248,N_14434,N_14092);
and U15249 (N_15249,N_14271,N_13636);
nor U15250 (N_15250,N_12806,N_12590);
xor U15251 (N_15251,N_13806,N_13050);
nand U15252 (N_15252,N_12102,N_10398);
and U15253 (N_15253,N_13285,N_14419);
nand U15254 (N_15254,N_10888,N_11850);
nand U15255 (N_15255,N_14727,N_11762);
nand U15256 (N_15256,N_14137,N_12957);
xnor U15257 (N_15257,N_14624,N_10117);
and U15258 (N_15258,N_11412,N_13405);
xnor U15259 (N_15259,N_14866,N_14956);
xor U15260 (N_15260,N_10309,N_10487);
or U15261 (N_15261,N_11281,N_14331);
nand U15262 (N_15262,N_10977,N_10970);
nand U15263 (N_15263,N_10189,N_10120);
or U15264 (N_15264,N_11997,N_13372);
xnor U15265 (N_15265,N_14159,N_10859);
nor U15266 (N_15266,N_12675,N_12014);
or U15267 (N_15267,N_12054,N_12674);
nand U15268 (N_15268,N_13529,N_10978);
and U15269 (N_15269,N_13960,N_11243);
xor U15270 (N_15270,N_13279,N_13327);
nor U15271 (N_15271,N_11624,N_12912);
and U15272 (N_15272,N_14763,N_10345);
nand U15273 (N_15273,N_13000,N_14824);
nand U15274 (N_15274,N_10229,N_14845);
nand U15275 (N_15275,N_13690,N_11244);
nor U15276 (N_15276,N_11860,N_13657);
nor U15277 (N_15277,N_11006,N_13509);
nand U15278 (N_15278,N_14383,N_14015);
or U15279 (N_15279,N_14709,N_11303);
nor U15280 (N_15280,N_11509,N_14604);
nand U15281 (N_15281,N_14902,N_10640);
or U15282 (N_15282,N_11080,N_10301);
xnor U15283 (N_15283,N_11727,N_10627);
nand U15284 (N_15284,N_14411,N_12798);
and U15285 (N_15285,N_11426,N_14988);
nand U15286 (N_15286,N_10082,N_10354);
or U15287 (N_15287,N_11067,N_13267);
and U15288 (N_15288,N_13428,N_11587);
nor U15289 (N_15289,N_12547,N_14728);
nand U15290 (N_15290,N_14224,N_12682);
nand U15291 (N_15291,N_10952,N_10499);
nand U15292 (N_15292,N_11712,N_12482);
xnor U15293 (N_15293,N_12228,N_14926);
and U15294 (N_15294,N_11029,N_11377);
or U15295 (N_15295,N_12535,N_13635);
or U15296 (N_15296,N_13754,N_13052);
nor U15297 (N_15297,N_13319,N_11481);
or U15298 (N_15298,N_10368,N_14592);
and U15299 (N_15299,N_14884,N_12977);
or U15300 (N_15300,N_11034,N_10913);
nand U15301 (N_15301,N_12091,N_13214);
nand U15302 (N_15302,N_14609,N_13536);
and U15303 (N_15303,N_14773,N_10830);
xor U15304 (N_15304,N_12690,N_12789);
or U15305 (N_15305,N_13234,N_14676);
and U15306 (N_15306,N_12730,N_13877);
and U15307 (N_15307,N_14648,N_13245);
nor U15308 (N_15308,N_10842,N_14507);
and U15309 (N_15309,N_12788,N_10591);
and U15310 (N_15310,N_11239,N_10033);
and U15311 (N_15311,N_14441,N_14220);
and U15312 (N_15312,N_14819,N_13366);
xor U15313 (N_15313,N_11781,N_13810);
xnor U15314 (N_15314,N_13827,N_13145);
nor U15315 (N_15315,N_12061,N_13104);
nor U15316 (N_15316,N_12577,N_10609);
nor U15317 (N_15317,N_13435,N_14666);
or U15318 (N_15318,N_11349,N_14966);
nor U15319 (N_15319,N_12585,N_13720);
and U15320 (N_15320,N_12727,N_11141);
nor U15321 (N_15321,N_13471,N_10441);
nor U15322 (N_15322,N_10312,N_10244);
xor U15323 (N_15323,N_14086,N_12233);
nand U15324 (N_15324,N_13805,N_10308);
nand U15325 (N_15325,N_13565,N_13561);
or U15326 (N_15326,N_11782,N_13530);
nor U15327 (N_15327,N_11825,N_11657);
xnor U15328 (N_15328,N_10392,N_10677);
or U15329 (N_15329,N_11699,N_14696);
nor U15330 (N_15330,N_14237,N_14284);
nor U15331 (N_15331,N_10936,N_12616);
nand U15332 (N_15332,N_11093,N_14858);
or U15333 (N_15333,N_12558,N_13158);
xor U15334 (N_15334,N_14934,N_14499);
and U15335 (N_15335,N_14713,N_12708);
nor U15336 (N_15336,N_13413,N_11101);
nand U15337 (N_15337,N_11511,N_13001);
or U15338 (N_15338,N_13522,N_11944);
or U15339 (N_15339,N_11083,N_10100);
and U15340 (N_15340,N_11328,N_10882);
or U15341 (N_15341,N_11645,N_12202);
and U15342 (N_15342,N_13641,N_13250);
nor U15343 (N_15343,N_12212,N_11374);
and U15344 (N_15344,N_12260,N_13573);
nor U15345 (N_15345,N_13220,N_13548);
nor U15346 (N_15346,N_12663,N_14582);
and U15347 (N_15347,N_13246,N_10824);
nand U15348 (N_15348,N_10147,N_14381);
or U15349 (N_15349,N_10972,N_14927);
nor U15350 (N_15350,N_11761,N_11601);
and U15351 (N_15351,N_10358,N_13603);
nand U15352 (N_15352,N_13626,N_13385);
nand U15353 (N_15353,N_10198,N_14929);
and U15354 (N_15354,N_10351,N_14883);
nand U15355 (N_15355,N_10178,N_14488);
nand U15356 (N_15356,N_14509,N_10203);
or U15357 (N_15357,N_12261,N_12040);
nor U15358 (N_15358,N_13688,N_11214);
and U15359 (N_15359,N_11200,N_13947);
nor U15360 (N_15360,N_13888,N_10850);
nand U15361 (N_15361,N_10848,N_14684);
or U15362 (N_15362,N_10019,N_12691);
nor U15363 (N_15363,N_12253,N_14321);
or U15364 (N_15364,N_11687,N_11070);
nand U15365 (N_15365,N_11421,N_12549);
nor U15366 (N_15366,N_14980,N_11545);
and U15367 (N_15367,N_14317,N_13785);
or U15368 (N_15368,N_13893,N_12216);
or U15369 (N_15369,N_12634,N_11917);
nor U15370 (N_15370,N_13840,N_12819);
nor U15371 (N_15371,N_13020,N_10819);
or U15372 (N_15372,N_13282,N_12767);
nor U15373 (N_15373,N_13919,N_11756);
and U15374 (N_15374,N_11724,N_13713);
and U15375 (N_15375,N_12684,N_14993);
nand U15376 (N_15376,N_10603,N_14277);
nor U15377 (N_15377,N_14390,N_12296);
nor U15378 (N_15378,N_14796,N_14665);
xor U15379 (N_15379,N_14402,N_12984);
nand U15380 (N_15380,N_14125,N_12215);
xnor U15381 (N_15381,N_10006,N_10960);
nor U15382 (N_15382,N_11642,N_10216);
nor U15383 (N_15383,N_10817,N_11822);
nor U15384 (N_15384,N_14749,N_13391);
nor U15385 (N_15385,N_12845,N_13367);
nand U15386 (N_15386,N_13606,N_13291);
and U15387 (N_15387,N_10426,N_10743);
or U15388 (N_15388,N_14898,N_10494);
nand U15389 (N_15389,N_12381,N_10085);
and U15390 (N_15390,N_14812,N_10995);
nor U15391 (N_15391,N_14860,N_10981);
nor U15392 (N_15392,N_14363,N_10649);
nand U15393 (N_15393,N_10797,N_12309);
nand U15394 (N_15394,N_14215,N_10729);
nand U15395 (N_15395,N_14954,N_10755);
xnor U15396 (N_15396,N_11746,N_13535);
nand U15397 (N_15397,N_13414,N_13080);
or U15398 (N_15398,N_11574,N_13227);
and U15399 (N_15399,N_10545,N_10849);
nor U15400 (N_15400,N_12306,N_13329);
nand U15401 (N_15401,N_14719,N_13571);
or U15402 (N_15402,N_10302,N_11983);
nor U15403 (N_15403,N_13855,N_13663);
xor U15404 (N_15404,N_11073,N_11017);
and U15405 (N_15405,N_13687,N_11773);
nand U15406 (N_15406,N_13342,N_14769);
nor U15407 (N_15407,N_14367,N_14459);
and U15408 (N_15408,N_14508,N_13989);
or U15409 (N_15409,N_10375,N_14362);
nand U15410 (N_15410,N_13630,N_10298);
and U15411 (N_15411,N_13186,N_13553);
and U15412 (N_15412,N_10377,N_12288);
xor U15413 (N_15413,N_13984,N_13229);
or U15414 (N_15414,N_13373,N_13418);
and U15415 (N_15415,N_12636,N_10841);
or U15416 (N_15416,N_13057,N_14223);
nor U15417 (N_15417,N_14098,N_14911);
or U15418 (N_15418,N_12827,N_14930);
and U15419 (N_15419,N_14463,N_13073);
nor U15420 (N_15420,N_10679,N_12157);
nor U15421 (N_15421,N_14073,N_13977);
xor U15422 (N_15422,N_14139,N_14058);
nor U15423 (N_15423,N_10518,N_10731);
nand U15424 (N_15424,N_14521,N_12981);
xor U15425 (N_15425,N_12893,N_13006);
or U15426 (N_15426,N_12480,N_14518);
xnor U15427 (N_15427,N_13510,N_13894);
nand U15428 (N_15428,N_12625,N_12935);
nand U15429 (N_15429,N_12970,N_14716);
nor U15430 (N_15430,N_14755,N_13583);
nor U15431 (N_15431,N_11414,N_11927);
nor U15432 (N_15432,N_14961,N_10990);
nor U15433 (N_15433,N_10152,N_14345);
or U15434 (N_15434,N_10174,N_11103);
or U15435 (N_15435,N_10226,N_11627);
or U15436 (N_15436,N_12398,N_13970);
and U15437 (N_15437,N_11120,N_11033);
nand U15438 (N_15438,N_14998,N_11282);
nand U15439 (N_15439,N_12668,N_13651);
nand U15440 (N_15440,N_14619,N_11921);
and U15441 (N_15441,N_11295,N_13699);
and U15442 (N_15442,N_13400,N_14742);
or U15443 (N_15443,N_13141,N_13394);
nand U15444 (N_15444,N_12133,N_10811);
nor U15445 (N_15445,N_14729,N_12487);
and U15446 (N_15446,N_11948,N_10110);
nor U15447 (N_15447,N_12136,N_12598);
or U15448 (N_15448,N_13381,N_12741);
nor U15449 (N_15449,N_13299,N_10013);
or U15450 (N_15450,N_10973,N_13352);
and U15451 (N_15451,N_10620,N_13454);
or U15452 (N_15452,N_10059,N_13268);
and U15453 (N_15453,N_14061,N_11286);
and U15454 (N_15454,N_13124,N_14401);
nor U15455 (N_15455,N_10886,N_14612);
nor U15456 (N_15456,N_11260,N_11183);
nand U15457 (N_15457,N_10321,N_11475);
xnor U15458 (N_15458,N_11664,N_10961);
or U15459 (N_15459,N_11052,N_13964);
and U15460 (N_15460,N_14739,N_10246);
nor U15461 (N_15461,N_14555,N_11250);
or U15462 (N_15462,N_14148,N_14001);
nor U15463 (N_15463,N_14193,N_12840);
xor U15464 (N_15464,N_12382,N_12150);
nand U15465 (N_15465,N_12265,N_11843);
or U15466 (N_15466,N_11592,N_12110);
nand U15467 (N_15467,N_11833,N_14562);
nand U15468 (N_15468,N_11406,N_10626);
xnor U15469 (N_15469,N_12994,N_13852);
nand U15470 (N_15470,N_11739,N_10526);
nor U15471 (N_15471,N_11911,N_11838);
nor U15472 (N_15472,N_12966,N_13361);
nor U15473 (N_15473,N_14206,N_11629);
nor U15474 (N_15474,N_10654,N_12046);
or U15475 (N_15475,N_13231,N_10918);
or U15476 (N_15476,N_11202,N_10877);
or U15477 (N_15477,N_13046,N_10653);
nand U15478 (N_15478,N_11916,N_14484);
or U15479 (N_15479,N_10386,N_11538);
and U15480 (N_15480,N_14782,N_12807);
nor U15481 (N_15481,N_13370,N_13783);
xnor U15482 (N_15482,N_12696,N_12861);
or U15483 (N_15483,N_10264,N_10118);
and U15484 (N_15484,N_12113,N_12195);
nor U15485 (N_15485,N_13797,N_12865);
or U15486 (N_15486,N_12906,N_14632);
nor U15487 (N_15487,N_10456,N_10781);
nand U15488 (N_15488,N_13114,N_13421);
nor U15489 (N_15489,N_14734,N_10472);
nand U15490 (N_15490,N_13388,N_14169);
nand U15491 (N_15491,N_10183,N_12364);
or U15492 (N_15492,N_12976,N_11265);
and U15493 (N_15493,N_13259,N_11388);
and U15494 (N_15494,N_13127,N_12553);
nor U15495 (N_15495,N_13420,N_10942);
nor U15496 (N_15496,N_14743,N_14520);
nand U15497 (N_15497,N_10370,N_13089);
or U15498 (N_15498,N_11300,N_14633);
nand U15499 (N_15499,N_12009,N_12600);
nand U15500 (N_15500,N_13646,N_13508);
nor U15501 (N_15501,N_10768,N_14583);
and U15502 (N_15502,N_10567,N_10634);
and U15503 (N_15503,N_12890,N_13774);
and U15504 (N_15504,N_11057,N_13684);
and U15505 (N_15505,N_12773,N_11126);
xor U15506 (N_15506,N_10201,N_13217);
or U15507 (N_15507,N_13676,N_13251);
nor U15508 (N_15508,N_10565,N_13788);
xor U15509 (N_15509,N_13110,N_14952);
nor U15510 (N_15510,N_11438,N_11700);
and U15511 (N_15511,N_14574,N_12315);
nand U15512 (N_15512,N_12705,N_13144);
nand U15513 (N_15513,N_11325,N_14029);
nand U15514 (N_15514,N_12412,N_11075);
or U15515 (N_15515,N_14646,N_13584);
nor U15516 (N_15516,N_14413,N_13578);
and U15517 (N_15517,N_11259,N_11345);
and U15518 (N_15518,N_11298,N_10955);
nand U15519 (N_15519,N_11512,N_12321);
nor U15520 (N_15520,N_10821,N_11723);
nor U15521 (N_15521,N_14685,N_10279);
nor U15522 (N_15522,N_11753,N_12162);
nand U15523 (N_15523,N_12479,N_11373);
nand U15524 (N_15524,N_10388,N_11975);
nand U15525 (N_15525,N_11868,N_14981);
nor U15526 (N_15526,N_10315,N_12645);
nor U15527 (N_15527,N_12495,N_14610);
nor U15528 (N_15528,N_12060,N_13937);
and U15529 (N_15529,N_12410,N_13596);
and U15530 (N_15530,N_12754,N_12978);
and U15531 (N_15531,N_14165,N_10860);
or U15532 (N_15532,N_14744,N_12622);
nand U15533 (N_15533,N_14937,N_14260);
or U15534 (N_15534,N_13972,N_11755);
nand U15535 (N_15535,N_14542,N_14551);
or U15536 (N_15536,N_14259,N_13835);
and U15537 (N_15537,N_12746,N_10151);
or U15538 (N_15538,N_13461,N_14393);
and U15539 (N_15539,N_10578,N_11293);
nand U15540 (N_15540,N_10055,N_13496);
or U15541 (N_15541,N_11873,N_11321);
nor U15542 (N_15542,N_11161,N_14008);
nand U15543 (N_15543,N_11430,N_13568);
or U15544 (N_15544,N_11100,N_14836);
and U15545 (N_15545,N_11251,N_13660);
nand U15546 (N_15546,N_10415,N_11456);
or U15547 (N_15547,N_13701,N_13277);
or U15548 (N_15548,N_11800,N_11102);
and U15549 (N_15549,N_13376,N_10148);
xor U15550 (N_15550,N_10812,N_14270);
nand U15551 (N_15551,N_14184,N_12312);
nor U15552 (N_15552,N_10215,N_13820);
or U15553 (N_15553,N_12948,N_13537);
or U15554 (N_15554,N_14995,N_12269);
and U15555 (N_15555,N_11937,N_13861);
nand U15556 (N_15556,N_12949,N_14496);
or U15557 (N_15557,N_12720,N_12494);
nor U15558 (N_15558,N_13570,N_12273);
xnor U15559 (N_15559,N_11178,N_13781);
or U15560 (N_15560,N_10460,N_13497);
and U15561 (N_15561,N_10748,N_13094);
and U15562 (N_15562,N_14392,N_11352);
nand U15563 (N_15563,N_10698,N_13880);
and U15564 (N_15564,N_10879,N_14853);
xnor U15565 (N_15565,N_14281,N_10138);
and U15566 (N_15566,N_11537,N_13514);
and U15567 (N_15567,N_13275,N_10457);
and U15568 (N_15568,N_12919,N_10396);
xor U15569 (N_15569,N_13230,N_13485);
nand U15570 (N_15570,N_10080,N_10208);
and U15571 (N_15571,N_11455,N_10419);
and U15572 (N_15572,N_12714,N_11151);
nand U15573 (N_15573,N_13940,N_12179);
or U15574 (N_15574,N_10774,N_10031);
nor U15575 (N_15575,N_10016,N_12752);
nor U15576 (N_15576,N_12947,N_10051);
and U15577 (N_15577,N_13812,N_12029);
or U15578 (N_15578,N_11935,N_12290);
or U15579 (N_15579,N_13574,N_13752);
nor U15580 (N_15580,N_11003,N_10758);
xnor U15581 (N_15581,N_13027,N_11518);
or U15582 (N_15582,N_12158,N_12884);
or U15583 (N_15583,N_14458,N_11112);
nor U15584 (N_15584,N_10307,N_13287);
nor U15585 (N_15585,N_14286,N_14765);
and U15586 (N_15586,N_10788,N_12766);
nor U15587 (N_15587,N_10721,N_11283);
nor U15588 (N_15588,N_12107,N_10746);
or U15589 (N_15589,N_13223,N_10765);
nor U15590 (N_15590,N_11717,N_13029);
and U15591 (N_15591,N_13368,N_11423);
nor U15592 (N_15592,N_14100,N_10865);
nand U15593 (N_15593,N_13064,N_10543);
nand U15594 (N_15594,N_11292,N_14847);
nor U15595 (N_15595,N_11600,N_13782);
nand U15596 (N_15596,N_11740,N_11468);
xor U15597 (N_15597,N_14686,N_11277);
nor U15598 (N_15598,N_10092,N_11764);
nand U15599 (N_15599,N_10437,N_10562);
and U15600 (N_15600,N_10466,N_11550);
or U15601 (N_15601,N_10237,N_11920);
or U15602 (N_15602,N_10500,N_14454);
nand U15603 (N_15603,N_10809,N_13233);
nand U15604 (N_15604,N_11846,N_11870);
or U15605 (N_15605,N_14118,N_11199);
nand U15606 (N_15606,N_11961,N_13807);
or U15607 (N_15607,N_11203,N_10590);
xor U15608 (N_15608,N_14817,N_11150);
and U15609 (N_15609,N_10831,N_14130);
nor U15610 (N_15610,N_10953,N_14815);
xor U15611 (N_15611,N_13176,N_11365);
or U15612 (N_15612,N_11718,N_10641);
and U15613 (N_15613,N_13710,N_14011);
nor U15614 (N_15614,N_10159,N_12047);
nor U15615 (N_15615,N_11180,N_12769);
nor U15616 (N_15616,N_11834,N_13343);
and U15617 (N_15617,N_10764,N_12028);
nor U15618 (N_15618,N_12768,N_13135);
nor U15619 (N_15619,N_12627,N_12137);
and U15620 (N_15620,N_14695,N_11138);
and U15621 (N_15621,N_11386,N_13321);
or U15622 (N_15622,N_10793,N_11750);
nand U15623 (N_15623,N_10221,N_14479);
nand U15624 (N_15624,N_11043,N_12287);
nor U15625 (N_15625,N_11088,N_10897);
or U15626 (N_15626,N_13870,N_14840);
nand U15627 (N_15627,N_14820,N_12041);
and U15628 (N_15628,N_11309,N_13825);
nand U15629 (N_15629,N_13741,N_13956);
nor U15630 (N_15630,N_11050,N_10858);
xor U15631 (N_15631,N_14528,N_14615);
or U15632 (N_15632,N_10618,N_14218);
xnor U15633 (N_15633,N_12071,N_10141);
or U15634 (N_15634,N_10699,N_10125);
nor U15635 (N_15635,N_13426,N_12559);
nand U15636 (N_15636,N_11949,N_10258);
nand U15637 (N_15637,N_12579,N_14505);
nor U15638 (N_15638,N_11165,N_10504);
nor U15639 (N_15639,N_14811,N_12350);
and U15640 (N_15640,N_11612,N_14057);
nand U15641 (N_15641,N_11284,N_11596);
and U15642 (N_15642,N_10311,N_12736);
or U15643 (N_15643,N_13928,N_14282);
or U15644 (N_15644,N_11235,N_10390);
or U15645 (N_15645,N_11646,N_12087);
or U15646 (N_15646,N_12596,N_12037);
and U15647 (N_15647,N_13666,N_11858);
nand U15648 (N_15648,N_13261,N_12950);
or U15649 (N_15649,N_12224,N_10667);
and U15650 (N_15650,N_11331,N_12219);
and U15651 (N_15651,N_11318,N_12867);
and U15652 (N_15652,N_14856,N_13475);
xnor U15653 (N_15653,N_13460,N_12771);
xor U15654 (N_15654,N_10124,N_11171);
nand U15655 (N_15655,N_11483,N_14654);
nor U15656 (N_15656,N_11354,N_11672);
or U15657 (N_15657,N_11849,N_13467);
nand U15658 (N_15658,N_12640,N_13716);
or U15659 (N_15659,N_13477,N_14672);
nand U15660 (N_15660,N_14570,N_12100);
nand U15661 (N_15661,N_10612,N_10624);
or U15662 (N_15662,N_14660,N_13211);
and U15663 (N_15663,N_14162,N_12408);
and U15664 (N_15664,N_11363,N_13002);
and U15665 (N_15665,N_14287,N_12504);
nor U15666 (N_15666,N_11992,N_13226);
or U15667 (N_15667,N_14560,N_10704);
nand U15668 (N_15668,N_11758,N_11960);
or U15669 (N_15669,N_11986,N_11338);
nor U15670 (N_15670,N_11759,N_12388);
or U15671 (N_15671,N_11176,N_14485);
and U15672 (N_15672,N_13856,N_12359);
nand U15673 (N_15673,N_13383,N_11784);
nor U15674 (N_15674,N_14945,N_10313);
or U15675 (N_15675,N_11398,N_14644);
nand U15676 (N_15676,N_12999,N_11394);
and U15677 (N_15677,N_11732,N_11765);
and U15678 (N_15678,N_14504,N_11744);
nor U15679 (N_15679,N_11113,N_12117);
and U15680 (N_15680,N_12820,N_12528);
or U15681 (N_15681,N_10894,N_13860);
nand U15682 (N_15682,N_13892,N_14000);
and U15683 (N_15683,N_12012,N_11527);
nand U15684 (N_15684,N_10920,N_12648);
or U15685 (N_15685,N_14872,N_14030);
or U15686 (N_15686,N_13550,N_14906);
xnor U15687 (N_15687,N_10316,N_14662);
or U15688 (N_15688,N_13766,N_13351);
or U15689 (N_15689,N_11173,N_12561);
and U15690 (N_15690,N_11836,N_10910);
nand U15691 (N_15691,N_14298,N_10574);
and U15692 (N_15692,N_13300,N_13469);
or U15693 (N_15693,N_13281,N_12659);
or U15694 (N_15694,N_10172,N_10642);
or U15695 (N_15695,N_13062,N_12426);
xnor U15696 (N_15696,N_12721,N_14412);
and U15697 (N_15697,N_11247,N_14792);
nand U15698 (N_15698,N_11131,N_12020);
nand U15699 (N_15699,N_11532,N_14473);
nor U15700 (N_15700,N_10856,N_13492);
or U15701 (N_15701,N_12490,N_14537);
and U15702 (N_15702,N_13256,N_14951);
or U15703 (N_15703,N_13890,N_12839);
or U15704 (N_15704,N_13118,N_11548);
nor U15705 (N_15705,N_14041,N_10335);
and U15706 (N_15706,N_13237,N_11933);
nand U15707 (N_15707,N_12712,N_12537);
and U15708 (N_15708,N_11790,N_11702);
xor U15709 (N_15709,N_10002,N_10822);
or U15710 (N_15710,N_12791,N_13488);
nor U15711 (N_15711,N_10436,N_10069);
and U15712 (N_15712,N_11094,N_10056);
or U15713 (N_15713,N_14154,N_12128);
or U15714 (N_15714,N_14584,N_13501);
nor U15715 (N_15715,N_11939,N_12974);
nor U15716 (N_15716,N_12834,N_10440);
nor U15717 (N_15717,N_12155,N_14667);
and U15718 (N_15718,N_13802,N_12583);
or U15719 (N_15719,N_14048,N_10608);
or U15720 (N_15720,N_12973,N_12774);
nand U15721 (N_15721,N_10224,N_10490);
nor U15722 (N_15722,N_14923,N_12238);
or U15723 (N_15723,N_11291,N_14040);
nor U15724 (N_15724,N_11585,N_13528);
or U15725 (N_15725,N_13991,N_12342);
or U15726 (N_15726,N_14017,N_13679);
nand U15727 (N_15727,N_10406,N_10757);
and U15728 (N_15728,N_14649,N_10883);
or U15729 (N_15729,N_11168,N_12749);
nor U15730 (N_15730,N_12399,N_10288);
or U15731 (N_15731,N_14885,N_13643);
nor U15732 (N_15732,N_12051,N_11495);
and U15733 (N_15733,N_14786,N_13930);
and U15734 (N_15734,N_12022,N_12278);
nor U15735 (N_15735,N_12591,N_10077);
nor U15736 (N_15736,N_11661,N_10365);
nor U15737 (N_15737,N_12015,N_12888);
and U15738 (N_15738,N_12082,N_13362);
nor U15739 (N_15739,N_14994,N_12325);
or U15740 (N_15740,N_11730,N_10064);
nor U15741 (N_15741,N_10303,N_13513);
nand U15742 (N_15742,N_13434,N_12166);
or U15743 (N_15743,N_14177,N_12914);
nor U15744 (N_15744,N_13452,N_13402);
and U15745 (N_15745,N_10360,N_13609);
nand U15746 (N_15746,N_11267,N_14530);
nand U15747 (N_15747,N_12863,N_11864);
nor U15748 (N_15748,N_14721,N_13273);
xor U15749 (N_15749,N_11053,N_10000);
xnor U15750 (N_15750,N_11697,N_12868);
and U15751 (N_15751,N_12709,N_12869);
nor U15752 (N_15752,N_12930,N_11375);
nor U15753 (N_15753,N_13816,N_10719);
nand U15754 (N_15754,N_11853,N_14826);
nor U15755 (N_15755,N_12274,N_11445);
xnor U15756 (N_15756,N_11163,N_13015);
and U15757 (N_15757,N_14910,N_10715);
and U15758 (N_15758,N_10863,N_10710);
nor U15759 (N_15759,N_14631,N_12817);
nand U15760 (N_15760,N_13150,N_10688);
or U15761 (N_15761,N_13932,N_10304);
xor U15762 (N_15762,N_13724,N_13714);
nor U15763 (N_15763,N_12623,N_12782);
and U15764 (N_15764,N_13119,N_11734);
and U15765 (N_15765,N_13204,N_11872);
nand U15766 (N_15766,N_12954,N_10026);
and U15767 (N_15767,N_13463,N_14349);
and U15768 (N_15768,N_14781,N_14494);
and U15769 (N_15769,N_12523,N_10692);
and U15770 (N_15770,N_14262,N_12647);
xnor U15771 (N_15771,N_12681,N_12814);
and U15772 (N_15772,N_12711,N_13677);
nand U15773 (N_15773,N_10182,N_14032);
or U15774 (N_15774,N_11233,N_14882);
or U15775 (N_15775,N_11348,N_12698);
nand U15776 (N_15776,N_13013,N_11851);
nand U15777 (N_15777,N_11107,N_11708);
and U15778 (N_15778,N_10691,N_14801);
xor U15779 (N_15779,N_11119,N_12610);
nor U15780 (N_15780,N_11774,N_14664);
nand U15781 (N_15781,N_11656,N_11658);
nor U15782 (N_15782,N_11787,N_11551);
and U15783 (N_15783,N_11329,N_11418);
or U15784 (N_15784,N_13443,N_13992);
nand U15785 (N_15785,N_13419,N_11169);
nor U15786 (N_15786,N_13854,N_11429);
nand U15787 (N_15787,N_10847,N_11319);
or U15788 (N_15788,N_14904,N_11659);
nor U15789 (N_15789,N_11114,N_11015);
xor U15790 (N_15790,N_14140,N_12843);
and U15791 (N_15791,N_10452,N_10636);
or U15792 (N_15792,N_10989,N_12624);
nor U15793 (N_15793,N_14449,N_12217);
or U15794 (N_15794,N_13210,N_12565);
and U15795 (N_15795,N_13047,N_13473);
nand U15796 (N_15796,N_13563,N_10291);
and U15797 (N_15797,N_11485,N_10593);
and U15798 (N_15798,N_10366,N_11639);
nor U15799 (N_15799,N_14372,N_10496);
or U15800 (N_15800,N_10123,N_11798);
or U15801 (N_15801,N_12609,N_13795);
nand U15802 (N_15802,N_10652,N_11496);
nor U15803 (N_15803,N_11662,N_11245);
nand U15804 (N_15804,N_10121,N_11899);
or U15805 (N_15805,N_14962,N_10434);
xnor U15806 (N_15806,N_10951,N_10648);
nand U15807 (N_15807,N_13215,N_13702);
or U15808 (N_15808,N_13472,N_14939);
or U15809 (N_15809,N_11140,N_10589);
or U15810 (N_15810,N_10628,N_10270);
xor U15811 (N_15811,N_11912,N_11181);
and U15812 (N_15812,N_10355,N_12203);
or U15813 (N_15813,N_10444,N_11258);
xnor U15814 (N_15814,N_12761,N_14155);
xor U15815 (N_15815,N_10592,N_12654);
nor U15816 (N_15816,N_14627,N_12126);
nand U15817 (N_15817,N_10572,N_10650);
nor U15818 (N_15818,N_13591,N_11816);
nand U15819 (N_15819,N_11488,N_11544);
xor U15820 (N_15820,N_14959,N_12436);
nand U15821 (N_15821,N_10061,N_10282);
nor U15822 (N_15822,N_13655,N_10011);
nor U15823 (N_15823,N_14854,N_12038);
nand U15824 (N_15824,N_13462,N_13133);
nand U15825 (N_15825,N_12170,N_11945);
nor U15826 (N_15826,N_10331,N_14265);
nand U15827 (N_15827,N_12924,N_14269);
nand U15828 (N_15828,N_14129,N_11419);
or U15829 (N_15829,N_11068,N_12729);
nor U15830 (N_15830,N_10890,N_11978);
or U15831 (N_15831,N_12540,N_13415);
nand U15832 (N_15832,N_12655,N_13585);
and U15833 (N_15833,N_11145,N_13294);
nor U15834 (N_15834,N_10079,N_13398);
or U15835 (N_15835,N_11137,N_12004);
nor U15836 (N_15836,N_12332,N_12560);
nand U15837 (N_15837,N_12220,N_11023);
or U15838 (N_15838,N_13173,N_14348);
and U15839 (N_15839,N_11317,N_14795);
xnor U15840 (N_15840,N_14813,N_11826);
xor U15841 (N_15841,N_14880,N_12095);
or U15842 (N_15842,N_14502,N_13909);
nand U15843 (N_15843,N_12064,N_14989);
nor U15844 (N_15844,N_10867,N_12106);
or U15845 (N_15845,N_11632,N_13773);
and U15846 (N_15846,N_14127,N_10933);
xnor U15847 (N_15847,N_12291,N_12434);
or U15848 (N_15848,N_13429,N_12246);
nor U15849 (N_15849,N_13380,N_12200);
and U15850 (N_15850,N_13406,N_14620);
xor U15851 (N_15851,N_12519,N_11618);
and U15852 (N_15852,N_12039,N_14731);
or U15853 (N_15853,N_13665,N_10815);
or U15854 (N_15854,N_11876,N_10658);
nor U15855 (N_15855,N_14843,N_13610);
nand U15856 (N_15856,N_12959,N_12149);
or U15857 (N_15857,N_12176,N_10529);
nor U15858 (N_15858,N_12237,N_11111);
nor U15859 (N_15859,N_11091,N_14387);
or U15860 (N_15860,N_14301,N_14578);
nor U15861 (N_15861,N_13876,N_11982);
nand U15862 (N_15862,N_12423,N_11820);
or U15863 (N_15863,N_13490,N_11540);
or U15864 (N_15864,N_10881,N_12193);
nor U15865 (N_15865,N_11256,N_12470);
nand U15866 (N_15866,N_10761,N_13090);
and U15867 (N_15867,N_12633,N_11002);
or U15868 (N_15868,N_13447,N_12473);
or U15869 (N_15869,N_14388,N_14775);
xor U15870 (N_15870,N_10619,N_12129);
or U15871 (N_15871,N_10602,N_10310);
xnor U15872 (N_15872,N_10336,N_12207);
xnor U15873 (N_15873,N_14766,N_12322);
and U15874 (N_15874,N_13389,N_13072);
nor U15875 (N_15875,N_14635,N_12152);
nor U15876 (N_15876,N_13734,N_11788);
xor U15877 (N_15877,N_12079,N_11821);
and U15878 (N_15878,N_12832,N_12351);
nor U15879 (N_15879,N_10747,N_12983);
xor U15880 (N_15880,N_10607,N_12837);
xnor U15881 (N_15881,N_14087,N_12103);
and U15882 (N_15882,N_13516,N_14586);
nand U15883 (N_15883,N_10616,N_10766);
nand U15884 (N_15884,N_12532,N_14572);
nand U15885 (N_15885,N_14236,N_11729);
xnor U15886 (N_15886,N_12205,N_14136);
and U15887 (N_15887,N_11886,N_13994);
or U15888 (N_15888,N_13209,N_11097);
nor U15889 (N_15889,N_11953,N_11380);
nand U15890 (N_15890,N_14096,N_14196);
nand U15891 (N_15891,N_14010,N_12448);
nand U15892 (N_15892,N_13975,N_14222);
xnor U15893 (N_15893,N_11990,N_12085);
or U15894 (N_15894,N_10435,N_14679);
or U15895 (N_15895,N_14947,N_10724);
and U15896 (N_15896,N_14421,N_13744);
nor U15897 (N_15897,N_11908,N_13161);
or U15898 (N_15898,N_14203,N_11617);
nor U15899 (N_15899,N_12883,N_12526);
or U15900 (N_15900,N_13945,N_10372);
and U15901 (N_15901,N_11799,N_10384);
or U15902 (N_15902,N_10488,N_10350);
nor U15903 (N_15903,N_11623,N_11615);
or U15904 (N_15904,N_14736,N_10241);
nor U15905 (N_15905,N_11275,N_10248);
xor U15906 (N_15906,N_10807,N_13430);
nor U15907 (N_15907,N_10674,N_13654);
nand U15908 (N_15908,N_11875,N_10694);
and U15909 (N_15909,N_14598,N_13562);
nand U15910 (N_15910,N_12415,N_11752);
and U15911 (N_15911,N_13465,N_13926);
nand U15912 (N_15912,N_14879,N_11595);
and U15913 (N_15913,N_14591,N_11358);
nor U15914 (N_15914,N_10114,N_13614);
and U15915 (N_15915,N_11128,N_13470);
or U15916 (N_15916,N_12138,N_10838);
and U15917 (N_15917,N_11508,N_13948);
nand U15918 (N_15918,N_14360,N_13091);
nor U15919 (N_15919,N_14707,N_13637);
and U15920 (N_15920,N_12008,N_12894);
xnor U15921 (N_15921,N_12283,N_12898);
and U15922 (N_15922,N_12165,N_10143);
nor U15923 (N_15923,N_11666,N_11311);
and U15924 (N_15924,N_14442,N_12175);
or U15925 (N_15925,N_13680,N_10617);
or U15926 (N_15926,N_10495,N_10352);
and U15927 (N_15927,N_11499,N_11542);
nor U15928 (N_15928,N_11560,N_10379);
xnor U15929 (N_15929,N_14151,N_12146);
and U15930 (N_15930,N_11972,N_10922);
nor U15931 (N_15931,N_12292,N_10786);
xnor U15932 (N_15932,N_11525,N_11271);
nand U15933 (N_15933,N_12310,N_11970);
or U15934 (N_15934,N_13958,N_11510);
nor U15935 (N_15935,N_14733,N_14268);
or U15936 (N_15936,N_11671,N_11725);
nand U15937 (N_15937,N_12057,N_14821);
and U15938 (N_15938,N_11783,N_11306);
nand U15939 (N_15939,N_10107,N_14279);
and U15940 (N_15940,N_14532,N_10359);
nor U15941 (N_15941,N_14830,N_14659);
nor U15942 (N_15942,N_10711,N_10866);
or U15943 (N_15943,N_14611,N_10035);
and U15944 (N_15944,N_13879,N_12568);
nor U15945 (N_15945,N_10794,N_14899);
and U15946 (N_15946,N_14673,N_12043);
nand U15947 (N_15947,N_11462,N_11172);
nand U15948 (N_15948,N_13152,N_12988);
nand U15949 (N_15949,N_10707,N_14354);
and U15950 (N_15950,N_10461,N_10186);
and U15951 (N_15951,N_10115,N_12951);
nand U15952 (N_15952,N_12998,N_14308);
or U15953 (N_15953,N_13599,N_10645);
nor U15954 (N_15954,N_12247,N_14506);
xor U15955 (N_15955,N_13081,N_14622);
nand U15956 (N_15956,N_10146,N_12718);
and U15957 (N_15957,N_12209,N_12083);
and U15958 (N_15958,N_11228,N_12460);
or U15959 (N_15959,N_14498,N_12181);
nand U15960 (N_15960,N_12432,N_11395);
or U15961 (N_15961,N_12464,N_11519);
or U15962 (N_15962,N_12467,N_14370);
nor U15963 (N_15963,N_12403,N_11400);
and U15964 (N_15964,N_13192,N_12088);
nand U15965 (N_15965,N_13266,N_14309);
nor U15966 (N_15966,N_14323,N_11737);
xor U15967 (N_15967,N_13564,N_13847);
or U15968 (N_15968,N_14095,N_10516);
or U15969 (N_15969,N_10919,N_13315);
and U15970 (N_15970,N_13726,N_12140);
and U15971 (N_15971,N_13450,N_10129);
nand U15972 (N_15972,N_10783,N_14453);
and U15973 (N_15973,N_10696,N_12075);
or U15974 (N_15974,N_14075,N_13151);
nand U15975 (N_15975,N_10991,N_14753);
xor U15976 (N_15976,N_12571,N_13622);
and U15977 (N_15977,N_11289,N_13725);
nor U15978 (N_15978,N_14754,N_11720);
nor U15979 (N_15979,N_14229,N_11272);
xnor U15980 (N_15980,N_13608,N_10928);
or U15981 (N_15981,N_10685,N_14616);
and U15982 (N_15982,N_11032,N_13236);
nor U15983 (N_15983,N_10739,N_14202);
xnor U15984 (N_15984,N_11189,N_14974);
and U15985 (N_15985,N_13815,N_12452);
nor U15986 (N_15986,N_14807,N_14149);
or U15987 (N_15987,N_14925,N_12862);
nand U15988 (N_15988,N_11249,N_11980);
and U15989 (N_15989,N_14917,N_11686);
nand U15990 (N_15990,N_12213,N_14629);
or U15991 (N_15991,N_11915,N_10191);
xor U15992 (N_15992,N_11217,N_12345);
nor U15993 (N_15993,N_12118,N_13061);
nand U15994 (N_15994,N_12324,N_11928);
or U15995 (N_15995,N_11852,N_12544);
nand U15996 (N_15996,N_14711,N_12904);
or U15997 (N_15997,N_13617,N_13953);
nand U15998 (N_15998,N_14232,N_13732);
or U15999 (N_15999,N_13917,N_10975);
and U16000 (N_16000,N_14128,N_10207);
nand U16001 (N_16001,N_13491,N_12453);
nor U16002 (N_16002,N_10332,N_14055);
nand U16003 (N_16003,N_11981,N_10997);
and U16004 (N_16004,N_13179,N_10344);
or U16005 (N_16005,N_10199,N_13786);
or U16006 (N_16006,N_10250,N_12725);
and U16007 (N_16007,N_13648,N_10508);
or U16008 (N_16008,N_11316,N_12353);
nand U16009 (N_16009,N_14777,N_12685);
nand U16010 (N_16010,N_11004,N_12847);
or U16011 (N_16011,N_10364,N_10853);
xnor U16012 (N_16012,N_13963,N_12844);
nor U16013 (N_16013,N_13913,N_13739);
nor U16014 (N_16014,N_10892,N_11824);
nor U16015 (N_16015,N_10733,N_12556);
xnor U16016 (N_16016,N_13750,N_13954);
nand U16017 (N_16017,N_14278,N_13598);
nor U16018 (N_16018,N_11692,N_12377);
xnor U16019 (N_16019,N_12795,N_10446);
and U16020 (N_16020,N_13408,N_12151);
or U16021 (N_16021,N_14567,N_11124);
and U16022 (N_16022,N_11344,N_13286);
nand U16023 (N_16023,N_12077,N_12927);
or U16024 (N_16024,N_11881,N_10062);
nand U16025 (N_16025,N_10004,N_10873);
nor U16026 (N_16026,N_11174,N_10644);
nand U16027 (N_16027,N_14642,N_14878);
nor U16028 (N_16028,N_13661,N_13177);
nor U16029 (N_16029,N_12911,N_13936);
nand U16030 (N_16030,N_10438,N_14698);
nand U16031 (N_16031,N_10959,N_11677);
and U16032 (N_16032,N_11742,N_12331);
or U16033 (N_16033,N_13182,N_14009);
nand U16034 (N_16034,N_10548,N_11336);
nor U16035 (N_16035,N_14703,N_13787);
or U16036 (N_16036,N_14386,N_11324);
and U16037 (N_16037,N_11207,N_12178);
nor U16038 (N_16038,N_11355,N_14464);
nor U16039 (N_16039,N_12344,N_12945);
nand U16040 (N_16040,N_11848,N_12042);
or U16041 (N_16041,N_14188,N_14398);
xnor U16042 (N_16042,N_14094,N_12450);
xnor U16043 (N_16043,N_12780,N_13107);
nand U16044 (N_16044,N_14798,N_13851);
and U16045 (N_16045,N_11628,N_11413);
nand U16046 (N_16046,N_10322,N_14046);
and U16047 (N_16047,N_11709,N_14233);
nor U16048 (N_16048,N_13205,N_10800);
and U16049 (N_16049,N_13853,N_10233);
nand U16050 (N_16050,N_14207,N_10582);
or U16051 (N_16051,N_14789,N_11923);
nor U16052 (N_16052,N_14045,N_10727);
and U16053 (N_16053,N_12454,N_14471);
or U16054 (N_16054,N_11399,N_13131);
or U16055 (N_16055,N_13358,N_11695);
nor U16056 (N_16056,N_10718,N_10614);
nor U16057 (N_16057,N_10278,N_11024);
nor U16058 (N_16058,N_12430,N_12227);
nand U16059 (N_16059,N_12469,N_14477);
xor U16060 (N_16060,N_13969,N_10037);
or U16061 (N_16061,N_11340,N_13532);
nor U16062 (N_16062,N_11583,N_12199);
xnor U16063 (N_16063,N_11768,N_11366);
and U16064 (N_16064,N_12429,N_11660);
xnor U16065 (N_16065,N_10160,N_12264);
and U16066 (N_16066,N_13602,N_11847);
and U16067 (N_16067,N_12327,N_11443);
and U16068 (N_16068,N_12231,N_14183);
or U16069 (N_16069,N_12431,N_11654);
nand U16070 (N_16070,N_13916,N_13875);
and U16071 (N_16071,N_10523,N_13770);
nor U16072 (N_16072,N_11210,N_13212);
xor U16073 (N_16073,N_10039,N_11472);
nand U16074 (N_16074,N_12631,N_12035);
or U16075 (N_16075,N_10007,N_13206);
or U16076 (N_16076,N_10098,N_10507);
xor U16077 (N_16077,N_11170,N_14688);
xor U16078 (N_16078,N_14957,N_12411);
and U16079 (N_16079,N_14022,N_10742);
nand U16080 (N_16080,N_14871,N_12355);
nand U16081 (N_16081,N_11794,N_12284);
nand U16082 (N_16082,N_11498,N_13931);
and U16083 (N_16083,N_14640,N_12441);
nor U16084 (N_16084,N_13221,N_12145);
nand U16085 (N_16085,N_14770,N_13541);
or U16086 (N_16086,N_10594,N_14867);
xor U16087 (N_16087,N_10551,N_13433);
and U16088 (N_16088,N_12045,N_13925);
xor U16089 (N_16089,N_14571,N_13034);
nand U16090 (N_16090,N_10528,N_10017);
nor U16091 (N_16091,N_10632,N_11840);
or U16092 (N_16092,N_12197,N_10261);
or U16093 (N_16093,N_11684,N_13427);
nor U16094 (N_16094,N_12853,N_13067);
nor U16095 (N_16095,N_13705,N_10140);
nand U16096 (N_16096,N_10916,N_13163);
or U16097 (N_16097,N_13500,N_12702);
and U16098 (N_16098,N_10214,N_11327);
and U16099 (N_16099,N_10655,N_14007);
or U16100 (N_16100,N_11584,N_12191);
and U16101 (N_16101,N_12011,N_12090);
or U16102 (N_16102,N_14174,N_11297);
xor U16103 (N_16103,N_12604,N_12686);
nand U16104 (N_16104,N_10818,N_14197);
nor U16105 (N_16105,N_12792,N_13041);
nor U16106 (N_16106,N_13762,N_13147);
nand U16107 (N_16107,N_13738,N_14849);
xor U16108 (N_16108,N_13946,N_14868);
nand U16109 (N_16109,N_12842,N_13850);
and U16110 (N_16110,N_10756,N_10714);
nor U16111 (N_16111,N_10253,N_10163);
nor U16112 (N_16112,N_12500,N_11404);
xor U16113 (N_16113,N_13554,N_11505);
xnor U16114 (N_16114,N_13035,N_13594);
nor U16115 (N_16115,N_12222,N_14102);
nor U16116 (N_16116,N_11432,N_12759);
nor U16117 (N_16117,N_11604,N_13729);
and U16118 (N_16118,N_10405,N_11493);
nand U16119 (N_16119,N_10341,N_11835);
xnor U16120 (N_16120,N_12533,N_13938);
or U16121 (N_16121,N_10181,N_12013);
xnor U16122 (N_16122,N_13518,N_11254);
or U16123 (N_16123,N_12081,N_14242);
nor U16124 (N_16124,N_11653,N_13867);
or U16125 (N_16125,N_14145,N_11607);
or U16126 (N_16126,N_14759,N_11268);
and U16127 (N_16127,N_12148,N_11706);
or U16128 (N_16128,N_11359,N_13728);
and U16129 (N_16129,N_13324,N_12676);
nor U16130 (N_16130,N_12692,N_10623);
nor U16131 (N_16131,N_10734,N_13017);
nor U16132 (N_16132,N_14838,N_14358);
nand U16133 (N_16133,N_11556,N_14706);
or U16134 (N_16134,N_12400,N_12551);
and U16135 (N_16135,N_13809,N_14536);
nand U16136 (N_16136,N_13301,N_10014);
or U16137 (N_16137,N_14462,N_14005);
and U16138 (N_16138,N_12534,N_14804);
or U16139 (N_16139,N_13922,N_14124);
and U16140 (N_16140,N_11269,N_10367);
nor U16141 (N_16141,N_10433,N_10709);
and U16142 (N_16142,N_14767,N_13955);
and U16143 (N_16143,N_12232,N_14566);
nand U16144 (N_16144,N_11007,N_13611);
nor U16145 (N_16145,N_14158,N_13625);
and U16146 (N_16146,N_11037,N_12608);
or U16147 (N_16147,N_13098,N_14888);
or U16148 (N_16148,N_11900,N_12941);
nand U16149 (N_16149,N_12225,N_10985);
or U16150 (N_16150,N_13834,N_12929);
nand U16151 (N_16151,N_14827,N_10868);
and U16152 (N_16152,N_11904,N_13831);
and U16153 (N_16153,N_10837,N_10763);
or U16154 (N_16154,N_14693,N_13924);
nor U16155 (N_16155,N_10965,N_11898);
or U16156 (N_16156,N_13038,N_13010);
and U16157 (N_16157,N_11326,N_13842);
or U16158 (N_16158,N_12543,N_12187);
and U16159 (N_16159,N_13878,N_14049);
or U16160 (N_16160,N_14784,N_13674);
xnor U16161 (N_16161,N_11048,N_10429);
xor U16162 (N_16162,N_10090,N_14913);
and U16163 (N_16163,N_11625,N_13102);
xnor U16164 (N_16164,N_14519,N_10483);
and U16165 (N_16165,N_12689,N_10491);
or U16166 (N_16166,N_14933,N_10103);
or U16167 (N_16167,N_11453,N_12594);
nor U16168 (N_16168,N_12688,N_12241);
or U16169 (N_16169,N_12070,N_11555);
and U16170 (N_16170,N_12765,N_14680);
or U16171 (N_16171,N_12606,N_14595);
xor U16172 (N_16172,N_10795,N_11893);
and U16173 (N_16173,N_13826,N_12779);
nand U16174 (N_16174,N_14576,N_14663);
and U16175 (N_16175,N_12527,N_12346);
xor U16176 (N_16176,N_14985,N_13422);
and U16177 (N_16177,N_10173,N_12650);
nand U16178 (N_16178,N_13123,N_11964);
or U16179 (N_16179,N_14231,N_14546);
or U16180 (N_16180,N_11839,N_10034);
or U16181 (N_16181,N_13228,N_12885);
xnor U16182 (N_16182,N_13547,N_12174);
nor U16183 (N_16183,N_10323,N_12651);
nor U16184 (N_16184,N_11313,N_12433);
nand U16185 (N_16185,N_14216,N_14164);
nor U16186 (N_16186,N_10802,N_11294);
nor U16187 (N_16187,N_12418,N_13957);
nand U16188 (N_16188,N_13138,N_11565);
nand U16189 (N_16189,N_13076,N_10380);
xor U16190 (N_16190,N_14436,N_13283);
and U16191 (N_16191,N_11296,N_12280);
nor U16192 (N_16192,N_10431,N_13566);
and U16193 (N_16193,N_13592,N_13801);
nor U16194 (N_16194,N_13448,N_11865);
nor U16195 (N_16195,N_11148,N_13239);
nand U16196 (N_16196,N_11440,N_13155);
or U16197 (N_16197,N_13316,N_10934);
and U16198 (N_16198,N_13187,N_11186);
nor U16199 (N_16199,N_11257,N_14745);
or U16200 (N_16200,N_12602,N_14714);
and U16201 (N_16201,N_14263,N_11482);
or U16202 (N_16202,N_10428,N_13142);
nand U16203 (N_16203,N_11597,N_14455);
nand U16204 (N_16204,N_12603,N_13743);
nand U16205 (N_16205,N_13658,N_14705);
xor U16206 (N_16206,N_12092,N_13355);
or U16207 (N_16207,N_13549,N_14292);
nand U16208 (N_16208,N_13525,N_14235);
and U16209 (N_16209,N_11909,N_14992);
and U16210 (N_16210,N_13423,N_14750);
and U16211 (N_16211,N_10086,N_10058);
xnor U16212 (N_16212,N_10682,N_13873);
or U16213 (N_16213,N_12122,N_10418);
nor U16214 (N_16214,N_12588,N_10912);
nor U16215 (N_16215,N_12667,N_11231);
and U16216 (N_16216,N_10993,N_10662);
and U16217 (N_16217,N_12573,N_14108);
nand U16218 (N_16218,N_11005,N_13999);
or U16219 (N_16219,N_14335,N_12142);
or U16220 (N_16220,N_10206,N_14738);
or U16221 (N_16221,N_11775,N_12267);
and U16222 (N_16222,N_12115,N_14920);
and U16223 (N_16223,N_11011,N_13691);
nand U16224 (N_16224,N_14643,N_11044);
nor U16225 (N_16225,N_11796,N_11451);
or U16226 (N_16226,N_14889,N_14589);
or U16227 (N_16227,N_11913,N_14967);
and U16228 (N_16228,N_12307,N_12093);
nor U16229 (N_16229,N_11652,N_14337);
xnor U16230 (N_16230,N_11401,N_12440);
xor U16231 (N_16231,N_13849,N_10078);
nor U16232 (N_16232,N_11407,N_13889);
xor U16233 (N_16233,N_10409,N_12135);
nand U16234 (N_16234,N_12569,N_10736);
nand U16235 (N_16235,N_11857,N_13456);
nand U16236 (N_16236,N_14150,N_10042);
nor U16237 (N_16237,N_14613,N_11109);
or U16238 (N_16238,N_11614,N_12266);
nor U16239 (N_16239,N_10421,N_14076);
nand U16240 (N_16240,N_13512,N_11143);
nand U16241 (N_16241,N_13779,N_14730);
nand U16242 (N_16242,N_10142,N_12809);
nor U16243 (N_16243,N_12120,N_13526);
nand U16244 (N_16244,N_12778,N_10665);
nand U16245 (N_16245,N_11342,N_10629);
nand U16246 (N_16246,N_10932,N_12986);
nor U16247 (N_16247,N_14973,N_14318);
and U16248 (N_16248,N_10505,N_10969);
nand U16249 (N_16249,N_14647,N_11710);
and U16250 (N_16250,N_14712,N_12067);
or U16251 (N_16251,N_12285,N_11929);
or U16252 (N_16252,N_12063,N_12548);
nor U16253 (N_16253,N_14905,N_14152);
or U16254 (N_16254,N_12255,N_10832);
nor U16255 (N_16255,N_10235,N_11305);
nor U16256 (N_16256,N_13322,N_14932);
nor U16257 (N_16257,N_10371,N_13401);
nor U16258 (N_16258,N_14683,N_11435);
nor U16259 (N_16259,N_12997,N_11497);
nor U16260 (N_16260,N_14580,N_10559);
nor U16261 (N_16261,N_10326,N_14395);
nand U16262 (N_16262,N_11335,N_14084);
xnor U16263 (N_16263,N_10683,N_12895);
and U16264 (N_16264,N_10043,N_10362);
xor U16265 (N_16265,N_11778,N_10647);
and U16266 (N_16266,N_11219,N_11942);
nor U16267 (N_16267,N_14912,N_11895);
or U16268 (N_16268,N_11288,N_13494);
nand U16269 (N_16269,N_11158,N_11998);
nand U16270 (N_16270,N_14556,N_10861);
xor U16271 (N_16271,N_11531,N_13943);
nor U16272 (N_16272,N_12263,N_14652);
nand U16273 (N_16273,N_10324,N_10726);
nor U16274 (N_16274,N_14511,N_12990);
or U16275 (N_16275,N_13284,N_11795);
xor U16276 (N_16276,N_11022,N_10782);
and U16277 (N_16277,N_10750,N_13683);
nor U16278 (N_16278,N_13318,N_10905);
or U16279 (N_16279,N_12518,N_10728);
or U16280 (N_16280,N_10760,N_11974);
and U16281 (N_16281,N_13445,N_10139);
nand U16282 (N_16282,N_11479,N_10656);
xnor U16283 (N_16283,N_10289,N_12513);
and U16284 (N_16284,N_11175,N_11722);
nor U16285 (N_16285,N_13241,N_14524);
and U16286 (N_16286,N_10534,N_10531);
nand U16287 (N_16287,N_10387,N_12328);
nor U16288 (N_16288,N_12793,N_12405);
and U16289 (N_16289,N_12920,N_11422);
or U16290 (N_16290,N_13431,N_13392);
nand U16291 (N_16291,N_11626,N_14093);
and U16292 (N_16292,N_10827,N_14214);
and U16293 (N_16293,N_13897,N_11786);
or U16294 (N_16294,N_13996,N_13753);
nand U16295 (N_16295,N_13776,N_13122);
or U16296 (N_16296,N_13664,N_13764);
and U16297 (N_16297,N_10519,N_11803);
or U16298 (N_16298,N_13437,N_13981);
and U16299 (N_16299,N_13264,N_14342);
xor U16300 (N_16300,N_12672,N_13546);
nand U16301 (N_16301,N_14873,N_11649);
nand U16302 (N_16302,N_11035,N_10536);
and U16303 (N_16303,N_10787,N_11529);
nor U16304 (N_16304,N_13757,N_14305);
or U16305 (N_16305,N_14944,N_11058);
or U16306 (N_16306,N_12656,N_14517);
nand U16307 (N_16307,N_13317,N_13959);
nor U16308 (N_16308,N_14245,N_14700);
or U16309 (N_16309,N_14178,N_13464);
or U16310 (N_16310,N_11559,N_12352);
or U16311 (N_16311,N_14818,N_14825);
nand U16312 (N_16312,N_12755,N_10382);
nand U16313 (N_16313,N_11061,N_13864);
and U16314 (N_16314,N_14564,N_14002);
nand U16315 (N_16315,N_14378,N_10568);
or U16316 (N_16316,N_11855,N_12562);
or U16317 (N_16317,N_14452,N_14928);
nand U16318 (N_16318,N_10353,N_12652);
xnor U16319 (N_16319,N_11402,N_10675);
or U16320 (N_16320,N_14435,N_14384);
and U16321 (N_16321,N_10880,N_13476);
and U16322 (N_16322,N_11640,N_11989);
xor U16323 (N_16323,N_13718,N_11831);
and U16324 (N_16324,N_10520,N_10430);
and U16325 (N_16325,N_13813,N_11648);
nand U16326 (N_16326,N_13911,N_11956);
nor U16327 (N_16327,N_10979,N_12946);
xnor U16328 (N_16328,N_10798,N_11397);
or U16329 (N_16329,N_13130,N_10722);
or U16330 (N_16330,N_13252,N_12743);
nand U16331 (N_16331,N_11159,N_10512);
or U16332 (N_16332,N_14290,N_10752);
or U16333 (N_16333,N_12979,N_13082);
or U16334 (N_16334,N_10631,N_11478);
and U16335 (N_16335,N_14423,N_12635);
nor U16336 (N_16336,N_12642,N_13511);
and U16337 (N_16337,N_14450,N_12800);
nor U16338 (N_16338,N_13695,N_10712);
xor U16339 (N_16339,N_11805,N_10911);
and U16340 (N_16340,N_14312,N_14857);
nand U16341 (N_16341,N_11698,N_10871);
or U16342 (N_16342,N_12738,N_11382);
or U16343 (N_16343,N_11135,N_11393);
xor U16344 (N_16344,N_10068,N_13105);
nand U16345 (N_16345,N_14587,N_11157);
nand U16346 (N_16346,N_13978,N_13749);
nor U16347 (N_16347,N_11049,N_10643);
nor U16348 (N_16348,N_14043,N_10732);
nor U16349 (N_16349,N_14250,N_13973);
and U16350 (N_16350,N_13332,N_13558);
nand U16351 (N_16351,N_11206,N_13843);
nand U16352 (N_16352,N_13671,N_13862);
nand U16353 (N_16353,N_11903,N_14355);
nor U16354 (N_16354,N_12343,N_13063);
nand U16355 (N_16355,N_10576,N_12073);
nor U16356 (N_16356,N_13615,N_13338);
nand U16357 (N_16357,N_14264,N_12892);
and U16358 (N_16358,N_14788,N_12938);
or U16359 (N_16359,N_12101,N_13837);
or U16360 (N_16360,N_13449,N_11558);
and U16361 (N_16361,N_14539,N_14588);
or U16362 (N_16362,N_12401,N_13884);
nand U16363 (N_16363,N_13707,N_14034);
xor U16364 (N_16364,N_12127,N_10799);
and U16365 (N_16365,N_10595,N_14977);
nand U16366 (N_16366,N_13159,N_10479);
nand U16367 (N_16367,N_10256,N_10378);
nand U16368 (N_16368,N_12491,N_10108);
nor U16369 (N_16369,N_11089,N_11714);
and U16370 (N_16370,N_12438,N_10188);
and U16371 (N_16371,N_13712,N_10779);
or U16372 (N_16372,N_11444,N_12742);
or U16373 (N_16373,N_11749,N_11667);
nand U16374 (N_16374,N_10762,N_10956);
nand U16375 (N_16375,N_13686,N_13883);
and U16376 (N_16376,N_13325,N_12514);
and U16377 (N_16377,N_12790,N_10530);
or U16378 (N_16378,N_14809,N_11491);
or U16379 (N_16379,N_12485,N_11090);
and U16380 (N_16380,N_13822,N_11602);
nor U16381 (N_16381,N_10547,N_13914);
and U16382 (N_16382,N_13481,N_13360);
nor U16383 (N_16383,N_12758,N_14751);
and U16384 (N_16384,N_11424,N_10935);
or U16385 (N_16385,N_11001,N_12096);
nor U16386 (N_16386,N_14172,N_13976);
xnor U16387 (N_16387,N_13735,N_12787);
nand U16388 (N_16388,N_12484,N_14243);
and U16389 (N_16389,N_10717,N_13058);
xnor U16390 (N_16390,N_12293,N_10455);
and U16391 (N_16391,N_12875,N_12049);
xnor U16392 (N_16392,N_12183,N_14208);
and U16393 (N_16393,N_13480,N_11930);
and U16394 (N_16394,N_12961,N_13297);
or U16395 (N_16395,N_10204,N_11549);
nor U16396 (N_16396,N_10363,N_14416);
nor U16397 (N_16397,N_14936,N_12601);
or U16398 (N_16398,N_12402,N_13742);
or U16399 (N_16399,N_12297,N_10982);
or U16400 (N_16400,N_12848,N_11827);
nand U16401 (N_16401,N_13804,N_11025);
nor U16402 (N_16402,N_14953,N_12972);
nor U16403 (N_16403,N_11763,N_12921);
and U16404 (N_16404,N_10703,N_10930);
or U16405 (N_16405,N_11963,N_10914);
nor U16406 (N_16406,N_11745,N_14437);
nand U16407 (N_16407,N_11371,N_13895);
and U16408 (N_16408,N_12078,N_12336);
or U16409 (N_16409,N_11967,N_14173);
and U16410 (N_16410,N_11155,N_11894);
or U16411 (N_16411,N_14079,N_10778);
nand U16412 (N_16412,N_10239,N_12048);
and U16413 (N_16413,N_10402,N_13662);
or U16414 (N_16414,N_12775,N_11019);
or U16415 (N_16415,N_13019,N_11428);
and U16416 (N_16416,N_11726,N_11780);
and U16417 (N_16417,N_11552,N_14239);
nand U16418 (N_16418,N_11689,N_13096);
nand U16419 (N_16419,N_14350,N_11829);
and U16420 (N_16420,N_13379,N_11117);
nor U16421 (N_16421,N_13715,N_13410);
or U16422 (N_16422,N_11477,N_13503);
or U16423 (N_16423,N_13650,N_10869);
nor U16424 (N_16424,N_11533,N_14021);
xor U16425 (N_16425,N_13863,N_12939);
and U16426 (N_16426,N_11791,N_10052);
xor U16427 (N_16427,N_13356,N_14779);
nand U16428 (N_16428,N_14352,N_12846);
and U16429 (N_16429,N_14082,N_11026);
and U16430 (N_16430,N_10983,N_11815);
and U16431 (N_16431,N_14315,N_13808);
xnor U16432 (N_16432,N_10539,N_13156);
or U16433 (N_16433,N_14255,N_12172);
nand U16434 (N_16434,N_10980,N_14418);
nand U16435 (N_16435,N_10903,N_12370);
nand U16436 (N_16436,N_12638,N_10950);
or U16437 (N_16437,N_14168,N_11877);
nand U16438 (N_16438,N_10403,N_13589);
or U16439 (N_16439,N_12605,N_14483);
nor U16440 (N_16440,N_12308,N_12161);
nand U16441 (N_16441,N_14448,N_13075);
nor U16442 (N_16442,N_13240,N_10813);
or U16443 (N_16443,N_11878,N_12953);
nand U16444 (N_16444,N_12903,N_13097);
nor U16445 (N_16445,N_11859,N_12770);
nor U16446 (N_16446,N_13349,N_10193);
nor U16447 (N_16447,N_13659,N_14190);
nor U16448 (N_16448,N_13891,N_14829);
and U16449 (N_16449,N_14131,N_12794);
or U16450 (N_16450,N_12335,N_10751);
nand U16451 (N_16451,N_12338,N_10070);
and U16452 (N_16452,N_11473,N_14787);
xnor U16453 (N_16453,N_13466,N_14495);
nor U16454 (N_16454,N_10265,N_14874);
and U16455 (N_16455,N_10305,N_12808);
xnor U16456 (N_16456,N_14275,N_11572);
or U16457 (N_16457,N_11869,N_10225);
xor U16458 (N_16458,N_11954,N_13310);
nor U16459 (N_16459,N_14313,N_14297);
or U16460 (N_16460,N_14031,N_12052);
nor U16461 (N_16461,N_14451,N_10564);
or U16462 (N_16462,N_13755,N_13498);
and U16463 (N_16463,N_14185,N_10047);
nor U16464 (N_16464,N_14861,N_12728);
nand U16465 (N_16465,N_12360,N_14195);
nand U16466 (N_16466,N_13706,N_14726);
and U16467 (N_16467,N_14960,N_14746);
xnor U16468 (N_16468,N_12831,N_10820);
or U16469 (N_16469,N_14267,N_14288);
or U16470 (N_16470,N_13045,N_10015);
nor U16471 (N_16471,N_13444,N_11074);
or U16472 (N_16472,N_10966,N_13397);
xor U16473 (N_16473,N_13248,N_11063);
nor U16474 (N_16474,N_10346,N_11302);
nand U16475 (N_16475,N_12428,N_11263);
or U16476 (N_16476,N_14373,N_13711);
nor U16477 (N_16477,N_12876,N_10134);
and U16478 (N_16478,N_12933,N_13028);
and U16479 (N_16479,N_14056,N_10588);
or U16480 (N_16480,N_13199,N_14984);
or U16481 (N_16481,N_13219,N_10775);
and U16482 (N_16482,N_11322,N_10468);
nand U16483 (N_16483,N_12958,N_12169);
nand U16484 (N_16484,N_11127,N_13830);
and U16485 (N_16485,N_14343,N_12733);
and U16486 (N_16486,N_10971,N_11253);
nand U16487 (N_16487,N_11030,N_14482);
nor U16488 (N_16488,N_12502,N_10509);
xor U16489 (N_16489,N_13331,N_14141);
xor U16490 (N_16490,N_11716,N_14116);
nor U16491 (N_16491,N_13190,N_13616);
or U16492 (N_16492,N_11590,N_13904);
and U16493 (N_16493,N_10369,N_10835);
or U16494 (N_16494,N_11226,N_11819);
or U16495 (N_16495,N_14274,N_14341);
xor U16496 (N_16496,N_14708,N_12854);
and U16497 (N_16497,N_13871,N_10071);
nand U16498 (N_16498,N_10805,N_10772);
and U16499 (N_16499,N_14590,N_12908);
nand U16500 (N_16500,N_13934,N_13771);
nor U16501 (N_16501,N_14379,N_12965);
nand U16502 (N_16502,N_11362,N_12422);
or U16503 (N_16503,N_12944,N_12517);
or U16504 (N_16504,N_13780,N_13577);
nor U16505 (N_16505,N_11062,N_12458);
and U16506 (N_16506,N_10826,N_14805);
nand U16507 (N_16507,N_13407,N_14409);
nor U16508 (N_16508,N_11579,N_14931);
nand U16509 (N_16509,N_13983,N_13059);
or U16510 (N_16510,N_14772,N_14114);
and U16511 (N_16511,N_10083,N_13269);
nand U16512 (N_16512,N_11501,N_10464);
nor U16513 (N_16513,N_12163,N_12372);
xor U16514 (N_16514,N_12182,N_12234);
nor U16515 (N_16515,N_10744,N_14533);
nor U16516 (N_16516,N_10194,N_12811);
and U16517 (N_16517,N_12838,N_14996);
nor U16518 (N_16518,N_11731,N_10197);
or U16519 (N_16519,N_13022,N_12159);
nor U16520 (N_16520,N_12389,N_13432);
nor U16521 (N_16521,N_10081,N_14403);
nor U16522 (N_16522,N_12361,N_12282);
nand U16523 (N_16523,N_11279,N_12937);
or U16524 (N_16524,N_12799,N_12031);
and U16525 (N_16525,N_13312,N_10740);
or U16526 (N_16526,N_11973,N_13117);
xor U16527 (N_16527,N_13865,N_14303);
or U16528 (N_16528,N_12021,N_13818);
or U16529 (N_16529,N_10889,N_14608);
nand U16530 (N_16530,N_14424,N_13579);
xnor U16531 (N_16531,N_14422,N_12572);
or U16532 (N_16532,N_10102,N_11046);
nand U16533 (N_16533,N_10716,N_14558);
or U16534 (N_16534,N_10395,N_10611);
nor U16535 (N_16535,N_13993,N_14460);
and U16536 (N_16536,N_10876,N_12210);
nor U16537 (N_16537,N_12753,N_13262);
nand U16538 (N_16538,N_10513,N_12478);
and U16539 (N_16539,N_11409,N_12618);
xor U16540 (N_16540,N_13590,N_11751);
xor U16541 (N_16541,N_12251,N_14979);
or U16542 (N_16542,N_14047,N_14491);
nor U16543 (N_16543,N_10939,N_10407);
or U16544 (N_16544,N_14111,N_13040);
or U16545 (N_16545,N_10801,N_10268);
nor U16546 (N_16546,N_14330,N_14066);
and U16547 (N_16547,N_14653,N_12801);
or U16548 (N_16548,N_14283,N_13078);
nor U16549 (N_16549,N_12417,N_10958);
nand U16550 (N_16550,N_11896,N_10840);
and U16551 (N_16551,N_10277,N_14440);
or U16552 (N_16552,N_10532,N_13556);
nand U16553 (N_16553,N_14780,N_10700);
nor U16554 (N_16554,N_12065,N_12962);
nor U16555 (N_16555,N_14553,N_10273);
and U16556 (N_16556,N_13942,N_13747);
and U16557 (N_16557,N_12230,N_12374);
and U16558 (N_16558,N_12097,N_13483);
nand U16559 (N_16559,N_10803,N_12488);
nand U16560 (N_16560,N_11770,N_10828);
or U16561 (N_16561,N_12337,N_11757);
nand U16562 (N_16562,N_12557,N_10075);
nor U16563 (N_16563,N_11060,N_13907);
nand U16564 (N_16564,N_10333,N_12276);
xnor U16565 (N_16565,N_13184,N_13545);
or U16566 (N_16566,N_10180,N_14147);
nand U16567 (N_16567,N_13411,N_10247);
or U16568 (N_16568,N_12516,N_14522);
or U16569 (N_16569,N_11152,N_11154);
nor U16570 (N_16570,N_10895,N_14014);
or U16571 (N_16571,N_10994,N_13727);
nor U16572 (N_16572,N_13597,N_10808);
and U16573 (N_16573,N_13887,N_14389);
and U16574 (N_16574,N_10777,N_14722);
nor U16575 (N_16575,N_14322,N_11312);
xor U16576 (N_16576,N_12874,N_14081);
nor U16577 (N_16577,N_10585,N_11008);
nand U16578 (N_16578,N_12563,N_10296);
or U16579 (N_16579,N_10045,N_14924);
nand U16580 (N_16580,N_12936,N_11078);
nand U16581 (N_16581,N_12649,N_14070);
and U16582 (N_16582,N_12570,N_10439);
xor U16583 (N_16583,N_14126,N_12185);
or U16584 (N_16584,N_12363,N_14426);
xnor U16585 (N_16585,N_12783,N_13772);
xor U16586 (N_16586,N_14657,N_11332);
and U16587 (N_16587,N_14153,N_14334);
or U16588 (N_16588,N_13140,N_14238);
and U16589 (N_16589,N_10864,N_10046);
nand U16590 (N_16590,N_14549,N_14490);
and U16591 (N_16591,N_10272,N_11887);
and U16592 (N_16592,N_14397,N_13274);
or U16593 (N_16593,N_14258,N_13247);
and U16594 (N_16594,N_11951,N_13638);
nor U16595 (N_16595,N_10621,N_11842);
or U16596 (N_16596,N_12314,N_14863);
nand U16597 (N_16597,N_10900,N_10637);
or U16598 (N_16598,N_14036,N_13552);
or U16599 (N_16599,N_14761,N_13272);
and U16600 (N_16600,N_10145,N_13364);
and U16601 (N_16601,N_14650,N_13627);
xor U16602 (N_16602,N_11056,N_12475);
xnor U16603 (N_16603,N_12918,N_12476);
nand U16604 (N_16604,N_12614,N_10854);
nor U16605 (N_16605,N_13748,N_14050);
and U16606 (N_16606,N_14603,N_12420);
nor U16607 (N_16607,N_13077,N_14291);
or U16608 (N_16608,N_12576,N_11735);
or U16609 (N_16609,N_11066,N_11638);
nand U16610 (N_16610,N_12619,N_13099);
and U16611 (N_16611,N_13165,N_12019);
nand U16612 (N_16612,N_10475,N_13908);
and U16613 (N_16613,N_14391,N_13693);
nor U16614 (N_16614,N_12271,N_14020);
nand U16615 (N_16615,N_11416,N_11405);
or U16616 (N_16616,N_11160,N_13520);
nor U16617 (N_16617,N_10697,N_14850);
or U16618 (N_16618,N_11576,N_13505);
or U16619 (N_16619,N_14489,N_12455);
and U16620 (N_16620,N_11940,N_14690);
or U16621 (N_16621,N_14121,N_13258);
xnor U16622 (N_16622,N_11806,N_12541);
xor U16623 (N_16623,N_13424,N_11118);
nor U16624 (N_16624,N_10024,N_14891);
and U16625 (N_16625,N_10689,N_14492);
nand U16626 (N_16626,N_13157,N_14841);
nand U16627 (N_16627,N_12940,N_11334);
nor U16628 (N_16628,N_10300,N_13723);
or U16629 (N_16629,N_14561,N_12992);
or U16630 (N_16630,N_14655,N_12879);
nor U16631 (N_16631,N_10478,N_12171);
nor U16632 (N_16632,N_12856,N_10659);
nand U16633 (N_16633,N_13121,N_12735);
nor U16634 (N_16634,N_13396,N_11077);
nand U16635 (N_16635,N_12024,N_14146);
or U16636 (N_16636,N_10032,N_12367);
xor U16637 (N_16637,N_11045,N_12786);
or U16638 (N_16638,N_13631,N_13921);
and U16639 (N_16639,N_10480,N_11156);
nor U16640 (N_16640,N_11808,N_10212);
and U16641 (N_16641,N_13278,N_11460);
and U16642 (N_16642,N_14552,N_11613);
xnor U16643 (N_16643,N_12724,N_13968);
and U16644 (N_16644,N_13334,N_10506);
nor U16645 (N_16645,N_10893,N_14563);
nor U16646 (N_16646,N_10546,N_12396);
or U16647 (N_16647,N_14192,N_12449);
nor U16648 (N_16648,N_13905,N_13016);
nor U16649 (N_16649,N_13515,N_11270);
xor U16650 (N_16650,N_14732,N_10144);
or U16651 (N_16651,N_11215,N_14697);
nand U16652 (N_16652,N_13793,N_10020);
and U16653 (N_16653,N_14068,N_14310);
or U16654 (N_16654,N_13775,N_13311);
nor U16655 (N_16655,N_14228,N_14329);
or U16656 (N_16656,N_14191,N_13791);
nor U16657 (N_16657,N_10393,N_13703);
or U16658 (N_16658,N_12982,N_14246);
nand U16659 (N_16659,N_10537,N_13486);
nor U16660 (N_16660,N_11925,N_10132);
and U16661 (N_16661,N_10839,N_12678);
or U16662 (N_16662,N_14901,N_13697);
or U16663 (N_16663,N_11663,N_11010);
and U16664 (N_16664,N_10878,N_13811);
nand U16665 (N_16665,N_10599,N_13828);
nor U16666 (N_16666,N_14080,N_11958);
and U16667 (N_16667,N_11036,N_10053);
nor U16668 (N_16668,N_10555,N_12575);
nand U16669 (N_16669,N_11465,N_12375);
or U16670 (N_16670,N_12910,N_14637);
and U16671 (N_16671,N_14078,N_12424);
nand U16672 (N_16672,N_12889,N_11095);
and U16673 (N_16673,N_10553,N_13350);
nand U16674 (N_16674,N_12507,N_11586);
nand U16675 (N_16675,N_11670,N_12520);
xor U16676 (N_16676,N_11914,N_12525);
xnor U16677 (N_16677,N_10486,N_14353);
or U16678 (N_16678,N_11553,N_10687);
nor U16679 (N_16679,N_11955,N_14077);
or U16680 (N_16680,N_11610,N_11212);
and U16681 (N_16681,N_14757,N_12385);
xnor U16682 (N_16682,N_13036,N_12289);
or U16683 (N_16683,N_10904,N_10467);
and U16684 (N_16684,N_13719,N_10074);
and U16685 (N_16685,N_10195,N_10130);
or U16686 (N_16686,N_13649,N_13845);
xor U16687 (N_16687,N_12913,N_14167);
or U16688 (N_16688,N_11804,N_12952);
or U16689 (N_16689,N_11837,N_11415);
nand U16690 (N_16690,N_13083,N_12386);
or U16691 (N_16691,N_14256,N_10785);
nand U16692 (N_16692,N_14396,N_14839);
nand U16693 (N_16693,N_10638,N_10522);
nand U16694 (N_16694,N_11216,N_14276);
nand U16695 (N_16695,N_11028,N_14634);
nor U16696 (N_16696,N_10394,N_10284);
and U16697 (N_16697,N_14332,N_14299);
or U16698 (N_16698,N_14895,N_10227);
nor U16699 (N_16699,N_10005,N_13271);
nand U16700 (N_16700,N_11086,N_12369);
and U16701 (N_16701,N_11262,N_14922);
xor U16702 (N_16702,N_14876,N_14316);
nand U16703 (N_16703,N_12751,N_13139);
nand U16704 (N_16704,N_11255,N_10260);
or U16705 (N_16705,N_11234,N_11534);
nand U16706 (N_16706,N_11356,N_13929);
nand U16707 (N_16707,N_12373,N_12317);
nor U16708 (N_16708,N_11232,N_13792);
xnor U16709 (N_16709,N_11743,N_10937);
nor U16710 (N_16710,N_14704,N_10945);
nor U16711 (N_16711,N_10330,N_11467);
and U16712 (N_16712,N_11598,N_14674);
nor U16713 (N_16713,N_10126,N_13009);
or U16714 (N_16714,N_12597,N_13799);
or U16715 (N_16715,N_12693,N_10622);
xnor U16716 (N_16716,N_12816,N_10556);
nand U16717 (N_16717,N_12406,N_12010);
nand U16718 (N_16718,N_11569,N_14382);
or U16719 (N_16719,N_12987,N_13257);
nand U16720 (N_16720,N_14802,N_12268);
nand U16721 (N_16721,N_13276,N_12922);
nand U16722 (N_16722,N_11016,N_10297);
and U16723 (N_16723,N_11516,N_13668);
and U16724 (N_16724,N_14415,N_10664);
and U16725 (N_16725,N_12123,N_12881);
and U16726 (N_16726,N_13962,N_12404);
nand U16727 (N_16727,N_13653,N_12719);
or U16728 (N_16728,N_11197,N_13768);
and U16729 (N_16729,N_10503,N_12901);
or U16730 (N_16730,N_12080,N_10635);
nor U16731 (N_16731,N_12368,N_10639);
and U16732 (N_16732,N_11469,N_14797);
xor U16733 (N_16733,N_11299,N_13069);
nand U16734 (N_16734,N_11208,N_11650);
xnor U16735 (N_16735,N_10218,N_14914);
nand U16736 (N_16736,N_12397,N_14892);
xor U16737 (N_16737,N_14107,N_14557);
or U16738 (N_16738,N_14417,N_11076);
and U16739 (N_16739,N_11458,N_10884);
nor U16740 (N_16740,N_11500,N_13923);
nand U16741 (N_16741,N_10668,N_13758);
nor U16742 (N_16742,N_14946,N_13021);
and U16743 (N_16743,N_11266,N_13390);
or U16744 (N_16744,N_11339,N_11728);
and U16745 (N_16745,N_12379,N_12340);
nand U16746 (N_16746,N_10222,N_11389);
or U16747 (N_16747,N_14950,N_11350);
nand U16748 (N_16748,N_10745,N_11330);
nor U16749 (N_16749,N_13323,N_14691);
nor U16750 (N_16750,N_12830,N_12621);
nand U16751 (N_16751,N_10054,N_12821);
or U16752 (N_16752,N_11069,N_14623);
nand U16753 (N_16753,N_14069,N_10862);
and U16754 (N_16754,N_14404,N_10948);
nor U16755 (N_16755,N_10941,N_13290);
nor U16756 (N_16756,N_13534,N_10684);
and U16757 (N_16757,N_11229,N_11065);
xor U16758 (N_16758,N_10767,N_13933);
or U16759 (N_16759,N_14806,N_14921);
nand U16760 (N_16760,N_14179,N_10334);
nand U16761 (N_16761,N_11442,N_12249);
nand U16762 (N_16762,N_13803,N_12301);
nand U16763 (N_16763,N_11828,N_11644);
and U16764 (N_16764,N_11906,N_13979);
and U16765 (N_16765,N_11630,N_12032);
nor U16766 (N_16766,N_10843,N_14219);
nor U16767 (N_16767,N_14266,N_14501);
nand U16768 (N_16768,N_12056,N_13990);
xnor U16769 (N_16769,N_14122,N_14968);
nor U16770 (N_16770,N_11691,N_11771);
and U16771 (N_16771,N_13821,N_10806);
xnor U16772 (N_16772,N_14249,N_14385);
nand U16773 (N_16773,N_12515,N_12044);
and U16774 (N_16774,N_14211,N_12822);
and U16775 (N_16775,N_14510,N_11707);
or U16776 (N_16776,N_14978,N_11643);
or U16777 (N_16777,N_14715,N_12757);
or U16778 (N_16778,N_12036,N_10067);
nand U16779 (N_16779,N_13436,N_14254);
and U16780 (N_16780,N_12144,N_11810);
nor U16781 (N_16781,N_14862,N_10404);
xnor U16782 (N_16782,N_13125,N_12437);
nand U16783 (N_16783,N_11669,N_10929);
or U16784 (N_16784,N_11213,N_14101);
and U16785 (N_16785,N_14581,N_10845);
and U16786 (N_16786,N_10511,N_10598);
and U16787 (N_16787,N_11952,N_10535);
nor U16788 (N_16788,N_11890,N_11224);
nor U16789 (N_16789,N_12007,N_10470);
nor U16790 (N_16790,N_10127,N_13185);
and U16791 (N_16791,N_11589,N_11000);
or U16792 (N_16792,N_10385,N_10701);
or U16793 (N_16793,N_14531,N_12915);
nand U16794 (N_16794,N_14699,N_14083);
or U16795 (N_16795,N_12916,N_11106);
nor U16796 (N_16796,N_10485,N_11227);
xor U16797 (N_16797,N_14347,N_10192);
nor U16798 (N_16798,N_13295,N_11620);
nand U16799 (N_16799,N_14368,N_13952);
nor U16800 (N_16800,N_13149,N_10476);
nor U16801 (N_16801,N_13129,N_10651);
or U16802 (N_16802,N_13800,N_11807);
or U16803 (N_16803,N_12644,N_10517);
and U16804 (N_16804,N_12483,N_10149);
nand U16805 (N_16805,N_12099,N_12365);
nand U16806 (N_16806,N_13692,N_13763);
nand U16807 (N_16807,N_12586,N_10663);
nor U16808 (N_16808,N_14013,N_10184);
nor U16809 (N_16809,N_12744,N_10257);
or U16810 (N_16810,N_11830,N_10769);
nand U16811 (N_16811,N_14803,N_13232);
and U16812 (N_16812,N_11674,N_11634);
nand U16813 (N_16813,N_14897,N_11897);
and U16814 (N_16814,N_12683,N_14351);
nand U16815 (N_16815,N_11179,N_13623);
and U16816 (N_16816,N_11882,N_14420);
and U16817 (N_16817,N_14194,N_13188);
nor U16818 (N_16818,N_10804,N_12076);
or U16819 (N_16819,N_14970,N_14625);
nand U16820 (N_16820,N_14645,N_14307);
nor U16821 (N_16821,N_13673,N_10458);
nor U16822 (N_16822,N_12991,N_14294);
xor U16823 (N_16823,N_10463,N_10738);
nor U16824 (N_16824,N_11314,N_14425);
and U16825 (N_16825,N_14251,N_11924);
and U16826 (N_16826,N_12699,N_11223);
xnor U16827 (N_16827,N_10561,N_11185);
and U16828 (N_16828,N_11241,N_13722);
nor U16829 (N_16829,N_13987,N_14443);
nand U16830 (N_16830,N_12859,N_12180);
nand U16831 (N_16831,N_12134,N_14257);
and U16832 (N_16832,N_13624,N_14143);
and U16833 (N_16833,N_11685,N_14289);
or U16834 (N_16834,N_13442,N_10606);
nor U16835 (N_16835,N_11315,N_11880);
or U16836 (N_16836,N_11320,N_14747);
and U16837 (N_16837,N_12339,N_11441);
or U16838 (N_16838,N_12304,N_12980);
or U16839 (N_16839,N_10170,N_13004);
nand U16840 (N_16840,N_13652,N_10112);
and U16841 (N_16841,N_13819,N_11713);
xnor U16842 (N_16842,N_13026,N_14810);
and U16843 (N_16843,N_14226,N_14142);
or U16844 (N_16844,N_12542,N_11570);
nor U16845 (N_16845,N_10030,N_11092);
nand U16846 (N_16846,N_11969,N_11931);
nand U16847 (N_16847,N_13740,N_12989);
or U16848 (N_16848,N_14099,N_11573);
nor U16849 (N_16849,N_14896,N_11125);
xor U16850 (N_16850,N_11577,N_10338);
nand U16851 (N_16851,N_10416,N_14682);
or U16852 (N_16852,N_13302,N_12812);
xnor U16853 (N_16853,N_12878,N_10274);
or U16854 (N_16854,N_11593,N_14336);
xnor U16855 (N_16855,N_12131,N_11448);
or U16856 (N_16856,N_14893,N_12395);
and U16857 (N_16857,N_14186,N_14375);
and U16858 (N_16858,N_13524,N_13384);
xnor U16859 (N_16859,N_14210,N_10425);
nand U16860 (N_16860,N_14791,N_14677);
and U16861 (N_16861,N_12852,N_14641);
nand U16862 (N_16862,N_13168,N_11513);
or U16863 (N_16863,N_13175,N_12713);
nor U16864 (N_16864,N_14306,N_12279);
nor U16865 (N_16865,N_11492,N_11947);
nor U16866 (N_16866,N_13639,N_14916);
or U16867 (N_16867,N_12211,N_11564);
nand U16868 (N_16868,N_14534,N_13482);
nor U16869 (N_16869,N_10730,N_12587);
nor U16870 (N_16870,N_14886,N_11085);
nand U16871 (N_16871,N_14955,N_11591);
and U16872 (N_16872,N_14112,N_12964);
nand U16873 (N_16873,N_10104,N_10153);
nand U16874 (N_16874,N_13644,N_10337);
nand U16875 (N_16875,N_12443,N_12223);
nand U16876 (N_16876,N_10583,N_14012);
or U16877 (N_16877,N_12677,N_13689);
or U16878 (N_16878,N_12810,N_13479);
or U16879 (N_16879,N_11844,N_11683);
and U16880 (N_16880,N_11054,N_11194);
or U16881 (N_16881,N_10091,N_14366);
or U16882 (N_16882,N_10187,N_12244);
nor U16883 (N_16883,N_10834,N_13313);
nor U16884 (N_16884,N_10964,N_10927);
and U16885 (N_16885,N_14429,N_14480);
nor U16886 (N_16886,N_11520,N_12068);
nor U16887 (N_16887,N_10164,N_13198);
xor U16888 (N_16888,N_10770,N_11031);
nand U16889 (N_16889,N_13538,N_11436);
nor U16890 (N_16890,N_13737,N_11099);
nor U16891 (N_16891,N_13559,N_13823);
nor U16892 (N_16892,N_14834,N_13507);
and U16893 (N_16893,N_11494,N_10759);
nand U16894 (N_16894,N_10157,N_13721);
and U16895 (N_16895,N_12632,N_12218);
and U16896 (N_16896,N_14400,N_11606);
or U16897 (N_16897,N_14325,N_10119);
nor U16898 (N_16898,N_12748,N_11301);
xnor U16899 (N_16899,N_12626,N_13066);
and U16900 (N_16900,N_14285,N_13270);
and U16901 (N_16901,N_12524,N_13733);
or U16902 (N_16902,N_10976,N_12841);
xor U16903 (N_16903,N_11861,N_12116);
nand U16904 (N_16904,N_13032,N_14406);
or U16905 (N_16905,N_11996,N_12026);
nand U16906 (N_16906,N_11701,N_10720);
or U16907 (N_16907,N_12427,N_10771);
nand U16908 (N_16908,N_12139,N_12098);
nor U16909 (N_16909,N_12000,N_13502);
and U16910 (N_16910,N_14364,N_14280);
or U16911 (N_16911,N_11310,N_11384);
and U16912 (N_16912,N_14204,N_13593);
nand U16913 (N_16913,N_10474,N_10735);
nand U16914 (N_16914,N_13093,N_11736);
nand U16915 (N_16915,N_11809,N_14760);
xor U16916 (N_16916,N_14940,N_14431);
nand U16917 (N_16917,N_13700,N_12492);
xnor U16918 (N_16918,N_12629,N_10737);
nand U16919 (N_16919,N_13838,N_13128);
nand U16920 (N_16920,N_10135,N_13070);
and U16921 (N_16921,N_13253,N_12665);
nand U16922 (N_16922,N_10515,N_11184);
nor U16923 (N_16923,N_11411,N_12072);
nor U16924 (N_16924,N_14293,N_10105);
nand U16925 (N_16925,N_12931,N_14569);
xnor U16926 (N_16926,N_12058,N_11588);
xnor U16927 (N_16927,N_12143,N_14067);
nand U16928 (N_16928,N_13560,N_12017);
nor U16929 (N_16929,N_12258,N_12124);
and U16930 (N_16930,N_14538,N_11979);
and U16931 (N_16931,N_13453,N_14975);
nand U16932 (N_16932,N_12380,N_14544);
and U16933 (N_16933,N_14523,N_12897);
nand U16934 (N_16934,N_13731,N_13495);
nor U16935 (N_16935,N_10596,N_10784);
xnor U16936 (N_16936,N_10560,N_14890);
nor U16937 (N_16937,N_10484,N_10870);
nand U16938 (N_16938,N_13971,N_13459);
or U16939 (N_16939,N_12687,N_13403);
and U16940 (N_16940,N_11474,N_14816);
nand U16941 (N_16941,N_11609,N_10836);
and U16942 (N_16942,N_10489,N_13619);
and U16943 (N_16943,N_11651,N_11343);
or U16944 (N_16944,N_12229,N_10946);
nor U16945 (N_16945,N_14176,N_11594);
nand U16946 (N_16946,N_11385,N_12554);
nor U16947 (N_16947,N_11201,N_13900);
and U16948 (N_16948,N_12700,N_11631);
nand U16949 (N_16949,N_13314,N_10240);
nand U16950 (N_16950,N_10449,N_11575);
nor U16951 (N_16951,N_11891,N_14300);
or U16952 (N_16952,N_11884,N_10943);
nor U16953 (N_16953,N_10400,N_13003);
nand U16954 (N_16954,N_12059,N_12313);
nor U16955 (N_16955,N_13374,N_13154);
nor U16956 (N_16956,N_14848,N_12776);
or U16957 (N_16957,N_13858,N_12993);
nor U16958 (N_16958,N_11987,N_14822);
nor U16959 (N_16959,N_10432,N_12489);
and U16960 (N_16960,N_14694,N_13717);
or U16961 (N_16961,N_13051,N_11425);
and U16962 (N_16962,N_14446,N_11563);
nand U16963 (N_16963,N_11693,N_11454);
nor U16964 (N_16964,N_11856,N_11883);
or U16965 (N_16965,N_12578,N_11676);
nor U16966 (N_16966,N_13293,N_11621);
nor U16967 (N_16967,N_14593,N_11139);
and U16968 (N_16968,N_14089,N_12531);
nor U16969 (N_16969,N_13794,N_13487);
nor U16970 (N_16970,N_10154,N_14038);
and U16971 (N_16971,N_14516,N_11567);
and U16972 (N_16972,N_14466,N_13519);
xnor U16973 (N_16973,N_12646,N_10066);
nand U16974 (N_16974,N_13308,N_11144);
nand U16975 (N_16975,N_13604,N_14027);
and U16976 (N_16976,N_10389,N_12731);
nand U16977 (N_16977,N_10205,N_14182);
nand U16978 (N_16978,N_10413,N_14253);
nand U16979 (N_16979,N_13704,N_11449);
and U16980 (N_16980,N_11237,N_12112);
or U16981 (N_16981,N_10003,N_12899);
nand U16982 (N_16982,N_12069,N_14832);
or U16983 (N_16983,N_10287,N_14512);
nand U16984 (N_16984,N_13698,N_13457);
nand U16985 (N_16985,N_10502,N_13193);
or U16986 (N_16986,N_13656,N_12326);
or U16987 (N_16987,N_13489,N_14630);
and U16988 (N_16988,N_12062,N_12960);
nor U16989 (N_16989,N_10065,N_10563);
xnor U16990 (N_16990,N_12034,N_11962);
or U16991 (N_16991,N_13033,N_14915);
nand U16992 (N_16992,N_10251,N_13200);
nand U16993 (N_16993,N_10923,N_13330);
nand U16994 (N_16994,N_14987,N_14374);
or U16995 (N_16995,N_11463,N_10493);
nand U16996 (N_16996,N_12245,N_12710);
nand U16997 (N_16997,N_11867,N_11536);
or U16998 (N_16998,N_11276,N_11814);
nand U16999 (N_16999,N_12356,N_10901);
xor U17000 (N_17000,N_11121,N_10996);
or U17001 (N_17001,N_12236,N_12239);
and U17002 (N_17002,N_13195,N_13306);
or U17003 (N_17003,N_12459,N_10179);
and U17004 (N_17004,N_14991,N_13642);
nor U17005 (N_17005,N_12486,N_12855);
nor U17006 (N_17006,N_14467,N_14133);
nor U17007 (N_17007,N_12186,N_13254);
or U17008 (N_17008,N_11447,N_13839);
and U17009 (N_17009,N_13326,N_12499);
or U17010 (N_17010,N_14535,N_10243);
nand U17011 (N_17011,N_13178,N_11547);
xnor U17012 (N_17012,N_11417,N_11182);
or U17013 (N_17013,N_11530,N_14132);
and U17014 (N_17014,N_13796,N_14110);
and U17015 (N_17015,N_12637,N_11889);
or U17016 (N_17016,N_13759,N_11918);
and U17017 (N_17017,N_14109,N_11910);
nand U17018 (N_17018,N_14444,N_11665);
nand U17019 (N_17019,N_13112,N_14776);
or U17020 (N_17020,N_13965,N_11177);
xnor U17021 (N_17021,N_12257,N_14687);
and U17022 (N_17022,N_14134,N_10318);
nand U17023 (N_17023,N_14577,N_14881);
nor U17024 (N_17024,N_10998,N_12955);
nand U17025 (N_17025,N_12242,N_11866);
nor U17026 (N_17026,N_12717,N_14428);
nand U17027 (N_17027,N_14042,N_14621);
nand U17028 (N_17028,N_13708,N_12184);
or U17029 (N_17029,N_11304,N_13409);
and U17030 (N_17030,N_10885,N_14983);
xnor U17031 (N_17031,N_12508,N_13126);
nor U17032 (N_17032,N_14756,N_11218);
and U17033 (N_17033,N_12550,N_10999);
nor U17034 (N_17034,N_11360,N_12926);
xnor U17035 (N_17035,N_12673,N_10514);
nor U17036 (N_17036,N_14302,N_12670);
nor U17037 (N_17037,N_12630,N_10899);
xor U17038 (N_17038,N_13967,N_14319);
or U17039 (N_17039,N_10525,N_12114);
nor U17040 (N_17040,N_10023,N_11506);
nand U17041 (N_17041,N_13395,N_10816);
nand U17042 (N_17042,N_12259,N_13798);
nand U17043 (N_17043,N_10223,N_13203);
and U17044 (N_17044,N_11040,N_13101);
nand U17045 (N_17045,N_13164,N_13543);
nand U17046 (N_17046,N_13336,N_12784);
and U17047 (N_17047,N_14500,N_12298);
or U17048 (N_17048,N_12457,N_14064);
or U17049 (N_17049,N_10725,N_12546);
nor U17050 (N_17050,N_10238,N_11561);
or U17051 (N_17051,N_11146,N_13335);
or U17052 (N_17052,N_12466,N_13980);
nor U17053 (N_17053,N_13371,N_11580);
or U17054 (N_17054,N_14230,N_10320);
nor U17055 (N_17055,N_12592,N_13309);
nor U17056 (N_17056,N_13049,N_13095);
nand U17057 (N_17057,N_13506,N_14718);
and U17058 (N_17058,N_13551,N_12628);
nand U17059 (N_17059,N_13647,N_11392);
or U17060 (N_17060,N_13265,N_14597);
or U17061 (N_17061,N_12445,N_12664);
or U17062 (N_17062,N_13814,N_13346);
or U17063 (N_17063,N_12005,N_14969);
and U17064 (N_17064,N_10544,N_13817);
or U17065 (N_17065,N_11985,N_13613);
nor U17066 (N_17066,N_12707,N_13756);
and U17067 (N_17067,N_13166,N_14198);
xor U17068 (N_17068,N_13425,N_12329);
or U17069 (N_17069,N_14091,N_14156);
nor U17070 (N_17070,N_10586,N_11222);
nand U17071 (N_17071,N_12221,N_12613);
or U17072 (N_17072,N_13446,N_12555);
and U17073 (N_17073,N_10255,N_14799);
and U17074 (N_17074,N_10554,N_12877);
and U17075 (N_17075,N_14617,N_10949);
nand U17076 (N_17076,N_13640,N_12704);
xnor U17077 (N_17077,N_12552,N_13504);
nand U17078 (N_17078,N_11811,N_11364);
or U17079 (N_17079,N_11608,N_14227);
nor U17080 (N_17080,N_10422,N_13170);
nor U17081 (N_17081,N_11523,N_10600);
or U17082 (N_17082,N_11905,N_13292);
nor U17083 (N_17083,N_13761,N_10510);
and U17084 (N_17084,N_14601,N_14606);
nand U17085 (N_17085,N_12167,N_11012);
nand U17086 (N_17086,N_11976,N_12813);
nor U17087 (N_17087,N_10281,N_12805);
nor U17088 (N_17088,N_13455,N_10376);
or U17089 (N_17089,N_14044,N_11486);
xor U17090 (N_17090,N_10217,N_12772);
or U17091 (N_17091,N_10266,N_14314);
nand U17092 (N_17092,N_14035,N_14958);
and U17093 (N_17093,N_12442,N_11919);
or U17094 (N_17094,N_14106,N_10533);
or U17095 (N_17095,N_13588,N_12074);
and U17096 (N_17096,N_12850,N_10171);
xor U17097 (N_17097,N_12737,N_12446);
nor U17098 (N_17098,N_10290,N_13100);
or U17099 (N_17099,N_10106,N_12909);
or U17100 (N_17100,N_10615,N_10150);
nor U17101 (N_17101,N_12750,N_10524);
nor U17102 (N_17102,N_14605,N_13023);
nand U17103 (N_17103,N_10944,N_11741);
or U17104 (N_17104,N_11290,N_13191);
or U17105 (N_17105,N_14244,N_14181);
nor U17106 (N_17106,N_12599,N_12870);
nor U17107 (N_17107,N_13451,N_13517);
or U17108 (N_17108,N_14003,N_13789);
and U17109 (N_17109,N_13912,N_12658);
and U17110 (N_17110,N_13458,N_12362);
and U17111 (N_17111,N_12703,N_10447);
and U17112 (N_17112,N_12316,N_10009);
or U17113 (N_17113,N_11087,N_10169);
nor U17114 (N_17114,N_12580,N_13054);
nand U17115 (N_17115,N_10175,N_13633);
and U17116 (N_17116,N_12252,N_11307);
and U17117 (N_17117,N_13103,N_12002);
xor U17118 (N_17118,N_13995,N_10166);
or U17119 (N_17119,N_12387,N_12905);
nand U17120 (N_17120,N_14359,N_13084);
and U17121 (N_17121,N_11507,N_12566);
nor U17122 (N_17122,N_12164,N_10176);
nor U17123 (N_17123,N_13790,N_13533);
nand U17124 (N_17124,N_10690,N_12094);
and U17125 (N_17125,N_14737,N_11147);
and U17126 (N_17126,N_14835,N_14938);
and U17127 (N_17127,N_12880,N_11504);
nor U17128 (N_17128,N_14380,N_10232);
nand U17129 (N_17129,N_11888,N_12121);
nor U17130 (N_17130,N_10587,N_11818);
nor U17131 (N_17131,N_14702,N_11351);
nand U17132 (N_17132,N_13567,N_11984);
and U17133 (N_17133,N_12456,N_14024);
nor U17134 (N_17134,N_14614,N_14723);
and U17135 (N_17135,N_12299,N_13113);
or U17136 (N_17136,N_12444,N_12545);
nor U17137 (N_17137,N_10672,N_12105);
and U17138 (N_17138,N_13527,N_12303);
nand U17139 (N_17139,N_12660,N_13218);
or U17140 (N_17140,N_12300,N_11115);
and U17141 (N_17141,N_10713,N_13760);
and U17142 (N_17142,N_14550,N_11059);
or U17143 (N_17143,N_12706,N_13160);
or U17144 (N_17144,N_14661,N_10968);
or U17145 (N_17145,N_12745,N_10314);
xor U17146 (N_17146,N_12593,N_10262);
nand U17147 (N_17147,N_13416,N_13375);
nor U17148 (N_17148,N_12498,N_13382);
and U17149 (N_17149,N_11096,N_13249);
or U17150 (N_17150,N_10292,N_12435);
nand U17151 (N_17151,N_11977,N_10347);
and U17152 (N_17152,N_12760,N_12349);
nor U17153 (N_17153,N_14771,N_10573);
nor U17154 (N_17154,N_11539,N_11221);
nand U17155 (N_17155,N_10269,N_14016);
nand U17156 (N_17156,N_13784,N_11195);
nand U17157 (N_17157,N_11116,N_12511);
nand U17158 (N_17158,N_12033,N_14618);
and U17159 (N_17159,N_12934,N_10947);
nand U17160 (N_17160,N_13745,N_13746);
or U17161 (N_17161,N_10605,N_14525);
xnor U17162 (N_17162,N_12383,N_13143);
or U17163 (N_17163,N_10038,N_12109);
and U17164 (N_17164,N_13183,N_10552);
and U17165 (N_17165,N_12160,N_10412);
nor U17166 (N_17166,N_13988,N_13478);
or U17167 (N_17167,N_14783,N_11965);
and U17168 (N_17168,N_14689,N_14774);
and U17169 (N_17169,N_12928,N_14748);
nand U17170 (N_17170,N_13542,N_10477);
and U17171 (N_17171,N_10158,N_13399);
nor U17172 (N_17172,N_14671,N_12777);
nor U17173 (N_17173,N_10498,N_11484);
nor U17174 (N_17174,N_11132,N_13576);
or U17175 (N_17175,N_14877,N_12887);
xor U17176 (N_17176,N_14346,N_14465);
or U17177 (N_17177,N_12530,N_14163);
and U17178 (N_17178,N_13868,N_14965);
nor U17179 (N_17179,N_14113,N_14855);
or U17180 (N_17180,N_11696,N_14470);
and U17181 (N_17181,N_13951,N_11039);
or U17182 (N_17182,N_12574,N_12732);
nand U17183 (N_17183,N_13288,N_11747);
nor U17184 (N_17184,N_14221,N_11950);
or U17185 (N_17185,N_14919,N_10613);
nor U17186 (N_17186,N_13043,N_11503);
or U17187 (N_17187,N_11081,N_11341);
nand U17188 (N_17188,N_13224,N_12529);
or U17189 (N_17189,N_10773,N_10391);
or U17190 (N_17190,N_12969,N_12333);
nor U17191 (N_17191,N_12740,N_10420);
and U17192 (N_17192,N_12521,N_12414);
nor U17193 (N_17193,N_12896,N_10678);
nor U17194 (N_17194,N_14543,N_14852);
or U17195 (N_17195,N_12564,N_10584);
nor U17196 (N_17196,N_14740,N_11703);
or U17197 (N_17197,N_10029,N_14311);
or U17198 (N_17198,N_13244,N_12815);
nor U17199 (N_17199,N_12824,N_14247);
or U17200 (N_17200,N_12620,N_12872);
xor U17201 (N_17201,N_11230,N_12468);
nand U17202 (N_17202,N_10161,N_12589);
or U17203 (N_17203,N_12825,N_10094);
nor U17204 (N_17204,N_12177,N_12286);
nor U17205 (N_17205,N_12722,N_11082);
or U17206 (N_17206,N_13874,N_14844);
nor U17207 (N_17207,N_10705,N_13263);
nor U17208 (N_17208,N_14717,N_12125);
nand U17209 (N_17209,N_10383,N_14019);
nand U17210 (N_17210,N_12173,N_11020);
nand U17211 (N_17211,N_12679,N_14785);
nor U17212 (N_17212,N_12835,N_13328);
and U17213 (N_17213,N_10349,N_11926);
or U17214 (N_17214,N_14865,N_10283);
nor U17215 (N_17215,N_12694,N_13108);
or U17216 (N_17216,N_10267,N_11308);
nand U17217 (N_17217,N_10113,N_10200);
nand U17218 (N_17218,N_12607,N_14710);
and U17219 (N_17219,N_10252,N_13601);
xnor U17220 (N_17220,N_11367,N_13011);
nand U17221 (N_17221,N_10492,N_13949);
or U17222 (N_17222,N_11162,N_10088);
nor U17223 (N_17223,N_10044,N_14540);
and U17224 (N_17224,N_14828,N_14548);
or U17225 (N_17225,N_10343,N_10230);
and U17226 (N_17226,N_11487,N_10575);
and U17227 (N_17227,N_13769,N_11738);
xor U17228 (N_17228,N_12505,N_14234);
nand U17229 (N_17229,N_11105,N_10902);
xor U17230 (N_17230,N_11211,N_12851);
or U17231 (N_17231,N_13213,N_12886);
and U17232 (N_17232,N_14658,N_14456);
or U17233 (N_17233,N_14942,N_14675);
or U17234 (N_17234,N_10018,N_14160);
xnor U17235 (N_17235,N_13386,N_10325);
xnor U17236 (N_17236,N_13910,N_12925);
xor U17237 (N_17237,N_13048,N_14851);
nor U17238 (N_17238,N_10597,N_14209);
or U17239 (N_17239,N_11264,N_10541);
and U17240 (N_17240,N_11522,N_13531);
or U17241 (N_17241,N_14117,N_13645);
and U17242 (N_17242,N_14941,N_10373);
nand U17243 (N_17243,N_14039,N_12697);
nand U17244 (N_17244,N_10984,N_13222);
and U17245 (N_17245,N_14526,N_14949);
nand U17246 (N_17246,N_13014,N_11995);
nor U17247 (N_17247,N_14894,N_13736);
nand U17248 (N_17248,N_10131,N_13137);
and U17249 (N_17249,N_13393,N_14900);
or U17250 (N_17250,N_11517,N_11142);
or U17251 (N_17251,N_11466,N_14607);
and U17252 (N_17252,N_10133,N_12243);
nor U17253 (N_17253,N_12726,N_14764);
or U17254 (N_17254,N_10823,N_11242);
and U17255 (N_17255,N_10342,N_11566);
and U17256 (N_17256,N_10604,N_13216);
or U17257 (N_17257,N_12119,N_13882);
nand U17258 (N_17258,N_14814,N_14559);
nand U17259 (N_17259,N_12923,N_13007);
nand U17260 (N_17260,N_10657,N_10521);
nor U17261 (N_17261,N_13678,N_14326);
nand U17262 (N_17262,N_12995,N_14399);
and U17263 (N_17263,N_10987,N_11789);
or U17264 (N_17264,N_12657,N_12154);
nor U17265 (N_17265,N_14692,N_10680);
and U17266 (N_17266,N_11041,N_12701);
nand U17267 (N_17267,N_11038,N_14943);
xnor U17268 (N_17268,N_14189,N_11637);
nand U17269 (N_17269,N_10550,N_13670);
and U17270 (N_17270,N_11252,N_12902);
and U17271 (N_17271,N_10925,N_10954);
or U17272 (N_17272,N_11287,N_11240);
xnor U17273 (N_17273,N_10887,N_12439);
nand U17274 (N_17274,N_12666,N_11812);
nand U17275 (N_17275,N_13056,N_11191);
nand U17276 (N_17276,N_12762,N_12023);
or U17277 (N_17277,N_13344,N_10669);
nand U17278 (N_17278,N_12956,N_11450);
xor U17279 (N_17279,N_12671,N_14371);
nand U17280 (N_17280,N_12472,N_12617);
nor U17281 (N_17281,N_12907,N_14123);
or U17282 (N_17282,N_13523,N_11018);
nand U17283 (N_17283,N_13832,N_11238);
or U17284 (N_17284,N_11932,N_10706);
nand U17285 (N_17285,N_10986,N_11841);
and U17286 (N_17286,N_12204,N_14724);
or U17287 (N_17287,N_10275,N_13341);
nor U17288 (N_17288,N_12639,N_12295);
nand U17289 (N_17289,N_14085,N_14602);
or U17290 (N_17290,N_11153,N_10137);
nand U17291 (N_17291,N_14074,N_10465);
xnor U17292 (N_17292,N_11568,N_10443);
and U17293 (N_17293,N_10962,N_12262);
xnor U17294 (N_17294,N_13025,N_11461);
and U17295 (N_17295,N_10177,N_12390);
or U17296 (N_17296,N_13181,N_14357);
or U17297 (N_17297,N_14628,N_11149);
xnor U17298 (N_17298,N_10280,N_13136);
nor U17299 (N_17299,N_13305,N_12323);
or U17300 (N_17300,N_10424,N_12715);
and U17301 (N_17301,N_14405,N_10242);
or U17302 (N_17302,N_14104,N_14859);
nor U17303 (N_17303,N_11378,N_10357);
nand U17304 (N_17304,N_12864,N_11104);
or U17305 (N_17305,N_13575,N_13377);
xnor U17306 (N_17306,N_14600,N_13243);
nor U17307 (N_17307,N_10319,N_11733);
xor U17308 (N_17308,N_14972,N_13024);
or U17309 (N_17309,N_14833,N_11526);
or U17310 (N_17310,N_13079,N_10286);
and U17311 (N_17311,N_11225,N_10190);
xor U17312 (N_17312,N_11187,N_12256);
and U17313 (N_17313,N_14846,N_14427);
nand U17314 (N_17314,N_10501,N_11236);
nor U17315 (N_17315,N_13751,N_12763);
or U17316 (N_17316,N_14472,N_14808);
nor U17317 (N_17317,N_10875,N_11546);
or U17318 (N_17318,N_11437,N_14361);
nor U17319 (N_17319,N_14908,N_13944);
or U17320 (N_17320,N_14161,N_12421);
nand U17321 (N_17321,N_13289,N_12804);
and U17322 (N_17322,N_10497,N_12612);
and U17323 (N_17323,N_12509,N_11769);
nand U17324 (N_17324,N_14272,N_11636);
nor U17325 (N_17325,N_12235,N_14515);
nand U17326 (N_17326,N_11907,N_13109);
xor U17327 (N_17327,N_10340,N_11133);
nor U17328 (N_17328,N_12003,N_12451);
nor U17329 (N_17329,N_14187,N_13824);
and U17330 (N_17330,N_11205,N_14295);
and U17331 (N_17331,N_11993,N_11368);
nor U17332 (N_17332,N_14842,N_13012);
nand U17333 (N_17333,N_12447,N_10259);
and U17334 (N_17334,N_12153,N_10057);
nor U17335 (N_17335,N_14365,N_10072);
nand U17336 (N_17336,N_12985,N_12669);
and U17337 (N_17337,N_14918,N_10540);
nor U17338 (N_17338,N_10317,N_11198);
nor U17339 (N_17339,N_10571,N_12168);
xor U17340 (N_17340,N_11129,N_12348);
nand U17341 (N_17341,N_11901,N_11879);
nor U17342 (N_17342,N_13886,N_10906);
nor U17343 (N_17343,N_11793,N_13685);
or U17344 (N_17344,N_10754,N_13918);
nor U17345 (N_17345,N_10294,N_10857);
nand U17346 (N_17346,N_14004,N_13848);
and U17347 (N_17347,N_14333,N_14432);
or U17348 (N_17348,N_11521,N_12510);
nor U17349 (N_17349,N_10356,N_13777);
and U17350 (N_17350,N_12302,N_14180);
nand U17351 (N_17351,N_14768,N_10299);
xnor U17352 (N_17352,N_13189,N_14051);
or U17353 (N_17353,N_14119,N_13607);
nor U17354 (N_17354,N_13071,N_12194);
nand U17355 (N_17355,N_14639,N_10459);
nor U17356 (N_17356,N_14052,N_10339);
nand U17357 (N_17357,N_14701,N_14033);
nor U17358 (N_17358,N_10401,N_14678);
nand U17359 (N_17359,N_12882,N_14793);
nor U17360 (N_17360,N_12584,N_14823);
xnor U17361 (N_17361,N_14241,N_11813);
nor U17362 (N_17362,N_11204,N_11502);
or U17363 (N_17363,N_11619,N_11524);
nor U17364 (N_17364,N_14596,N_13767);
and U17365 (N_17365,N_13620,N_13201);
or U17366 (N_17366,N_14296,N_12053);
nor U17367 (N_17367,N_10814,N_11383);
and U17368 (N_17368,N_11108,N_10907);
nand U17369 (N_17369,N_11136,N_14599);
nor U17370 (N_17370,N_11854,N_11446);
or U17371 (N_17371,N_11871,N_10661);
xnor U17372 (N_17372,N_10136,N_13132);
or U17373 (N_17373,N_10625,N_14545);
or U17374 (N_17374,N_10087,N_14026);
xor U17375 (N_17375,N_10796,N_11541);
nand U17376 (N_17376,N_12354,N_12371);
and U17377 (N_17377,N_14547,N_13225);
or U17378 (N_17378,N_13581,N_12192);
xnor U17379 (N_17379,N_13901,N_10451);
nor U17380 (N_17380,N_12462,N_11387);
nor U17381 (N_17381,N_11071,N_10220);
and U17382 (N_17382,N_14474,N_11452);
xor U17383 (N_17383,N_10695,N_14870);
and U17384 (N_17384,N_10789,N_10099);
or U17385 (N_17385,N_10708,N_11014);
and U17386 (N_17386,N_11874,N_12394);
nand U17387 (N_17387,N_10361,N_13694);
and U17388 (N_17388,N_11557,N_14157);
or U17389 (N_17389,N_10254,N_11480);
or U17390 (N_17390,N_12723,N_12833);
xnor U17391 (N_17391,N_11946,N_11166);
nand U17392 (N_17392,N_11785,N_11459);
nand U17393 (N_17393,N_12967,N_10101);
nor U17394 (N_17394,N_13521,N_13539);
nand U17395 (N_17395,N_14175,N_10162);
xnor U17396 (N_17396,N_11704,N_12496);
nand U17397 (N_17397,N_10963,N_10462);
and U17398 (N_17398,N_13961,N_11991);
or U17399 (N_17399,N_13065,N_11682);
and U17400 (N_17400,N_13836,N_12857);
or U17401 (N_17401,N_13053,N_13092);
xor U17402 (N_17402,N_10234,N_10915);
nor U17403 (N_17403,N_10780,N_10855);
nand U17404 (N_17404,N_13208,N_11323);
and U17405 (N_17405,N_12250,N_11966);
or U17406 (N_17406,N_14831,N_13634);
or U17407 (N_17407,N_11832,N_14430);
nor U17408 (N_17408,N_13174,N_10988);
nor U17409 (N_17409,N_12582,N_14948);
or U17410 (N_17410,N_14407,N_13180);
nor U17411 (N_17411,N_10285,N_12272);
nor U17412 (N_17412,N_11528,N_13030);
nand U17413 (N_17413,N_13675,N_11439);
xnor U17414 (N_17414,N_14997,N_10825);
or U17415 (N_17415,N_10093,N_12506);
and U17416 (N_17416,N_13841,N_10050);
or U17417 (N_17417,N_10454,N_12497);
and U17418 (N_17418,N_13974,N_10957);
nand U17419 (N_17419,N_10931,N_10028);
and U17420 (N_17420,N_12818,N_11376);
or U17421 (N_17421,N_12341,N_13885);
or U17422 (N_17422,N_11248,N_11802);
and U17423 (N_17423,N_14568,N_12975);
or U17424 (N_17424,N_13569,N_11390);
or U17425 (N_17425,N_13986,N_12226);
or U17426 (N_17426,N_11892,N_12376);
xor U17427 (N_17427,N_11633,N_14059);
or U17428 (N_17428,N_14681,N_11760);
nor U17429 (N_17429,N_13387,N_13347);
nand U17430 (N_17430,N_10938,N_14668);
nor U17431 (N_17431,N_13363,N_12188);
and U17432 (N_17432,N_12086,N_14115);
xor U17433 (N_17433,N_12214,N_10329);
nor U17434 (N_17434,N_13881,N_10471);
nand U17435 (N_17435,N_10791,N_13235);
xor U17436 (N_17436,N_13068,N_14097);
or U17437 (N_17437,N_12147,N_11021);
xnor U17438 (N_17438,N_14573,N_12823);
nand U17439 (N_17439,N_12662,N_13586);
nor U17440 (N_17440,N_10040,N_13260);
or U17441 (N_17441,N_12828,N_11434);
or U17442 (N_17442,N_14071,N_12190);
and U17443 (N_17443,N_11064,N_12996);
nor U17444 (N_17444,N_12581,N_10073);
xor U17445 (N_17445,N_10926,N_11605);
or U17446 (N_17446,N_14324,N_10445);
or U17447 (N_17447,N_11754,N_13872);
or U17448 (N_17448,N_13982,N_10646);
and U17449 (N_17449,N_11379,N_13337);
nand U17450 (N_17450,N_10469,N_11681);
nor U17451 (N_17451,N_12030,N_13339);
nand U17452 (N_17452,N_10021,N_10063);
or U17453 (N_17453,N_12481,N_13345);
nor U17454 (N_17454,N_11164,N_12643);
nor U17455 (N_17455,N_13365,N_14875);
or U17456 (N_17456,N_10601,N_10427);
nor U17457 (N_17457,N_10577,N_10686);
nand U17458 (N_17458,N_14669,N_13985);
nand U17459 (N_17459,N_10185,N_12797);
nor U17460 (N_17460,N_11673,N_14636);
or U17461 (N_17461,N_14438,N_12615);
or U17462 (N_17462,N_13595,N_12391);
or U17463 (N_17463,N_11110,N_10676);
nor U17464 (N_17464,N_10295,N_13669);
and U17465 (N_17465,N_13672,N_12538);
and U17466 (N_17466,N_10049,N_13044);
or U17467 (N_17467,N_13008,N_13031);
nor U17468 (N_17468,N_13896,N_12392);
nor U17469 (N_17469,N_10219,N_14273);
or U17470 (N_17470,N_13116,N_12425);
nor U17471 (N_17471,N_14439,N_10549);
nor U17472 (N_17472,N_13087,N_12001);
nor U17473 (N_17473,N_12461,N_11767);
nand U17474 (N_17474,N_10833,N_14261);
and U17475 (N_17475,N_12104,N_11042);
xor U17476 (N_17476,N_14565,N_12873);
nand U17477 (N_17477,N_14023,N_14120);
xor U17478 (N_17478,N_12305,N_10723);
and U17479 (N_17479,N_13681,N_14338);
nand U17480 (N_17480,N_13153,N_12089);
nand U17481 (N_17481,N_12347,N_13730);
nand U17482 (N_17482,N_13582,N_11941);
and U17483 (N_17483,N_12084,N_14135);
or U17484 (N_17484,N_14964,N_14461);
nor U17485 (N_17485,N_10673,N_12006);
nand U17486 (N_17486,N_11420,N_14344);
nor U17487 (N_17487,N_12294,N_11192);
nand U17488 (N_17488,N_11817,N_13628);
nor U17489 (N_17489,N_13440,N_11027);
nor U17490 (N_17490,N_13438,N_13088);
nand U17491 (N_17491,N_11721,N_13242);
nand U17492 (N_17492,N_14638,N_11719);
and U17493 (N_17493,N_11622,N_12311);
xnor U17494 (N_17494,N_12378,N_13540);
or U17495 (N_17495,N_13833,N_14377);
nand U17496 (N_17496,N_11777,N_11009);
nor U17497 (N_17497,N_12018,N_13709);
nor U17498 (N_17498,N_11679,N_10702);
or U17499 (N_17499,N_11988,N_14758);
nand U17500 (N_17500,N_13921,N_13412);
xnor U17501 (N_17501,N_10009,N_13842);
and U17502 (N_17502,N_10306,N_11786);
and U17503 (N_17503,N_12053,N_11607);
nor U17504 (N_17504,N_14211,N_12703);
or U17505 (N_17505,N_10991,N_12426);
or U17506 (N_17506,N_13577,N_10271);
nor U17507 (N_17507,N_14140,N_11936);
and U17508 (N_17508,N_10103,N_11785);
nand U17509 (N_17509,N_11604,N_13172);
nand U17510 (N_17510,N_10119,N_12806);
or U17511 (N_17511,N_13604,N_12731);
and U17512 (N_17512,N_12610,N_13747);
nor U17513 (N_17513,N_14113,N_14448);
xor U17514 (N_17514,N_10478,N_12710);
nand U17515 (N_17515,N_12937,N_12279);
nand U17516 (N_17516,N_11929,N_13909);
nor U17517 (N_17517,N_14687,N_14016);
and U17518 (N_17518,N_12271,N_10732);
nor U17519 (N_17519,N_13244,N_10225);
nor U17520 (N_17520,N_12171,N_12445);
nor U17521 (N_17521,N_13935,N_12820);
xnor U17522 (N_17522,N_10883,N_12497);
and U17523 (N_17523,N_14243,N_11692);
xnor U17524 (N_17524,N_11939,N_12487);
nor U17525 (N_17525,N_12737,N_13522);
nand U17526 (N_17526,N_12345,N_10196);
or U17527 (N_17527,N_11935,N_13066);
or U17528 (N_17528,N_10558,N_14811);
or U17529 (N_17529,N_13635,N_11576);
xor U17530 (N_17530,N_10678,N_12624);
xor U17531 (N_17531,N_10552,N_11513);
and U17532 (N_17532,N_14139,N_13374);
xnor U17533 (N_17533,N_10601,N_14129);
nor U17534 (N_17534,N_13919,N_14593);
xnor U17535 (N_17535,N_14946,N_12966);
and U17536 (N_17536,N_12380,N_11215);
nand U17537 (N_17537,N_10536,N_14882);
and U17538 (N_17538,N_14177,N_10911);
and U17539 (N_17539,N_11969,N_12256);
nand U17540 (N_17540,N_13312,N_11736);
nand U17541 (N_17541,N_12712,N_10501);
nor U17542 (N_17542,N_12119,N_10242);
nor U17543 (N_17543,N_10203,N_14312);
nor U17544 (N_17544,N_13569,N_14713);
xor U17545 (N_17545,N_11595,N_11458);
nand U17546 (N_17546,N_10143,N_14243);
nand U17547 (N_17547,N_10710,N_12365);
and U17548 (N_17548,N_12661,N_11905);
xor U17549 (N_17549,N_14855,N_12141);
nor U17550 (N_17550,N_13403,N_13435);
nor U17551 (N_17551,N_11125,N_13569);
or U17552 (N_17552,N_14519,N_12657);
nand U17553 (N_17553,N_10150,N_11252);
nand U17554 (N_17554,N_11128,N_10577);
nand U17555 (N_17555,N_13498,N_12044);
and U17556 (N_17556,N_14927,N_11866);
or U17557 (N_17557,N_12699,N_10062);
and U17558 (N_17558,N_10792,N_10350);
or U17559 (N_17559,N_14682,N_14167);
nor U17560 (N_17560,N_10294,N_12718);
nand U17561 (N_17561,N_14415,N_13381);
and U17562 (N_17562,N_14481,N_13331);
nor U17563 (N_17563,N_13182,N_12856);
nand U17564 (N_17564,N_12661,N_12303);
or U17565 (N_17565,N_13647,N_14960);
xnor U17566 (N_17566,N_12006,N_10285);
nor U17567 (N_17567,N_13745,N_14870);
or U17568 (N_17568,N_10751,N_12278);
nand U17569 (N_17569,N_11485,N_13016);
and U17570 (N_17570,N_13166,N_10848);
nor U17571 (N_17571,N_11055,N_11922);
xor U17572 (N_17572,N_11858,N_11258);
or U17573 (N_17573,N_10742,N_14681);
and U17574 (N_17574,N_11405,N_10321);
or U17575 (N_17575,N_11573,N_14502);
nor U17576 (N_17576,N_11398,N_14594);
and U17577 (N_17577,N_14156,N_11090);
and U17578 (N_17578,N_10595,N_13950);
nand U17579 (N_17579,N_11323,N_11339);
nand U17580 (N_17580,N_10633,N_14184);
nand U17581 (N_17581,N_13942,N_10841);
and U17582 (N_17582,N_12056,N_14938);
nand U17583 (N_17583,N_14270,N_12664);
xor U17584 (N_17584,N_10557,N_11475);
nand U17585 (N_17585,N_10475,N_13851);
nor U17586 (N_17586,N_13843,N_13235);
and U17587 (N_17587,N_12835,N_11043);
nand U17588 (N_17588,N_11938,N_13709);
nand U17589 (N_17589,N_13872,N_14574);
and U17590 (N_17590,N_11188,N_11315);
nor U17591 (N_17591,N_12634,N_10630);
nand U17592 (N_17592,N_13729,N_13883);
nand U17593 (N_17593,N_13709,N_10811);
nor U17594 (N_17594,N_13770,N_13792);
and U17595 (N_17595,N_11226,N_11884);
nor U17596 (N_17596,N_13434,N_11707);
xnor U17597 (N_17597,N_12152,N_11480);
xor U17598 (N_17598,N_11358,N_14461);
nor U17599 (N_17599,N_14392,N_13258);
nand U17600 (N_17600,N_13127,N_12114);
xor U17601 (N_17601,N_11571,N_14320);
or U17602 (N_17602,N_13598,N_12102);
xnor U17603 (N_17603,N_12523,N_13254);
nor U17604 (N_17604,N_11326,N_14057);
or U17605 (N_17605,N_11061,N_10658);
xnor U17606 (N_17606,N_12869,N_10133);
xor U17607 (N_17607,N_10890,N_11929);
and U17608 (N_17608,N_14935,N_14612);
xnor U17609 (N_17609,N_13901,N_11743);
and U17610 (N_17610,N_12115,N_14652);
nand U17611 (N_17611,N_10844,N_11385);
nor U17612 (N_17612,N_10013,N_10715);
nor U17613 (N_17613,N_13239,N_14537);
and U17614 (N_17614,N_14708,N_12218);
nor U17615 (N_17615,N_13047,N_11860);
nor U17616 (N_17616,N_14358,N_11088);
or U17617 (N_17617,N_14107,N_11475);
nand U17618 (N_17618,N_12350,N_10645);
or U17619 (N_17619,N_11732,N_13650);
and U17620 (N_17620,N_13697,N_10836);
nor U17621 (N_17621,N_10390,N_14927);
and U17622 (N_17622,N_13813,N_14875);
and U17623 (N_17623,N_12696,N_14645);
or U17624 (N_17624,N_12225,N_14594);
and U17625 (N_17625,N_11391,N_11702);
and U17626 (N_17626,N_11609,N_10203);
or U17627 (N_17627,N_13398,N_13708);
or U17628 (N_17628,N_10523,N_14048);
nor U17629 (N_17629,N_13071,N_10872);
nor U17630 (N_17630,N_12260,N_12619);
and U17631 (N_17631,N_13676,N_13941);
nor U17632 (N_17632,N_12355,N_13707);
nand U17633 (N_17633,N_14339,N_14869);
or U17634 (N_17634,N_10262,N_10425);
nor U17635 (N_17635,N_11012,N_10459);
nor U17636 (N_17636,N_13023,N_11024);
nand U17637 (N_17637,N_11148,N_10291);
and U17638 (N_17638,N_12765,N_13515);
nand U17639 (N_17639,N_11788,N_11031);
nand U17640 (N_17640,N_13322,N_13122);
nand U17641 (N_17641,N_12150,N_11085);
nand U17642 (N_17642,N_12287,N_12262);
nand U17643 (N_17643,N_12535,N_11039);
and U17644 (N_17644,N_11070,N_10979);
or U17645 (N_17645,N_14223,N_11722);
xnor U17646 (N_17646,N_12337,N_12759);
and U17647 (N_17647,N_14732,N_11914);
and U17648 (N_17648,N_10900,N_13447);
and U17649 (N_17649,N_11664,N_14220);
nor U17650 (N_17650,N_13986,N_10728);
or U17651 (N_17651,N_13773,N_13980);
nor U17652 (N_17652,N_13925,N_11291);
nor U17653 (N_17653,N_12269,N_12076);
or U17654 (N_17654,N_14860,N_12968);
or U17655 (N_17655,N_12220,N_11686);
and U17656 (N_17656,N_10138,N_13994);
nand U17657 (N_17657,N_12778,N_11491);
nor U17658 (N_17658,N_11385,N_11099);
and U17659 (N_17659,N_14564,N_13609);
and U17660 (N_17660,N_10794,N_13271);
nand U17661 (N_17661,N_14543,N_12582);
or U17662 (N_17662,N_11082,N_11100);
or U17663 (N_17663,N_10648,N_12713);
nand U17664 (N_17664,N_10291,N_12017);
and U17665 (N_17665,N_14109,N_13935);
nor U17666 (N_17666,N_12487,N_14888);
and U17667 (N_17667,N_10282,N_11790);
nor U17668 (N_17668,N_14436,N_10794);
and U17669 (N_17669,N_11600,N_10804);
nor U17670 (N_17670,N_14609,N_11971);
nor U17671 (N_17671,N_11545,N_14933);
and U17672 (N_17672,N_11982,N_12379);
and U17673 (N_17673,N_12767,N_12708);
nor U17674 (N_17674,N_10957,N_12322);
or U17675 (N_17675,N_12641,N_14485);
or U17676 (N_17676,N_13987,N_10891);
nor U17677 (N_17677,N_14454,N_13556);
nand U17678 (N_17678,N_12743,N_11336);
nand U17679 (N_17679,N_12846,N_14589);
or U17680 (N_17680,N_14244,N_11488);
and U17681 (N_17681,N_14609,N_11041);
nand U17682 (N_17682,N_11675,N_12107);
nand U17683 (N_17683,N_11316,N_13750);
nor U17684 (N_17684,N_11883,N_11539);
and U17685 (N_17685,N_11700,N_10995);
nor U17686 (N_17686,N_13825,N_12114);
and U17687 (N_17687,N_14511,N_10499);
nor U17688 (N_17688,N_10272,N_13851);
nand U17689 (N_17689,N_11456,N_13723);
nand U17690 (N_17690,N_10591,N_11447);
xnor U17691 (N_17691,N_14911,N_12438);
or U17692 (N_17692,N_14111,N_14054);
and U17693 (N_17693,N_13033,N_12145);
nor U17694 (N_17694,N_10107,N_11150);
and U17695 (N_17695,N_12290,N_14553);
nor U17696 (N_17696,N_10000,N_11433);
xnor U17697 (N_17697,N_12735,N_14175);
xnor U17698 (N_17698,N_13222,N_12066);
nand U17699 (N_17699,N_12148,N_14704);
nor U17700 (N_17700,N_10057,N_12582);
nor U17701 (N_17701,N_11523,N_13755);
nand U17702 (N_17702,N_14527,N_12432);
nor U17703 (N_17703,N_12535,N_12985);
or U17704 (N_17704,N_14283,N_13903);
or U17705 (N_17705,N_13491,N_13089);
nor U17706 (N_17706,N_10043,N_13388);
nor U17707 (N_17707,N_13280,N_12459);
nor U17708 (N_17708,N_10470,N_12290);
nand U17709 (N_17709,N_13853,N_10096);
and U17710 (N_17710,N_10272,N_14691);
nand U17711 (N_17711,N_11710,N_11102);
xnor U17712 (N_17712,N_14402,N_12878);
and U17713 (N_17713,N_12099,N_11456);
or U17714 (N_17714,N_11596,N_12635);
nor U17715 (N_17715,N_12299,N_12055);
or U17716 (N_17716,N_13389,N_14241);
or U17717 (N_17717,N_14884,N_13785);
nand U17718 (N_17718,N_10674,N_10968);
nor U17719 (N_17719,N_12620,N_12639);
xor U17720 (N_17720,N_10251,N_10354);
or U17721 (N_17721,N_13159,N_10733);
or U17722 (N_17722,N_12597,N_10658);
nor U17723 (N_17723,N_13243,N_10452);
and U17724 (N_17724,N_12165,N_12881);
and U17725 (N_17725,N_12914,N_11271);
and U17726 (N_17726,N_10058,N_14442);
and U17727 (N_17727,N_12600,N_14658);
and U17728 (N_17728,N_10244,N_11410);
and U17729 (N_17729,N_10293,N_14691);
nand U17730 (N_17730,N_11865,N_13238);
nor U17731 (N_17731,N_13063,N_13952);
nand U17732 (N_17732,N_13514,N_14509);
and U17733 (N_17733,N_11032,N_12893);
nand U17734 (N_17734,N_13614,N_13860);
nor U17735 (N_17735,N_11641,N_14203);
nand U17736 (N_17736,N_11652,N_14019);
and U17737 (N_17737,N_13274,N_12562);
xor U17738 (N_17738,N_11781,N_13314);
or U17739 (N_17739,N_10475,N_14815);
and U17740 (N_17740,N_12908,N_12039);
or U17741 (N_17741,N_14260,N_13776);
or U17742 (N_17742,N_13021,N_12671);
xnor U17743 (N_17743,N_11271,N_11613);
or U17744 (N_17744,N_14209,N_13192);
and U17745 (N_17745,N_10389,N_10167);
nand U17746 (N_17746,N_13609,N_13548);
or U17747 (N_17747,N_14451,N_12987);
and U17748 (N_17748,N_12631,N_13607);
or U17749 (N_17749,N_10278,N_11493);
nor U17750 (N_17750,N_13227,N_13946);
or U17751 (N_17751,N_10816,N_11713);
and U17752 (N_17752,N_12277,N_14117);
and U17753 (N_17753,N_11415,N_12010);
and U17754 (N_17754,N_14604,N_11915);
and U17755 (N_17755,N_10926,N_13230);
or U17756 (N_17756,N_10387,N_13783);
or U17757 (N_17757,N_11287,N_12939);
xor U17758 (N_17758,N_12552,N_13540);
xor U17759 (N_17759,N_10316,N_12633);
and U17760 (N_17760,N_14911,N_14356);
or U17761 (N_17761,N_11850,N_14215);
and U17762 (N_17762,N_13632,N_11357);
nand U17763 (N_17763,N_10737,N_12924);
and U17764 (N_17764,N_12588,N_10132);
nand U17765 (N_17765,N_13334,N_14407);
xor U17766 (N_17766,N_12129,N_12111);
or U17767 (N_17767,N_14756,N_11405);
nand U17768 (N_17768,N_11194,N_10171);
nand U17769 (N_17769,N_12259,N_11775);
or U17770 (N_17770,N_12512,N_11623);
and U17771 (N_17771,N_12141,N_10988);
or U17772 (N_17772,N_13578,N_13831);
or U17773 (N_17773,N_12299,N_10555);
or U17774 (N_17774,N_12897,N_12328);
nor U17775 (N_17775,N_10085,N_13031);
nor U17776 (N_17776,N_10483,N_13444);
nand U17777 (N_17777,N_14614,N_11287);
or U17778 (N_17778,N_14646,N_13396);
nor U17779 (N_17779,N_11745,N_10218);
nand U17780 (N_17780,N_13215,N_11790);
and U17781 (N_17781,N_11299,N_12396);
or U17782 (N_17782,N_10435,N_12833);
nor U17783 (N_17783,N_11317,N_13084);
xor U17784 (N_17784,N_10662,N_11191);
or U17785 (N_17785,N_12777,N_11338);
and U17786 (N_17786,N_12789,N_10192);
nor U17787 (N_17787,N_12967,N_14097);
or U17788 (N_17788,N_12725,N_10653);
xnor U17789 (N_17789,N_14214,N_11686);
xnor U17790 (N_17790,N_13146,N_10040);
nand U17791 (N_17791,N_13977,N_11863);
xor U17792 (N_17792,N_12406,N_12216);
and U17793 (N_17793,N_12755,N_10021);
or U17794 (N_17794,N_14031,N_14739);
nor U17795 (N_17795,N_10302,N_10131);
or U17796 (N_17796,N_12694,N_13853);
nor U17797 (N_17797,N_11507,N_12890);
nor U17798 (N_17798,N_12612,N_13323);
or U17799 (N_17799,N_12330,N_11447);
xor U17800 (N_17800,N_10548,N_10780);
and U17801 (N_17801,N_12374,N_11341);
nor U17802 (N_17802,N_14348,N_10238);
nand U17803 (N_17803,N_14020,N_14584);
or U17804 (N_17804,N_11955,N_14257);
or U17805 (N_17805,N_14783,N_11178);
nor U17806 (N_17806,N_13331,N_10955);
or U17807 (N_17807,N_12224,N_14085);
nor U17808 (N_17808,N_11965,N_11211);
nor U17809 (N_17809,N_13808,N_12710);
nand U17810 (N_17810,N_13873,N_10328);
nand U17811 (N_17811,N_13840,N_11414);
and U17812 (N_17812,N_12531,N_12766);
and U17813 (N_17813,N_11155,N_13119);
nor U17814 (N_17814,N_11189,N_10485);
nand U17815 (N_17815,N_11577,N_13949);
nor U17816 (N_17816,N_12349,N_14722);
nand U17817 (N_17817,N_13121,N_12887);
or U17818 (N_17818,N_10428,N_11919);
xnor U17819 (N_17819,N_13924,N_11395);
nand U17820 (N_17820,N_12537,N_12858);
or U17821 (N_17821,N_11175,N_14421);
and U17822 (N_17822,N_12669,N_14678);
nand U17823 (N_17823,N_14951,N_14472);
or U17824 (N_17824,N_12214,N_10345);
nand U17825 (N_17825,N_11464,N_13908);
nor U17826 (N_17826,N_11064,N_10822);
nor U17827 (N_17827,N_12661,N_14490);
and U17828 (N_17828,N_11030,N_12386);
nor U17829 (N_17829,N_13245,N_13504);
nor U17830 (N_17830,N_13312,N_10348);
nand U17831 (N_17831,N_11377,N_12863);
nor U17832 (N_17832,N_12457,N_11354);
nor U17833 (N_17833,N_10101,N_10001);
nor U17834 (N_17834,N_12090,N_10275);
nand U17835 (N_17835,N_11020,N_13622);
or U17836 (N_17836,N_13109,N_13626);
nand U17837 (N_17837,N_10914,N_12597);
nor U17838 (N_17838,N_10976,N_13569);
and U17839 (N_17839,N_11843,N_12867);
nand U17840 (N_17840,N_11481,N_14421);
or U17841 (N_17841,N_14673,N_14426);
nand U17842 (N_17842,N_10831,N_14694);
nor U17843 (N_17843,N_13190,N_13268);
nand U17844 (N_17844,N_13480,N_12225);
nor U17845 (N_17845,N_10173,N_11250);
or U17846 (N_17846,N_13874,N_13370);
nand U17847 (N_17847,N_11502,N_14024);
xor U17848 (N_17848,N_10552,N_12600);
or U17849 (N_17849,N_13034,N_11632);
or U17850 (N_17850,N_11787,N_13526);
xor U17851 (N_17851,N_13762,N_11644);
and U17852 (N_17852,N_12312,N_12735);
xnor U17853 (N_17853,N_10185,N_13440);
and U17854 (N_17854,N_13863,N_11392);
nor U17855 (N_17855,N_12240,N_14802);
and U17856 (N_17856,N_12760,N_13305);
nor U17857 (N_17857,N_12868,N_10982);
nand U17858 (N_17858,N_12042,N_10863);
or U17859 (N_17859,N_12017,N_14346);
or U17860 (N_17860,N_10800,N_10035);
and U17861 (N_17861,N_14386,N_13550);
nor U17862 (N_17862,N_13217,N_11941);
nor U17863 (N_17863,N_14344,N_14422);
or U17864 (N_17864,N_12393,N_10125);
or U17865 (N_17865,N_10570,N_12181);
or U17866 (N_17866,N_11531,N_14181);
nand U17867 (N_17867,N_13520,N_14202);
nor U17868 (N_17868,N_12733,N_13153);
and U17869 (N_17869,N_12989,N_14686);
and U17870 (N_17870,N_10702,N_12058);
and U17871 (N_17871,N_11425,N_12330);
nand U17872 (N_17872,N_11655,N_11738);
nand U17873 (N_17873,N_10529,N_13873);
and U17874 (N_17874,N_11574,N_10610);
or U17875 (N_17875,N_13702,N_11948);
nor U17876 (N_17876,N_13679,N_14851);
and U17877 (N_17877,N_13437,N_10799);
nor U17878 (N_17878,N_10960,N_14876);
nor U17879 (N_17879,N_13326,N_12544);
and U17880 (N_17880,N_10551,N_14829);
xor U17881 (N_17881,N_13089,N_11983);
nand U17882 (N_17882,N_12133,N_12096);
nor U17883 (N_17883,N_12534,N_12850);
xor U17884 (N_17884,N_14920,N_10501);
nand U17885 (N_17885,N_11270,N_11536);
nand U17886 (N_17886,N_11831,N_14634);
or U17887 (N_17887,N_14240,N_12607);
or U17888 (N_17888,N_11503,N_13012);
nor U17889 (N_17889,N_10273,N_10097);
nand U17890 (N_17890,N_12023,N_13416);
xor U17891 (N_17891,N_11274,N_11539);
and U17892 (N_17892,N_10028,N_12171);
nor U17893 (N_17893,N_12684,N_14353);
nand U17894 (N_17894,N_13729,N_14699);
nand U17895 (N_17895,N_12062,N_13969);
xor U17896 (N_17896,N_11772,N_10832);
or U17897 (N_17897,N_13977,N_14335);
nand U17898 (N_17898,N_11821,N_13090);
or U17899 (N_17899,N_13190,N_11601);
or U17900 (N_17900,N_11472,N_12544);
nand U17901 (N_17901,N_10375,N_10582);
and U17902 (N_17902,N_13529,N_14407);
or U17903 (N_17903,N_10100,N_11778);
or U17904 (N_17904,N_12910,N_14716);
or U17905 (N_17905,N_12280,N_14059);
nand U17906 (N_17906,N_12819,N_11870);
and U17907 (N_17907,N_13935,N_14847);
and U17908 (N_17908,N_10905,N_10899);
nand U17909 (N_17909,N_10084,N_12113);
xor U17910 (N_17910,N_14735,N_11217);
and U17911 (N_17911,N_14355,N_13666);
and U17912 (N_17912,N_14825,N_13077);
or U17913 (N_17913,N_12744,N_10326);
nand U17914 (N_17914,N_13033,N_13152);
and U17915 (N_17915,N_13920,N_10739);
or U17916 (N_17916,N_12406,N_10915);
xnor U17917 (N_17917,N_12540,N_10216);
or U17918 (N_17918,N_14812,N_14708);
or U17919 (N_17919,N_14236,N_13433);
and U17920 (N_17920,N_12498,N_11992);
nor U17921 (N_17921,N_12389,N_10721);
nor U17922 (N_17922,N_11474,N_14971);
nor U17923 (N_17923,N_14768,N_12628);
and U17924 (N_17924,N_13131,N_10470);
or U17925 (N_17925,N_14817,N_10318);
nor U17926 (N_17926,N_13798,N_10680);
nor U17927 (N_17927,N_14114,N_10126);
or U17928 (N_17928,N_13013,N_12952);
nor U17929 (N_17929,N_11289,N_10071);
xor U17930 (N_17930,N_14189,N_10606);
nor U17931 (N_17931,N_12977,N_13932);
nor U17932 (N_17932,N_11938,N_14510);
or U17933 (N_17933,N_11081,N_11347);
nand U17934 (N_17934,N_12818,N_12285);
nor U17935 (N_17935,N_14639,N_11598);
nand U17936 (N_17936,N_14141,N_10600);
or U17937 (N_17937,N_10868,N_12566);
nand U17938 (N_17938,N_11007,N_10179);
nand U17939 (N_17939,N_12594,N_12620);
and U17940 (N_17940,N_12313,N_14457);
and U17941 (N_17941,N_12857,N_12425);
nand U17942 (N_17942,N_10538,N_10731);
and U17943 (N_17943,N_13563,N_13965);
nor U17944 (N_17944,N_13501,N_14650);
and U17945 (N_17945,N_11530,N_14524);
nand U17946 (N_17946,N_11439,N_13209);
nor U17947 (N_17947,N_12491,N_11026);
xnor U17948 (N_17948,N_12272,N_11815);
and U17949 (N_17949,N_13700,N_12333);
nand U17950 (N_17950,N_13018,N_11327);
and U17951 (N_17951,N_11055,N_13345);
and U17952 (N_17952,N_10614,N_12579);
and U17953 (N_17953,N_12865,N_13478);
and U17954 (N_17954,N_11609,N_12167);
and U17955 (N_17955,N_13480,N_14932);
xor U17956 (N_17956,N_11343,N_13199);
nor U17957 (N_17957,N_14290,N_13412);
or U17958 (N_17958,N_12927,N_13973);
xor U17959 (N_17959,N_11922,N_13050);
and U17960 (N_17960,N_14712,N_11224);
nor U17961 (N_17961,N_11297,N_13796);
and U17962 (N_17962,N_14219,N_13744);
nor U17963 (N_17963,N_13868,N_14002);
nand U17964 (N_17964,N_12228,N_14648);
nand U17965 (N_17965,N_10346,N_13148);
or U17966 (N_17966,N_14109,N_12863);
nand U17967 (N_17967,N_11038,N_12591);
and U17968 (N_17968,N_10563,N_11039);
nand U17969 (N_17969,N_11466,N_13186);
and U17970 (N_17970,N_14877,N_14296);
nor U17971 (N_17971,N_10736,N_14101);
nor U17972 (N_17972,N_11775,N_12308);
nor U17973 (N_17973,N_10236,N_12001);
nor U17974 (N_17974,N_12263,N_14392);
nor U17975 (N_17975,N_12950,N_10717);
nor U17976 (N_17976,N_12734,N_10961);
nor U17977 (N_17977,N_10327,N_11575);
nor U17978 (N_17978,N_13957,N_13855);
xor U17979 (N_17979,N_13356,N_12319);
nand U17980 (N_17980,N_12799,N_10278);
nor U17981 (N_17981,N_14022,N_12659);
xnor U17982 (N_17982,N_14648,N_10199);
nand U17983 (N_17983,N_12506,N_14614);
nor U17984 (N_17984,N_14803,N_14359);
xor U17985 (N_17985,N_12110,N_10860);
nor U17986 (N_17986,N_12841,N_11275);
nor U17987 (N_17987,N_14916,N_13004);
nor U17988 (N_17988,N_13945,N_14003);
and U17989 (N_17989,N_10894,N_13773);
and U17990 (N_17990,N_14168,N_11532);
nor U17991 (N_17991,N_13505,N_13977);
or U17992 (N_17992,N_13864,N_12396);
and U17993 (N_17993,N_13131,N_13723);
nand U17994 (N_17994,N_12560,N_11368);
nand U17995 (N_17995,N_11262,N_11535);
or U17996 (N_17996,N_14603,N_11653);
and U17997 (N_17997,N_10253,N_10864);
and U17998 (N_17998,N_11843,N_14653);
and U17999 (N_17999,N_14694,N_13675);
nand U18000 (N_18000,N_12478,N_10042);
and U18001 (N_18001,N_14862,N_10829);
nor U18002 (N_18002,N_13584,N_14768);
nor U18003 (N_18003,N_12953,N_10620);
and U18004 (N_18004,N_13599,N_11798);
or U18005 (N_18005,N_14531,N_13110);
and U18006 (N_18006,N_14290,N_11115);
or U18007 (N_18007,N_14152,N_12695);
nand U18008 (N_18008,N_11156,N_13831);
and U18009 (N_18009,N_11596,N_13442);
xnor U18010 (N_18010,N_14032,N_12864);
nand U18011 (N_18011,N_10904,N_13587);
or U18012 (N_18012,N_13996,N_14496);
nor U18013 (N_18013,N_13483,N_11505);
and U18014 (N_18014,N_14602,N_11438);
nor U18015 (N_18015,N_12524,N_11982);
and U18016 (N_18016,N_10154,N_11455);
xnor U18017 (N_18017,N_13744,N_14791);
nor U18018 (N_18018,N_10985,N_14002);
nor U18019 (N_18019,N_10218,N_12426);
nand U18020 (N_18020,N_12524,N_11980);
and U18021 (N_18021,N_13140,N_10764);
and U18022 (N_18022,N_11752,N_13604);
nand U18023 (N_18023,N_14053,N_12222);
nand U18024 (N_18024,N_13536,N_12483);
or U18025 (N_18025,N_10117,N_12181);
xor U18026 (N_18026,N_11751,N_10683);
or U18027 (N_18027,N_11897,N_14683);
and U18028 (N_18028,N_11262,N_14663);
or U18029 (N_18029,N_12247,N_14309);
and U18030 (N_18030,N_12741,N_10591);
xor U18031 (N_18031,N_11471,N_12332);
and U18032 (N_18032,N_11700,N_10417);
nor U18033 (N_18033,N_12222,N_11090);
nand U18034 (N_18034,N_13113,N_12206);
and U18035 (N_18035,N_13934,N_11925);
nand U18036 (N_18036,N_13517,N_13655);
or U18037 (N_18037,N_11324,N_11867);
nand U18038 (N_18038,N_14915,N_10676);
or U18039 (N_18039,N_10677,N_10708);
xor U18040 (N_18040,N_11138,N_14455);
and U18041 (N_18041,N_14596,N_14680);
nor U18042 (N_18042,N_14917,N_13705);
and U18043 (N_18043,N_14468,N_13955);
and U18044 (N_18044,N_11838,N_11092);
or U18045 (N_18045,N_11880,N_14872);
nor U18046 (N_18046,N_13670,N_11062);
nor U18047 (N_18047,N_13457,N_14338);
or U18048 (N_18048,N_12862,N_12534);
nor U18049 (N_18049,N_13972,N_13555);
or U18050 (N_18050,N_10776,N_14468);
and U18051 (N_18051,N_13342,N_14706);
and U18052 (N_18052,N_11995,N_11233);
nor U18053 (N_18053,N_12502,N_11376);
nand U18054 (N_18054,N_11409,N_10689);
or U18055 (N_18055,N_14577,N_10819);
nand U18056 (N_18056,N_14550,N_11679);
and U18057 (N_18057,N_11549,N_14672);
nand U18058 (N_18058,N_11445,N_12422);
or U18059 (N_18059,N_11095,N_11713);
or U18060 (N_18060,N_12103,N_10831);
nand U18061 (N_18061,N_11918,N_10305);
nand U18062 (N_18062,N_13024,N_13306);
nor U18063 (N_18063,N_12458,N_12394);
nor U18064 (N_18064,N_13069,N_12179);
xor U18065 (N_18065,N_14062,N_10648);
or U18066 (N_18066,N_10505,N_12000);
or U18067 (N_18067,N_13016,N_13023);
nand U18068 (N_18068,N_12264,N_10756);
nor U18069 (N_18069,N_14656,N_12295);
nand U18070 (N_18070,N_14245,N_13081);
or U18071 (N_18071,N_10910,N_12144);
nor U18072 (N_18072,N_11262,N_12092);
or U18073 (N_18073,N_12355,N_13200);
nor U18074 (N_18074,N_12937,N_10634);
or U18075 (N_18075,N_12973,N_13879);
or U18076 (N_18076,N_10793,N_14465);
or U18077 (N_18077,N_10762,N_13737);
or U18078 (N_18078,N_13501,N_13212);
or U18079 (N_18079,N_10702,N_12589);
nor U18080 (N_18080,N_12068,N_14193);
nand U18081 (N_18081,N_14159,N_13537);
xnor U18082 (N_18082,N_12365,N_14641);
and U18083 (N_18083,N_13078,N_12323);
and U18084 (N_18084,N_11321,N_12585);
nor U18085 (N_18085,N_13541,N_10987);
xor U18086 (N_18086,N_10841,N_14335);
nor U18087 (N_18087,N_10431,N_10947);
or U18088 (N_18088,N_14271,N_14452);
or U18089 (N_18089,N_13129,N_14380);
or U18090 (N_18090,N_12500,N_11145);
and U18091 (N_18091,N_12157,N_10791);
nand U18092 (N_18092,N_12413,N_14982);
or U18093 (N_18093,N_12391,N_10420);
nor U18094 (N_18094,N_11266,N_11570);
nor U18095 (N_18095,N_10794,N_11421);
nor U18096 (N_18096,N_13004,N_13148);
nand U18097 (N_18097,N_13624,N_12227);
nand U18098 (N_18098,N_13986,N_11463);
nor U18099 (N_18099,N_10125,N_14641);
and U18100 (N_18100,N_14757,N_13864);
nor U18101 (N_18101,N_14761,N_14604);
or U18102 (N_18102,N_10418,N_14890);
xor U18103 (N_18103,N_14733,N_11895);
nor U18104 (N_18104,N_12998,N_10470);
or U18105 (N_18105,N_10870,N_11135);
xor U18106 (N_18106,N_10468,N_14823);
or U18107 (N_18107,N_13248,N_11850);
xnor U18108 (N_18108,N_14767,N_14441);
nor U18109 (N_18109,N_10116,N_11442);
nand U18110 (N_18110,N_13396,N_13149);
or U18111 (N_18111,N_11880,N_14198);
xor U18112 (N_18112,N_14375,N_10970);
nor U18113 (N_18113,N_14541,N_13537);
or U18114 (N_18114,N_13737,N_11050);
and U18115 (N_18115,N_11201,N_10476);
and U18116 (N_18116,N_12691,N_13046);
or U18117 (N_18117,N_11695,N_11462);
nor U18118 (N_18118,N_14201,N_10129);
or U18119 (N_18119,N_10246,N_14421);
nand U18120 (N_18120,N_10720,N_13376);
nand U18121 (N_18121,N_12193,N_14463);
or U18122 (N_18122,N_14973,N_14751);
or U18123 (N_18123,N_11735,N_11437);
nand U18124 (N_18124,N_10614,N_14621);
nand U18125 (N_18125,N_12943,N_11662);
nor U18126 (N_18126,N_10896,N_14513);
nand U18127 (N_18127,N_13171,N_10761);
xor U18128 (N_18128,N_11643,N_10257);
xnor U18129 (N_18129,N_13763,N_11086);
nand U18130 (N_18130,N_11350,N_13149);
nor U18131 (N_18131,N_10388,N_12650);
xnor U18132 (N_18132,N_13856,N_13718);
xnor U18133 (N_18133,N_10047,N_12537);
nor U18134 (N_18134,N_12786,N_11841);
nor U18135 (N_18135,N_13742,N_12541);
xor U18136 (N_18136,N_12126,N_14808);
or U18137 (N_18137,N_14781,N_13328);
or U18138 (N_18138,N_12881,N_12128);
or U18139 (N_18139,N_10806,N_13010);
and U18140 (N_18140,N_11755,N_14534);
nor U18141 (N_18141,N_11774,N_12965);
and U18142 (N_18142,N_12752,N_13903);
nor U18143 (N_18143,N_11477,N_14769);
nor U18144 (N_18144,N_11962,N_10916);
nor U18145 (N_18145,N_11500,N_10100);
xnor U18146 (N_18146,N_11607,N_12352);
and U18147 (N_18147,N_13698,N_12065);
or U18148 (N_18148,N_10228,N_14167);
and U18149 (N_18149,N_13078,N_14209);
and U18150 (N_18150,N_11562,N_12419);
nand U18151 (N_18151,N_11203,N_10426);
nor U18152 (N_18152,N_14668,N_11137);
and U18153 (N_18153,N_13657,N_12632);
xnor U18154 (N_18154,N_14452,N_13313);
nand U18155 (N_18155,N_14896,N_10020);
or U18156 (N_18156,N_11363,N_14235);
nand U18157 (N_18157,N_13715,N_10603);
nand U18158 (N_18158,N_10730,N_11015);
or U18159 (N_18159,N_12522,N_10363);
and U18160 (N_18160,N_10775,N_11769);
and U18161 (N_18161,N_12959,N_10084);
and U18162 (N_18162,N_13844,N_13519);
nor U18163 (N_18163,N_14635,N_13901);
or U18164 (N_18164,N_12125,N_12001);
nand U18165 (N_18165,N_11244,N_14987);
nor U18166 (N_18166,N_10479,N_13762);
or U18167 (N_18167,N_13845,N_12533);
nor U18168 (N_18168,N_11277,N_14781);
or U18169 (N_18169,N_10889,N_13581);
nand U18170 (N_18170,N_12343,N_12002);
nand U18171 (N_18171,N_12834,N_13505);
nand U18172 (N_18172,N_11950,N_13524);
nand U18173 (N_18173,N_12486,N_13076);
and U18174 (N_18174,N_13614,N_10268);
and U18175 (N_18175,N_12996,N_10099);
and U18176 (N_18176,N_12481,N_11684);
or U18177 (N_18177,N_10780,N_14779);
nand U18178 (N_18178,N_14007,N_11577);
nand U18179 (N_18179,N_10281,N_14201);
xnor U18180 (N_18180,N_14873,N_12712);
nand U18181 (N_18181,N_13950,N_11370);
or U18182 (N_18182,N_12198,N_14435);
xor U18183 (N_18183,N_11584,N_14417);
or U18184 (N_18184,N_12110,N_10600);
and U18185 (N_18185,N_10503,N_13322);
nand U18186 (N_18186,N_13588,N_14008);
or U18187 (N_18187,N_13398,N_14459);
nor U18188 (N_18188,N_13932,N_11404);
or U18189 (N_18189,N_13880,N_13493);
nor U18190 (N_18190,N_14565,N_11126);
xnor U18191 (N_18191,N_13419,N_12787);
or U18192 (N_18192,N_11132,N_10035);
or U18193 (N_18193,N_13329,N_13688);
nand U18194 (N_18194,N_10477,N_13788);
and U18195 (N_18195,N_11391,N_13925);
and U18196 (N_18196,N_12666,N_14585);
or U18197 (N_18197,N_12630,N_13557);
and U18198 (N_18198,N_14655,N_11624);
nor U18199 (N_18199,N_14650,N_13378);
and U18200 (N_18200,N_13235,N_13682);
nand U18201 (N_18201,N_12537,N_12734);
and U18202 (N_18202,N_13567,N_11899);
nor U18203 (N_18203,N_12332,N_12823);
and U18204 (N_18204,N_12083,N_10212);
nand U18205 (N_18205,N_13190,N_10936);
nand U18206 (N_18206,N_13609,N_14693);
nor U18207 (N_18207,N_13114,N_10324);
nand U18208 (N_18208,N_10058,N_11109);
or U18209 (N_18209,N_10845,N_11945);
nand U18210 (N_18210,N_10167,N_14361);
nand U18211 (N_18211,N_13344,N_11074);
nand U18212 (N_18212,N_11438,N_14604);
nor U18213 (N_18213,N_11651,N_10548);
or U18214 (N_18214,N_10254,N_10434);
nor U18215 (N_18215,N_11715,N_10457);
nand U18216 (N_18216,N_11737,N_10732);
nand U18217 (N_18217,N_11549,N_10380);
and U18218 (N_18218,N_14025,N_14300);
or U18219 (N_18219,N_10495,N_10977);
and U18220 (N_18220,N_10366,N_12757);
or U18221 (N_18221,N_12317,N_12662);
nand U18222 (N_18222,N_11186,N_14890);
and U18223 (N_18223,N_10404,N_11402);
nor U18224 (N_18224,N_13471,N_11750);
nor U18225 (N_18225,N_10980,N_11028);
or U18226 (N_18226,N_14910,N_12648);
and U18227 (N_18227,N_12050,N_10138);
nand U18228 (N_18228,N_14706,N_11608);
or U18229 (N_18229,N_10747,N_14905);
nor U18230 (N_18230,N_12646,N_12773);
nor U18231 (N_18231,N_13817,N_12600);
and U18232 (N_18232,N_10864,N_14643);
nand U18233 (N_18233,N_13441,N_11562);
nor U18234 (N_18234,N_12221,N_14307);
nand U18235 (N_18235,N_10619,N_14112);
and U18236 (N_18236,N_11466,N_10722);
nor U18237 (N_18237,N_11392,N_10106);
nand U18238 (N_18238,N_13628,N_11891);
and U18239 (N_18239,N_10335,N_13890);
xnor U18240 (N_18240,N_10882,N_12665);
and U18241 (N_18241,N_10819,N_14325);
nand U18242 (N_18242,N_14216,N_14443);
nor U18243 (N_18243,N_14623,N_13764);
or U18244 (N_18244,N_13645,N_11061);
nor U18245 (N_18245,N_10566,N_11093);
and U18246 (N_18246,N_11654,N_10468);
or U18247 (N_18247,N_10149,N_10988);
nand U18248 (N_18248,N_10980,N_12992);
nor U18249 (N_18249,N_11211,N_10354);
nand U18250 (N_18250,N_13660,N_11885);
nor U18251 (N_18251,N_11012,N_10982);
nand U18252 (N_18252,N_11170,N_14031);
nor U18253 (N_18253,N_12355,N_14307);
or U18254 (N_18254,N_13595,N_12902);
nand U18255 (N_18255,N_10278,N_14374);
xor U18256 (N_18256,N_13235,N_11811);
nor U18257 (N_18257,N_14730,N_13406);
nand U18258 (N_18258,N_13948,N_12275);
nand U18259 (N_18259,N_14113,N_13148);
nand U18260 (N_18260,N_10256,N_12684);
and U18261 (N_18261,N_12602,N_14594);
nor U18262 (N_18262,N_10119,N_10219);
or U18263 (N_18263,N_13908,N_12341);
nor U18264 (N_18264,N_13670,N_10842);
and U18265 (N_18265,N_13080,N_14962);
xnor U18266 (N_18266,N_12326,N_12830);
xnor U18267 (N_18267,N_11817,N_11007);
and U18268 (N_18268,N_13865,N_13351);
or U18269 (N_18269,N_12635,N_13478);
nand U18270 (N_18270,N_12116,N_14253);
or U18271 (N_18271,N_12746,N_13548);
nand U18272 (N_18272,N_12555,N_12232);
and U18273 (N_18273,N_12791,N_14952);
nor U18274 (N_18274,N_11843,N_13814);
or U18275 (N_18275,N_13058,N_10999);
nand U18276 (N_18276,N_10954,N_13501);
or U18277 (N_18277,N_14310,N_11244);
nor U18278 (N_18278,N_14589,N_12614);
nand U18279 (N_18279,N_12263,N_12732);
nor U18280 (N_18280,N_14965,N_12302);
nor U18281 (N_18281,N_14995,N_11218);
xnor U18282 (N_18282,N_14266,N_14899);
or U18283 (N_18283,N_14681,N_11254);
or U18284 (N_18284,N_11876,N_10215);
and U18285 (N_18285,N_14794,N_11777);
nand U18286 (N_18286,N_10117,N_14800);
nor U18287 (N_18287,N_10103,N_14381);
or U18288 (N_18288,N_14117,N_12954);
nor U18289 (N_18289,N_14238,N_10986);
xnor U18290 (N_18290,N_14933,N_13852);
and U18291 (N_18291,N_14529,N_14892);
xor U18292 (N_18292,N_11348,N_14064);
and U18293 (N_18293,N_14881,N_13235);
and U18294 (N_18294,N_10418,N_11911);
and U18295 (N_18295,N_11468,N_12572);
nor U18296 (N_18296,N_13591,N_14588);
nand U18297 (N_18297,N_10867,N_10089);
xnor U18298 (N_18298,N_14719,N_10829);
or U18299 (N_18299,N_13068,N_14944);
nor U18300 (N_18300,N_13901,N_13561);
and U18301 (N_18301,N_12252,N_10994);
nor U18302 (N_18302,N_12713,N_14723);
and U18303 (N_18303,N_11669,N_11824);
or U18304 (N_18304,N_13279,N_11429);
and U18305 (N_18305,N_10908,N_12837);
nor U18306 (N_18306,N_14651,N_10902);
and U18307 (N_18307,N_10020,N_10884);
nand U18308 (N_18308,N_14023,N_14621);
or U18309 (N_18309,N_11891,N_10213);
nor U18310 (N_18310,N_13518,N_13440);
nor U18311 (N_18311,N_11882,N_10767);
or U18312 (N_18312,N_14826,N_12227);
and U18313 (N_18313,N_14198,N_10826);
and U18314 (N_18314,N_13604,N_10066);
nor U18315 (N_18315,N_12534,N_11474);
xor U18316 (N_18316,N_10208,N_14520);
nand U18317 (N_18317,N_13063,N_10149);
nand U18318 (N_18318,N_10515,N_12921);
nand U18319 (N_18319,N_10650,N_10740);
nand U18320 (N_18320,N_12162,N_11834);
xnor U18321 (N_18321,N_13904,N_13224);
nor U18322 (N_18322,N_10314,N_10393);
and U18323 (N_18323,N_10805,N_10018);
xnor U18324 (N_18324,N_13518,N_14726);
and U18325 (N_18325,N_11966,N_14461);
nand U18326 (N_18326,N_10073,N_11201);
nor U18327 (N_18327,N_13384,N_11451);
nor U18328 (N_18328,N_13619,N_11537);
xor U18329 (N_18329,N_11969,N_11800);
or U18330 (N_18330,N_12396,N_13904);
and U18331 (N_18331,N_10580,N_10317);
or U18332 (N_18332,N_10935,N_11243);
nand U18333 (N_18333,N_10269,N_13388);
and U18334 (N_18334,N_10018,N_11734);
xor U18335 (N_18335,N_14898,N_13562);
nand U18336 (N_18336,N_12585,N_11717);
nor U18337 (N_18337,N_11683,N_14418);
and U18338 (N_18338,N_12981,N_13530);
nor U18339 (N_18339,N_12793,N_14311);
xnor U18340 (N_18340,N_11200,N_10436);
nand U18341 (N_18341,N_11976,N_12071);
nand U18342 (N_18342,N_13984,N_13162);
xnor U18343 (N_18343,N_13143,N_12238);
nand U18344 (N_18344,N_11304,N_10256);
or U18345 (N_18345,N_11384,N_10584);
nor U18346 (N_18346,N_14901,N_13878);
nor U18347 (N_18347,N_10903,N_10609);
and U18348 (N_18348,N_12660,N_13247);
nand U18349 (N_18349,N_12386,N_13997);
and U18350 (N_18350,N_10071,N_10773);
nor U18351 (N_18351,N_12877,N_14220);
or U18352 (N_18352,N_12015,N_10415);
nor U18353 (N_18353,N_11234,N_12901);
nor U18354 (N_18354,N_14765,N_13153);
nand U18355 (N_18355,N_13812,N_13939);
or U18356 (N_18356,N_13983,N_13362);
nand U18357 (N_18357,N_10969,N_14993);
and U18358 (N_18358,N_10805,N_13049);
nor U18359 (N_18359,N_11969,N_13546);
xor U18360 (N_18360,N_11891,N_14885);
and U18361 (N_18361,N_14237,N_13056);
nand U18362 (N_18362,N_10274,N_10657);
and U18363 (N_18363,N_10498,N_14422);
or U18364 (N_18364,N_11433,N_13003);
and U18365 (N_18365,N_12068,N_10069);
xor U18366 (N_18366,N_13460,N_11701);
and U18367 (N_18367,N_13998,N_12221);
nor U18368 (N_18368,N_13221,N_10620);
xnor U18369 (N_18369,N_11936,N_14599);
xor U18370 (N_18370,N_14827,N_12437);
or U18371 (N_18371,N_13282,N_13437);
nor U18372 (N_18372,N_10373,N_14497);
and U18373 (N_18373,N_10469,N_11804);
nor U18374 (N_18374,N_11072,N_14654);
or U18375 (N_18375,N_12326,N_10344);
nor U18376 (N_18376,N_10611,N_11085);
nor U18377 (N_18377,N_12776,N_11674);
and U18378 (N_18378,N_13157,N_11229);
nor U18379 (N_18379,N_12811,N_13453);
and U18380 (N_18380,N_10593,N_11912);
or U18381 (N_18381,N_11840,N_11102);
and U18382 (N_18382,N_11885,N_13198);
or U18383 (N_18383,N_10756,N_10142);
nand U18384 (N_18384,N_12496,N_13457);
nand U18385 (N_18385,N_12369,N_14973);
nand U18386 (N_18386,N_12803,N_10658);
and U18387 (N_18387,N_11822,N_14450);
or U18388 (N_18388,N_11949,N_12481);
and U18389 (N_18389,N_14322,N_10891);
or U18390 (N_18390,N_13736,N_11171);
xnor U18391 (N_18391,N_14601,N_10290);
and U18392 (N_18392,N_13280,N_11444);
or U18393 (N_18393,N_14296,N_10988);
or U18394 (N_18394,N_13332,N_11549);
or U18395 (N_18395,N_13634,N_12756);
or U18396 (N_18396,N_12738,N_11179);
nor U18397 (N_18397,N_12871,N_10539);
nand U18398 (N_18398,N_11325,N_10244);
nand U18399 (N_18399,N_13001,N_12494);
nor U18400 (N_18400,N_14093,N_11978);
or U18401 (N_18401,N_12864,N_12583);
nor U18402 (N_18402,N_14832,N_10810);
nand U18403 (N_18403,N_14902,N_12146);
nor U18404 (N_18404,N_14479,N_13490);
and U18405 (N_18405,N_14010,N_10227);
or U18406 (N_18406,N_11721,N_14550);
and U18407 (N_18407,N_14798,N_13215);
nor U18408 (N_18408,N_12280,N_13305);
nor U18409 (N_18409,N_14209,N_10554);
xor U18410 (N_18410,N_13919,N_11901);
xnor U18411 (N_18411,N_11725,N_10293);
or U18412 (N_18412,N_11345,N_10067);
nand U18413 (N_18413,N_14049,N_14439);
and U18414 (N_18414,N_14968,N_13922);
and U18415 (N_18415,N_14954,N_10214);
xnor U18416 (N_18416,N_13052,N_11168);
nand U18417 (N_18417,N_11895,N_12731);
or U18418 (N_18418,N_11626,N_14972);
xnor U18419 (N_18419,N_10374,N_14660);
nand U18420 (N_18420,N_10692,N_11536);
nand U18421 (N_18421,N_12822,N_13520);
and U18422 (N_18422,N_13209,N_11164);
or U18423 (N_18423,N_13366,N_12124);
nand U18424 (N_18424,N_14936,N_13651);
or U18425 (N_18425,N_10092,N_14500);
or U18426 (N_18426,N_14808,N_14805);
and U18427 (N_18427,N_12739,N_10723);
and U18428 (N_18428,N_11235,N_13046);
nand U18429 (N_18429,N_14174,N_11501);
and U18430 (N_18430,N_10463,N_12119);
nand U18431 (N_18431,N_13830,N_14619);
and U18432 (N_18432,N_13874,N_14482);
and U18433 (N_18433,N_12414,N_11841);
and U18434 (N_18434,N_13123,N_11442);
nor U18435 (N_18435,N_14984,N_10719);
nor U18436 (N_18436,N_10360,N_10136);
and U18437 (N_18437,N_13251,N_11206);
and U18438 (N_18438,N_14257,N_14358);
nor U18439 (N_18439,N_14888,N_14179);
xor U18440 (N_18440,N_12839,N_13962);
and U18441 (N_18441,N_11985,N_13502);
nor U18442 (N_18442,N_10535,N_12080);
or U18443 (N_18443,N_11550,N_13549);
xor U18444 (N_18444,N_12865,N_10538);
nand U18445 (N_18445,N_13838,N_10557);
xor U18446 (N_18446,N_14590,N_12699);
nor U18447 (N_18447,N_13450,N_10263);
nand U18448 (N_18448,N_14553,N_11510);
and U18449 (N_18449,N_12951,N_12735);
nand U18450 (N_18450,N_11213,N_10698);
or U18451 (N_18451,N_13212,N_13923);
nor U18452 (N_18452,N_12631,N_12388);
nor U18453 (N_18453,N_12656,N_14126);
or U18454 (N_18454,N_12618,N_11952);
and U18455 (N_18455,N_10202,N_12435);
nor U18456 (N_18456,N_12083,N_14189);
or U18457 (N_18457,N_14125,N_14470);
and U18458 (N_18458,N_14038,N_10686);
and U18459 (N_18459,N_14926,N_14702);
and U18460 (N_18460,N_13281,N_14428);
and U18461 (N_18461,N_13840,N_11380);
or U18462 (N_18462,N_11790,N_12998);
nor U18463 (N_18463,N_10443,N_11303);
and U18464 (N_18464,N_10548,N_11013);
and U18465 (N_18465,N_10588,N_12740);
and U18466 (N_18466,N_11646,N_10665);
nor U18467 (N_18467,N_13292,N_11901);
xor U18468 (N_18468,N_10743,N_11056);
nand U18469 (N_18469,N_13961,N_10080);
xnor U18470 (N_18470,N_10614,N_12834);
or U18471 (N_18471,N_12526,N_13183);
or U18472 (N_18472,N_12438,N_13761);
and U18473 (N_18473,N_13653,N_14201);
nand U18474 (N_18474,N_10169,N_14581);
and U18475 (N_18475,N_12108,N_11013);
nor U18476 (N_18476,N_14607,N_11864);
nor U18477 (N_18477,N_10121,N_12105);
nand U18478 (N_18478,N_11611,N_10784);
nand U18479 (N_18479,N_12953,N_13803);
or U18480 (N_18480,N_13789,N_14164);
and U18481 (N_18481,N_12912,N_11202);
xnor U18482 (N_18482,N_11508,N_13456);
and U18483 (N_18483,N_14217,N_14694);
and U18484 (N_18484,N_11353,N_14003);
and U18485 (N_18485,N_12932,N_11130);
and U18486 (N_18486,N_14359,N_13190);
nand U18487 (N_18487,N_11810,N_12507);
nand U18488 (N_18488,N_12318,N_11661);
and U18489 (N_18489,N_13448,N_11538);
nand U18490 (N_18490,N_10751,N_14658);
xnor U18491 (N_18491,N_13888,N_11688);
nor U18492 (N_18492,N_14836,N_12658);
nor U18493 (N_18493,N_14307,N_13772);
nor U18494 (N_18494,N_12410,N_12716);
or U18495 (N_18495,N_10293,N_14338);
xor U18496 (N_18496,N_10180,N_13171);
or U18497 (N_18497,N_12786,N_10837);
or U18498 (N_18498,N_11740,N_12798);
and U18499 (N_18499,N_11178,N_13698);
nand U18500 (N_18500,N_11196,N_13994);
or U18501 (N_18501,N_10685,N_11696);
nor U18502 (N_18502,N_12838,N_11055);
nand U18503 (N_18503,N_11288,N_12945);
nor U18504 (N_18504,N_14901,N_10799);
nor U18505 (N_18505,N_10736,N_14002);
nor U18506 (N_18506,N_12546,N_13496);
and U18507 (N_18507,N_11868,N_12466);
xor U18508 (N_18508,N_14849,N_11154);
or U18509 (N_18509,N_14121,N_11898);
nand U18510 (N_18510,N_10885,N_12993);
and U18511 (N_18511,N_12703,N_13562);
nor U18512 (N_18512,N_14790,N_14554);
or U18513 (N_18513,N_10098,N_12549);
and U18514 (N_18514,N_14598,N_14486);
or U18515 (N_18515,N_12632,N_11367);
or U18516 (N_18516,N_13181,N_11555);
or U18517 (N_18517,N_13309,N_14599);
xnor U18518 (N_18518,N_12365,N_14080);
nor U18519 (N_18519,N_10008,N_11579);
nand U18520 (N_18520,N_14007,N_10272);
nor U18521 (N_18521,N_14920,N_13929);
nand U18522 (N_18522,N_12755,N_14772);
nor U18523 (N_18523,N_10718,N_13213);
xor U18524 (N_18524,N_11249,N_13082);
nand U18525 (N_18525,N_12645,N_11422);
or U18526 (N_18526,N_14048,N_13440);
nor U18527 (N_18527,N_11300,N_10624);
nor U18528 (N_18528,N_11245,N_14216);
nor U18529 (N_18529,N_14509,N_11078);
or U18530 (N_18530,N_12949,N_13506);
nor U18531 (N_18531,N_12476,N_14705);
xor U18532 (N_18532,N_13444,N_11175);
nand U18533 (N_18533,N_11549,N_11827);
or U18534 (N_18534,N_11411,N_11889);
and U18535 (N_18535,N_12396,N_10592);
nand U18536 (N_18536,N_11692,N_13421);
nor U18537 (N_18537,N_11057,N_14419);
or U18538 (N_18538,N_14943,N_11577);
and U18539 (N_18539,N_12181,N_13223);
nor U18540 (N_18540,N_13144,N_11704);
or U18541 (N_18541,N_12469,N_13365);
nand U18542 (N_18542,N_14225,N_12972);
xnor U18543 (N_18543,N_14777,N_13114);
nand U18544 (N_18544,N_12232,N_14955);
and U18545 (N_18545,N_11594,N_11588);
nand U18546 (N_18546,N_12654,N_14595);
nor U18547 (N_18547,N_14466,N_12860);
and U18548 (N_18548,N_12836,N_13088);
nor U18549 (N_18549,N_13238,N_10550);
xor U18550 (N_18550,N_12501,N_10770);
and U18551 (N_18551,N_10333,N_13158);
nor U18552 (N_18552,N_14183,N_11801);
and U18553 (N_18553,N_14604,N_13313);
and U18554 (N_18554,N_12496,N_12754);
nor U18555 (N_18555,N_13014,N_10950);
and U18556 (N_18556,N_10739,N_14447);
or U18557 (N_18557,N_13025,N_11438);
or U18558 (N_18558,N_10674,N_11001);
nor U18559 (N_18559,N_11110,N_12398);
nor U18560 (N_18560,N_12210,N_13703);
or U18561 (N_18561,N_13340,N_12794);
nor U18562 (N_18562,N_10145,N_14681);
and U18563 (N_18563,N_11184,N_10476);
and U18564 (N_18564,N_10604,N_14621);
and U18565 (N_18565,N_14791,N_14889);
and U18566 (N_18566,N_10970,N_10416);
nor U18567 (N_18567,N_10509,N_11988);
and U18568 (N_18568,N_10719,N_10651);
nor U18569 (N_18569,N_10983,N_14364);
and U18570 (N_18570,N_11635,N_11458);
and U18571 (N_18571,N_10601,N_13681);
xor U18572 (N_18572,N_12891,N_14308);
nor U18573 (N_18573,N_11699,N_10120);
and U18574 (N_18574,N_12306,N_13327);
or U18575 (N_18575,N_13123,N_10745);
nor U18576 (N_18576,N_13918,N_13411);
nand U18577 (N_18577,N_12004,N_14693);
and U18578 (N_18578,N_11842,N_10749);
nor U18579 (N_18579,N_12254,N_10145);
nand U18580 (N_18580,N_11232,N_12014);
nand U18581 (N_18581,N_11850,N_14682);
nand U18582 (N_18582,N_12734,N_11961);
nor U18583 (N_18583,N_14992,N_11382);
and U18584 (N_18584,N_11129,N_14914);
or U18585 (N_18585,N_11542,N_14025);
xor U18586 (N_18586,N_12810,N_14599);
and U18587 (N_18587,N_14465,N_12278);
and U18588 (N_18588,N_14708,N_13208);
nor U18589 (N_18589,N_12476,N_12222);
nor U18590 (N_18590,N_11127,N_13557);
nand U18591 (N_18591,N_13126,N_10240);
nand U18592 (N_18592,N_12758,N_10046);
nand U18593 (N_18593,N_14553,N_11801);
nor U18594 (N_18594,N_13399,N_13864);
and U18595 (N_18595,N_12152,N_13376);
nand U18596 (N_18596,N_10264,N_11596);
xor U18597 (N_18597,N_13655,N_10056);
xnor U18598 (N_18598,N_10138,N_14928);
nor U18599 (N_18599,N_10201,N_11159);
and U18600 (N_18600,N_13500,N_13631);
or U18601 (N_18601,N_10020,N_13732);
nand U18602 (N_18602,N_10760,N_12470);
and U18603 (N_18603,N_12147,N_14641);
nor U18604 (N_18604,N_10891,N_12179);
or U18605 (N_18605,N_13644,N_11260);
nor U18606 (N_18606,N_13632,N_10428);
xnor U18607 (N_18607,N_10875,N_14906);
nand U18608 (N_18608,N_10928,N_10285);
nor U18609 (N_18609,N_12508,N_13906);
or U18610 (N_18610,N_12417,N_11744);
or U18611 (N_18611,N_13302,N_14451);
nand U18612 (N_18612,N_13631,N_13446);
or U18613 (N_18613,N_12467,N_14426);
and U18614 (N_18614,N_10205,N_10355);
nand U18615 (N_18615,N_14669,N_12461);
and U18616 (N_18616,N_12699,N_13513);
or U18617 (N_18617,N_12423,N_12353);
or U18618 (N_18618,N_14529,N_10306);
nor U18619 (N_18619,N_10190,N_12300);
and U18620 (N_18620,N_13871,N_12866);
nor U18621 (N_18621,N_11339,N_10110);
or U18622 (N_18622,N_12272,N_13751);
nand U18623 (N_18623,N_11287,N_10566);
or U18624 (N_18624,N_12775,N_10978);
or U18625 (N_18625,N_14105,N_10341);
nor U18626 (N_18626,N_10547,N_13734);
and U18627 (N_18627,N_13717,N_10013);
nand U18628 (N_18628,N_14078,N_14267);
nand U18629 (N_18629,N_13136,N_11126);
nor U18630 (N_18630,N_13411,N_13795);
nor U18631 (N_18631,N_14546,N_13891);
or U18632 (N_18632,N_10667,N_10959);
nor U18633 (N_18633,N_14812,N_12808);
or U18634 (N_18634,N_13766,N_13889);
nor U18635 (N_18635,N_14415,N_11840);
nor U18636 (N_18636,N_13199,N_10161);
xor U18637 (N_18637,N_11797,N_13687);
nand U18638 (N_18638,N_11574,N_11391);
xor U18639 (N_18639,N_13080,N_12350);
and U18640 (N_18640,N_10502,N_11552);
or U18641 (N_18641,N_12315,N_14965);
and U18642 (N_18642,N_11646,N_13957);
nand U18643 (N_18643,N_12821,N_14039);
nand U18644 (N_18644,N_14825,N_11748);
nor U18645 (N_18645,N_10351,N_12292);
or U18646 (N_18646,N_10106,N_13599);
and U18647 (N_18647,N_10276,N_10694);
nor U18648 (N_18648,N_12185,N_13751);
and U18649 (N_18649,N_13266,N_11951);
nand U18650 (N_18650,N_12366,N_11606);
nand U18651 (N_18651,N_14325,N_12284);
nand U18652 (N_18652,N_12524,N_12886);
nor U18653 (N_18653,N_10493,N_12724);
or U18654 (N_18654,N_11743,N_11798);
nand U18655 (N_18655,N_10938,N_11306);
xnor U18656 (N_18656,N_14624,N_14910);
and U18657 (N_18657,N_13993,N_14747);
and U18658 (N_18658,N_12317,N_14942);
or U18659 (N_18659,N_12957,N_14259);
or U18660 (N_18660,N_12152,N_11326);
and U18661 (N_18661,N_10092,N_12112);
and U18662 (N_18662,N_13574,N_11085);
or U18663 (N_18663,N_11219,N_14614);
and U18664 (N_18664,N_14139,N_10828);
nand U18665 (N_18665,N_10343,N_14914);
xnor U18666 (N_18666,N_13590,N_10794);
nand U18667 (N_18667,N_14365,N_10075);
nand U18668 (N_18668,N_12460,N_11286);
and U18669 (N_18669,N_14103,N_13202);
and U18670 (N_18670,N_10052,N_12231);
nand U18671 (N_18671,N_11781,N_13288);
nand U18672 (N_18672,N_14250,N_14584);
and U18673 (N_18673,N_11945,N_12387);
or U18674 (N_18674,N_13360,N_11418);
nor U18675 (N_18675,N_10809,N_14802);
nor U18676 (N_18676,N_11725,N_12014);
or U18677 (N_18677,N_11087,N_11228);
nor U18678 (N_18678,N_14959,N_12800);
xnor U18679 (N_18679,N_11386,N_10617);
nor U18680 (N_18680,N_11293,N_13682);
and U18681 (N_18681,N_14307,N_10199);
nor U18682 (N_18682,N_10010,N_11446);
and U18683 (N_18683,N_12979,N_12314);
and U18684 (N_18684,N_10817,N_13940);
nand U18685 (N_18685,N_13377,N_13876);
and U18686 (N_18686,N_13888,N_12051);
nand U18687 (N_18687,N_14897,N_14964);
or U18688 (N_18688,N_10477,N_13979);
nor U18689 (N_18689,N_13119,N_14977);
nor U18690 (N_18690,N_12476,N_12984);
and U18691 (N_18691,N_13098,N_14588);
nand U18692 (N_18692,N_11958,N_13984);
nor U18693 (N_18693,N_13091,N_11674);
or U18694 (N_18694,N_13342,N_10964);
or U18695 (N_18695,N_14902,N_10959);
nand U18696 (N_18696,N_12988,N_10944);
nor U18697 (N_18697,N_13337,N_13321);
nand U18698 (N_18698,N_11676,N_12689);
or U18699 (N_18699,N_11560,N_13564);
or U18700 (N_18700,N_12016,N_11712);
and U18701 (N_18701,N_12302,N_14248);
and U18702 (N_18702,N_14877,N_11416);
and U18703 (N_18703,N_10745,N_11560);
nand U18704 (N_18704,N_13206,N_12751);
and U18705 (N_18705,N_12716,N_11885);
nand U18706 (N_18706,N_14790,N_12101);
and U18707 (N_18707,N_11946,N_14592);
or U18708 (N_18708,N_10636,N_10414);
nand U18709 (N_18709,N_13538,N_11623);
and U18710 (N_18710,N_12272,N_13342);
and U18711 (N_18711,N_13313,N_10361);
nor U18712 (N_18712,N_10194,N_13297);
xor U18713 (N_18713,N_11031,N_12102);
or U18714 (N_18714,N_11806,N_11475);
nand U18715 (N_18715,N_10854,N_14502);
nor U18716 (N_18716,N_14762,N_12260);
or U18717 (N_18717,N_10915,N_13900);
xnor U18718 (N_18718,N_12340,N_12776);
xor U18719 (N_18719,N_12993,N_13823);
and U18720 (N_18720,N_12062,N_12037);
or U18721 (N_18721,N_13588,N_13081);
xor U18722 (N_18722,N_14284,N_10488);
and U18723 (N_18723,N_10060,N_14274);
nand U18724 (N_18724,N_10476,N_10832);
nand U18725 (N_18725,N_13847,N_12346);
and U18726 (N_18726,N_14193,N_14683);
nor U18727 (N_18727,N_12809,N_14549);
nor U18728 (N_18728,N_13810,N_14040);
nand U18729 (N_18729,N_13381,N_12542);
nand U18730 (N_18730,N_10421,N_11362);
xnor U18731 (N_18731,N_11688,N_11842);
and U18732 (N_18732,N_11024,N_14564);
or U18733 (N_18733,N_11303,N_10347);
and U18734 (N_18734,N_10501,N_12149);
nand U18735 (N_18735,N_14808,N_11944);
and U18736 (N_18736,N_13039,N_12287);
nor U18737 (N_18737,N_12475,N_14658);
xor U18738 (N_18738,N_11058,N_12162);
xnor U18739 (N_18739,N_10517,N_12629);
and U18740 (N_18740,N_14072,N_13156);
nor U18741 (N_18741,N_14339,N_10911);
xnor U18742 (N_18742,N_11637,N_13258);
and U18743 (N_18743,N_13651,N_14202);
and U18744 (N_18744,N_12919,N_10278);
nand U18745 (N_18745,N_11362,N_13161);
and U18746 (N_18746,N_13135,N_11809);
xnor U18747 (N_18747,N_14296,N_12768);
nand U18748 (N_18748,N_10740,N_14731);
nor U18749 (N_18749,N_11271,N_10410);
nand U18750 (N_18750,N_10464,N_11891);
nand U18751 (N_18751,N_10795,N_11991);
nor U18752 (N_18752,N_11125,N_12657);
and U18753 (N_18753,N_10805,N_12017);
nor U18754 (N_18754,N_14899,N_10443);
or U18755 (N_18755,N_11496,N_14523);
nor U18756 (N_18756,N_14976,N_14349);
or U18757 (N_18757,N_11039,N_13545);
or U18758 (N_18758,N_10872,N_12563);
nand U18759 (N_18759,N_12100,N_14534);
nand U18760 (N_18760,N_14137,N_13210);
nand U18761 (N_18761,N_12690,N_11840);
and U18762 (N_18762,N_10313,N_14875);
and U18763 (N_18763,N_12783,N_12450);
or U18764 (N_18764,N_12613,N_10350);
nand U18765 (N_18765,N_13795,N_10993);
nor U18766 (N_18766,N_10894,N_10216);
xnor U18767 (N_18767,N_12696,N_11405);
nor U18768 (N_18768,N_13569,N_12258);
xor U18769 (N_18769,N_11086,N_12889);
xor U18770 (N_18770,N_10862,N_10767);
nand U18771 (N_18771,N_13117,N_12781);
and U18772 (N_18772,N_14615,N_11757);
and U18773 (N_18773,N_13431,N_14821);
nand U18774 (N_18774,N_13446,N_12673);
nand U18775 (N_18775,N_13051,N_10078);
nand U18776 (N_18776,N_12120,N_10641);
or U18777 (N_18777,N_12717,N_11589);
nand U18778 (N_18778,N_12424,N_12162);
and U18779 (N_18779,N_11633,N_13236);
or U18780 (N_18780,N_11476,N_10551);
or U18781 (N_18781,N_14530,N_10667);
and U18782 (N_18782,N_13051,N_10954);
and U18783 (N_18783,N_12286,N_10493);
xor U18784 (N_18784,N_12264,N_13670);
and U18785 (N_18785,N_14018,N_12051);
nand U18786 (N_18786,N_11339,N_12289);
nand U18787 (N_18787,N_12100,N_13921);
and U18788 (N_18788,N_11722,N_14197);
nor U18789 (N_18789,N_10753,N_13827);
xnor U18790 (N_18790,N_13468,N_11983);
nand U18791 (N_18791,N_14248,N_10463);
and U18792 (N_18792,N_10161,N_10465);
and U18793 (N_18793,N_14768,N_12376);
or U18794 (N_18794,N_10417,N_14141);
nor U18795 (N_18795,N_11607,N_14147);
or U18796 (N_18796,N_14214,N_11852);
nand U18797 (N_18797,N_13657,N_12501);
nand U18798 (N_18798,N_10300,N_12057);
nor U18799 (N_18799,N_13810,N_10046);
or U18800 (N_18800,N_14218,N_13270);
and U18801 (N_18801,N_12529,N_10942);
xor U18802 (N_18802,N_13116,N_14907);
and U18803 (N_18803,N_10093,N_11157);
nor U18804 (N_18804,N_10352,N_14616);
and U18805 (N_18805,N_13892,N_11060);
or U18806 (N_18806,N_12636,N_10217);
nand U18807 (N_18807,N_12334,N_10582);
nor U18808 (N_18808,N_11160,N_12115);
or U18809 (N_18809,N_14144,N_12680);
nor U18810 (N_18810,N_14705,N_10611);
nor U18811 (N_18811,N_12868,N_13046);
and U18812 (N_18812,N_13880,N_11696);
nor U18813 (N_18813,N_10190,N_10852);
nand U18814 (N_18814,N_10288,N_14688);
nand U18815 (N_18815,N_13076,N_13185);
or U18816 (N_18816,N_10116,N_14483);
or U18817 (N_18817,N_12822,N_14464);
nor U18818 (N_18818,N_10497,N_14367);
nor U18819 (N_18819,N_14823,N_14812);
nor U18820 (N_18820,N_14290,N_14678);
nand U18821 (N_18821,N_11255,N_13775);
nand U18822 (N_18822,N_12667,N_11571);
nand U18823 (N_18823,N_12890,N_12860);
nand U18824 (N_18824,N_12095,N_14729);
xor U18825 (N_18825,N_12807,N_10297);
xor U18826 (N_18826,N_14117,N_11671);
nand U18827 (N_18827,N_13115,N_11249);
nand U18828 (N_18828,N_12724,N_10859);
and U18829 (N_18829,N_12365,N_14634);
xnor U18830 (N_18830,N_11247,N_13706);
and U18831 (N_18831,N_10944,N_11264);
and U18832 (N_18832,N_13522,N_12529);
or U18833 (N_18833,N_13057,N_12838);
or U18834 (N_18834,N_11584,N_11897);
nor U18835 (N_18835,N_14053,N_11199);
nand U18836 (N_18836,N_10244,N_14437);
and U18837 (N_18837,N_14665,N_13003);
nand U18838 (N_18838,N_12171,N_13145);
xnor U18839 (N_18839,N_11826,N_13796);
nor U18840 (N_18840,N_14594,N_12042);
and U18841 (N_18841,N_13420,N_11382);
and U18842 (N_18842,N_12302,N_10241);
nand U18843 (N_18843,N_14779,N_14674);
xnor U18844 (N_18844,N_14248,N_10434);
nor U18845 (N_18845,N_12538,N_12007);
nor U18846 (N_18846,N_11173,N_12880);
nor U18847 (N_18847,N_11934,N_13626);
xnor U18848 (N_18848,N_14811,N_14434);
and U18849 (N_18849,N_13705,N_11884);
or U18850 (N_18850,N_11407,N_13166);
or U18851 (N_18851,N_14300,N_13161);
or U18852 (N_18852,N_13711,N_12714);
nor U18853 (N_18853,N_14232,N_12887);
xor U18854 (N_18854,N_13789,N_13700);
xor U18855 (N_18855,N_13807,N_14941);
and U18856 (N_18856,N_13909,N_14921);
or U18857 (N_18857,N_10822,N_14946);
xnor U18858 (N_18858,N_13978,N_12006);
nor U18859 (N_18859,N_14701,N_13233);
and U18860 (N_18860,N_14787,N_12313);
nor U18861 (N_18861,N_11701,N_14419);
and U18862 (N_18862,N_12869,N_11940);
or U18863 (N_18863,N_11808,N_14973);
or U18864 (N_18864,N_11215,N_12158);
nand U18865 (N_18865,N_10424,N_13122);
or U18866 (N_18866,N_13888,N_13843);
and U18867 (N_18867,N_14398,N_10755);
xnor U18868 (N_18868,N_12514,N_13796);
and U18869 (N_18869,N_13299,N_10429);
nor U18870 (N_18870,N_14607,N_13161);
and U18871 (N_18871,N_11792,N_14162);
or U18872 (N_18872,N_14716,N_11969);
nand U18873 (N_18873,N_11441,N_12061);
nor U18874 (N_18874,N_14220,N_12722);
and U18875 (N_18875,N_10341,N_10953);
nor U18876 (N_18876,N_12376,N_10691);
xor U18877 (N_18877,N_14950,N_11701);
nand U18878 (N_18878,N_12013,N_13607);
and U18879 (N_18879,N_10364,N_10733);
and U18880 (N_18880,N_11807,N_12677);
and U18881 (N_18881,N_12991,N_13069);
nor U18882 (N_18882,N_14800,N_12566);
nor U18883 (N_18883,N_11993,N_12442);
or U18884 (N_18884,N_14245,N_13064);
nor U18885 (N_18885,N_13959,N_12507);
xor U18886 (N_18886,N_10722,N_11498);
nor U18887 (N_18887,N_11253,N_13739);
or U18888 (N_18888,N_13921,N_10221);
nor U18889 (N_18889,N_12371,N_11248);
nor U18890 (N_18890,N_12218,N_10600);
nand U18891 (N_18891,N_13923,N_11458);
nor U18892 (N_18892,N_11615,N_12859);
or U18893 (N_18893,N_10049,N_12235);
or U18894 (N_18894,N_11365,N_13823);
nor U18895 (N_18895,N_14195,N_13892);
nand U18896 (N_18896,N_13421,N_10383);
nand U18897 (N_18897,N_14514,N_10002);
and U18898 (N_18898,N_14268,N_14994);
and U18899 (N_18899,N_11646,N_14290);
xnor U18900 (N_18900,N_12797,N_12806);
and U18901 (N_18901,N_10887,N_10909);
and U18902 (N_18902,N_14650,N_11594);
and U18903 (N_18903,N_12664,N_12639);
or U18904 (N_18904,N_10292,N_12635);
and U18905 (N_18905,N_11858,N_11075);
nand U18906 (N_18906,N_14664,N_14785);
nand U18907 (N_18907,N_10281,N_13978);
nand U18908 (N_18908,N_14418,N_14032);
and U18909 (N_18909,N_10168,N_13610);
and U18910 (N_18910,N_12206,N_14265);
and U18911 (N_18911,N_11742,N_14976);
or U18912 (N_18912,N_11595,N_12269);
nand U18913 (N_18913,N_12090,N_12906);
nor U18914 (N_18914,N_13731,N_13159);
and U18915 (N_18915,N_10714,N_12948);
and U18916 (N_18916,N_14366,N_10694);
and U18917 (N_18917,N_14579,N_12602);
nor U18918 (N_18918,N_13702,N_14137);
nor U18919 (N_18919,N_14686,N_12840);
and U18920 (N_18920,N_14219,N_11398);
and U18921 (N_18921,N_14022,N_13184);
nand U18922 (N_18922,N_13145,N_13181);
or U18923 (N_18923,N_13159,N_13328);
nand U18924 (N_18924,N_14903,N_14831);
and U18925 (N_18925,N_12753,N_12856);
nand U18926 (N_18926,N_10355,N_10356);
and U18927 (N_18927,N_14514,N_14311);
nor U18928 (N_18928,N_14356,N_10752);
nor U18929 (N_18929,N_10365,N_14766);
nand U18930 (N_18930,N_13265,N_14500);
nor U18931 (N_18931,N_14842,N_11732);
nand U18932 (N_18932,N_11957,N_11045);
xnor U18933 (N_18933,N_10831,N_10557);
xnor U18934 (N_18934,N_13856,N_10819);
or U18935 (N_18935,N_10039,N_13638);
and U18936 (N_18936,N_12210,N_11049);
nor U18937 (N_18937,N_13395,N_10964);
or U18938 (N_18938,N_10937,N_14004);
nor U18939 (N_18939,N_14075,N_10953);
nor U18940 (N_18940,N_10243,N_12755);
and U18941 (N_18941,N_11053,N_14585);
xnor U18942 (N_18942,N_14756,N_14125);
and U18943 (N_18943,N_10354,N_12790);
and U18944 (N_18944,N_10794,N_11684);
nand U18945 (N_18945,N_13075,N_14034);
nor U18946 (N_18946,N_13245,N_10523);
nor U18947 (N_18947,N_11601,N_10825);
nor U18948 (N_18948,N_14858,N_11248);
nand U18949 (N_18949,N_14292,N_12917);
and U18950 (N_18950,N_13443,N_10581);
or U18951 (N_18951,N_13522,N_10799);
nand U18952 (N_18952,N_14914,N_12082);
nor U18953 (N_18953,N_10190,N_12739);
nor U18954 (N_18954,N_12494,N_13293);
and U18955 (N_18955,N_11286,N_10324);
and U18956 (N_18956,N_12051,N_14856);
or U18957 (N_18957,N_14173,N_14905);
and U18958 (N_18958,N_12188,N_11267);
or U18959 (N_18959,N_13212,N_13245);
or U18960 (N_18960,N_12856,N_10487);
and U18961 (N_18961,N_13760,N_11092);
nor U18962 (N_18962,N_13565,N_10029);
nor U18963 (N_18963,N_12018,N_14839);
xnor U18964 (N_18964,N_13854,N_11608);
and U18965 (N_18965,N_12965,N_14505);
and U18966 (N_18966,N_10420,N_10486);
and U18967 (N_18967,N_10361,N_11466);
xnor U18968 (N_18968,N_14123,N_13398);
and U18969 (N_18969,N_13264,N_14210);
nor U18970 (N_18970,N_10550,N_11038);
nor U18971 (N_18971,N_12779,N_11874);
nor U18972 (N_18972,N_13586,N_11316);
or U18973 (N_18973,N_14311,N_10290);
or U18974 (N_18974,N_13008,N_13802);
nand U18975 (N_18975,N_11551,N_11745);
nor U18976 (N_18976,N_13112,N_13037);
or U18977 (N_18977,N_12232,N_12692);
and U18978 (N_18978,N_11209,N_10158);
nor U18979 (N_18979,N_11218,N_10532);
or U18980 (N_18980,N_12967,N_14922);
or U18981 (N_18981,N_11279,N_12188);
and U18982 (N_18982,N_12797,N_13073);
xnor U18983 (N_18983,N_11611,N_12679);
and U18984 (N_18984,N_11320,N_13395);
or U18985 (N_18985,N_11438,N_11032);
nor U18986 (N_18986,N_14233,N_14611);
nand U18987 (N_18987,N_10397,N_10549);
and U18988 (N_18988,N_12518,N_12881);
or U18989 (N_18989,N_10618,N_10559);
nand U18990 (N_18990,N_10019,N_11142);
and U18991 (N_18991,N_14157,N_12158);
nand U18992 (N_18992,N_13159,N_14891);
or U18993 (N_18993,N_11028,N_10478);
nor U18994 (N_18994,N_12203,N_14036);
nand U18995 (N_18995,N_10491,N_11308);
xnor U18996 (N_18996,N_13635,N_13685);
and U18997 (N_18997,N_10944,N_14036);
and U18998 (N_18998,N_11965,N_13643);
nor U18999 (N_18999,N_12134,N_10588);
nor U19000 (N_19000,N_14427,N_14429);
xnor U19001 (N_19001,N_14759,N_11218);
nor U19002 (N_19002,N_12193,N_12973);
nand U19003 (N_19003,N_12084,N_10051);
and U19004 (N_19004,N_13642,N_10131);
or U19005 (N_19005,N_13499,N_10900);
or U19006 (N_19006,N_11389,N_10180);
xor U19007 (N_19007,N_14746,N_11993);
nand U19008 (N_19008,N_12048,N_10417);
or U19009 (N_19009,N_11961,N_10590);
nor U19010 (N_19010,N_11501,N_14839);
nand U19011 (N_19011,N_13733,N_13406);
nand U19012 (N_19012,N_10610,N_12119);
and U19013 (N_19013,N_10820,N_11810);
and U19014 (N_19014,N_14040,N_13022);
or U19015 (N_19015,N_11061,N_11071);
and U19016 (N_19016,N_11733,N_12626);
and U19017 (N_19017,N_11647,N_11092);
or U19018 (N_19018,N_11054,N_14597);
or U19019 (N_19019,N_12761,N_12579);
nand U19020 (N_19020,N_12624,N_11404);
or U19021 (N_19021,N_14512,N_12611);
and U19022 (N_19022,N_10156,N_14932);
xor U19023 (N_19023,N_10473,N_13121);
and U19024 (N_19024,N_11970,N_12053);
nor U19025 (N_19025,N_11839,N_11915);
and U19026 (N_19026,N_10947,N_10737);
nor U19027 (N_19027,N_14140,N_10223);
nand U19028 (N_19028,N_10594,N_10147);
or U19029 (N_19029,N_12321,N_13889);
nand U19030 (N_19030,N_14873,N_14153);
and U19031 (N_19031,N_12658,N_12527);
or U19032 (N_19032,N_12749,N_11296);
or U19033 (N_19033,N_12609,N_10099);
nor U19034 (N_19034,N_14612,N_10681);
nor U19035 (N_19035,N_13673,N_12416);
nor U19036 (N_19036,N_13151,N_13585);
or U19037 (N_19037,N_12908,N_11583);
nor U19038 (N_19038,N_11758,N_10755);
nor U19039 (N_19039,N_13821,N_14592);
xor U19040 (N_19040,N_12253,N_10772);
xor U19041 (N_19041,N_14578,N_12380);
nand U19042 (N_19042,N_14565,N_13851);
and U19043 (N_19043,N_13529,N_13910);
or U19044 (N_19044,N_11642,N_13480);
xor U19045 (N_19045,N_14877,N_12514);
xnor U19046 (N_19046,N_11509,N_13216);
and U19047 (N_19047,N_11120,N_10920);
nor U19048 (N_19048,N_13418,N_13923);
and U19049 (N_19049,N_13968,N_10115);
and U19050 (N_19050,N_14905,N_12416);
nand U19051 (N_19051,N_14804,N_11372);
or U19052 (N_19052,N_12115,N_14867);
or U19053 (N_19053,N_11377,N_10994);
and U19054 (N_19054,N_12969,N_10838);
nand U19055 (N_19055,N_10423,N_11070);
or U19056 (N_19056,N_11290,N_12977);
or U19057 (N_19057,N_14221,N_13107);
nor U19058 (N_19058,N_12344,N_12556);
nor U19059 (N_19059,N_13351,N_11164);
or U19060 (N_19060,N_12807,N_12112);
nand U19061 (N_19061,N_13461,N_11351);
or U19062 (N_19062,N_13521,N_11141);
xor U19063 (N_19063,N_10007,N_13372);
xnor U19064 (N_19064,N_10694,N_11147);
and U19065 (N_19065,N_10511,N_13843);
xor U19066 (N_19066,N_14181,N_11513);
nand U19067 (N_19067,N_11746,N_10892);
nand U19068 (N_19068,N_13873,N_11263);
or U19069 (N_19069,N_11804,N_12563);
nor U19070 (N_19070,N_14737,N_10319);
and U19071 (N_19071,N_13710,N_11437);
nor U19072 (N_19072,N_12974,N_13107);
or U19073 (N_19073,N_14174,N_10718);
and U19074 (N_19074,N_12479,N_10047);
or U19075 (N_19075,N_11847,N_11677);
and U19076 (N_19076,N_11210,N_11641);
nand U19077 (N_19077,N_12979,N_13325);
xnor U19078 (N_19078,N_10193,N_13485);
xor U19079 (N_19079,N_10505,N_12823);
and U19080 (N_19080,N_13772,N_12819);
or U19081 (N_19081,N_14416,N_12199);
and U19082 (N_19082,N_11374,N_12763);
nor U19083 (N_19083,N_11002,N_11093);
nand U19084 (N_19084,N_13235,N_10191);
or U19085 (N_19085,N_10685,N_13759);
nand U19086 (N_19086,N_11842,N_14938);
and U19087 (N_19087,N_11197,N_14884);
nor U19088 (N_19088,N_12097,N_10935);
xor U19089 (N_19089,N_14379,N_11964);
or U19090 (N_19090,N_13332,N_10788);
and U19091 (N_19091,N_11509,N_11391);
nand U19092 (N_19092,N_10142,N_11816);
or U19093 (N_19093,N_10819,N_12210);
nor U19094 (N_19094,N_13930,N_11261);
nand U19095 (N_19095,N_14961,N_14506);
nand U19096 (N_19096,N_12356,N_14814);
xnor U19097 (N_19097,N_12698,N_14349);
and U19098 (N_19098,N_14922,N_14092);
or U19099 (N_19099,N_12030,N_10127);
and U19100 (N_19100,N_12526,N_10858);
nand U19101 (N_19101,N_10771,N_10329);
and U19102 (N_19102,N_14685,N_12110);
and U19103 (N_19103,N_11939,N_11301);
nor U19104 (N_19104,N_10902,N_10908);
or U19105 (N_19105,N_11391,N_10430);
nor U19106 (N_19106,N_11080,N_12522);
or U19107 (N_19107,N_12505,N_14506);
nor U19108 (N_19108,N_12618,N_11835);
nor U19109 (N_19109,N_11351,N_13264);
and U19110 (N_19110,N_12518,N_10528);
and U19111 (N_19111,N_14167,N_10943);
and U19112 (N_19112,N_13746,N_13287);
or U19113 (N_19113,N_11854,N_14080);
nand U19114 (N_19114,N_13588,N_10139);
or U19115 (N_19115,N_12342,N_13533);
nor U19116 (N_19116,N_10733,N_10777);
and U19117 (N_19117,N_13165,N_10693);
or U19118 (N_19118,N_10547,N_12549);
and U19119 (N_19119,N_14318,N_10332);
nand U19120 (N_19120,N_11963,N_14082);
and U19121 (N_19121,N_10572,N_12091);
nand U19122 (N_19122,N_13418,N_13238);
xor U19123 (N_19123,N_10619,N_11508);
or U19124 (N_19124,N_12121,N_12516);
nand U19125 (N_19125,N_11139,N_13049);
xnor U19126 (N_19126,N_14810,N_12508);
nand U19127 (N_19127,N_12928,N_13993);
or U19128 (N_19128,N_13395,N_13630);
and U19129 (N_19129,N_10119,N_13974);
and U19130 (N_19130,N_10660,N_14803);
nor U19131 (N_19131,N_12920,N_13736);
and U19132 (N_19132,N_13188,N_13810);
and U19133 (N_19133,N_14410,N_13889);
nand U19134 (N_19134,N_12777,N_10258);
xnor U19135 (N_19135,N_14806,N_13698);
or U19136 (N_19136,N_13757,N_11854);
nor U19137 (N_19137,N_11220,N_13516);
nand U19138 (N_19138,N_10910,N_10287);
nor U19139 (N_19139,N_11156,N_10604);
or U19140 (N_19140,N_11046,N_13865);
and U19141 (N_19141,N_11666,N_11688);
nor U19142 (N_19142,N_12422,N_12341);
xor U19143 (N_19143,N_13880,N_10489);
nand U19144 (N_19144,N_10304,N_13328);
and U19145 (N_19145,N_13424,N_11149);
and U19146 (N_19146,N_14487,N_12451);
nor U19147 (N_19147,N_12765,N_11208);
nand U19148 (N_19148,N_14685,N_11137);
and U19149 (N_19149,N_11343,N_14059);
or U19150 (N_19150,N_13307,N_12293);
or U19151 (N_19151,N_13510,N_12871);
nand U19152 (N_19152,N_14142,N_14760);
or U19153 (N_19153,N_10191,N_12295);
nand U19154 (N_19154,N_10608,N_11175);
and U19155 (N_19155,N_14982,N_11845);
and U19156 (N_19156,N_10150,N_12134);
nor U19157 (N_19157,N_12188,N_12428);
nor U19158 (N_19158,N_12870,N_14076);
nand U19159 (N_19159,N_14561,N_12402);
nor U19160 (N_19160,N_13130,N_14093);
nor U19161 (N_19161,N_13722,N_14764);
and U19162 (N_19162,N_10744,N_13451);
nand U19163 (N_19163,N_10478,N_11275);
or U19164 (N_19164,N_12224,N_10745);
or U19165 (N_19165,N_12382,N_10644);
nand U19166 (N_19166,N_11571,N_10157);
and U19167 (N_19167,N_11949,N_11158);
or U19168 (N_19168,N_12832,N_14018);
nand U19169 (N_19169,N_10564,N_13648);
and U19170 (N_19170,N_11642,N_13859);
and U19171 (N_19171,N_13280,N_13095);
or U19172 (N_19172,N_10513,N_14089);
and U19173 (N_19173,N_13287,N_11906);
nand U19174 (N_19174,N_12825,N_12901);
xnor U19175 (N_19175,N_12293,N_14584);
xnor U19176 (N_19176,N_12075,N_10644);
and U19177 (N_19177,N_13476,N_12577);
nor U19178 (N_19178,N_13956,N_11880);
xor U19179 (N_19179,N_10028,N_12919);
nor U19180 (N_19180,N_13120,N_12087);
or U19181 (N_19181,N_12241,N_14111);
xnor U19182 (N_19182,N_10098,N_13017);
nand U19183 (N_19183,N_14059,N_10464);
nor U19184 (N_19184,N_12368,N_11904);
nor U19185 (N_19185,N_13718,N_13590);
or U19186 (N_19186,N_12505,N_12882);
and U19187 (N_19187,N_10237,N_12314);
nand U19188 (N_19188,N_13328,N_12628);
nand U19189 (N_19189,N_10747,N_12492);
and U19190 (N_19190,N_12707,N_12474);
nand U19191 (N_19191,N_11154,N_10886);
xor U19192 (N_19192,N_11873,N_11616);
nand U19193 (N_19193,N_12902,N_11876);
or U19194 (N_19194,N_13449,N_11661);
nor U19195 (N_19195,N_12349,N_12359);
nor U19196 (N_19196,N_12357,N_13672);
and U19197 (N_19197,N_14110,N_12003);
xor U19198 (N_19198,N_14058,N_13192);
or U19199 (N_19199,N_14570,N_10299);
nand U19200 (N_19200,N_11437,N_13065);
and U19201 (N_19201,N_13096,N_10617);
nor U19202 (N_19202,N_12199,N_10123);
nor U19203 (N_19203,N_14978,N_13658);
nand U19204 (N_19204,N_14519,N_13965);
or U19205 (N_19205,N_14131,N_13472);
or U19206 (N_19206,N_10408,N_11468);
or U19207 (N_19207,N_14996,N_10288);
or U19208 (N_19208,N_11029,N_13260);
and U19209 (N_19209,N_13896,N_14167);
nor U19210 (N_19210,N_14264,N_10363);
or U19211 (N_19211,N_13778,N_14171);
nor U19212 (N_19212,N_12847,N_12731);
nor U19213 (N_19213,N_11477,N_13568);
nand U19214 (N_19214,N_12918,N_14779);
nand U19215 (N_19215,N_12728,N_11571);
nand U19216 (N_19216,N_11986,N_11961);
and U19217 (N_19217,N_14755,N_11522);
nor U19218 (N_19218,N_14769,N_11214);
or U19219 (N_19219,N_13412,N_12692);
xor U19220 (N_19220,N_12620,N_12642);
nand U19221 (N_19221,N_10937,N_12652);
nor U19222 (N_19222,N_10587,N_13101);
or U19223 (N_19223,N_13363,N_10053);
or U19224 (N_19224,N_13819,N_13021);
and U19225 (N_19225,N_14308,N_10373);
nor U19226 (N_19226,N_11668,N_12700);
nor U19227 (N_19227,N_12590,N_10375);
and U19228 (N_19228,N_13770,N_13584);
nand U19229 (N_19229,N_11919,N_11581);
and U19230 (N_19230,N_10524,N_14831);
or U19231 (N_19231,N_12428,N_11465);
xor U19232 (N_19232,N_13012,N_12665);
nor U19233 (N_19233,N_12633,N_11298);
nand U19234 (N_19234,N_10087,N_13606);
and U19235 (N_19235,N_13936,N_14100);
xor U19236 (N_19236,N_14880,N_13110);
nand U19237 (N_19237,N_10134,N_12751);
or U19238 (N_19238,N_14200,N_13148);
xnor U19239 (N_19239,N_12004,N_13917);
nor U19240 (N_19240,N_11782,N_14227);
xor U19241 (N_19241,N_13792,N_13825);
and U19242 (N_19242,N_10265,N_12683);
nand U19243 (N_19243,N_14411,N_13417);
and U19244 (N_19244,N_11201,N_10798);
nand U19245 (N_19245,N_14546,N_14171);
nor U19246 (N_19246,N_12399,N_12325);
or U19247 (N_19247,N_13991,N_12597);
or U19248 (N_19248,N_12683,N_10430);
nor U19249 (N_19249,N_13585,N_14460);
nand U19250 (N_19250,N_13516,N_14399);
and U19251 (N_19251,N_13116,N_12468);
nand U19252 (N_19252,N_12317,N_13374);
nor U19253 (N_19253,N_11679,N_10226);
or U19254 (N_19254,N_13388,N_10611);
nand U19255 (N_19255,N_12371,N_10643);
and U19256 (N_19256,N_12142,N_12325);
nand U19257 (N_19257,N_10984,N_14760);
nor U19258 (N_19258,N_12485,N_13874);
xnor U19259 (N_19259,N_10833,N_12916);
or U19260 (N_19260,N_13206,N_13200);
nor U19261 (N_19261,N_14422,N_13336);
and U19262 (N_19262,N_12174,N_10465);
or U19263 (N_19263,N_11376,N_11666);
and U19264 (N_19264,N_10065,N_13951);
and U19265 (N_19265,N_13673,N_14500);
and U19266 (N_19266,N_13749,N_13623);
xnor U19267 (N_19267,N_10897,N_10935);
nor U19268 (N_19268,N_10859,N_12024);
or U19269 (N_19269,N_11128,N_13297);
or U19270 (N_19270,N_12041,N_10528);
nor U19271 (N_19271,N_11214,N_11182);
xor U19272 (N_19272,N_12405,N_13075);
nand U19273 (N_19273,N_13146,N_13596);
nor U19274 (N_19274,N_11104,N_11679);
and U19275 (N_19275,N_13111,N_10795);
and U19276 (N_19276,N_12255,N_14868);
nand U19277 (N_19277,N_10513,N_11271);
nand U19278 (N_19278,N_13671,N_11070);
nand U19279 (N_19279,N_12532,N_13224);
and U19280 (N_19280,N_14637,N_10649);
or U19281 (N_19281,N_10399,N_13944);
and U19282 (N_19282,N_14605,N_10157);
nor U19283 (N_19283,N_10336,N_13361);
nor U19284 (N_19284,N_10349,N_10622);
and U19285 (N_19285,N_11390,N_12685);
nor U19286 (N_19286,N_11535,N_13511);
nand U19287 (N_19287,N_11979,N_14507);
nor U19288 (N_19288,N_11909,N_12447);
nand U19289 (N_19289,N_14676,N_13826);
or U19290 (N_19290,N_12445,N_13228);
or U19291 (N_19291,N_12902,N_11095);
nor U19292 (N_19292,N_10692,N_10472);
nor U19293 (N_19293,N_11938,N_14608);
nand U19294 (N_19294,N_12699,N_12899);
nor U19295 (N_19295,N_13255,N_10164);
nor U19296 (N_19296,N_10159,N_10871);
nor U19297 (N_19297,N_10185,N_14254);
xnor U19298 (N_19298,N_12492,N_10628);
and U19299 (N_19299,N_10842,N_11835);
and U19300 (N_19300,N_12914,N_10176);
or U19301 (N_19301,N_14188,N_11106);
xor U19302 (N_19302,N_10071,N_12731);
or U19303 (N_19303,N_12411,N_13286);
or U19304 (N_19304,N_11845,N_11943);
nand U19305 (N_19305,N_13798,N_10378);
nand U19306 (N_19306,N_10987,N_11501);
or U19307 (N_19307,N_10171,N_13089);
nand U19308 (N_19308,N_13946,N_13870);
and U19309 (N_19309,N_12381,N_13793);
xor U19310 (N_19310,N_10642,N_12670);
nor U19311 (N_19311,N_12259,N_11730);
nand U19312 (N_19312,N_12588,N_10036);
nand U19313 (N_19313,N_14770,N_10554);
or U19314 (N_19314,N_13780,N_11197);
and U19315 (N_19315,N_11685,N_13482);
and U19316 (N_19316,N_13381,N_13235);
nand U19317 (N_19317,N_13081,N_14052);
nand U19318 (N_19318,N_11034,N_14825);
xor U19319 (N_19319,N_11564,N_12265);
xor U19320 (N_19320,N_11579,N_14000);
nand U19321 (N_19321,N_12514,N_14737);
nand U19322 (N_19322,N_10903,N_14931);
nor U19323 (N_19323,N_12839,N_12329);
nor U19324 (N_19324,N_12689,N_13055);
nor U19325 (N_19325,N_14809,N_14321);
and U19326 (N_19326,N_14964,N_10970);
nor U19327 (N_19327,N_14869,N_13756);
nand U19328 (N_19328,N_11506,N_13847);
or U19329 (N_19329,N_12819,N_11878);
or U19330 (N_19330,N_12601,N_13326);
nor U19331 (N_19331,N_14634,N_10267);
or U19332 (N_19332,N_11749,N_12533);
or U19333 (N_19333,N_14425,N_10902);
nor U19334 (N_19334,N_14711,N_14308);
and U19335 (N_19335,N_12468,N_11086);
nand U19336 (N_19336,N_10812,N_11077);
and U19337 (N_19337,N_14834,N_13042);
nor U19338 (N_19338,N_14508,N_10737);
nor U19339 (N_19339,N_12095,N_11282);
or U19340 (N_19340,N_10261,N_12966);
and U19341 (N_19341,N_12597,N_10982);
or U19342 (N_19342,N_11739,N_10277);
nand U19343 (N_19343,N_12912,N_10577);
xor U19344 (N_19344,N_13276,N_10017);
or U19345 (N_19345,N_13296,N_11986);
nand U19346 (N_19346,N_10439,N_10093);
nor U19347 (N_19347,N_12244,N_12895);
nand U19348 (N_19348,N_12987,N_11342);
nand U19349 (N_19349,N_12739,N_13620);
xnor U19350 (N_19350,N_13096,N_14157);
or U19351 (N_19351,N_13167,N_11192);
or U19352 (N_19352,N_14684,N_10458);
xor U19353 (N_19353,N_13730,N_10838);
xnor U19354 (N_19354,N_12249,N_10418);
and U19355 (N_19355,N_10153,N_10228);
nand U19356 (N_19356,N_11688,N_12574);
or U19357 (N_19357,N_11735,N_14808);
nand U19358 (N_19358,N_12076,N_10258);
nor U19359 (N_19359,N_13450,N_10794);
nand U19360 (N_19360,N_11723,N_14873);
and U19361 (N_19361,N_11407,N_14616);
and U19362 (N_19362,N_11593,N_10372);
or U19363 (N_19363,N_13668,N_12695);
nand U19364 (N_19364,N_11009,N_10537);
nand U19365 (N_19365,N_10315,N_11667);
nand U19366 (N_19366,N_11689,N_13158);
xnor U19367 (N_19367,N_13377,N_13046);
nand U19368 (N_19368,N_12860,N_14106);
or U19369 (N_19369,N_14001,N_14118);
nand U19370 (N_19370,N_10529,N_14968);
nand U19371 (N_19371,N_13176,N_10808);
and U19372 (N_19372,N_10690,N_12032);
or U19373 (N_19373,N_13544,N_12044);
nor U19374 (N_19374,N_11804,N_11523);
or U19375 (N_19375,N_14483,N_12852);
or U19376 (N_19376,N_13712,N_14164);
xor U19377 (N_19377,N_12068,N_12168);
nor U19378 (N_19378,N_14780,N_14839);
nand U19379 (N_19379,N_12958,N_12045);
nand U19380 (N_19380,N_11743,N_14837);
or U19381 (N_19381,N_10664,N_12619);
and U19382 (N_19382,N_13044,N_11880);
nor U19383 (N_19383,N_13380,N_12826);
nand U19384 (N_19384,N_10776,N_10758);
nand U19385 (N_19385,N_13363,N_11820);
and U19386 (N_19386,N_13791,N_11598);
nand U19387 (N_19387,N_12560,N_12246);
nor U19388 (N_19388,N_12553,N_12081);
and U19389 (N_19389,N_12470,N_12528);
nand U19390 (N_19390,N_12258,N_10845);
nand U19391 (N_19391,N_13267,N_11656);
and U19392 (N_19392,N_10029,N_12749);
or U19393 (N_19393,N_13431,N_13473);
nand U19394 (N_19394,N_13881,N_14335);
and U19395 (N_19395,N_11236,N_10594);
nand U19396 (N_19396,N_12609,N_14083);
or U19397 (N_19397,N_10480,N_11052);
nand U19398 (N_19398,N_13262,N_13079);
nand U19399 (N_19399,N_14063,N_12064);
or U19400 (N_19400,N_10496,N_10325);
and U19401 (N_19401,N_14125,N_10358);
nand U19402 (N_19402,N_11067,N_11197);
nor U19403 (N_19403,N_12398,N_14608);
and U19404 (N_19404,N_13936,N_12309);
nand U19405 (N_19405,N_14421,N_11678);
nand U19406 (N_19406,N_11531,N_14093);
nor U19407 (N_19407,N_10264,N_10279);
nand U19408 (N_19408,N_12052,N_13954);
and U19409 (N_19409,N_12387,N_10337);
and U19410 (N_19410,N_11299,N_10221);
nor U19411 (N_19411,N_10491,N_12257);
or U19412 (N_19412,N_14254,N_12059);
nand U19413 (N_19413,N_14674,N_10034);
or U19414 (N_19414,N_11277,N_10235);
xnor U19415 (N_19415,N_11307,N_10411);
nor U19416 (N_19416,N_10789,N_13817);
or U19417 (N_19417,N_12378,N_10201);
nand U19418 (N_19418,N_14080,N_14772);
nor U19419 (N_19419,N_10156,N_14195);
and U19420 (N_19420,N_10821,N_10133);
nor U19421 (N_19421,N_10153,N_11613);
nor U19422 (N_19422,N_12137,N_10588);
and U19423 (N_19423,N_11803,N_10324);
nand U19424 (N_19424,N_12380,N_11613);
and U19425 (N_19425,N_10268,N_13393);
and U19426 (N_19426,N_14300,N_12467);
nor U19427 (N_19427,N_12256,N_14804);
nand U19428 (N_19428,N_14043,N_10985);
or U19429 (N_19429,N_14229,N_10264);
and U19430 (N_19430,N_12534,N_11557);
or U19431 (N_19431,N_14136,N_11057);
and U19432 (N_19432,N_14069,N_13968);
nor U19433 (N_19433,N_14699,N_11327);
xnor U19434 (N_19434,N_13645,N_13171);
and U19435 (N_19435,N_14277,N_10541);
or U19436 (N_19436,N_13437,N_13502);
nand U19437 (N_19437,N_14277,N_13875);
or U19438 (N_19438,N_11079,N_14789);
or U19439 (N_19439,N_12682,N_13003);
and U19440 (N_19440,N_11594,N_11892);
and U19441 (N_19441,N_10619,N_12816);
nand U19442 (N_19442,N_10795,N_12266);
nand U19443 (N_19443,N_13846,N_10398);
and U19444 (N_19444,N_14179,N_11607);
nor U19445 (N_19445,N_10639,N_14220);
xnor U19446 (N_19446,N_13047,N_11064);
nand U19447 (N_19447,N_10101,N_10126);
or U19448 (N_19448,N_10236,N_11461);
nand U19449 (N_19449,N_14504,N_14676);
and U19450 (N_19450,N_12622,N_10709);
nor U19451 (N_19451,N_14920,N_14356);
nor U19452 (N_19452,N_11008,N_10225);
nor U19453 (N_19453,N_10452,N_10776);
nand U19454 (N_19454,N_14598,N_12338);
nand U19455 (N_19455,N_10138,N_13940);
nor U19456 (N_19456,N_12786,N_13259);
and U19457 (N_19457,N_11359,N_14315);
and U19458 (N_19458,N_12385,N_10831);
nand U19459 (N_19459,N_11500,N_10257);
xor U19460 (N_19460,N_14736,N_14579);
or U19461 (N_19461,N_10774,N_12981);
and U19462 (N_19462,N_13869,N_11160);
nand U19463 (N_19463,N_12990,N_10386);
nand U19464 (N_19464,N_13033,N_14762);
nor U19465 (N_19465,N_12697,N_10405);
nor U19466 (N_19466,N_10929,N_11249);
and U19467 (N_19467,N_12465,N_12627);
or U19468 (N_19468,N_13972,N_10120);
nand U19469 (N_19469,N_10283,N_14372);
nor U19470 (N_19470,N_10037,N_14696);
nand U19471 (N_19471,N_10674,N_11354);
and U19472 (N_19472,N_12479,N_13728);
nor U19473 (N_19473,N_11759,N_14166);
and U19474 (N_19474,N_10068,N_12552);
or U19475 (N_19475,N_10519,N_14387);
nand U19476 (N_19476,N_10615,N_13305);
nand U19477 (N_19477,N_12832,N_10846);
nand U19478 (N_19478,N_12488,N_12686);
or U19479 (N_19479,N_11584,N_10379);
nor U19480 (N_19480,N_10626,N_14632);
nor U19481 (N_19481,N_14273,N_12766);
nand U19482 (N_19482,N_12785,N_10463);
nor U19483 (N_19483,N_10230,N_10290);
nor U19484 (N_19484,N_11164,N_12092);
or U19485 (N_19485,N_11185,N_14183);
nor U19486 (N_19486,N_14102,N_13661);
or U19487 (N_19487,N_12558,N_12137);
and U19488 (N_19488,N_14431,N_11733);
nor U19489 (N_19489,N_11590,N_14367);
nand U19490 (N_19490,N_14293,N_14434);
or U19491 (N_19491,N_11300,N_13741);
and U19492 (N_19492,N_10341,N_10347);
or U19493 (N_19493,N_14643,N_12333);
or U19494 (N_19494,N_14559,N_10175);
xor U19495 (N_19495,N_12117,N_12240);
nor U19496 (N_19496,N_13761,N_11644);
and U19497 (N_19497,N_14695,N_10585);
xor U19498 (N_19498,N_10353,N_10662);
or U19499 (N_19499,N_10208,N_14008);
nor U19500 (N_19500,N_12965,N_11095);
xor U19501 (N_19501,N_14808,N_11710);
and U19502 (N_19502,N_14437,N_11380);
nor U19503 (N_19503,N_11067,N_13737);
or U19504 (N_19504,N_12335,N_10750);
nor U19505 (N_19505,N_14721,N_11002);
nand U19506 (N_19506,N_10501,N_13870);
nand U19507 (N_19507,N_10238,N_13514);
or U19508 (N_19508,N_12299,N_12387);
and U19509 (N_19509,N_14496,N_10840);
nor U19510 (N_19510,N_13197,N_11686);
nor U19511 (N_19511,N_11641,N_14545);
nand U19512 (N_19512,N_10079,N_12913);
and U19513 (N_19513,N_11279,N_10575);
or U19514 (N_19514,N_12019,N_11154);
nand U19515 (N_19515,N_11449,N_10545);
and U19516 (N_19516,N_12676,N_14485);
nand U19517 (N_19517,N_10644,N_12202);
xor U19518 (N_19518,N_13341,N_13808);
nor U19519 (N_19519,N_11770,N_14591);
nor U19520 (N_19520,N_13870,N_13564);
nand U19521 (N_19521,N_13033,N_14756);
nand U19522 (N_19522,N_10771,N_12062);
and U19523 (N_19523,N_13471,N_14032);
nand U19524 (N_19524,N_10393,N_12885);
nand U19525 (N_19525,N_12286,N_12952);
xor U19526 (N_19526,N_14398,N_11182);
nor U19527 (N_19527,N_11887,N_12473);
or U19528 (N_19528,N_10662,N_12782);
nand U19529 (N_19529,N_12538,N_14837);
nor U19530 (N_19530,N_13767,N_13279);
and U19531 (N_19531,N_13997,N_11869);
nor U19532 (N_19532,N_11543,N_14250);
nand U19533 (N_19533,N_14751,N_13842);
and U19534 (N_19534,N_12346,N_14858);
nor U19535 (N_19535,N_13613,N_11754);
nor U19536 (N_19536,N_14948,N_10333);
and U19537 (N_19537,N_13972,N_12237);
xnor U19538 (N_19538,N_10542,N_12789);
xor U19539 (N_19539,N_11991,N_11066);
and U19540 (N_19540,N_10121,N_10925);
xor U19541 (N_19541,N_10025,N_11671);
or U19542 (N_19542,N_14040,N_11449);
xor U19543 (N_19543,N_13537,N_12612);
nor U19544 (N_19544,N_12110,N_12322);
and U19545 (N_19545,N_10420,N_13320);
nand U19546 (N_19546,N_14335,N_11646);
nand U19547 (N_19547,N_10869,N_10548);
or U19548 (N_19548,N_12058,N_13158);
xnor U19549 (N_19549,N_14569,N_10002);
and U19550 (N_19550,N_12649,N_10321);
and U19551 (N_19551,N_10663,N_12695);
and U19552 (N_19552,N_10780,N_13550);
xor U19553 (N_19553,N_12493,N_10513);
nand U19554 (N_19554,N_14950,N_11531);
or U19555 (N_19555,N_13697,N_11938);
or U19556 (N_19556,N_12466,N_12005);
xor U19557 (N_19557,N_10829,N_13460);
nor U19558 (N_19558,N_14076,N_12839);
and U19559 (N_19559,N_13557,N_12991);
nor U19560 (N_19560,N_13299,N_10470);
nand U19561 (N_19561,N_14197,N_12000);
or U19562 (N_19562,N_14590,N_12632);
and U19563 (N_19563,N_13100,N_12013);
nor U19564 (N_19564,N_14227,N_11126);
or U19565 (N_19565,N_11350,N_11644);
and U19566 (N_19566,N_13492,N_13497);
and U19567 (N_19567,N_13692,N_14359);
or U19568 (N_19568,N_11324,N_12021);
and U19569 (N_19569,N_11772,N_11478);
xor U19570 (N_19570,N_13949,N_10408);
nand U19571 (N_19571,N_13446,N_12182);
nand U19572 (N_19572,N_13984,N_12017);
or U19573 (N_19573,N_11588,N_12872);
nand U19574 (N_19574,N_14697,N_10000);
xor U19575 (N_19575,N_12966,N_10403);
or U19576 (N_19576,N_13439,N_13398);
nand U19577 (N_19577,N_11262,N_14933);
and U19578 (N_19578,N_12822,N_11193);
xor U19579 (N_19579,N_13667,N_12464);
or U19580 (N_19580,N_14858,N_10382);
or U19581 (N_19581,N_11797,N_11728);
and U19582 (N_19582,N_11658,N_14619);
or U19583 (N_19583,N_13313,N_11773);
or U19584 (N_19584,N_13458,N_14430);
nand U19585 (N_19585,N_10206,N_12107);
and U19586 (N_19586,N_10368,N_10103);
nor U19587 (N_19587,N_11672,N_14892);
or U19588 (N_19588,N_14781,N_12652);
or U19589 (N_19589,N_11545,N_12576);
and U19590 (N_19590,N_10530,N_11607);
or U19591 (N_19591,N_11620,N_10737);
xnor U19592 (N_19592,N_14294,N_11036);
and U19593 (N_19593,N_10240,N_11311);
and U19594 (N_19594,N_11581,N_13660);
nand U19595 (N_19595,N_10915,N_11361);
or U19596 (N_19596,N_14939,N_13265);
nor U19597 (N_19597,N_10292,N_11313);
and U19598 (N_19598,N_10226,N_13137);
nor U19599 (N_19599,N_13443,N_10887);
xnor U19600 (N_19600,N_13868,N_11153);
or U19601 (N_19601,N_13386,N_12902);
nor U19602 (N_19602,N_11029,N_14647);
or U19603 (N_19603,N_12596,N_10719);
xnor U19604 (N_19604,N_11652,N_14313);
xor U19605 (N_19605,N_12256,N_13421);
xnor U19606 (N_19606,N_14175,N_11431);
or U19607 (N_19607,N_14061,N_13717);
and U19608 (N_19608,N_10798,N_11031);
xor U19609 (N_19609,N_13849,N_14490);
and U19610 (N_19610,N_12878,N_12612);
and U19611 (N_19611,N_12898,N_11848);
and U19612 (N_19612,N_12964,N_13830);
or U19613 (N_19613,N_14751,N_11350);
or U19614 (N_19614,N_11941,N_14422);
and U19615 (N_19615,N_11161,N_10835);
nor U19616 (N_19616,N_12529,N_10110);
xnor U19617 (N_19617,N_12482,N_12959);
nor U19618 (N_19618,N_12363,N_12475);
nor U19619 (N_19619,N_14779,N_12936);
or U19620 (N_19620,N_10203,N_12548);
nand U19621 (N_19621,N_11048,N_14815);
and U19622 (N_19622,N_13136,N_13668);
nor U19623 (N_19623,N_10682,N_14653);
and U19624 (N_19624,N_13103,N_13878);
and U19625 (N_19625,N_13969,N_13880);
and U19626 (N_19626,N_12540,N_14144);
nor U19627 (N_19627,N_11571,N_14265);
nand U19628 (N_19628,N_14823,N_10400);
nor U19629 (N_19629,N_10072,N_14858);
nor U19630 (N_19630,N_11590,N_12735);
nor U19631 (N_19631,N_12235,N_12089);
nand U19632 (N_19632,N_14776,N_14026);
nor U19633 (N_19633,N_11673,N_14273);
nand U19634 (N_19634,N_12103,N_10257);
xnor U19635 (N_19635,N_10018,N_12452);
and U19636 (N_19636,N_13448,N_13037);
nand U19637 (N_19637,N_10859,N_14959);
nor U19638 (N_19638,N_12487,N_14071);
nor U19639 (N_19639,N_13257,N_14653);
or U19640 (N_19640,N_14579,N_14650);
nand U19641 (N_19641,N_11950,N_14657);
nand U19642 (N_19642,N_14157,N_12334);
nor U19643 (N_19643,N_11924,N_11042);
xnor U19644 (N_19644,N_12394,N_13492);
nor U19645 (N_19645,N_13000,N_12074);
xor U19646 (N_19646,N_11331,N_12750);
or U19647 (N_19647,N_10989,N_10933);
or U19648 (N_19648,N_14878,N_13909);
nor U19649 (N_19649,N_11404,N_13052);
or U19650 (N_19650,N_14831,N_10992);
nor U19651 (N_19651,N_12215,N_12313);
or U19652 (N_19652,N_10597,N_14605);
or U19653 (N_19653,N_10529,N_13515);
xor U19654 (N_19654,N_10547,N_12597);
or U19655 (N_19655,N_12899,N_10923);
nor U19656 (N_19656,N_10706,N_13165);
nor U19657 (N_19657,N_14522,N_12061);
nand U19658 (N_19658,N_12176,N_13844);
nand U19659 (N_19659,N_10424,N_10792);
nand U19660 (N_19660,N_11906,N_13054);
nor U19661 (N_19661,N_12327,N_10707);
nor U19662 (N_19662,N_11689,N_10990);
and U19663 (N_19663,N_12107,N_10693);
or U19664 (N_19664,N_14551,N_10325);
and U19665 (N_19665,N_13439,N_14483);
nor U19666 (N_19666,N_11605,N_11120);
or U19667 (N_19667,N_13383,N_13785);
xor U19668 (N_19668,N_13485,N_14849);
nor U19669 (N_19669,N_14850,N_14042);
or U19670 (N_19670,N_13652,N_11439);
and U19671 (N_19671,N_11408,N_10136);
nor U19672 (N_19672,N_11104,N_14463);
nand U19673 (N_19673,N_10555,N_12455);
nor U19674 (N_19674,N_11535,N_10978);
nand U19675 (N_19675,N_10992,N_14151);
and U19676 (N_19676,N_11825,N_10908);
or U19677 (N_19677,N_14868,N_10374);
nor U19678 (N_19678,N_10959,N_12016);
and U19679 (N_19679,N_10860,N_13616);
nand U19680 (N_19680,N_10224,N_10273);
nor U19681 (N_19681,N_11241,N_10960);
nor U19682 (N_19682,N_10634,N_12561);
nand U19683 (N_19683,N_11828,N_10577);
or U19684 (N_19684,N_11521,N_11352);
and U19685 (N_19685,N_12979,N_13978);
or U19686 (N_19686,N_14292,N_13499);
or U19687 (N_19687,N_14109,N_13891);
nor U19688 (N_19688,N_14375,N_11939);
or U19689 (N_19689,N_11457,N_13570);
or U19690 (N_19690,N_12460,N_13816);
or U19691 (N_19691,N_14952,N_11180);
nand U19692 (N_19692,N_13123,N_11314);
nand U19693 (N_19693,N_10676,N_11339);
or U19694 (N_19694,N_11262,N_10803);
nor U19695 (N_19695,N_14390,N_11396);
nand U19696 (N_19696,N_13921,N_12812);
nand U19697 (N_19697,N_11362,N_10677);
and U19698 (N_19698,N_12063,N_14879);
or U19699 (N_19699,N_11323,N_13045);
nor U19700 (N_19700,N_12926,N_12782);
and U19701 (N_19701,N_14442,N_12468);
xnor U19702 (N_19702,N_10615,N_11516);
and U19703 (N_19703,N_13636,N_13256);
nor U19704 (N_19704,N_12646,N_12339);
xor U19705 (N_19705,N_10261,N_10999);
nor U19706 (N_19706,N_10956,N_10138);
nor U19707 (N_19707,N_12335,N_14546);
and U19708 (N_19708,N_10181,N_12527);
and U19709 (N_19709,N_12414,N_11754);
and U19710 (N_19710,N_13563,N_14870);
and U19711 (N_19711,N_14230,N_11335);
or U19712 (N_19712,N_14935,N_11670);
nand U19713 (N_19713,N_10106,N_11082);
nand U19714 (N_19714,N_11926,N_12865);
nand U19715 (N_19715,N_11604,N_13778);
nand U19716 (N_19716,N_12661,N_13317);
nor U19717 (N_19717,N_11327,N_14051);
and U19718 (N_19718,N_12747,N_14698);
and U19719 (N_19719,N_14611,N_11773);
nand U19720 (N_19720,N_14159,N_12135);
nor U19721 (N_19721,N_10445,N_11005);
nor U19722 (N_19722,N_13588,N_10321);
or U19723 (N_19723,N_11691,N_11110);
nor U19724 (N_19724,N_13135,N_11761);
nand U19725 (N_19725,N_10476,N_13569);
or U19726 (N_19726,N_13108,N_10684);
and U19727 (N_19727,N_10339,N_10239);
and U19728 (N_19728,N_12396,N_12282);
nand U19729 (N_19729,N_12368,N_10157);
or U19730 (N_19730,N_12161,N_10512);
nor U19731 (N_19731,N_12670,N_14122);
nand U19732 (N_19732,N_14765,N_12664);
xor U19733 (N_19733,N_12497,N_10351);
or U19734 (N_19734,N_13044,N_13126);
nor U19735 (N_19735,N_10017,N_14237);
nand U19736 (N_19736,N_13584,N_13338);
xnor U19737 (N_19737,N_13179,N_12528);
or U19738 (N_19738,N_10277,N_11693);
nand U19739 (N_19739,N_10422,N_12161);
nand U19740 (N_19740,N_11728,N_12373);
nor U19741 (N_19741,N_11264,N_12963);
nor U19742 (N_19742,N_13816,N_11627);
or U19743 (N_19743,N_14425,N_12795);
nor U19744 (N_19744,N_11431,N_12745);
nand U19745 (N_19745,N_12391,N_12078);
nor U19746 (N_19746,N_14468,N_14336);
nand U19747 (N_19747,N_10567,N_14412);
nor U19748 (N_19748,N_13878,N_10267);
nand U19749 (N_19749,N_10582,N_12257);
xnor U19750 (N_19750,N_14480,N_10162);
and U19751 (N_19751,N_10675,N_10713);
nand U19752 (N_19752,N_13499,N_14454);
and U19753 (N_19753,N_10973,N_11807);
or U19754 (N_19754,N_13830,N_12492);
or U19755 (N_19755,N_13892,N_14654);
nor U19756 (N_19756,N_11791,N_11132);
xnor U19757 (N_19757,N_10458,N_14364);
and U19758 (N_19758,N_11849,N_13404);
or U19759 (N_19759,N_12024,N_10720);
and U19760 (N_19760,N_11533,N_11627);
and U19761 (N_19761,N_14449,N_10995);
and U19762 (N_19762,N_14451,N_12358);
and U19763 (N_19763,N_13420,N_11781);
or U19764 (N_19764,N_14528,N_10544);
and U19765 (N_19765,N_14082,N_12967);
nand U19766 (N_19766,N_14771,N_11379);
and U19767 (N_19767,N_12616,N_13886);
or U19768 (N_19768,N_13439,N_11728);
or U19769 (N_19769,N_13558,N_11068);
nand U19770 (N_19770,N_10569,N_14548);
xor U19771 (N_19771,N_13793,N_10833);
and U19772 (N_19772,N_13004,N_10546);
nor U19773 (N_19773,N_10772,N_13989);
nand U19774 (N_19774,N_13688,N_12307);
nor U19775 (N_19775,N_14132,N_14011);
or U19776 (N_19776,N_10364,N_10949);
and U19777 (N_19777,N_13992,N_10228);
xnor U19778 (N_19778,N_14312,N_10103);
nor U19779 (N_19779,N_12208,N_14389);
and U19780 (N_19780,N_14447,N_13542);
nor U19781 (N_19781,N_14960,N_12356);
and U19782 (N_19782,N_14514,N_12100);
nand U19783 (N_19783,N_11963,N_13408);
nand U19784 (N_19784,N_14173,N_14550);
nor U19785 (N_19785,N_11483,N_14689);
xor U19786 (N_19786,N_11687,N_11136);
nand U19787 (N_19787,N_14218,N_13609);
nand U19788 (N_19788,N_12135,N_11548);
nand U19789 (N_19789,N_10330,N_10259);
nand U19790 (N_19790,N_11105,N_11145);
xnor U19791 (N_19791,N_11129,N_14322);
nor U19792 (N_19792,N_10315,N_11603);
nor U19793 (N_19793,N_10658,N_11496);
nand U19794 (N_19794,N_12373,N_14134);
and U19795 (N_19795,N_12172,N_14639);
nor U19796 (N_19796,N_10949,N_12825);
xnor U19797 (N_19797,N_14853,N_10079);
nand U19798 (N_19798,N_14626,N_11751);
nand U19799 (N_19799,N_10961,N_11875);
or U19800 (N_19800,N_12939,N_13597);
and U19801 (N_19801,N_12639,N_13311);
nor U19802 (N_19802,N_12597,N_14161);
and U19803 (N_19803,N_11391,N_11032);
and U19804 (N_19804,N_14187,N_14855);
or U19805 (N_19805,N_14067,N_12861);
nand U19806 (N_19806,N_14431,N_11536);
or U19807 (N_19807,N_14461,N_12637);
or U19808 (N_19808,N_13703,N_13432);
and U19809 (N_19809,N_13099,N_10513);
or U19810 (N_19810,N_14791,N_11624);
xnor U19811 (N_19811,N_10876,N_12487);
nand U19812 (N_19812,N_10468,N_10743);
or U19813 (N_19813,N_13512,N_12566);
and U19814 (N_19814,N_11188,N_11849);
and U19815 (N_19815,N_13873,N_12441);
or U19816 (N_19816,N_12352,N_12191);
and U19817 (N_19817,N_12288,N_14836);
and U19818 (N_19818,N_12512,N_11099);
and U19819 (N_19819,N_13658,N_11808);
and U19820 (N_19820,N_10999,N_12159);
or U19821 (N_19821,N_11754,N_11776);
or U19822 (N_19822,N_14399,N_13988);
and U19823 (N_19823,N_14799,N_12456);
nand U19824 (N_19824,N_14252,N_11163);
and U19825 (N_19825,N_14909,N_14034);
and U19826 (N_19826,N_14338,N_11795);
nor U19827 (N_19827,N_14926,N_10829);
xor U19828 (N_19828,N_12179,N_13313);
and U19829 (N_19829,N_13610,N_12251);
or U19830 (N_19830,N_13270,N_13057);
and U19831 (N_19831,N_14802,N_11690);
or U19832 (N_19832,N_11235,N_12333);
and U19833 (N_19833,N_10760,N_14162);
nor U19834 (N_19834,N_14447,N_10045);
nor U19835 (N_19835,N_11521,N_10569);
nand U19836 (N_19836,N_13556,N_14785);
xor U19837 (N_19837,N_10549,N_11891);
or U19838 (N_19838,N_13162,N_11784);
nand U19839 (N_19839,N_14791,N_14751);
nand U19840 (N_19840,N_14047,N_14691);
nor U19841 (N_19841,N_14371,N_12619);
or U19842 (N_19842,N_12005,N_14706);
nand U19843 (N_19843,N_12282,N_12824);
and U19844 (N_19844,N_10733,N_14190);
and U19845 (N_19845,N_13374,N_13749);
nand U19846 (N_19846,N_11370,N_14349);
and U19847 (N_19847,N_11723,N_10514);
nor U19848 (N_19848,N_11283,N_11781);
nor U19849 (N_19849,N_11566,N_14885);
and U19850 (N_19850,N_10908,N_14257);
or U19851 (N_19851,N_14232,N_11120);
xor U19852 (N_19852,N_13149,N_11605);
and U19853 (N_19853,N_14379,N_10984);
xor U19854 (N_19854,N_10635,N_13872);
and U19855 (N_19855,N_12351,N_12235);
nor U19856 (N_19856,N_11390,N_11883);
nor U19857 (N_19857,N_11544,N_10540);
and U19858 (N_19858,N_13066,N_13381);
nor U19859 (N_19859,N_12579,N_12241);
and U19860 (N_19860,N_14814,N_12324);
or U19861 (N_19861,N_14895,N_10427);
and U19862 (N_19862,N_10111,N_12509);
or U19863 (N_19863,N_12793,N_11731);
nand U19864 (N_19864,N_12316,N_14034);
and U19865 (N_19865,N_12268,N_13665);
and U19866 (N_19866,N_14012,N_12707);
or U19867 (N_19867,N_13092,N_11951);
xnor U19868 (N_19868,N_14920,N_12914);
or U19869 (N_19869,N_11117,N_14515);
nor U19870 (N_19870,N_14941,N_10017);
nand U19871 (N_19871,N_13652,N_12596);
or U19872 (N_19872,N_14577,N_10698);
nor U19873 (N_19873,N_10021,N_11500);
or U19874 (N_19874,N_12781,N_14818);
and U19875 (N_19875,N_12379,N_13506);
and U19876 (N_19876,N_11934,N_12582);
xnor U19877 (N_19877,N_12268,N_12479);
nor U19878 (N_19878,N_13269,N_13018);
nor U19879 (N_19879,N_13591,N_10103);
nand U19880 (N_19880,N_13246,N_14905);
and U19881 (N_19881,N_12754,N_12105);
and U19882 (N_19882,N_10121,N_12489);
and U19883 (N_19883,N_10323,N_10845);
nand U19884 (N_19884,N_11855,N_14344);
nand U19885 (N_19885,N_10400,N_14418);
and U19886 (N_19886,N_14729,N_11958);
nor U19887 (N_19887,N_14306,N_14991);
nor U19888 (N_19888,N_10759,N_13271);
nand U19889 (N_19889,N_13774,N_11687);
nand U19890 (N_19890,N_10832,N_13390);
nor U19891 (N_19891,N_11610,N_10172);
nand U19892 (N_19892,N_10355,N_13973);
or U19893 (N_19893,N_10534,N_12757);
nand U19894 (N_19894,N_11634,N_10479);
nand U19895 (N_19895,N_11266,N_14452);
or U19896 (N_19896,N_10892,N_11633);
or U19897 (N_19897,N_14415,N_13717);
xnor U19898 (N_19898,N_11080,N_12469);
nand U19899 (N_19899,N_14815,N_14486);
nand U19900 (N_19900,N_10686,N_13990);
or U19901 (N_19901,N_13615,N_10546);
or U19902 (N_19902,N_13358,N_10279);
nor U19903 (N_19903,N_13487,N_14712);
xnor U19904 (N_19904,N_13622,N_12876);
nor U19905 (N_19905,N_10781,N_12276);
xor U19906 (N_19906,N_12578,N_13290);
or U19907 (N_19907,N_14457,N_13826);
or U19908 (N_19908,N_11119,N_14217);
and U19909 (N_19909,N_13443,N_10373);
or U19910 (N_19910,N_14627,N_14235);
and U19911 (N_19911,N_13395,N_12053);
nand U19912 (N_19912,N_10778,N_14269);
or U19913 (N_19913,N_14458,N_11956);
and U19914 (N_19914,N_14525,N_14808);
nand U19915 (N_19915,N_13711,N_11238);
and U19916 (N_19916,N_14227,N_14362);
or U19917 (N_19917,N_10181,N_13329);
and U19918 (N_19918,N_10221,N_13357);
xnor U19919 (N_19919,N_12986,N_10705);
and U19920 (N_19920,N_14382,N_10152);
nor U19921 (N_19921,N_13832,N_14187);
or U19922 (N_19922,N_14806,N_14533);
and U19923 (N_19923,N_12127,N_13935);
nand U19924 (N_19924,N_10096,N_12940);
nor U19925 (N_19925,N_14959,N_11808);
or U19926 (N_19926,N_10560,N_13915);
or U19927 (N_19927,N_14486,N_13405);
or U19928 (N_19928,N_12697,N_12514);
nand U19929 (N_19929,N_11455,N_12324);
and U19930 (N_19930,N_10396,N_13619);
nor U19931 (N_19931,N_12994,N_10513);
nand U19932 (N_19932,N_12749,N_13368);
nand U19933 (N_19933,N_10075,N_13835);
and U19934 (N_19934,N_10701,N_10089);
nor U19935 (N_19935,N_11352,N_12637);
nor U19936 (N_19936,N_12017,N_13616);
xnor U19937 (N_19937,N_10261,N_11154);
xor U19938 (N_19938,N_12237,N_12982);
nor U19939 (N_19939,N_11318,N_10657);
nand U19940 (N_19940,N_10274,N_13678);
nor U19941 (N_19941,N_13822,N_10396);
or U19942 (N_19942,N_11504,N_11400);
or U19943 (N_19943,N_10835,N_11421);
nand U19944 (N_19944,N_13713,N_12620);
or U19945 (N_19945,N_11847,N_13956);
nor U19946 (N_19946,N_14142,N_11874);
nor U19947 (N_19947,N_13318,N_10122);
or U19948 (N_19948,N_11937,N_12878);
nand U19949 (N_19949,N_10858,N_11474);
and U19950 (N_19950,N_11493,N_10935);
or U19951 (N_19951,N_11129,N_12068);
nand U19952 (N_19952,N_13582,N_12546);
nor U19953 (N_19953,N_11076,N_13181);
xor U19954 (N_19954,N_14519,N_13315);
and U19955 (N_19955,N_13183,N_13711);
or U19956 (N_19956,N_10767,N_12236);
nor U19957 (N_19957,N_14822,N_12236);
xor U19958 (N_19958,N_13451,N_13523);
nand U19959 (N_19959,N_11858,N_10503);
nor U19960 (N_19960,N_13058,N_10755);
or U19961 (N_19961,N_10307,N_12854);
or U19962 (N_19962,N_14272,N_14837);
nor U19963 (N_19963,N_10743,N_14456);
or U19964 (N_19964,N_14256,N_13686);
nor U19965 (N_19965,N_13490,N_12859);
nor U19966 (N_19966,N_11021,N_12528);
nand U19967 (N_19967,N_13284,N_12568);
and U19968 (N_19968,N_13088,N_13981);
or U19969 (N_19969,N_14550,N_14439);
nand U19970 (N_19970,N_11608,N_10602);
xor U19971 (N_19971,N_13317,N_10045);
nand U19972 (N_19972,N_12490,N_14793);
and U19973 (N_19973,N_11860,N_10182);
nor U19974 (N_19974,N_12243,N_12045);
xnor U19975 (N_19975,N_12998,N_14538);
nor U19976 (N_19976,N_13999,N_11267);
and U19977 (N_19977,N_11202,N_10549);
nor U19978 (N_19978,N_11261,N_13205);
and U19979 (N_19979,N_10171,N_14990);
and U19980 (N_19980,N_12326,N_11480);
xor U19981 (N_19981,N_13821,N_11151);
nor U19982 (N_19982,N_12133,N_10694);
and U19983 (N_19983,N_13741,N_12339);
nand U19984 (N_19984,N_11307,N_10297);
and U19985 (N_19985,N_10333,N_11768);
nand U19986 (N_19986,N_13251,N_12652);
nand U19987 (N_19987,N_14722,N_10252);
and U19988 (N_19988,N_10742,N_12168);
and U19989 (N_19989,N_13397,N_10753);
nor U19990 (N_19990,N_14062,N_12474);
nor U19991 (N_19991,N_11030,N_13882);
or U19992 (N_19992,N_12262,N_12768);
nand U19993 (N_19993,N_11344,N_13724);
and U19994 (N_19994,N_14918,N_14993);
or U19995 (N_19995,N_10114,N_11104);
and U19996 (N_19996,N_14144,N_14788);
nor U19997 (N_19997,N_11216,N_11599);
nor U19998 (N_19998,N_10650,N_11324);
or U19999 (N_19999,N_10992,N_11547);
nor UO_0 (O_0,N_18939,N_18267);
nor UO_1 (O_1,N_15536,N_15126);
nand UO_2 (O_2,N_18041,N_19322);
or UO_3 (O_3,N_15311,N_15990);
nor UO_4 (O_4,N_17375,N_16513);
and UO_5 (O_5,N_17119,N_15969);
nor UO_6 (O_6,N_17090,N_17561);
and UO_7 (O_7,N_17577,N_19469);
nor UO_8 (O_8,N_16050,N_17579);
and UO_9 (O_9,N_19804,N_16441);
and UO_10 (O_10,N_17804,N_18929);
and UO_11 (O_11,N_15222,N_17947);
nor UO_12 (O_12,N_18729,N_15602);
nand UO_13 (O_13,N_17792,N_15179);
nand UO_14 (O_14,N_15260,N_17278);
or UO_15 (O_15,N_15957,N_17843);
and UO_16 (O_16,N_19766,N_18578);
nand UO_17 (O_17,N_19512,N_18030);
nor UO_18 (O_18,N_16867,N_18474);
nand UO_19 (O_19,N_15944,N_18935);
and UO_20 (O_20,N_17930,N_16192);
nand UO_21 (O_21,N_16484,N_19857);
and UO_22 (O_22,N_15510,N_15921);
or UO_23 (O_23,N_16187,N_16585);
xor UO_24 (O_24,N_17621,N_18287);
nand UO_25 (O_25,N_17218,N_17258);
nor UO_26 (O_26,N_17607,N_17370);
and UO_27 (O_27,N_16046,N_19896);
nand UO_28 (O_28,N_18228,N_19984);
nand UO_29 (O_29,N_15976,N_17540);
or UO_30 (O_30,N_15670,N_19286);
or UO_31 (O_31,N_15967,N_16219);
and UO_32 (O_32,N_19131,N_15011);
xor UO_33 (O_33,N_15893,N_15088);
nor UO_34 (O_34,N_19256,N_17536);
nand UO_35 (O_35,N_18317,N_17475);
nor UO_36 (O_36,N_15265,N_16234);
nor UO_37 (O_37,N_18015,N_15672);
and UO_38 (O_38,N_19353,N_17864);
or UO_39 (O_39,N_15569,N_17973);
and UO_40 (O_40,N_18523,N_16641);
nor UO_41 (O_41,N_15859,N_15480);
or UO_42 (O_42,N_18011,N_19452);
or UO_43 (O_43,N_15800,N_15711);
and UO_44 (O_44,N_15550,N_17886);
nand UO_45 (O_45,N_19156,N_16105);
nand UO_46 (O_46,N_19468,N_15201);
nand UO_47 (O_47,N_18167,N_18599);
or UO_48 (O_48,N_15357,N_15185);
or UO_49 (O_49,N_17147,N_19513);
nand UO_50 (O_50,N_16727,N_17632);
or UO_51 (O_51,N_18942,N_17593);
or UO_52 (O_52,N_16753,N_18581);
xor UO_53 (O_53,N_19503,N_17360);
nor UO_54 (O_54,N_19532,N_15530);
nor UO_55 (O_55,N_15429,N_16704);
nor UO_56 (O_56,N_17736,N_18674);
nor UO_57 (O_57,N_18473,N_18520);
or UO_58 (O_58,N_17247,N_17677);
or UO_59 (O_59,N_16266,N_15998);
or UO_60 (O_60,N_18428,N_16025);
or UO_61 (O_61,N_19367,N_17458);
nand UO_62 (O_62,N_19166,N_18535);
and UO_63 (O_63,N_19244,N_18824);
nor UO_64 (O_64,N_18651,N_19902);
and UO_65 (O_65,N_17887,N_18441);
and UO_66 (O_66,N_16583,N_18775);
or UO_67 (O_67,N_17958,N_15726);
xnor UO_68 (O_68,N_17266,N_16568);
or UO_69 (O_69,N_15235,N_16560);
nand UO_70 (O_70,N_17639,N_19006);
nand UO_71 (O_71,N_19790,N_17200);
or UO_72 (O_72,N_15060,N_15558);
nor UO_73 (O_73,N_18237,N_19674);
and UO_74 (O_74,N_16558,N_18903);
nor UO_75 (O_75,N_19253,N_18146);
and UO_76 (O_76,N_15432,N_17584);
nand UO_77 (O_77,N_16353,N_15067);
nor UO_78 (O_78,N_17707,N_17866);
and UO_79 (O_79,N_17211,N_19356);
and UO_80 (O_80,N_16196,N_16685);
nand UO_81 (O_81,N_19888,N_17327);
nor UO_82 (O_82,N_18077,N_15952);
nand UO_83 (O_83,N_18958,N_15239);
and UO_84 (O_84,N_19912,N_17062);
and UO_85 (O_85,N_17397,N_17992);
xnor UO_86 (O_86,N_19575,N_18984);
and UO_87 (O_87,N_17782,N_16902);
or UO_88 (O_88,N_18005,N_19341);
or UO_89 (O_89,N_18685,N_16162);
nor UO_90 (O_90,N_16080,N_15254);
nand UO_91 (O_91,N_19147,N_19934);
nor UO_92 (O_92,N_17559,N_19894);
nor UO_93 (O_93,N_16709,N_18629);
nand UO_94 (O_94,N_15621,N_18117);
nor UO_95 (O_95,N_19613,N_17869);
and UO_96 (O_96,N_18879,N_16775);
and UO_97 (O_97,N_17092,N_17322);
nor UO_98 (O_98,N_16909,N_16799);
or UO_99 (O_99,N_17784,N_17028);
or UO_100 (O_100,N_17925,N_19714);
or UO_101 (O_101,N_16765,N_17021);
or UO_102 (O_102,N_17957,N_16516);
and UO_103 (O_103,N_16041,N_15308);
and UO_104 (O_104,N_19499,N_15870);
and UO_105 (O_105,N_17588,N_19737);
or UO_106 (O_106,N_17800,N_16414);
and UO_107 (O_107,N_16602,N_18300);
nor UO_108 (O_108,N_15358,N_18573);
or UO_109 (O_109,N_19635,N_15160);
xor UO_110 (O_110,N_19853,N_18512);
or UO_111 (O_111,N_19397,N_15050);
nor UO_112 (O_112,N_19652,N_15001);
or UO_113 (O_113,N_18332,N_18008);
nor UO_114 (O_114,N_19366,N_16142);
nor UO_115 (O_115,N_16331,N_18564);
nor UO_116 (O_116,N_16153,N_19535);
or UO_117 (O_117,N_15455,N_16437);
nor UO_118 (O_118,N_15457,N_15072);
nor UO_119 (O_119,N_16675,N_16169);
nor UO_120 (O_120,N_19660,N_16475);
or UO_121 (O_121,N_16688,N_16469);
nand UO_122 (O_122,N_19205,N_16949);
or UO_123 (O_123,N_18388,N_18736);
or UO_124 (O_124,N_19507,N_16536);
nand UO_125 (O_125,N_15167,N_18088);
nand UO_126 (O_126,N_15137,N_19667);
nand UO_127 (O_127,N_17451,N_15722);
and UO_128 (O_128,N_16999,N_18427);
or UO_129 (O_129,N_19296,N_19325);
nor UO_130 (O_130,N_15594,N_19377);
or UO_131 (O_131,N_19510,N_15792);
and UO_132 (O_132,N_15042,N_17171);
nor UO_133 (O_133,N_15778,N_19424);
xor UO_134 (O_134,N_18432,N_18524);
or UO_135 (O_135,N_17259,N_15400);
and UO_136 (O_136,N_15494,N_18014);
or UO_137 (O_137,N_15693,N_18424);
xor UO_138 (O_138,N_17306,N_15826);
and UO_139 (O_139,N_15350,N_19076);
nor UO_140 (O_140,N_19569,N_17951);
nor UO_141 (O_141,N_19594,N_19907);
and UO_142 (O_142,N_18928,N_19062);
or UO_143 (O_143,N_18807,N_19181);
nor UO_144 (O_144,N_19648,N_19277);
or UO_145 (O_145,N_17042,N_17516);
nor UO_146 (O_146,N_15213,N_19379);
nor UO_147 (O_147,N_16336,N_15718);
or UO_148 (O_148,N_16817,N_17931);
or UO_149 (O_149,N_16600,N_18546);
xnor UO_150 (O_150,N_19347,N_16708);
or UO_151 (O_151,N_16757,N_18101);
nand UO_152 (O_152,N_19772,N_17648);
nor UO_153 (O_153,N_15922,N_17441);
or UO_154 (O_154,N_16253,N_17618);
nor UO_155 (O_155,N_18589,N_19375);
or UO_156 (O_156,N_18197,N_17201);
nor UO_157 (O_157,N_15811,N_17891);
and UO_158 (O_158,N_19485,N_15227);
and UO_159 (O_159,N_19640,N_19793);
nand UO_160 (O_160,N_18349,N_16945);
xor UO_161 (O_161,N_17236,N_16334);
nor UO_162 (O_162,N_19068,N_19935);
nand UO_163 (O_163,N_16029,N_19722);
xor UO_164 (O_164,N_15977,N_15995);
or UO_165 (O_165,N_17146,N_16835);
or UO_166 (O_166,N_15296,N_15272);
xnor UO_167 (O_167,N_18991,N_15393);
xor UO_168 (O_168,N_16185,N_16917);
xor UO_169 (O_169,N_16498,N_17733);
or UO_170 (O_170,N_17275,N_16391);
nand UO_171 (O_171,N_19111,N_15119);
nor UO_172 (O_172,N_19255,N_15698);
nor UO_173 (O_173,N_19559,N_17675);
or UO_174 (O_174,N_15192,N_16190);
and UO_175 (O_175,N_18183,N_18856);
nor UO_176 (O_176,N_18190,N_19762);
and UO_177 (O_177,N_16188,N_19928);
nand UO_178 (O_178,N_17576,N_15053);
and UO_179 (O_179,N_19232,N_16923);
nor UO_180 (O_180,N_16845,N_19583);
nand UO_181 (O_181,N_16718,N_16210);
or UO_182 (O_182,N_18061,N_18464);
nor UO_183 (O_183,N_17606,N_16034);
nand UO_184 (O_184,N_18418,N_18967);
xnor UO_185 (O_185,N_18602,N_16822);
or UO_186 (O_186,N_17646,N_19556);
or UO_187 (O_187,N_15159,N_16309);
or UO_188 (O_188,N_19663,N_18141);
or UO_189 (O_189,N_19415,N_19936);
and UO_190 (O_190,N_15301,N_19291);
or UO_191 (O_191,N_19658,N_18431);
and UO_192 (O_192,N_17603,N_16514);
or UO_193 (O_193,N_18628,N_16293);
nand UO_194 (O_194,N_17227,N_16120);
or UO_195 (O_195,N_18838,N_17741);
and UO_196 (O_196,N_16487,N_19702);
nor UO_197 (O_197,N_16296,N_15626);
nand UO_198 (O_198,N_15405,N_19779);
xnor UO_199 (O_199,N_19701,N_19630);
or UO_200 (O_200,N_19226,N_16150);
nor UO_201 (O_201,N_18849,N_15030);
nor UO_202 (O_202,N_17273,N_17487);
nand UO_203 (O_203,N_18012,N_16154);
and UO_204 (O_204,N_17706,N_16642);
or UO_205 (O_205,N_19242,N_15127);
nand UO_206 (O_206,N_17356,N_18145);
or UO_207 (O_207,N_18569,N_18102);
nand UO_208 (O_208,N_19211,N_18483);
nand UO_209 (O_209,N_16624,N_18983);
or UO_210 (O_210,N_15741,N_18627);
or UO_211 (O_211,N_19519,N_19798);
and UO_212 (O_212,N_17769,N_18703);
and UO_213 (O_213,N_16938,N_18105);
or UO_214 (O_214,N_16399,N_15907);
and UO_215 (O_215,N_17323,N_16337);
or UO_216 (O_216,N_16865,N_18761);
or UO_217 (O_217,N_18953,N_19363);
nor UO_218 (O_218,N_17000,N_18742);
or UO_219 (O_219,N_16065,N_19725);
nor UO_220 (O_220,N_17031,N_18846);
nor UO_221 (O_221,N_18282,N_19267);
nand UO_222 (O_222,N_15679,N_15439);
nor UO_223 (O_223,N_15526,N_17783);
and UO_224 (O_224,N_16995,N_17143);
nor UO_225 (O_225,N_17971,N_15233);
and UO_226 (O_226,N_18710,N_15194);
or UO_227 (O_227,N_17474,N_17043);
nor UO_228 (O_228,N_18809,N_19236);
nor UO_229 (O_229,N_17751,N_19593);
or UO_230 (O_230,N_15568,N_17387);
nand UO_231 (O_231,N_16049,N_18894);
or UO_232 (O_232,N_17531,N_18676);
and UO_233 (O_233,N_16305,N_15168);
and UO_234 (O_234,N_19158,N_16397);
and UO_235 (O_235,N_19830,N_16850);
or UO_236 (O_236,N_19453,N_18469);
or UO_237 (O_237,N_18510,N_15318);
nand UO_238 (O_238,N_16179,N_19838);
or UO_239 (O_239,N_18471,N_18071);
nand UO_240 (O_240,N_18618,N_15292);
nor UO_241 (O_241,N_16117,N_16417);
or UO_242 (O_242,N_18301,N_18962);
nor UO_243 (O_243,N_16479,N_15057);
and UO_244 (O_244,N_19653,N_19247);
or UO_245 (O_245,N_16425,N_16198);
or UO_246 (O_246,N_17354,N_18978);
and UO_247 (O_247,N_18160,N_19116);
and UO_248 (O_248,N_17248,N_15054);
xor UO_249 (O_249,N_19600,N_18611);
nor UO_250 (O_250,N_18373,N_19360);
and UO_251 (O_251,N_17668,N_15863);
or UO_252 (O_252,N_15485,N_15342);
or UO_253 (O_253,N_18749,N_18671);
and UO_254 (O_254,N_19438,N_17877);
nand UO_255 (O_255,N_16904,N_18293);
xnor UO_256 (O_256,N_18539,N_19390);
or UO_257 (O_257,N_17066,N_17312);
nor UO_258 (O_258,N_19066,N_19029);
nor UO_259 (O_259,N_15305,N_18173);
or UO_260 (O_260,N_18166,N_17320);
and UO_261 (O_261,N_15066,N_16956);
nand UO_262 (O_262,N_17009,N_19228);
or UO_263 (O_263,N_15516,N_19125);
and UO_264 (O_264,N_17976,N_16075);
nand UO_265 (O_265,N_17902,N_18188);
and UO_266 (O_266,N_15573,N_19478);
nand UO_267 (O_267,N_17546,N_18501);
or UO_268 (O_268,N_19549,N_16690);
and UO_269 (O_269,N_15195,N_19713);
xnor UO_270 (O_270,N_19840,N_19812);
nor UO_271 (O_271,N_15496,N_19140);
and UO_272 (O_272,N_16459,N_18247);
nor UO_273 (O_273,N_17609,N_18971);
nand UO_274 (O_274,N_15158,N_16400);
nor UO_275 (O_275,N_18381,N_15096);
and UO_276 (O_276,N_18229,N_19774);
nand UO_277 (O_277,N_18369,N_17983);
and UO_278 (O_278,N_18837,N_15788);
or UO_279 (O_279,N_16091,N_19107);
nand UO_280 (O_280,N_17870,N_17928);
or UO_281 (O_281,N_15383,N_16227);
or UO_282 (O_282,N_17879,N_18679);
or UO_283 (O_283,N_17033,N_16106);
nor UO_284 (O_284,N_15370,N_16357);
and UO_285 (O_285,N_16385,N_16355);
nand UO_286 (O_286,N_17113,N_18647);
and UO_287 (O_287,N_18920,N_15263);
nor UO_288 (O_288,N_16754,N_18492);
or UO_289 (O_289,N_16571,N_19686);
and UO_290 (O_290,N_15020,N_19188);
xor UO_291 (O_291,N_15097,N_19588);
nand UO_292 (O_292,N_18205,N_17257);
nand UO_293 (O_293,N_16665,N_17269);
xnor UO_294 (O_294,N_15304,N_18993);
nor UO_295 (O_295,N_19515,N_19173);
nor UO_296 (O_296,N_18514,N_18162);
xor UO_297 (O_297,N_16540,N_19005);
or UO_298 (O_298,N_15970,N_15850);
and UO_299 (O_299,N_19218,N_15356);
xor UO_300 (O_300,N_16032,N_15899);
and UO_301 (O_301,N_19099,N_18482);
nor UO_302 (O_302,N_19446,N_18415);
and UO_303 (O_303,N_19486,N_16736);
nand UO_304 (O_304,N_15106,N_17127);
or UO_305 (O_305,N_19179,N_15047);
nand UO_306 (O_306,N_18147,N_17539);
and UO_307 (O_307,N_19570,N_15366);
nand UO_308 (O_308,N_18495,N_18808);
and UO_309 (O_309,N_15361,N_16705);
nand UO_310 (O_310,N_16378,N_16450);
nand UO_311 (O_311,N_19333,N_19248);
nand UO_312 (O_312,N_15117,N_16166);
nor UO_313 (O_313,N_15663,N_18734);
nor UO_314 (O_314,N_18669,N_15489);
nand UO_315 (O_315,N_16746,N_17328);
and UO_316 (O_316,N_16742,N_19698);
xor UO_317 (O_317,N_16054,N_18263);
and UO_318 (O_318,N_15327,N_18092);
nand UO_319 (O_319,N_19350,N_17154);
nand UO_320 (O_320,N_17221,N_15996);
or UO_321 (O_321,N_16729,N_17348);
nand UO_322 (O_322,N_18989,N_18236);
or UO_323 (O_323,N_18318,N_16647);
nor UO_324 (O_324,N_18787,N_19448);
and UO_325 (O_325,N_18810,N_17187);
and UO_326 (O_326,N_19237,N_18038);
xor UO_327 (O_327,N_17486,N_16189);
and UO_328 (O_328,N_19430,N_17704);
and UO_329 (O_329,N_17595,N_15412);
nor UO_330 (O_330,N_16788,N_15545);
nor UO_331 (O_331,N_16841,N_15759);
xnor UO_332 (O_332,N_15810,N_15680);
nand UO_333 (O_333,N_15343,N_19688);
or UO_334 (O_334,N_18754,N_18766);
nand UO_335 (O_335,N_15593,N_17802);
and UO_336 (O_336,N_18410,N_15026);
or UO_337 (O_337,N_17742,N_16332);
nand UO_338 (O_338,N_17319,N_17903);
and UO_339 (O_339,N_19871,N_15801);
nand UO_340 (O_340,N_16860,N_19887);
nand UO_341 (O_341,N_16934,N_18259);
xnor UO_342 (O_342,N_15320,N_18897);
nand UO_343 (O_343,N_16152,N_17857);
xnor UO_344 (O_344,N_15796,N_16340);
nor UO_345 (O_345,N_18901,N_16930);
nand UO_346 (O_346,N_18299,N_17270);
nor UO_347 (O_347,N_16526,N_19069);
and UO_348 (O_348,N_17461,N_19715);
nand UO_349 (O_349,N_15938,N_15837);
or UO_350 (O_350,N_15328,N_16392);
or UO_351 (O_351,N_18968,N_16172);
nor UO_352 (O_352,N_18047,N_19923);
and UO_353 (O_353,N_18003,N_17238);
nand UO_354 (O_354,N_17940,N_18306);
or UO_355 (O_355,N_15785,N_18178);
and UO_356 (O_356,N_16660,N_18890);
or UO_357 (O_357,N_16952,N_19335);
or UO_358 (O_358,N_15084,N_15075);
nor UO_359 (O_359,N_18574,N_15107);
or UO_360 (O_360,N_16725,N_17768);
nor UO_361 (O_361,N_18600,N_19862);
xnor UO_362 (O_362,N_16456,N_18877);
and UO_363 (O_363,N_18798,N_15755);
nand UO_364 (O_364,N_19345,N_19605);
or UO_365 (O_365,N_17393,N_16766);
and UO_366 (O_366,N_18768,N_16711);
and UO_367 (O_367,N_16460,N_15856);
and UO_368 (O_368,N_18295,N_16001);
nand UO_369 (O_369,N_15184,N_16656);
or UO_370 (O_370,N_15341,N_15884);
and UO_371 (O_371,N_16377,N_18490);
and UO_372 (O_372,N_16070,N_17465);
xnor UO_373 (O_373,N_16100,N_15476);
xor UO_374 (O_374,N_15662,N_19966);
nor UO_375 (O_375,N_17614,N_15094);
and UO_376 (O_376,N_15849,N_15465);
and UO_377 (O_377,N_16811,N_19699);
and UO_378 (O_378,N_19032,N_17206);
or UO_379 (O_379,N_16370,N_17485);
nand UO_380 (O_380,N_18632,N_18379);
or UO_381 (O_381,N_19436,N_16321);
and UO_382 (O_382,N_15068,N_15716);
nand UO_383 (O_383,N_17183,N_18079);
or UO_384 (O_384,N_17529,N_15453);
or UO_385 (O_385,N_16026,N_16300);
or UO_386 (O_386,N_15939,N_15677);
nor UO_387 (O_387,N_17335,N_16416);
or UO_388 (O_388,N_16174,N_19233);
or UO_389 (O_389,N_17608,N_18530);
and UO_390 (O_390,N_17100,N_17933);
or UO_391 (O_391,N_16792,N_17695);
nand UO_392 (O_392,N_19419,N_15620);
and UO_393 (O_393,N_17426,N_18116);
nor UO_394 (O_394,N_17083,N_16202);
nor UO_395 (O_395,N_17845,N_15266);
or UO_396 (O_396,N_16576,N_15157);
or UO_397 (O_397,N_17712,N_18401);
or UO_398 (O_398,N_19839,N_18241);
and UO_399 (O_399,N_17728,N_16206);
and UO_400 (O_400,N_16474,N_15063);
or UO_401 (O_401,N_15277,N_19372);
or UO_402 (O_402,N_16719,N_16243);
or UO_403 (O_403,N_19744,N_19975);
nor UO_404 (O_404,N_15808,N_18653);
and UO_405 (O_405,N_19252,N_18119);
nor UO_406 (O_406,N_18394,N_18786);
nor UO_407 (O_407,N_16298,N_19551);
nor UO_408 (O_408,N_17049,N_17209);
nor UO_409 (O_409,N_17883,N_19500);
or UO_410 (O_410,N_18944,N_15003);
nor UO_411 (O_411,N_18608,N_16078);
nand UO_412 (O_412,N_15388,N_17553);
or UO_413 (O_413,N_18278,N_15232);
xor UO_414 (O_414,N_19108,N_16177);
nand UO_415 (O_415,N_17219,N_18719);
and UO_416 (O_416,N_19059,N_16407);
xor UO_417 (O_417,N_19297,N_15392);
nor UO_418 (O_418,N_19985,N_17650);
nor UO_419 (O_419,N_15431,N_18872);
or UO_420 (O_420,N_17523,N_19691);
nand UO_421 (O_421,N_19773,N_15668);
nor UO_422 (O_422,N_18350,N_15177);
or UO_423 (O_423,N_17024,N_18888);
nor UO_424 (O_424,N_17839,N_16413);
and UO_425 (O_425,N_18018,N_16255);
or UO_426 (O_426,N_19019,N_17509);
nor UO_427 (O_427,N_15210,N_18209);
and UO_428 (O_428,N_19346,N_17019);
or UO_429 (O_429,N_17967,N_17210);
or UO_430 (O_430,N_19796,N_17405);
nor UO_431 (O_431,N_16241,N_17184);
and UO_432 (O_432,N_16804,N_17331);
nor UO_433 (O_433,N_18806,N_15659);
and UO_434 (O_434,N_17350,N_15842);
and UO_435 (O_435,N_16648,N_19083);
and UO_436 (O_436,N_19824,N_17310);
nand UO_437 (O_437,N_15460,N_15614);
or UO_438 (O_438,N_18123,N_17010);
nor UO_439 (O_439,N_15902,N_15943);
nand UO_440 (O_440,N_18399,N_15840);
nor UO_441 (O_441,N_17231,N_16491);
xor UO_442 (O_442,N_16922,N_16988);
and UO_443 (O_443,N_15867,N_17308);
or UO_444 (O_444,N_15329,N_16247);
nor UO_445 (O_445,N_17956,N_19901);
nor UO_446 (O_446,N_16423,N_17084);
and UO_447 (O_447,N_18156,N_15724);
nand UO_448 (O_448,N_15256,N_18334);
nand UO_449 (O_449,N_19842,N_15259);
nand UO_450 (O_450,N_17311,N_15701);
and UO_451 (O_451,N_17916,N_16869);
nand UO_452 (O_452,N_17252,N_16856);
nand UO_453 (O_453,N_19012,N_16424);
or UO_454 (O_454,N_16836,N_16014);
and UO_455 (O_455,N_17108,N_15830);
nand UO_456 (O_456,N_15517,N_16268);
nor UO_457 (O_457,N_19403,N_18750);
nand UO_458 (O_458,N_16489,N_17449);
nor UO_459 (O_459,N_18034,N_18716);
or UO_460 (O_460,N_16135,N_15942);
xor UO_461 (O_461,N_19983,N_16833);
nand UO_462 (O_462,N_18817,N_17279);
nor UO_463 (O_463,N_19542,N_15487);
or UO_464 (O_464,N_18982,N_15686);
nor UO_465 (O_465,N_16104,N_18131);
nand UO_466 (O_466,N_18681,N_19329);
xnor UO_467 (O_467,N_17496,N_15484);
nand UO_468 (O_468,N_19183,N_16477);
or UO_469 (O_469,N_19628,N_18091);
nor UO_470 (O_470,N_15841,N_17798);
nor UO_471 (O_471,N_18276,N_17199);
or UO_472 (O_472,N_18780,N_19293);
or UO_473 (O_473,N_17409,N_18498);
nand UO_474 (O_474,N_19175,N_19268);
nand UO_475 (O_475,N_15869,N_17400);
and UO_476 (O_476,N_17203,N_18743);
nand UO_477 (O_477,N_16567,N_18286);
nor UO_478 (O_478,N_17796,N_19860);
nor UO_479 (O_479,N_18931,N_16672);
xor UO_480 (O_480,N_19023,N_16270);
nand UO_481 (O_481,N_19411,N_16131);
nand UO_482 (O_482,N_18974,N_18258);
nor UO_483 (O_483,N_19258,N_16012);
and UO_484 (O_484,N_15048,N_18217);
nor UO_485 (O_485,N_19449,N_19938);
nand UO_486 (O_486,N_17093,N_16093);
nand UO_487 (O_487,N_18172,N_16271);
nand UO_488 (O_488,N_19201,N_19604);
nor UO_489 (O_489,N_19200,N_17657);
or UO_490 (O_490,N_19475,N_19843);
xnor UO_491 (O_491,N_19127,N_15598);
or UO_492 (O_492,N_16303,N_17503);
or UO_493 (O_493,N_16180,N_19048);
and UO_494 (O_494,N_19877,N_19101);
nor UO_495 (O_495,N_15228,N_17726);
nor UO_496 (O_496,N_19434,N_17686);
nand UO_497 (O_497,N_19321,N_16519);
and UO_498 (O_498,N_19817,N_18717);
nor UO_499 (O_499,N_19493,N_18138);
nand UO_500 (O_500,N_16589,N_19084);
nor UO_501 (O_501,N_17655,N_16073);
and UO_502 (O_502,N_19885,N_19548);
or UO_503 (O_503,N_16452,N_17039);
or UO_504 (O_504,N_16146,N_16318);
nor UO_505 (O_505,N_16593,N_17568);
nand UO_506 (O_506,N_18829,N_16480);
and UO_507 (O_507,N_19882,N_17340);
and UO_508 (O_508,N_17478,N_19832);
or UO_509 (O_509,N_16242,N_18227);
and UO_510 (O_510,N_16977,N_19792);
xor UO_511 (O_511,N_18239,N_17263);
nand UO_512 (O_512,N_18272,N_16927);
and UO_513 (O_513,N_16971,N_17212);
and UO_514 (O_514,N_15171,N_18044);
nor UO_515 (O_515,N_16828,N_18221);
or UO_516 (O_516,N_15139,N_18828);
nand UO_517 (O_517,N_19884,N_15150);
and UO_518 (O_518,N_17790,N_19065);
nor UO_519 (O_519,N_15482,N_19522);
and UO_520 (O_520,N_16992,N_18827);
or UO_521 (O_521,N_16114,N_17388);
nand UO_522 (O_522,N_19903,N_15717);
and UO_523 (O_523,N_17929,N_15447);
nand UO_524 (O_524,N_18916,N_16525);
and UO_525 (O_525,N_18475,N_15984);
or UO_526 (O_526,N_17477,N_19566);
nor UO_527 (O_527,N_19889,N_19310);
and UO_528 (O_528,N_18715,N_15631);
or UO_529 (O_529,N_18556,N_17027);
nor UO_530 (O_530,N_16465,N_18985);
xor UO_531 (O_531,N_18056,N_15008);
and UO_532 (O_532,N_18774,N_19913);
xor UO_533 (O_533,N_16857,N_15086);
nor UO_534 (O_534,N_17437,N_17906);
or UO_535 (O_535,N_19892,N_16053);
or UO_536 (O_536,N_18923,N_18892);
xnor UO_537 (O_537,N_17801,N_15448);
or UO_538 (O_538,N_17109,N_15634);
and UO_539 (O_539,N_15322,N_16249);
and UO_540 (O_540,N_15153,N_18839);
and UO_541 (O_541,N_15035,N_16607);
nand UO_542 (O_542,N_17999,N_17134);
and UO_543 (O_543,N_17436,N_17432);
nor UO_544 (O_544,N_16755,N_15678);
nor UO_545 (O_545,N_17690,N_17394);
or UO_546 (O_546,N_17885,N_18195);
nor UO_547 (O_547,N_18289,N_15622);
xnor UO_548 (O_548,N_19825,N_16699);
and UO_549 (O_549,N_15381,N_15844);
xor UO_550 (O_550,N_17234,N_18850);
nand UO_551 (O_551,N_15949,N_18347);
nor UO_552 (O_552,N_17767,N_17277);
nor UO_553 (O_553,N_18635,N_19137);
nand UO_554 (O_554,N_17589,N_16778);
nand UO_555 (O_555,N_15493,N_15567);
and UO_556 (O_556,N_15860,N_17865);
or UO_557 (O_557,N_18351,N_15131);
or UO_558 (O_558,N_15403,N_15806);
nand UO_559 (O_559,N_16597,N_15528);
nor UO_560 (O_560,N_15772,N_19526);
and UO_561 (O_561,N_18692,N_16052);
nor UO_562 (O_562,N_19965,N_15839);
or UO_563 (O_563,N_15225,N_17103);
and UO_564 (O_564,N_15733,N_15791);
or UO_565 (O_565,N_17991,N_19245);
nand UO_566 (O_566,N_17750,N_19251);
nand UO_567 (O_567,N_16191,N_15878);
xnor UO_568 (O_568,N_18551,N_16214);
nor UO_569 (O_569,N_17285,N_19805);
and UO_570 (O_570,N_17551,N_19246);
nand UO_571 (O_571,N_16329,N_19278);
nand UO_572 (O_572,N_17440,N_18650);
and UO_573 (O_573,N_18057,N_15783);
or UO_574 (O_574,N_17821,N_18438);
nand UO_575 (O_575,N_18848,N_19178);
and UO_576 (O_576,N_19326,N_19053);
or UO_577 (O_577,N_19909,N_16693);
or UO_578 (O_578,N_17452,N_15498);
and UO_579 (O_579,N_18862,N_17734);
and UO_580 (O_580,N_16634,N_16557);
nor UO_581 (O_581,N_17156,N_18112);
xnor UO_582 (O_582,N_17878,N_17274);
nor UO_583 (O_583,N_17115,N_19197);
xnor UO_584 (O_584,N_17402,N_18446);
and UO_585 (O_585,N_15789,N_15348);
nand UO_586 (O_586,N_19868,N_19204);
nor UO_587 (O_587,N_19064,N_17158);
nor UO_588 (O_588,N_19741,N_17890);
nor UO_589 (O_589,N_19481,N_17601);
or UO_590 (O_590,N_15214,N_15803);
or UO_591 (O_591,N_15955,N_17756);
nand UO_592 (O_592,N_19213,N_16295);
and UO_593 (O_593,N_16274,N_18368);
nor UO_594 (O_594,N_19898,N_18309);
nand UO_595 (O_595,N_16759,N_16047);
or UO_596 (O_596,N_17545,N_16269);
nor UO_597 (O_597,N_15339,N_19285);
or UO_598 (O_598,N_15038,N_17052);
and UO_599 (O_599,N_19707,N_16681);
or UO_600 (O_600,N_17046,N_16819);
nand UO_601 (O_601,N_18214,N_17729);
or UO_602 (O_602,N_16712,N_18595);
nor UO_603 (O_603,N_17121,N_18255);
or UO_604 (O_604,N_19539,N_17454);
or UO_605 (O_605,N_16914,N_15190);
nor UO_606 (O_606,N_15845,N_15641);
nand UO_607 (O_607,N_16750,N_16387);
or UO_608 (O_608,N_16854,N_18649);
or UO_609 (O_609,N_18756,N_15317);
or UO_610 (O_610,N_15963,N_18610);
nand UO_611 (O_611,N_16458,N_19269);
nand UO_612 (O_612,N_16967,N_15466);
and UO_613 (O_613,N_18997,N_17223);
and UO_614 (O_614,N_17137,N_19524);
nand UO_615 (O_615,N_18507,N_17722);
nand UO_616 (O_616,N_18323,N_16045);
nand UO_617 (O_617,N_16862,N_17423);
or UO_618 (O_618,N_17530,N_17691);
nor UO_619 (O_619,N_17316,N_18893);
or UO_620 (O_620,N_15384,N_15099);
nor UO_621 (O_621,N_16159,N_19152);
nor UO_622 (O_622,N_17816,N_15876);
or UO_623 (O_623,N_17245,N_19937);
nor UO_624 (O_624,N_18095,N_16211);
and UO_625 (O_625,N_15833,N_19501);
nand UO_626 (O_626,N_18932,N_17989);
nor UO_627 (O_627,N_18238,N_19704);
nor UO_628 (O_628,N_19562,N_17153);
nand UO_629 (O_629,N_18759,N_18840);
or UO_630 (O_630,N_15648,N_18009);
and UO_631 (O_631,N_16530,N_18995);
nor UO_632 (O_632,N_16584,N_18891);
or UO_633 (O_633,N_17959,N_18576);
and UO_634 (O_634,N_19413,N_16731);
nor UO_635 (O_635,N_18370,N_18346);
xor UO_636 (O_636,N_19624,N_18883);
or UO_637 (O_637,N_18531,N_17182);
and UO_638 (O_638,N_17180,N_17721);
nor UO_639 (O_639,N_17372,N_16827);
and UO_640 (O_640,N_18338,N_15278);
nand UO_641 (O_641,N_16951,N_19726);
and UO_642 (O_642,N_18290,N_18362);
and UO_643 (O_643,N_17411,N_16194);
and UO_644 (O_644,N_18555,N_17725);
xnor UO_645 (O_645,N_18051,N_19437);
and UO_646 (O_646,N_19133,N_16622);
and UO_647 (O_647,N_19525,N_17761);
nor UO_648 (O_648,N_15580,N_15290);
or UO_649 (O_649,N_19946,N_18752);
or UO_650 (O_650,N_17280,N_19141);
xor UO_651 (O_651,N_17494,N_18860);
or UO_652 (O_652,N_19564,N_15514);
nand UO_653 (O_653,N_16851,N_19264);
nand UO_654 (O_654,N_19121,N_15694);
nand UO_655 (O_655,N_18665,N_15426);
and UO_656 (O_656,N_17597,N_16082);
or UO_657 (O_657,N_17346,N_16373);
or UO_658 (O_658,N_18284,N_15502);
and UO_659 (O_659,N_19599,N_19775);
nor UO_660 (O_660,N_18517,N_18788);
and UO_661 (O_661,N_16215,N_19915);
xnor UO_662 (O_662,N_18296,N_16145);
or UO_663 (O_663,N_16950,N_16763);
nand UO_664 (O_664,N_15874,N_16698);
and UO_665 (O_665,N_16116,N_15597);
nand UO_666 (O_666,N_16134,N_17057);
xor UO_667 (O_667,N_17949,N_16842);
nand UO_668 (O_668,N_17442,N_17484);
xnor UO_669 (O_669,N_15972,N_18212);
and UO_670 (O_670,N_15832,N_17235);
nor UO_671 (O_671,N_16156,N_17082);
nor UO_672 (O_672,N_15243,N_19785);
or UO_673 (O_673,N_18181,N_17829);
or UO_674 (O_674,N_18782,N_15034);
nor UO_675 (O_675,N_17631,N_18853);
and UO_676 (O_676,N_19122,N_18082);
nor UO_677 (O_677,N_19727,N_19060);
nand UO_678 (O_678,N_16734,N_19550);
or UO_679 (O_679,N_17177,N_15334);
nor UO_680 (O_680,N_16982,N_16533);
xor UO_681 (O_681,N_17538,N_19011);
and UO_682 (O_682,N_18733,N_16896);
or UO_683 (O_683,N_16535,N_15182);
and UO_684 (O_684,N_19738,N_15111);
nand UO_685 (O_685,N_19948,N_15398);
nand UO_686 (O_686,N_19344,N_19338);
or UO_687 (O_687,N_16733,N_16216);
nand UO_688 (O_688,N_16859,N_16954);
or UO_689 (O_689,N_15461,N_16010);
or UO_690 (O_690,N_19459,N_15611);
and UO_691 (O_691,N_16879,N_15234);
nand UO_692 (O_692,N_17026,N_19135);
or UO_693 (O_693,N_17242,N_15275);
and UO_694 (O_694,N_19638,N_16148);
and UO_695 (O_695,N_19052,N_15113);
nor UO_696 (O_696,N_16259,N_15414);
xnor UO_697 (O_697,N_17634,N_17667);
and UO_698 (O_698,N_17995,N_18367);
or UO_699 (O_699,N_15515,N_19538);
or UO_700 (O_700,N_16651,N_18330);
or UO_701 (O_701,N_19088,N_19279);
nor UO_702 (O_702,N_17993,N_15492);
or UO_703 (O_703,N_16668,N_18244);
nor UO_704 (O_704,N_17016,N_18233);
nor UO_705 (O_705,N_19180,N_18844);
nor UO_706 (O_706,N_17738,N_16640);
nand UO_707 (O_707,N_16213,N_18407);
nor UO_708 (O_708,N_15617,N_16611);
xnor UO_709 (O_709,N_15813,N_16072);
nand UO_710 (O_710,N_18084,N_18053);
and UO_711 (O_711,N_18478,N_19273);
or UO_712 (O_712,N_15787,N_15572);
and UO_713 (O_713,N_17944,N_17382);
and UO_714 (O_714,N_15653,N_17481);
and UO_715 (O_715,N_18508,N_19890);
or UO_716 (O_716,N_19646,N_17564);
or UO_717 (O_717,N_19138,N_19846);
or UO_718 (O_718,N_15959,N_17264);
and UO_719 (O_719,N_17915,N_17166);
nor UO_720 (O_720,N_15206,N_17932);
nor UO_721 (O_721,N_19040,N_19466);
xor UO_722 (O_722,N_18880,N_15240);
or UO_723 (O_723,N_17445,N_18680);
or UO_724 (O_724,N_16101,N_18143);
and UO_725 (O_725,N_17367,N_18919);
nor UO_726 (O_726,N_17169,N_17662);
and UO_727 (O_727,N_19378,N_15186);
or UO_728 (O_728,N_18273,N_16591);
nor UO_729 (O_729,N_17378,N_17291);
nor UO_730 (O_730,N_15121,N_19159);
and UO_731 (O_731,N_19465,N_19261);
nor UO_732 (O_732,N_16825,N_16898);
or UO_733 (O_733,N_19536,N_15851);
nand UO_734 (O_734,N_16223,N_15132);
nor UO_735 (O_735,N_19708,N_18500);
nand UO_736 (O_736,N_18857,N_19754);
or UO_737 (O_737,N_15176,N_16657);
or UO_738 (O_738,N_17731,N_18909);
nand UO_739 (O_739,N_16884,N_18193);
nor UO_740 (O_740,N_16590,N_16887);
or UO_741 (O_741,N_17600,N_17532);
nor UO_742 (O_742,N_19953,N_16881);
nor UO_743 (O_743,N_15422,N_16885);
or UO_744 (O_744,N_18460,N_19852);
nor UO_745 (O_745,N_15689,N_15207);
or UO_746 (O_746,N_16615,N_19129);
and UO_747 (O_747,N_16261,N_16979);
or UO_748 (O_748,N_15401,N_18470);
or UO_749 (O_749,N_18072,N_18966);
and UO_750 (O_750,N_15760,N_16931);
or UO_751 (O_751,N_17427,N_18873);
or UO_752 (O_752,N_19456,N_18922);
and UO_753 (O_753,N_19308,N_18662);
nand UO_754 (O_754,N_17766,N_17840);
nor UO_755 (O_755,N_16126,N_17665);
and UO_756 (O_756,N_17927,N_15005);
and UO_757 (O_757,N_18972,N_17160);
xor UO_758 (O_758,N_15781,N_15574);
nor UO_759 (O_759,N_16451,N_16312);
and UO_760 (O_760,N_15525,N_16447);
nor UO_761 (O_761,N_15604,N_18973);
nand UO_762 (O_762,N_16273,N_17628);
nor UO_763 (O_763,N_16960,N_15032);
nor UO_764 (O_764,N_16978,N_18876);
nand UO_765 (O_765,N_15793,N_16741);
or UO_766 (O_766,N_17806,N_17110);
nand UO_767 (O_767,N_19949,N_19093);
or UO_768 (O_768,N_17926,N_16511);
xnor UO_769 (O_769,N_15576,N_16411);
nand UO_770 (O_770,N_15377,N_19492);
nand UO_771 (O_771,N_19899,N_17699);
or UO_772 (O_772,N_16092,N_15188);
nand UO_773 (O_773,N_18636,N_18176);
nor UO_774 (O_774,N_17168,N_19970);
or UO_775 (O_775,N_15421,N_16044);
nand UO_776 (O_776,N_16360,N_17975);
nor UO_777 (O_777,N_15387,N_16028);
nand UO_778 (O_778,N_18479,N_18693);
or UO_779 (O_779,N_17172,N_18675);
or UO_780 (O_780,N_18663,N_18519);
or UO_781 (O_781,N_19835,N_16412);
or UO_782 (O_782,N_18220,N_18961);
nand UO_783 (O_783,N_19078,N_16311);
nor UO_784 (O_784,N_15506,N_18792);
nor UO_785 (O_785,N_16015,N_18121);
and UO_786 (O_786,N_17643,N_17313);
and UO_787 (O_787,N_18938,N_16575);
nor UO_788 (O_788,N_15173,N_18137);
xnor UO_789 (O_789,N_15581,N_15989);
nor UO_790 (O_790,N_18136,N_19304);
or UO_791 (O_791,N_15202,N_19607);
nor UO_792 (O_792,N_19495,N_19855);
xor UO_793 (O_793,N_18593,N_17611);
nor UO_794 (O_794,N_16061,N_19900);
xor UO_795 (O_795,N_18385,N_19747);
nor UO_796 (O_796,N_15051,N_19721);
xor UO_797 (O_797,N_16715,N_17626);
nor UO_798 (O_798,N_17048,N_15508);
and UO_799 (O_799,N_15960,N_18887);
nand UO_800 (O_800,N_15036,N_17735);
nand UO_801 (O_801,N_16383,N_19540);
or UO_802 (O_802,N_17988,N_15671);
or UO_803 (O_803,N_19886,N_17408);
nor UO_804 (O_804,N_18731,N_17353);
and UO_805 (O_805,N_15300,N_17953);
nand UO_806 (O_806,N_16739,N_16663);
nand UO_807 (O_807,N_16779,N_18924);
or UO_808 (O_808,N_17703,N_17747);
and UO_809 (O_809,N_18250,N_17006);
and UO_810 (O_810,N_16201,N_15913);
and UO_811 (O_811,N_15299,N_18561);
and UO_812 (O_812,N_15865,N_18818);
and UO_813 (O_813,N_16580,N_15843);
or UO_814 (O_814,N_19207,N_17471);
nand UO_815 (O_815,N_15436,N_15782);
nand UO_816 (O_816,N_18527,N_18403);
or UO_817 (O_817,N_16024,N_16007);
and UO_818 (O_818,N_19265,N_15091);
or UO_819 (O_819,N_17102,N_17262);
nor UO_820 (O_820,N_18843,N_15479);
nand UO_821 (O_821,N_18149,N_17661);
nor UO_822 (O_822,N_17326,N_17364);
nand UO_823 (O_823,N_19621,N_18398);
nor UO_824 (O_824,N_15629,N_17900);
and UO_825 (O_825,N_19417,N_19553);
or UO_826 (O_826,N_19927,N_19637);
xnor UO_827 (O_827,N_16097,N_15979);
xnor UO_828 (O_828,N_17499,N_17142);
and UO_829 (O_829,N_19401,N_17041);
and UO_830 (O_830,N_17068,N_17345);
and UO_831 (O_831,N_15561,N_18869);
nor UO_832 (O_832,N_18965,N_19429);
and UO_833 (O_833,N_19447,N_19420);
nand UO_834 (O_834,N_17811,N_17076);
nand UO_835 (O_835,N_19893,N_16434);
nor UO_836 (O_836,N_16351,N_15002);
and UO_837 (O_837,N_18712,N_15340);
or UO_838 (O_838,N_16791,N_17910);
or UO_839 (O_839,N_17133,N_19933);
nor UO_840 (O_840,N_15566,N_15014);
and UO_841 (O_841,N_17760,N_16504);
nand UO_842 (O_842,N_18525,N_17012);
nor UO_843 (O_843,N_19314,N_15413);
nor UO_844 (O_844,N_15537,N_18025);
nand UO_845 (O_845,N_16359,N_15746);
nor UO_846 (O_846,N_18337,N_15238);
nand UO_847 (O_847,N_15258,N_16144);
and UO_848 (O_848,N_15083,N_15302);
and UO_849 (O_849,N_17859,N_16631);
and UO_850 (O_850,N_17164,N_19193);
xor UO_851 (O_851,N_15993,N_17254);
nor UO_852 (O_852,N_16022,N_16740);
and UO_853 (O_853,N_17085,N_16772);
nor UO_854 (O_854,N_17038,N_18819);
xnor UO_855 (O_855,N_16846,N_18981);
nand UO_856 (O_856,N_16390,N_16366);
nor UO_857 (O_857,N_17619,N_16524);
or UO_858 (O_858,N_17265,N_19306);
nand UO_859 (O_859,N_18702,N_18861);
nand UO_860 (O_860,N_17309,N_17620);
or UO_861 (O_861,N_19262,N_18927);
nand UO_862 (O_862,N_18537,N_19027);
or UO_863 (O_863,N_15438,N_15369);
xor UO_864 (O_864,N_17352,N_19216);
or UO_865 (O_865,N_16071,N_16866);
nor UO_866 (O_866,N_18764,N_19581);
and UO_867 (O_867,N_19826,N_19587);
or UO_868 (O_868,N_17613,N_18055);
and UO_869 (O_869,N_17053,N_18324);
nor UO_870 (O_870,N_15070,N_15090);
xnor UO_871 (O_871,N_18040,N_15122);
nand UO_872 (O_872,N_19263,N_16232);
nor UO_873 (O_873,N_15244,N_19491);
nand UO_874 (O_874,N_18421,N_17193);
or UO_875 (O_875,N_18592,N_16356);
and UO_876 (O_876,N_15293,N_19557);
and UO_877 (O_877,N_16111,N_17519);
or UO_878 (O_878,N_17851,N_16875);
nor UO_879 (O_879,N_15471,N_19412);
xnor UO_880 (O_880,N_18128,N_17457);
or UO_881 (O_881,N_19971,N_15961);
nor UO_882 (O_882,N_15615,N_17863);
or UO_883 (O_883,N_15805,N_17963);
or UO_884 (O_884,N_15064,N_15100);
xor UO_885 (O_885,N_19117,N_18127);
and UO_886 (O_886,N_15916,N_16448);
nor UO_887 (O_887,N_19967,N_16581);
nand UO_888 (O_888,N_17152,N_19608);
and UO_889 (O_889,N_19703,N_16031);
nand UO_890 (O_890,N_17939,N_19545);
xnor UO_891 (O_891,N_16774,N_17037);
or UO_892 (O_892,N_15822,N_16962);
nand UO_893 (O_893,N_15149,N_18579);
or UO_894 (O_894,N_17842,N_15868);
nor UO_895 (O_895,N_19324,N_19003);
or UO_896 (O_896,N_19631,N_15284);
nor UO_897 (O_897,N_19103,N_18387);
nand UO_898 (O_898,N_16601,N_18371);
nand UO_899 (O_899,N_15740,N_16522);
and UO_900 (O_900,N_19656,N_18670);
or UO_901 (O_901,N_17497,N_19739);
or UO_902 (O_902,N_17054,N_16803);
nand UO_903 (O_903,N_16816,N_18226);
nand UO_904 (O_904,N_16129,N_19736);
nor UO_905 (O_905,N_17656,N_17466);
nor UO_906 (O_906,N_19845,N_16900);
and UO_907 (O_907,N_19655,N_16807);
nand UO_908 (O_908,N_18312,N_15468);
and UO_909 (O_909,N_16421,N_18557);
nand UO_910 (O_910,N_18080,N_18455);
or UO_911 (O_911,N_15777,N_15910);
nor UO_912 (O_912,N_17293,N_19085);
and UO_913 (O_913,N_18686,N_19471);
nand UO_914 (O_914,N_16067,N_16937);
or UO_915 (O_915,N_16002,N_16362);
nand UO_916 (O_916,N_15853,N_18090);
nand UO_917 (O_917,N_18447,N_16810);
nor UO_918 (O_918,N_16762,N_19482);
xor UO_919 (O_919,N_19870,N_18397);
nand UO_920 (O_920,N_16652,N_15497);
or UO_921 (O_921,N_17094,N_18165);
nor UO_922 (O_922,N_16163,N_17982);
or UO_923 (O_923,N_19765,N_19488);
nand UO_924 (O_924,N_19982,N_17758);
xor UO_925 (O_925,N_16785,N_19298);
nor UO_926 (O_926,N_19844,N_17174);
and UO_927 (O_927,N_16099,N_17089);
nand UO_928 (O_928,N_19235,N_18654);
and UO_929 (O_929,N_17654,N_18821);
nor UO_930 (O_930,N_19786,N_15028);
or UO_931 (O_931,N_17954,N_18245);
nor UO_932 (O_932,N_15434,N_17913);
or UO_933 (O_933,N_18321,N_18687);
nand UO_934 (O_934,N_19756,N_19386);
or UO_935 (O_935,N_16471,N_17711);
nand UO_936 (O_936,N_15344,N_16770);
and UO_937 (O_937,N_16798,N_15773);
nor UO_938 (O_938,N_19091,N_18776);
or UO_939 (O_939,N_19561,N_15061);
or UO_940 (O_940,N_16673,N_19171);
and UO_941 (O_941,N_17856,N_19584);
and UO_942 (O_942,N_16409,N_15307);
nand UO_943 (O_943,N_18964,N_19976);
nand UO_944 (O_944,N_18035,N_16051);
nor UO_945 (O_945,N_19502,N_17622);
or UO_946 (O_946,N_17424,N_17398);
nor UO_947 (O_947,N_15691,N_19506);
nor UO_948 (O_948,N_18210,N_15221);
and UO_949 (O_949,N_15744,N_18718);
nor UO_950 (O_950,N_15565,N_17329);
or UO_951 (O_951,N_18078,N_17379);
nor UO_952 (O_952,N_15303,N_17687);
nor UO_953 (O_953,N_19941,N_17482);
and UO_954 (O_954,N_15128,N_15769);
or UO_955 (O_955,N_18074,N_16874);
nand UO_956 (O_956,N_18601,N_18148);
nor UO_957 (O_957,N_16199,N_16961);
xor UO_958 (O_958,N_19980,N_19911);
nor UO_959 (O_959,N_17923,N_18449);
and UO_960 (O_960,N_17197,N_15347);
nand UO_961 (O_961,N_19611,N_17087);
and UO_962 (O_962,N_17537,N_18322);
nor UO_963 (O_963,N_19645,N_18913);
nor UO_964 (O_964,N_18832,N_15282);
or UO_965 (O_965,N_17765,N_17443);
xnor UO_966 (O_966,N_15660,N_19051);
or UO_967 (O_967,N_16604,N_16569);
nand UO_968 (O_968,N_18187,N_17159);
xor UO_969 (O_969,N_15987,N_15423);
and UO_970 (O_970,N_15854,N_18307);
or UO_971 (O_971,N_17222,N_17501);
nor UO_972 (O_972,N_18831,N_18115);
and UO_973 (O_973,N_16292,N_18185);
nor UO_974 (O_974,N_16928,N_19977);
or UO_975 (O_975,N_18028,N_16280);
nand UO_976 (O_976,N_17853,N_17363);
and UO_977 (O_977,N_18643,N_16861);
nand UO_978 (O_978,N_17091,N_17753);
and UO_979 (O_979,N_18534,N_16710);
or UO_980 (O_980,N_17938,N_18700);
or UO_981 (O_981,N_18484,N_19187);
xnor UO_982 (O_982,N_16908,N_18615);
nor UO_983 (O_983,N_18936,N_18854);
nand UO_984 (O_984,N_15473,N_16468);
or UO_985 (O_985,N_19202,N_16218);
or UO_986 (O_986,N_15931,N_15991);
or UO_987 (O_987,N_16103,N_19167);
and UO_988 (O_988,N_16233,N_16574);
and UO_989 (O_989,N_16855,N_17895);
nand UO_990 (O_990,N_15080,N_15009);
and UO_991 (O_991,N_19633,N_17435);
or UO_992 (O_992,N_16618,N_19579);
or UO_993 (O_993,N_18256,N_15872);
or UO_994 (O_994,N_15864,N_17841);
or UO_995 (O_995,N_18660,N_15105);
and UO_996 (O_996,N_16496,N_19661);
and UO_997 (O_997,N_15021,N_15951);
nor UO_998 (O_998,N_18915,N_19283);
and UO_999 (O_999,N_18157,N_19874);
nand UO_1000 (O_1000,N_18728,N_16130);
nand UO_1001 (O_1001,N_17521,N_17852);
and UO_1002 (O_1002,N_18815,N_17749);
and UO_1003 (O_1003,N_15390,N_15603);
nand UO_1004 (O_1004,N_17799,N_16614);
nand UO_1005 (O_1005,N_19063,N_17253);
or UO_1006 (O_1006,N_15973,N_18029);
nor UO_1007 (O_1007,N_17653,N_16443);
nor UO_1008 (O_1008,N_18667,N_18572);
or UO_1009 (O_1009,N_15948,N_17128);
or UO_1010 (O_1010,N_18100,N_16445);
nand UO_1011 (O_1011,N_16483,N_15950);
nor UO_1012 (O_1012,N_15203,N_19381);
and UO_1013 (O_1013,N_18956,N_19476);
and UO_1014 (O_1014,N_15470,N_17190);
nand UO_1015 (O_1015,N_18885,N_17566);
nor UO_1016 (O_1016,N_19694,N_18992);
nand UO_1017 (O_1017,N_18170,N_16283);
nor UO_1018 (O_1018,N_15607,N_18213);
or UO_1019 (O_1019,N_17506,N_19816);
xor UO_1020 (O_1020,N_17381,N_19473);
nor UO_1021 (O_1021,N_17846,N_17934);
nor UO_1022 (O_1022,N_17358,N_19305);
or UO_1023 (O_1023,N_19119,N_16876);
xnor UO_1024 (O_1024,N_17649,N_18277);
and UO_1025 (O_1025,N_19879,N_19533);
nand UO_1026 (O_1026,N_17255,N_15015);
and UO_1027 (O_1027,N_19730,N_18243);
nor UO_1028 (O_1028,N_19568,N_18594);
nand UO_1029 (O_1029,N_16771,N_18232);
nor UO_1030 (O_1030,N_16911,N_18159);
or UO_1031 (O_1031,N_16905,N_16840);
or UO_1032 (O_1032,N_19384,N_15481);
nor UO_1033 (O_1033,N_19861,N_15505);
nor UO_1034 (O_1034,N_19172,N_19169);
xor UO_1035 (O_1035,N_16784,N_18262);
nand UO_1036 (O_1036,N_16888,N_17535);
nand UO_1037 (O_1037,N_17698,N_17357);
or UO_1038 (O_1038,N_15041,N_18358);
nor UO_1039 (O_1039,N_17120,N_15823);
xor UO_1040 (O_1040,N_16780,N_19990);
nand UO_1041 (O_1041,N_17826,N_17338);
or UO_1042 (O_1042,N_16848,N_16873);
or UO_1043 (O_1043,N_16358,N_18563);
and UO_1044 (O_1044,N_18467,N_18779);
nor UO_1045 (O_1045,N_19209,N_19951);
or UO_1046 (O_1046,N_19385,N_19734);
nand UO_1047 (O_1047,N_19394,N_19102);
and UO_1048 (O_1048,N_15966,N_18491);
nand UO_1049 (O_1049,N_18253,N_15136);
xor UO_1050 (O_1050,N_15601,N_16981);
nand UO_1051 (O_1051,N_15108,N_18158);
and UO_1052 (O_1052,N_15046,N_18739);
nand UO_1053 (O_1053,N_18658,N_17779);
and UO_1054 (O_1054,N_19398,N_19257);
or UO_1055 (O_1055,N_17237,N_19170);
nor UO_1056 (O_1056,N_19644,N_16003);
nor UO_1057 (O_1057,N_16683,N_16493);
nor UO_1058 (O_1058,N_16212,N_18612);
nand UO_1059 (O_1059,N_19259,N_16346);
nand UO_1060 (O_1060,N_18976,N_19778);
nor UO_1061 (O_1061,N_19272,N_16700);
nand UO_1062 (O_1062,N_19072,N_19497);
xor UO_1063 (O_1063,N_19318,N_18225);
and UO_1064 (O_1064,N_17610,N_18544);
nor UO_1065 (O_1065,N_17542,N_19336);
xnor UO_1066 (O_1066,N_18999,N_16619);
nor UO_1067 (O_1067,N_19602,N_18064);
nand UO_1068 (O_1068,N_18722,N_19511);
or UO_1069 (O_1069,N_18582,N_19303);
and UO_1070 (O_1070,N_16320,N_15512);
nand UO_1071 (O_1071,N_17283,N_15467);
xnor UO_1072 (O_1072,N_17290,N_19595);
or UO_1073 (O_1073,N_16069,N_19837);
and UO_1074 (O_1074,N_19368,N_17463);
or UO_1075 (O_1075,N_15695,N_19120);
or UO_1076 (O_1076,N_19742,N_17456);
or UO_1077 (O_1077,N_16815,N_15591);
or UO_1078 (O_1078,N_19797,N_18625);
nand UO_1079 (O_1079,N_19254,N_19388);
or UO_1080 (O_1080,N_16279,N_19565);
or UO_1081 (O_1081,N_19761,N_19460);
and UO_1082 (O_1082,N_17702,N_18437);
or UO_1083 (O_1083,N_17544,N_16124);
nor UO_1084 (O_1084,N_18814,N_18395);
and UO_1085 (O_1085,N_17230,N_16276);
nand UO_1086 (O_1086,N_16363,N_17685);
nor UO_1087 (O_1087,N_19225,N_16847);
nor UO_1088 (O_1088,N_17970,N_17630);
and UO_1089 (O_1089,N_17555,N_16983);
nand UO_1090 (O_1090,N_16349,N_19618);
nor UO_1091 (O_1091,N_15650,N_17145);
nor UO_1092 (O_1092,N_18292,N_19030);
nor UO_1093 (O_1093,N_19361,N_15273);
xnor UO_1094 (O_1094,N_17696,N_15555);
or UO_1095 (O_1095,N_15940,N_15287);
nand UO_1096 (O_1096,N_18746,N_16401);
nand UO_1097 (O_1097,N_19528,N_19319);
or UO_1098 (O_1098,N_17965,N_16208);
and UO_1099 (O_1099,N_19118,N_18949);
or UO_1100 (O_1100,N_15045,N_19036);
or UO_1101 (O_1101,N_19109,N_17151);
or UO_1102 (O_1102,N_17228,N_15682);
nor UO_1103 (O_1103,N_17605,N_16327);
nor UO_1104 (O_1104,N_19718,N_19710);
nor UO_1105 (O_1105,N_15771,N_19044);
nand UO_1106 (O_1106,N_15352,N_19355);
nand UO_1107 (O_1107,N_15335,N_17977);
and UO_1108 (O_1108,N_15135,N_18314);
or UO_1109 (O_1109,N_16630,N_16786);
nand UO_1110 (O_1110,N_15880,N_18269);
or UO_1111 (O_1111,N_16714,N_17148);
nor UO_1112 (O_1112,N_15151,N_15570);
nand UO_1113 (O_1113,N_17583,N_16863);
xor UO_1114 (O_1114,N_18777,N_17179);
nor UO_1115 (O_1115,N_19589,N_16143);
and UO_1116 (O_1116,N_15205,N_15669);
nor UO_1117 (O_1117,N_19776,N_17762);
or UO_1118 (O_1118,N_15495,N_19794);
nor UO_1119 (O_1119,N_15640,N_17717);
or UO_1120 (O_1120,N_17492,N_15885);
and UO_1121 (O_1121,N_15606,N_15799);
nand UO_1122 (O_1122,N_16546,N_17590);
nand UO_1123 (O_1123,N_16467,N_15123);
nor UO_1124 (O_1124,N_15013,N_17410);
and UO_1125 (O_1125,N_16415,N_16616);
xor UO_1126 (O_1126,N_16079,N_15037);
nor UO_1127 (O_1127,N_15587,N_19294);
nor UO_1128 (O_1128,N_15163,N_18450);
nand UO_1129 (O_1129,N_17421,N_17414);
and UO_1130 (O_1130,N_15786,N_15719);
nor UO_1131 (O_1131,N_15862,N_15827);
nand UO_1132 (O_1132,N_19194,N_18357);
and UO_1133 (O_1133,N_17337,N_16564);
nor UO_1134 (O_1134,N_19827,N_15418);
and UO_1135 (O_1135,N_16021,N_15198);
and UO_1136 (O_1136,N_17663,N_19657);
and UO_1137 (O_1137,N_19537,N_17061);
and UO_1138 (O_1138,N_17282,N_17292);
and UO_1139 (O_1139,N_15816,N_18083);
nor UO_1140 (O_1140,N_16226,N_18881);
nand UO_1141 (O_1141,N_18476,N_19978);
xnor UO_1142 (O_1142,N_18930,N_17528);
or UO_1143 (O_1143,N_17808,N_19477);
nor UO_1144 (O_1144,N_15349,N_18753);
or UO_1145 (O_1145,N_16446,N_19800);
or UO_1146 (O_1146,N_18740,N_17476);
or UO_1147 (O_1147,N_16793,N_19523);
xor UO_1148 (O_1148,N_17377,N_16543);
nor UO_1149 (O_1149,N_17838,N_18032);
nand UO_1150 (O_1150,N_15743,N_15824);
and UO_1151 (O_1151,N_18865,N_19625);
and UO_1152 (O_1152,N_15217,N_16882);
or UO_1153 (O_1153,N_16402,N_17905);
nand UO_1154 (O_1154,N_16666,N_18230);
nand UO_1155 (O_1155,N_18585,N_15655);
or UO_1156 (O_1156,N_15204,N_16674);
or UO_1157 (O_1157,N_17683,N_15118);
xnor UO_1158 (O_1158,N_16453,N_18070);
or UO_1159 (O_1159,N_19328,N_15742);
nor UO_1160 (O_1160,N_18094,N_16702);
nand UO_1161 (O_1161,N_17718,N_18355);
nor UO_1162 (O_1162,N_16997,N_17395);
nand UO_1163 (O_1163,N_19028,N_16586);
nor UO_1164 (O_1164,N_15410,N_19757);
and UO_1165 (O_1165,N_16545,N_19994);
xnor UO_1166 (O_1166,N_18354,N_19190);
nand UO_1167 (O_1167,N_18639,N_19664);
nand UO_1168 (O_1168,N_18058,N_17719);
or UO_1169 (O_1169,N_15714,N_19284);
nand UO_1170 (O_1170,N_15642,N_19639);
or UO_1171 (O_1171,N_15483,N_18462);
or UO_1172 (O_1172,N_19567,N_17256);
nor UO_1173 (O_1173,N_15533,N_19461);
xor UO_1174 (O_1174,N_16935,N_16095);
nand UO_1175 (O_1175,N_15624,N_15676);
and UO_1176 (O_1176,N_15802,N_16537);
and UO_1177 (O_1177,N_15115,N_17155);
or UO_1178 (O_1178,N_15855,N_17195);
nor UO_1179 (O_1179,N_18360,N_18313);
nor UO_1180 (O_1180,N_19416,N_18619);
nand UO_1181 (O_1181,N_19791,N_17961);
nand UO_1182 (O_1182,N_18506,N_19910);
nor UO_1183 (O_1183,N_18098,N_18445);
xor UO_1184 (O_1184,N_15720,N_15362);
nor UO_1185 (O_1185,N_17889,N_16921);
nor UO_1186 (O_1186,N_16433,N_15231);
and UO_1187 (O_1187,N_16039,N_19441);
and UO_1188 (O_1188,N_16542,N_18270);
and UO_1189 (O_1189,N_19208,N_17185);
or UO_1190 (O_1190,N_19196,N_17070);
or UO_1191 (O_1191,N_16431,N_17640);
nor UO_1192 (O_1192,N_16203,N_17510);
and UO_1193 (O_1193,N_17772,N_16244);
nand UO_1194 (O_1194,N_15215,N_18004);
and UO_1195 (O_1195,N_18023,N_15945);
nor UO_1196 (O_1196,N_19856,N_16167);
nand UO_1197 (O_1197,N_17815,N_17918);
nand UO_1198 (O_1198,N_15723,N_18603);
nor UO_1199 (O_1199,N_17480,N_16588);
nand UO_1200 (O_1200,N_19299,N_15029);
or UO_1201 (O_1201,N_18908,N_16508);
nand UO_1202 (O_1202,N_15911,N_15252);
nand UO_1203 (O_1203,N_19153,N_15351);
and UO_1204 (O_1204,N_18198,N_15557);
nor UO_1205 (O_1205,N_18565,N_18336);
or UO_1206 (O_1206,N_18513,N_19365);
xor UO_1207 (O_1207,N_15763,N_15459);
nor UO_1208 (O_1208,N_16181,N_16968);
and UO_1209 (O_1209,N_17596,N_17533);
and UO_1210 (O_1210,N_18713,N_19222);
nor UO_1211 (O_1211,N_16991,N_19300);
and UO_1212 (O_1212,N_15968,N_18024);
nor UO_1213 (O_1213,N_17260,N_17888);
or UO_1214 (O_1214,N_17994,N_18043);
nand UO_1215 (O_1215,N_19875,N_19391);
and UO_1216 (O_1216,N_15588,N_16472);
nand UO_1217 (O_1217,N_16787,N_17462);
nor UO_1218 (O_1218,N_17178,N_19918);
or UO_1219 (O_1219,N_16209,N_17937);
or UO_1220 (O_1220,N_16517,N_16238);
nor UO_1221 (O_1221,N_15404,N_18502);
or UO_1222 (O_1222,N_19315,N_18268);
and UO_1223 (O_1223,N_15129,N_18863);
nor UO_1224 (O_1224,N_16565,N_18580);
or UO_1225 (O_1225,N_18553,N_16752);
and UO_1226 (O_1226,N_19115,N_18652);
and UO_1227 (O_1227,N_15897,N_15437);
nor UO_1228 (O_1228,N_15656,N_18182);
nor UO_1229 (O_1229,N_18103,N_16119);
and UO_1230 (O_1230,N_16654,N_15109);
nand UO_1231 (O_1231,N_18027,N_19867);
nor UO_1232 (O_1232,N_16379,N_19709);
nor UO_1233 (O_1233,N_17448,N_16371);
and UO_1234 (O_1234,N_18677,N_19920);
nor UO_1235 (O_1235,N_18408,N_18532);
and UO_1236 (O_1236,N_18917,N_15541);
nand UO_1237 (O_1237,N_19097,N_17715);
and UO_1238 (O_1238,N_17612,N_17518);
xor UO_1239 (O_1239,N_18720,N_19212);
or UO_1240 (O_1240,N_18216,N_17406);
or UO_1241 (O_1241,N_18106,N_18708);
nor UO_1242 (O_1242,N_19067,N_19128);
or UO_1243 (O_1243,N_15059,N_19444);
nand UO_1244 (O_1244,N_16128,N_17666);
or UO_1245 (O_1245,N_17602,N_17688);
xnor UO_1246 (O_1246,N_18404,N_15062);
nand UO_1247 (O_1247,N_18076,N_17380);
nand UO_1248 (O_1248,N_17101,N_16403);
xnor UO_1249 (O_1249,N_19929,N_15666);
xor UO_1250 (O_1250,N_18201,N_15102);
and UO_1251 (O_1251,N_17986,N_16396);
or UO_1252 (O_1252,N_19162,N_19290);
and UO_1253 (O_1253,N_15148,N_19282);
and UO_1254 (O_1254,N_18741,N_16388);
nor UO_1255 (O_1255,N_19496,N_15551);
nor UO_1256 (O_1256,N_19770,N_16669);
nand UO_1257 (O_1257,N_15651,N_15039);
and UO_1258 (O_1258,N_17095,N_16947);
nor UO_1259 (O_1259,N_16659,N_18633);
xor UO_1260 (O_1260,N_16482,N_17267);
and UO_1261 (O_1261,N_18448,N_19224);
nand UO_1262 (O_1262,N_15690,N_17775);
nor UO_1263 (O_1263,N_17303,N_18867);
xor UO_1264 (O_1264,N_19126,N_19677);
or UO_1265 (O_1265,N_15764,N_15274);
nand UO_1266 (O_1266,N_16419,N_17921);
or UO_1267 (O_1267,N_17571,N_18191);
nand UO_1268 (O_1268,N_18659,N_17192);
or UO_1269 (O_1269,N_17261,N_17582);
nand UO_1270 (O_1270,N_16969,N_19574);
or UO_1271 (O_1271,N_17342,N_19719);
or UO_1272 (O_1272,N_19487,N_19732);
nand UO_1273 (O_1273,N_18979,N_18918);
or UO_1274 (O_1274,N_16677,N_15031);
nor UO_1275 (O_1275,N_17483,N_17040);
nor UO_1276 (O_1276,N_17823,N_16497);
or UO_1277 (O_1277,N_18036,N_15715);
or UO_1278 (O_1278,N_17371,N_17055);
nand UO_1279 (O_1279,N_15074,N_17813);
nand UO_1280 (O_1280,N_17207,N_15372);
nor UO_1281 (O_1281,N_17777,N_16547);
nor UO_1282 (O_1282,N_17764,N_16764);
or UO_1283 (O_1283,N_18021,N_17399);
nor UO_1284 (O_1284,N_15224,N_19400);
or UO_1285 (O_1285,N_16577,N_17373);
or UO_1286 (O_1286,N_19706,N_16240);
or UO_1287 (O_1287,N_17468,N_19666);
and UO_1288 (O_1288,N_19505,N_19818);
nor UO_1289 (O_1289,N_17810,N_18900);
and UO_1290 (O_1290,N_17880,N_17984);
and UO_1291 (O_1291,N_16864,N_16794);
or UO_1292 (O_1292,N_19380,N_19470);
xor UO_1293 (O_1293,N_15016,N_16760);
or UO_1294 (O_1294,N_18826,N_18122);
nand UO_1295 (O_1295,N_15915,N_16084);
or UO_1296 (O_1296,N_15216,N_15078);
and UO_1297 (O_1297,N_19474,N_17709);
xor UO_1298 (O_1298,N_19331,N_19820);
nor UO_1299 (O_1299,N_19376,N_16347);
nand UO_1300 (O_1300,N_16802,N_15276);
nand UO_1301 (O_1301,N_17943,N_16090);
nor UO_1302 (O_1302,N_15608,N_15435);
or UO_1303 (O_1303,N_17872,N_18783);
xor UO_1304 (O_1304,N_16380,N_16628);
nor UO_1305 (O_1305,N_16094,N_16264);
xnor UO_1306 (O_1306,N_17946,N_18911);
and UO_1307 (O_1307,N_19642,N_19650);
nor UO_1308 (O_1308,N_15994,N_17876);
and UO_1309 (O_1309,N_16823,N_19395);
and UO_1310 (O_1310,N_16127,N_16749);
xor UO_1311 (O_1311,N_16136,N_18315);
or UO_1312 (O_1312,N_15325,N_17008);
or UO_1313 (O_1313,N_17225,N_19174);
or UO_1314 (O_1314,N_15920,N_18797);
nor UO_1315 (O_1315,N_17652,N_15033);
or UO_1316 (O_1316,N_18737,N_18329);
or UO_1317 (O_1317,N_15052,N_18656);
xor UO_1318 (O_1318,N_19275,N_18219);
or UO_1319 (O_1319,N_15532,N_16661);
nor UO_1320 (O_1320,N_17162,N_17748);
or UO_1321 (O_1321,N_16033,N_17489);
nor UO_1322 (O_1322,N_15583,N_17822);
and UO_1323 (O_1323,N_15578,N_16532);
xnor UO_1324 (O_1324,N_16118,N_18305);
and UO_1325 (O_1325,N_17324,N_16550);
or UO_1326 (O_1326,N_15903,N_15661);
or UO_1327 (O_1327,N_15752,N_16176);
nand UO_1328 (O_1328,N_15120,N_16060);
xnor UO_1329 (O_1329,N_17317,N_17479);
and UO_1330 (O_1330,N_17924,N_15270);
nor UO_1331 (O_1331,N_19221,N_19780);
nand UO_1332 (O_1332,N_18934,N_15451);
nor UO_1333 (O_1333,N_17332,N_18111);
and UO_1334 (O_1334,N_18242,N_18211);
nor UO_1335 (O_1335,N_16228,N_16996);
nand UO_1336 (O_1336,N_19323,N_19679);
or UO_1337 (O_1337,N_19146,N_15323);
xor UO_1338 (O_1338,N_18266,N_15181);
or UO_1339 (O_1339,N_16687,N_15486);
and UO_1340 (O_1340,N_15605,N_16929);
and UO_1341 (O_1341,N_18130,N_16110);
and UO_1342 (O_1342,N_19348,N_17776);
and UO_1343 (O_1343,N_18588,N_15399);
and UO_1344 (O_1344,N_19696,N_19807);
xor UO_1345 (O_1345,N_16043,N_15223);
xnor UO_1346 (O_1346,N_16697,N_16506);
nor UO_1347 (O_1347,N_19972,N_16137);
nand UO_1348 (O_1348,N_19629,N_18771);
or UO_1349 (O_1349,N_18135,N_15664);
xnor UO_1350 (O_1350,N_19123,N_18914);
nor UO_1351 (O_1351,N_17077,N_15076);
xnor UO_1352 (O_1352,N_18550,N_16306);
nand UO_1353 (O_1353,N_19833,N_18279);
nand UO_1354 (O_1354,N_18598,N_19087);
nand UO_1355 (O_1355,N_15600,N_19266);
or UO_1356 (O_1356,N_16368,N_18002);
nand UO_1357 (O_1357,N_19428,N_19454);
and UO_1358 (O_1358,N_16844,N_18529);
and UO_1359 (O_1359,N_17167,N_17368);
xnor UO_1360 (O_1360,N_16367,N_18142);
nand UO_1361 (O_1361,N_15835,N_18017);
nor UO_1362 (O_1362,N_15776,N_17135);
or UO_1363 (O_1363,N_18505,N_15848);
xnor UO_1364 (O_1364,N_18735,N_16680);
or UO_1365 (O_1365,N_18144,N_19320);
nand UO_1366 (O_1366,N_16473,N_17627);
nor UO_1367 (O_1367,N_16394,N_16936);
nand UO_1368 (O_1368,N_18794,N_15125);
or UO_1369 (O_1369,N_17990,N_15440);
and UO_1370 (O_1370,N_18841,N_19165);
and UO_1371 (O_1371,N_15395,N_16561);
nor UO_1372 (O_1372,N_16670,N_15360);
xnor UO_1373 (O_1373,N_15081,N_15784);
nor UO_1374 (O_1374,N_19327,N_15389);
or UO_1375 (O_1375,N_17797,N_16364);
nor UO_1376 (O_1376,N_18606,N_17587);
nor UO_1377 (O_1377,N_15006,N_18234);
or UO_1378 (O_1378,N_18714,N_18039);
and UO_1379 (O_1379,N_16728,N_16813);
or UO_1380 (O_1380,N_15609,N_19932);
xor UO_1381 (O_1381,N_15958,N_18655);
or UO_1382 (O_1382,N_18457,N_16643);
nand UO_1383 (O_1383,N_16286,N_19547);
or UO_1384 (O_1384,N_17365,N_18488);
xnor UO_1385 (O_1385,N_16829,N_15134);
or UO_1386 (O_1386,N_19164,N_17565);
or UO_1387 (O_1387,N_15330,N_16085);
or UO_1388 (O_1388,N_19219,N_15582);
nor UO_1389 (O_1389,N_18947,N_16986);
nor UO_1390 (O_1390,N_15522,N_17508);
or UO_1391 (O_1391,N_17420,N_18383);
nand UO_1392 (O_1392,N_15376,N_17955);
xor UO_1393 (O_1393,N_16064,N_16314);
or UO_1394 (O_1394,N_19926,N_18452);
or UO_1395 (O_1395,N_16457,N_19782);
xnor UO_1396 (O_1396,N_15478,N_15589);
and UO_1397 (O_1397,N_16973,N_18405);
and UO_1398 (O_1398,N_19623,N_15043);
nand UO_1399 (O_1399,N_15584,N_15962);
and UO_1400 (O_1400,N_18664,N_16133);
nor UO_1401 (O_1401,N_18150,N_18327);
nand UO_1402 (O_1402,N_16231,N_18781);
or UO_1403 (O_1403,N_16230,N_15643);
or UO_1404 (O_1404,N_16325,N_16806);
and UO_1405 (O_1405,N_18905,N_19405);
and UO_1406 (O_1406,N_16341,N_15262);
xor UO_1407 (O_1407,N_19243,N_18060);
or UO_1408 (O_1408,N_17030,N_18294);
or UO_1409 (O_1409,N_19802,N_18801);
nand UO_1410 (O_1410,N_17705,N_18541);
and UO_1411 (O_1411,N_16880,N_19010);
and UO_1412 (O_1412,N_17304,N_18069);
or UO_1413 (O_1413,N_15632,N_16987);
and UO_1414 (O_1414,N_17343,N_18925);
xor UO_1415 (O_1415,N_18522,N_18026);
or UO_1416 (O_1416,N_19406,N_18097);
xnor UO_1417 (O_1417,N_16515,N_16494);
or UO_1418 (O_1418,N_17513,N_16891);
or UO_1419 (O_1419,N_18696,N_15751);
nor UO_1420 (O_1420,N_18689,N_17391);
or UO_1421 (O_1421,N_17881,N_15219);
nand UO_1422 (O_1422,N_16323,N_18439);
and UO_1423 (O_1423,N_17467,N_18085);
nand UO_1424 (O_1424,N_17635,N_19295);
and UO_1425 (O_1425,N_19073,N_18486);
nor UO_1426 (O_1426,N_17693,N_18264);
xor UO_1427 (O_1427,N_16289,N_17286);
nor UO_1428 (O_1428,N_17296,N_19301);
nand UO_1429 (O_1429,N_15477,N_15018);
nand UO_1430 (O_1430,N_18683,N_18393);
xor UO_1431 (O_1431,N_18586,N_17198);
nand UO_1432 (O_1432,N_18348,N_16613);
nand UO_1433 (O_1433,N_16592,N_15886);
or UO_1434 (O_1434,N_19472,N_15739);
and UO_1435 (O_1435,N_15441,N_19945);
nand UO_1436 (O_1436,N_18802,N_16186);
and UO_1437 (O_1437,N_18955,N_18235);
nor UO_1438 (O_1438,N_17460,N_15754);
nor UO_1439 (O_1439,N_17828,N_16157);
or UO_1440 (O_1440,N_17415,N_19819);
nor UO_1441 (O_1441,N_19399,N_17567);
and UO_1442 (O_1442,N_19079,N_19781);
or UO_1443 (O_1443,N_18745,N_15056);
or UO_1444 (O_1444,N_17131,N_18013);
nor UO_1445 (O_1445,N_15542,N_16809);
or UO_1446 (O_1446,N_16566,N_16098);
nor UO_1447 (O_1447,N_17359,N_16639);
and UO_1448 (O_1448,N_15548,N_19641);
and UO_1449 (O_1449,N_17447,N_15658);
and UO_1450 (O_1450,N_19408,N_16030);
nand UO_1451 (O_1451,N_15986,N_16994);
xor UO_1452 (O_1452,N_17157,N_17780);
nand UO_1453 (O_1453,N_18657,N_18882);
and UO_1454 (O_1454,N_15732,N_19527);
and UO_1455 (O_1455,N_17522,N_15881);
or UO_1456 (O_1456,N_18542,N_19480);
nor UO_1457 (O_1457,N_18113,N_16518);
nor UO_1458 (O_1458,N_19422,N_19143);
nand UO_1459 (O_1459,N_16789,N_19964);
nor UO_1460 (O_1460,N_19026,N_17572);
and UO_1461 (O_1461,N_15133,N_17898);
nor UO_1462 (O_1462,N_19803,N_18970);
nand UO_1463 (O_1463,N_19572,N_15169);
or UO_1464 (O_1464,N_17336,N_15708);
or UO_1465 (O_1465,N_19801,N_15396);
nand UO_1466 (O_1466,N_19086,N_18926);
or UO_1467 (O_1467,N_16554,N_17325);
and UO_1468 (O_1468,N_15531,N_16326);
and UO_1469 (O_1469,N_16655,N_19811);
nand UO_1470 (O_1470,N_16076,N_17557);
nand UO_1471 (O_1471,N_15748,N_16361);
or UO_1472 (O_1472,N_15428,N_17299);
and UO_1473 (O_1473,N_19340,N_19829);
nand UO_1474 (O_1474,N_17334,N_19517);
and UO_1475 (O_1475,N_17321,N_19878);
and UO_1476 (O_1476,N_15337,N_17239);
or UO_1477 (O_1477,N_19577,N_16382);
or UO_1478 (O_1478,N_16272,N_19684);
or UO_1479 (O_1479,N_17150,N_18207);
or UO_1480 (O_1480,N_17130,N_17014);
nand UO_1481 (O_1481,N_16985,N_17403);
and UO_1482 (O_1482,N_16919,N_15463);
or UO_1483 (O_1483,N_15456,N_15563);
nand UO_1484 (O_1484,N_15616,N_18001);
xor UO_1485 (O_1485,N_19914,N_19145);
and UO_1486 (O_1486,N_17907,N_19897);
nand UO_1487 (O_1487,N_18584,N_16948);
nand UO_1488 (O_1488,N_19760,N_17770);
xor UO_1489 (O_1489,N_19598,N_15071);
or UO_1490 (O_1490,N_18800,N_18132);
or UO_1491 (O_1491,N_18874,N_16701);
and UO_1492 (O_1492,N_18723,N_16288);
nor UO_1493 (O_1493,N_15625,N_17029);
nor UO_1494 (O_1494,N_15896,N_16042);
nor UO_1495 (O_1495,N_16161,N_18114);
or UO_1496 (O_1496,N_17059,N_17060);
xor UO_1497 (O_1497,N_15734,N_15385);
and UO_1498 (O_1498,N_15143,N_15721);
and UO_1499 (O_1499,N_16495,N_17912);
or UO_1500 (O_1500,N_16222,N_18118);
or UO_1501 (O_1501,N_17974,N_15175);
and UO_1502 (O_1502,N_18748,N_18376);
nor UO_1503 (O_1503,N_18328,N_18548);
xnor UO_1504 (O_1504,N_15562,N_18378);
and UO_1505 (O_1505,N_19015,N_16430);
and UO_1506 (O_1506,N_18963,N_17669);
nand UO_1507 (O_1507,N_19943,N_17616);
nand UO_1508 (O_1508,N_15758,N_16436);
and UO_1509 (O_1509,N_18489,N_16671);
or UO_1510 (O_1510,N_19665,N_18414);
xor UO_1511 (O_1511,N_17985,N_18204);
nor UO_1512 (O_1512,N_18049,N_19203);
or UO_1513 (O_1513,N_17629,N_19230);
nand UO_1514 (O_1514,N_19443,N_17556);
and UO_1515 (O_1515,N_17063,N_15082);
xnor UO_1516 (O_1516,N_18697,N_18596);
or UO_1517 (O_1517,N_18353,N_17922);
nand UO_1518 (O_1518,N_16004,N_15946);
and UO_1519 (O_1519,N_18066,N_15596);
nor UO_1520 (O_1520,N_18271,N_15331);
nand UO_1521 (O_1521,N_17035,N_15647);
or UO_1522 (O_1522,N_17805,N_18770);
and UO_1523 (O_1523,N_16205,N_18994);
nand UO_1524 (O_1524,N_18046,N_18842);
xnor UO_1525 (O_1525,N_16529,N_15319);
nand UO_1526 (O_1526,N_18521,N_16173);
or UO_1527 (O_1527,N_17251,N_18020);
nand UO_1528 (O_1528,N_18310,N_19302);
and UO_1529 (O_1529,N_18960,N_18583);
nor UO_1530 (O_1530,N_15556,N_18855);
xor UO_1531 (O_1531,N_17697,N_17713);
xnor UO_1532 (O_1532,N_17138,N_18174);
or UO_1533 (O_1533,N_16510,N_18392);
nand UO_1534 (O_1534,N_16893,N_16872);
or UO_1535 (O_1535,N_17339,N_18820);
xor UO_1536 (O_1536,N_17658,N_16706);
or UO_1537 (O_1537,N_17302,N_19440);
and UO_1538 (O_1538,N_16435,N_16625);
nor UO_1539 (O_1539,N_17287,N_18419);
nand UO_1540 (O_1540,N_16141,N_15761);
and UO_1541 (O_1541,N_16265,N_17674);
nand UO_1542 (O_1542,N_17689,N_19810);
nor UO_1543 (O_1543,N_15288,N_15538);
and UO_1544 (O_1544,N_15236,N_16877);
nor UO_1545 (O_1545,N_16782,N_19521);
or UO_1546 (O_1546,N_19450,N_18545);
nand UO_1547 (O_1547,N_15639,N_17868);
nor UO_1548 (O_1548,N_18587,N_17835);
xnor UO_1549 (O_1549,N_16966,N_19463);
nand UO_1550 (O_1550,N_15683,N_16277);
and UO_1551 (O_1551,N_18822,N_17795);
nand UO_1552 (O_1552,N_18884,N_18342);
nand UO_1553 (O_1553,N_19541,N_15247);
and UO_1554 (O_1554,N_19759,N_19859);
or UO_1555 (O_1555,N_19788,N_15753);
or UO_1556 (O_1556,N_17117,N_19070);
or UO_1557 (O_1557,N_19606,N_19908);
xor UO_1558 (O_1558,N_18730,N_16892);
nor UO_1559 (O_1559,N_19260,N_16998);
and UO_1560 (O_1560,N_16499,N_16330);
nand UO_1561 (O_1561,N_16924,N_18790);
nor UO_1562 (O_1562,N_15750,N_15543);
nand UO_1563 (O_1563,N_16108,N_19239);
or UO_1564 (O_1564,N_18179,N_15544);
nand UO_1565 (O_1565,N_19215,N_17241);
and UO_1566 (O_1566,N_18104,N_16113);
and UO_1567 (O_1567,N_19132,N_15474);
nor UO_1568 (O_1568,N_19784,N_19150);
and UO_1569 (O_1569,N_17315,N_19716);
and UO_1570 (O_1570,N_18751,N_18200);
or UO_1571 (O_1571,N_16374,N_18308);
or UO_1572 (O_1572,N_15879,N_16527);
and UO_1573 (O_1573,N_18799,N_15712);
nor UO_1574 (O_1574,N_17097,N_19711);
and UO_1575 (O_1575,N_18081,N_17307);
nor UO_1576 (O_1576,N_18285,N_15971);
xnor UO_1577 (O_1577,N_15397,N_18411);
nand UO_1578 (O_1578,N_18375,N_16139);
nand UO_1579 (O_1579,N_17018,N_15965);
and UO_1580 (O_1580,N_18192,N_18605);
nor UO_1581 (O_1581,N_18481,N_16972);
or UO_1582 (O_1582,N_18154,N_16649);
nor UO_1583 (O_1583,N_18068,N_16913);
nand UO_1584 (O_1584,N_19457,N_16299);
nor UO_1585 (O_1585,N_17105,N_17874);
or UO_1586 (O_1586,N_16258,N_15571);
nand UO_1587 (O_1587,N_16814,N_15933);
and UO_1588 (O_1588,N_19922,N_17438);
or UO_1589 (O_1589,N_18496,N_17344);
nor UO_1590 (O_1590,N_17968,N_17431);
or UO_1591 (O_1591,N_16426,N_15992);
and UO_1592 (O_1592,N_17112,N_17047);
nand UO_1593 (O_1593,N_16553,N_18384);
nor UO_1594 (O_1594,N_19695,N_19479);
nor UO_1595 (O_1595,N_16501,N_17744);
nor UO_1596 (O_1596,N_17730,N_16916);
or UO_1597 (O_1597,N_15934,N_17268);
nor UO_1598 (O_1598,N_17909,N_16692);
nor UO_1599 (O_1599,N_19382,N_16716);
nor UO_1600 (O_1600,N_18007,N_19136);
nand UO_1601 (O_1601,N_18990,N_18769);
nand UO_1602 (O_1602,N_15747,N_16197);
xor UO_1603 (O_1603,N_16901,N_19697);
nor UO_1604 (O_1604,N_18062,N_17390);
nor UO_1605 (O_1605,N_15187,N_18335);
xnor UO_1606 (O_1606,N_16089,N_19956);
nand UO_1607 (O_1607,N_15923,N_18151);
nand UO_1608 (O_1608,N_15831,N_16957);
and UO_1609 (O_1609,N_17740,N_17773);
and UO_1610 (O_1610,N_19045,N_19149);
nor UO_1611 (O_1611,N_17893,N_15040);
or UO_1612 (O_1612,N_19182,N_15980);
xor UO_1613 (O_1613,N_19038,N_17670);
or UO_1614 (O_1614,N_18511,N_15828);
or UO_1615 (O_1615,N_16906,N_18791);
or UO_1616 (O_1616,N_19620,N_18878);
and UO_1617 (O_1617,N_15114,N_18133);
and UO_1618 (O_1618,N_19940,N_17681);
xor UO_1619 (O_1619,N_15380,N_19081);
or UO_1620 (O_1620,N_16870,N_16171);
nor UO_1621 (O_1621,N_17114,N_16633);
and UO_1622 (O_1622,N_15928,N_15630);
or UO_1623 (O_1623,N_18644,N_19752);
nand UO_1624 (O_1624,N_18459,N_17470);
nand UO_1625 (O_1625,N_17598,N_19047);
and UO_1626 (O_1626,N_19410,N_18356);
and UO_1627 (O_1627,N_17139,N_19514);
or UO_1628 (O_1628,N_17554,N_17894);
nor UO_1629 (O_1629,N_18343,N_17288);
nor UO_1630 (O_1630,N_18222,N_16747);
nor UO_1631 (O_1631,N_15095,N_18630);
nand UO_1632 (O_1632,N_16849,N_15501);
nor UO_1633 (O_1633,N_18509,N_19000);
and UO_1634 (O_1634,N_15162,N_15089);
or UO_1635 (O_1635,N_18444,N_18249);
nor UO_1636 (O_1636,N_18171,N_18823);
nor UO_1637 (O_1637,N_17882,N_17617);
nand UO_1638 (O_1638,N_16682,N_19359);
nor UO_1639 (O_1639,N_19157,N_19808);
and UO_1640 (O_1640,N_18016,N_16335);
or UO_1641 (O_1641,N_15692,N_17960);
nor UO_1642 (O_1642,N_19206,N_18297);
nor UO_1643 (O_1643,N_15518,N_19414);
nand UO_1644 (O_1644,N_17837,N_17074);
nand UO_1645 (O_1645,N_17830,N_16717);
nand UO_1646 (O_1646,N_15073,N_18331);
xnor UO_1647 (O_1647,N_18946,N_16008);
nand UO_1648 (O_1648,N_19374,N_17330);
or UO_1649 (O_1649,N_17818,N_18666);
nor UO_1650 (O_1650,N_19082,N_19590);
nor UO_1651 (O_1651,N_17096,N_18812);
and UO_1652 (O_1652,N_19134,N_16703);
or UO_1653 (O_1653,N_17642,N_18194);
nor UO_1654 (O_1654,N_18785,N_18613);
nand UO_1655 (O_1655,N_16959,N_15449);
and UO_1656 (O_1656,N_16404,N_17204);
nand UO_1657 (O_1657,N_17936,N_19831);
or UO_1658 (O_1658,N_15183,N_16492);
nor UO_1659 (O_1659,N_15704,N_17069);
or UO_1660 (O_1660,N_15757,N_17434);
xor UO_1661 (O_1661,N_16831,N_17716);
and UO_1662 (O_1662,N_15394,N_15610);
xnor UO_1663 (O_1663,N_16262,N_15382);
nand UO_1664 (O_1664,N_15391,N_16626);
nand UO_1665 (O_1665,N_16509,N_19404);
or UO_1666 (O_1666,N_16664,N_19467);
and UO_1667 (O_1667,N_19229,N_18252);
xor UO_1668 (O_1668,N_17025,N_16440);
and UO_1669 (O_1669,N_17429,N_15673);
xor UO_1670 (O_1670,N_18558,N_16686);
and UO_1671 (O_1671,N_18215,N_19168);
or UO_1672 (O_1672,N_17592,N_17072);
and UO_1673 (O_1673,N_19585,N_16463);
xnor UO_1674 (O_1674,N_19683,N_17036);
nand UO_1675 (O_1675,N_19809,N_19676);
and UO_1676 (O_1676,N_16695,N_18678);
nand UO_1677 (O_1677,N_15147,N_15069);
nand UO_1678 (O_1678,N_19021,N_19979);
and UO_1679 (O_1679,N_18833,N_18836);
nor UO_1680 (O_1680,N_16427,N_17604);
xor UO_1681 (O_1681,N_18937,N_16838);
nand UO_1682 (O_1682,N_19271,N_18607);
nor UO_1683 (O_1683,N_18518,N_19037);
xnor UO_1684 (O_1684,N_15775,N_19603);
or UO_1685 (O_1685,N_19270,N_17163);
nand UO_1686 (O_1686,N_17392,N_19498);
nor UO_1687 (O_1687,N_19671,N_19113);
nor UO_1688 (O_1688,N_15675,N_16942);
and UO_1689 (O_1689,N_16620,N_17809);
nor UO_1690 (O_1690,N_17032,N_16795);
and UO_1691 (O_1691,N_18326,N_17563);
nor UO_1692 (O_1692,N_16016,N_19917);
xnor UO_1693 (O_1693,N_15914,N_15306);
and UO_1694 (O_1694,N_18886,N_18417);
nor UO_1695 (O_1695,N_18948,N_16048);
or UO_1696 (O_1696,N_18240,N_19074);
and UO_1697 (O_1697,N_18319,N_15779);
or UO_1698 (O_1698,N_15674,N_16317);
and UO_1699 (O_1699,N_15092,N_19582);
and UO_1700 (O_1700,N_16812,N_19924);
nand UO_1701 (O_1701,N_19634,N_18000);
or UO_1702 (O_1702,N_17575,N_15745);
or UO_1703 (O_1703,N_18793,N_15241);
nor UO_1704 (O_1704,N_19442,N_16783);
nand UO_1705 (O_1705,N_19439,N_19576);
nand UO_1706 (O_1706,N_17710,N_19210);
nor UO_1707 (O_1707,N_17430,N_16605);
nor UO_1708 (O_1708,N_19371,N_16200);
or UO_1709 (O_1709,N_18206,N_18180);
xor UO_1710 (O_1710,N_16006,N_15326);
or UO_1711 (O_1711,N_16290,N_16907);
or UO_1712 (O_1712,N_15725,N_16886);
nand UO_1713 (O_1713,N_19992,N_17401);
or UO_1714 (O_1714,N_15924,N_15314);
xnor UO_1715 (O_1715,N_18864,N_18538);
xnor UO_1716 (O_1716,N_16235,N_17013);
nor UO_1717 (O_1717,N_16748,N_19354);
nand UO_1718 (O_1718,N_17056,N_16342);
nand UO_1719 (O_1719,N_17366,N_17979);
nor UO_1720 (O_1720,N_18504,N_18805);
nor UO_1721 (O_1721,N_16745,N_16393);
xnor UO_1722 (O_1722,N_17785,N_15586);
nor UO_1723 (O_1723,N_16738,N_16662);
nor UO_1724 (O_1724,N_19883,N_17803);
and UO_1725 (O_1725,N_16797,N_17224);
and UO_1726 (O_1726,N_15638,N_19337);
nor UO_1727 (O_1727,N_17226,N_15577);
xor UO_1728 (O_1728,N_17873,N_18795);
and UO_1729 (O_1729,N_15709,N_18540);
xnor UO_1730 (O_1730,N_15649,N_16023);
and UO_1731 (O_1731,N_19649,N_16899);
xnor UO_1732 (O_1732,N_17136,N_16345);
and UO_1733 (O_1733,N_15646,N_19614);
xor UO_1734 (O_1734,N_17250,N_18621);
xor UO_1735 (O_1735,N_15023,N_16595);
nand UO_1736 (O_1736,N_17746,N_16406);
nor UO_1737 (O_1737,N_19795,N_16470);
and UO_1738 (O_1738,N_18661,N_15652);
xnor UO_1739 (O_1739,N_15912,N_15226);
nand UO_1740 (O_1740,N_19020,N_16297);
nand UO_1741 (O_1741,N_19240,N_18552);
nor UO_1742 (O_1742,N_15310,N_19071);
nor UO_1743 (O_1743,N_19509,N_17099);
and UO_1744 (O_1744,N_18725,N_17599);
and UO_1745 (O_1745,N_16920,N_19049);
and UO_1746 (O_1746,N_18364,N_17098);
and UO_1747 (O_1747,N_18784,N_17220);
nor UO_1748 (O_1748,N_17490,N_17700);
or UO_1749 (O_1749,N_15579,N_15929);
or UO_1750 (O_1750,N_15685,N_15964);
and UO_1751 (O_1751,N_15513,N_16552);
and UO_1752 (O_1752,N_17500,N_18339);
nor UO_1753 (O_1753,N_19104,N_15124);
and UO_1754 (O_1754,N_17578,N_19124);
xor UO_1755 (O_1755,N_19451,N_16313);
or UO_1756 (O_1756,N_18688,N_17952);
nor UO_1757 (O_1757,N_19192,N_18089);
nand UO_1758 (O_1758,N_19351,N_16790);
nor UO_1759 (O_1759,N_15941,N_19724);
xnor UO_1760 (O_1760,N_15367,N_19863);
nand UO_1761 (O_1761,N_19851,N_17071);
nor UO_1762 (O_1762,N_17413,N_15756);
nand UO_1763 (O_1763,N_17723,N_17743);
xor UO_1764 (O_1764,N_17439,N_18648);
nand UO_1765 (O_1765,N_19009,N_17297);
nor UO_1766 (O_1766,N_15985,N_17787);
or UO_1767 (O_1767,N_16319,N_17794);
nor UO_1768 (O_1768,N_16852,N_19728);
or UO_1769 (O_1769,N_16225,N_16037);
or UO_1770 (O_1770,N_15130,N_16333);
or UO_1771 (O_1771,N_15269,N_17058);
nand UO_1772 (O_1772,N_17644,N_18772);
or UO_1773 (O_1773,N_18396,N_15294);
nor UO_1774 (O_1774,N_19669,N_17065);
nor UO_1775 (O_1775,N_16389,N_16976);
and UO_1776 (O_1776,N_16737,N_18231);
nor UO_1777 (O_1777,N_18075,N_17660);
and UO_1778 (O_1778,N_19998,N_17807);
and UO_1779 (O_1779,N_18765,N_18037);
nand UO_1780 (O_1780,N_16207,N_16758);
or UO_1781 (O_1781,N_15873,N_19176);
and UO_1782 (O_1782,N_16500,N_19092);
nand UO_1783 (O_1783,N_15155,N_17385);
xor UO_1784 (O_1784,N_18952,N_15645);
nand UO_1785 (O_1785,N_16348,N_19735);
and UO_1786 (O_1786,N_16534,N_19001);
or UO_1787 (O_1787,N_16121,N_18704);
nor UO_1788 (O_1788,N_16933,N_16013);
nor UO_1789 (O_1789,N_17233,N_16439);
nor UO_1790 (O_1790,N_19961,N_18726);
nand UO_1791 (O_1791,N_15475,N_18758);
nand UO_1792 (O_1792,N_15575,N_16691);
or UO_1793 (O_1793,N_15371,N_19392);
xor UO_1794 (O_1794,N_19280,N_18458);
or UO_1795 (O_1795,N_18898,N_19687);
or UO_1796 (O_1796,N_15904,N_16096);
and UO_1797 (O_1797,N_18223,N_17945);
and UO_1798 (O_1798,N_19407,N_17701);
or UO_1799 (O_1799,N_16503,N_19955);
nand UO_1800 (O_1800,N_18311,N_18010);
or UO_1801 (O_1801,N_15359,N_19075);
and UO_1802 (O_1802,N_16578,N_17786);
or UO_1803 (O_1803,N_19057,N_15248);
or UO_1804 (O_1804,N_15699,N_18134);
and UO_1805 (O_1805,N_18699,N_19191);
nor UO_1806 (O_1806,N_18834,N_19643);
nand UO_1807 (O_1807,N_17418,N_15315);
nand UO_1808 (O_1808,N_19651,N_15332);
nand UO_1809 (O_1809,N_15887,N_19891);
nor UO_1810 (O_1810,N_16310,N_17123);
and UO_1811 (O_1811,N_16112,N_16800);
nand UO_1812 (O_1812,N_17050,N_17512);
nand UO_1813 (O_1813,N_18340,N_15988);
and UO_1814 (O_1814,N_15454,N_18048);
xnor UO_1815 (O_1815,N_16587,N_18562);
nor UO_1816 (O_1816,N_19580,N_19342);
nand UO_1817 (O_1817,N_15815,N_17527);
and UO_1818 (O_1818,N_18954,N_18528);
and UO_1819 (O_1819,N_15500,N_16005);
nand UO_1820 (O_1820,N_15281,N_18304);
and UO_1821 (O_1821,N_19925,N_18682);
nand UO_1822 (O_1822,N_17088,N_15424);
and UO_1823 (O_1823,N_16889,N_15925);
or UO_1824 (O_1824,N_17472,N_19672);
nand UO_1825 (O_1825,N_16221,N_17078);
nor UO_1826 (O_1826,N_16521,N_18577);
or UO_1827 (O_1827,N_17935,N_16087);
nor UO_1828 (O_1828,N_15918,N_18570);
nand UO_1829 (O_1829,N_18261,N_17848);
xor UO_1830 (O_1830,N_15450,N_18406);
nor UO_1831 (O_1831,N_16528,N_18487);
nor UO_1832 (O_1832,N_16068,N_19534);
and UO_1833 (O_1833,N_15166,N_18218);
nor UO_1834 (O_1834,N_17004,N_17361);
or UO_1835 (O_1835,N_19362,N_16808);
or UO_1836 (O_1836,N_17491,N_19947);
xor UO_1837 (O_1837,N_17281,N_17651);
xor UO_1838 (O_1838,N_16562,N_16572);
xor UO_1839 (O_1839,N_16038,N_15055);
nand UO_1840 (O_1840,N_15706,N_16678);
or UO_1841 (O_1841,N_15926,N_17679);
xor UO_1842 (O_1842,N_19876,N_18412);
nand UO_1843 (O_1843,N_15427,N_18033);
or UO_1844 (O_1844,N_18998,N_18045);
xnor UO_1845 (O_1845,N_17011,N_19544);
nand UO_1846 (O_1846,N_15511,N_18341);
and UO_1847 (O_1847,N_17362,N_16160);
or UO_1848 (O_1848,N_19199,N_17176);
nand UO_1849 (O_1849,N_19311,N_17969);
or UO_1850 (O_1850,N_18566,N_19033);
or UO_1851 (O_1851,N_16598,N_16989);
nand UO_1852 (O_1852,N_18468,N_19733);
or UO_1853 (O_1853,N_16505,N_16743);
xnor UO_1854 (O_1854,N_16939,N_15834);
nand UO_1855 (O_1855,N_17140,N_19681);
nand UO_1856 (O_1856,N_17560,N_19996);
or UO_1857 (O_1857,N_17170,N_19058);
and UO_1858 (O_1858,N_18904,N_15524);
nor UO_1859 (O_1859,N_19723,N_18617);
or UO_1860 (O_1860,N_16442,N_15883);
and UO_1861 (O_1861,N_17517,N_16890);
or UO_1862 (O_1862,N_16868,N_15138);
and UO_1863 (O_1863,N_18830,N_16858);
nor UO_1864 (O_1864,N_17708,N_16147);
or UO_1865 (O_1865,N_18463,N_19617);
and UO_1866 (O_1866,N_18709,N_19627);
or UO_1867 (O_1867,N_19034,N_15560);
and UO_1868 (O_1868,N_19276,N_15794);
or UO_1869 (O_1869,N_16432,N_19025);
nor UO_1870 (O_1870,N_18155,N_17122);
or UO_1871 (O_1871,N_17724,N_19227);
xnor UO_1872 (O_1872,N_16170,N_18762);
nor UO_1873 (O_1873,N_15368,N_16372);
and UO_1874 (O_1874,N_18153,N_15336);
nand UO_1875 (O_1875,N_18291,N_16184);
and UO_1876 (O_1876,N_15246,N_17817);
nand UO_1877 (O_1877,N_19195,N_19516);
xnor UO_1878 (O_1878,N_18059,N_16478);
nand UO_1879 (O_1879,N_18435,N_15321);
nand UO_1880 (O_1880,N_19822,N_16386);
or UO_1881 (O_1881,N_16000,N_17757);
and UO_1882 (O_1882,N_18325,N_16897);
or UO_1883 (O_1883,N_16843,N_15797);
and UO_1884 (O_1884,N_19555,N_17126);
and UO_1885 (O_1885,N_18456,N_15895);
xor UO_1886 (O_1886,N_16107,N_17820);
or UO_1887 (O_1887,N_16539,N_18196);
nor UO_1888 (O_1888,N_19332,N_16726);
xor UO_1889 (O_1889,N_15430,N_19110);
nand UO_1890 (O_1890,N_19312,N_15590);
nor UO_1891 (O_1891,N_15521,N_16195);
and UO_1892 (O_1892,N_19950,N_18988);
nand UO_1893 (O_1893,N_15618,N_17899);
nor UO_1894 (O_1894,N_19995,N_16975);
or UO_1895 (O_1895,N_17896,N_16236);
and UO_1896 (O_1896,N_18851,N_16246);
nor UO_1897 (O_1897,N_19352,N_19986);
or UO_1898 (O_1898,N_18169,N_16767);
nand UO_1899 (O_1899,N_18895,N_16895);
or UO_1900 (O_1900,N_19464,N_15022);
and UO_1901 (O_1901,N_15103,N_17574);
nand UO_1902 (O_1902,N_16287,N_17417);
nand UO_1903 (O_1903,N_17911,N_15297);
nor UO_1904 (O_1904,N_15623,N_17289);
nor UO_1905 (O_1905,N_16548,N_18480);
nand UO_1906 (O_1906,N_18695,N_19989);
and UO_1907 (O_1907,N_16964,N_16796);
or UO_1908 (O_1908,N_19418,N_16418);
nand UO_1909 (O_1909,N_16158,N_15554);
nor UO_1910 (O_1910,N_17834,N_17997);
nor UO_1911 (O_1911,N_16556,N_18477);
and UO_1912 (O_1912,N_18691,N_19921);
xnor UO_1913 (O_1913,N_16926,N_15200);
nor UO_1914 (O_1914,N_19906,N_16444);
nand UO_1915 (O_1915,N_16428,N_17673);
nand UO_1916 (O_1916,N_16821,N_19931);
nor UO_1917 (O_1917,N_17672,N_17349);
or UO_1918 (O_1918,N_19930,N_15619);
and UO_1919 (O_1919,N_19007,N_18616);
nand UO_1920 (O_1920,N_16260,N_17534);
xnor UO_1921 (O_1921,N_18902,N_18986);
and UO_1922 (O_1922,N_17645,N_15935);
nand UO_1923 (O_1923,N_19409,N_19031);
nand UO_1924 (O_1924,N_17732,N_18120);
or UO_1925 (O_1925,N_15229,N_19905);
nand UO_1926 (O_1926,N_16338,N_19189);
or UO_1927 (O_1927,N_19177,N_15553);
nor UO_1928 (O_1928,N_17355,N_16339);
xor UO_1929 (O_1929,N_19016,N_16707);
nor UO_1930 (O_1930,N_16941,N_15657);
xnor UO_1931 (O_1931,N_18516,N_18189);
or UO_1932 (O_1932,N_17847,N_18443);
xor UO_1933 (O_1933,N_17941,N_17081);
nand UO_1934 (O_1934,N_15378,N_19330);
or UO_1935 (O_1935,N_15937,N_17573);
nor UO_1936 (O_1936,N_15145,N_15890);
nor UO_1937 (O_1937,N_18899,N_15464);
and UO_1938 (O_1938,N_18707,N_16599);
nand UO_1939 (O_1939,N_19973,N_18673);
xor UO_1940 (O_1940,N_19682,N_16563);
or UO_1941 (O_1941,N_15196,N_16291);
and UO_1942 (O_1942,N_17919,N_18969);
or UO_1943 (O_1943,N_15906,N_15539);
and UO_1944 (O_1944,N_15534,N_15809);
nand UO_1945 (O_1945,N_16304,N_19597);
or UO_1946 (O_1946,N_18945,N_16538);
nand UO_1947 (O_1947,N_15900,N_16871);
nand UO_1948 (O_1948,N_15313,N_17149);
nor UO_1949 (O_1949,N_16020,N_18208);
nor UO_1950 (O_1950,N_15164,N_18454);
or UO_1951 (O_1951,N_15289,N_18871);
nor UO_1952 (O_1952,N_17972,N_15774);
nor UO_1953 (O_1953,N_18727,N_15975);
nand UO_1954 (O_1954,N_17901,N_15255);
and UO_1955 (O_1955,N_18175,N_15093);
and UO_1956 (O_1956,N_16132,N_19114);
nor UO_1957 (O_1957,N_16155,N_17664);
nor UO_1958 (O_1958,N_19154,N_15846);
or UO_1959 (O_1959,N_18465,N_19685);
nor UO_1960 (O_1960,N_15445,N_16773);
xnor UO_1961 (O_1961,N_19287,N_19586);
nand UO_1962 (O_1962,N_19435,N_17625);
and UO_1963 (O_1963,N_15165,N_16744);
and UO_1964 (O_1964,N_18672,N_17020);
and UO_1965 (O_1965,N_19130,N_17249);
nor UO_1966 (O_1966,N_17213,N_18859);
and UO_1967 (O_1967,N_16653,N_19094);
nand UO_1968 (O_1968,N_17591,N_15101);
and UO_1969 (O_1969,N_17789,N_19763);
xor UO_1970 (O_1970,N_16307,N_17570);
nor UO_1971 (O_1971,N_16834,N_17832);
or UO_1972 (O_1972,N_17444,N_19421);
nand UO_1973 (O_1973,N_17550,N_15978);
or UO_1974 (O_1974,N_18124,N_18912);
nand UO_1975 (O_1975,N_17416,N_16629);
or UO_1976 (O_1976,N_17981,N_17964);
and UO_1977 (O_1977,N_17520,N_18280);
or UO_1978 (O_1978,N_19987,N_19895);
nor UO_1979 (O_1979,N_15633,N_16057);
nor UO_1980 (O_1980,N_17676,N_15770);
nor UO_1981 (O_1981,N_17386,N_17752);
or UO_1982 (O_1982,N_15298,N_19858);
xor UO_1983 (O_1983,N_15956,N_15353);
nor UO_1984 (O_1984,N_18423,N_19238);
and UO_1985 (O_1985,N_17594,N_17867);
and UO_1986 (O_1986,N_16912,N_17549);
nor UO_1987 (O_1987,N_18352,N_16138);
nand UO_1988 (O_1988,N_16011,N_17624);
xor UO_1989 (O_1989,N_19748,N_19749);
nand UO_1990 (O_1990,N_16281,N_16369);
nor UO_1991 (O_1991,N_19349,N_17196);
nand UO_1992 (O_1992,N_19745,N_18461);
and UO_1993 (O_1993,N_16405,N_19999);
nand UO_1994 (O_1994,N_15857,N_16220);
or UO_1995 (O_1995,N_17585,N_16667);
or UO_1996 (O_1996,N_15098,N_16102);
and UO_1997 (O_1997,N_16832,N_16993);
and UO_1998 (O_1998,N_17511,N_17781);
nand UO_1999 (O_1999,N_18497,N_15599);
nor UO_2000 (O_2000,N_16623,N_18126);
or UO_2001 (O_2001,N_18638,N_16980);
nand UO_2002 (O_2002,N_16263,N_15087);
or UO_2003 (O_2003,N_18637,N_19198);
or UO_2004 (O_2004,N_17871,N_19560);
xor UO_2005 (O_2005,N_15407,N_17045);
or UO_2006 (O_2006,N_16818,N_15324);
nand UO_2007 (O_2007,N_19334,N_16636);
nor UO_2008 (O_2008,N_18620,N_15829);
xor UO_2009 (O_2009,N_16603,N_17727);
and UO_2010 (O_2010,N_19962,N_16544);
or UO_2011 (O_2011,N_17548,N_17473);
or UO_2012 (O_2012,N_17633,N_15152);
nand UO_2013 (O_2013,N_19750,N_17547);
or UO_2014 (O_2014,N_19777,N_17892);
nand UO_2015 (O_2015,N_17111,N_15710);
nand UO_2016 (O_2016,N_19530,N_18164);
nand UO_2017 (O_2017,N_19872,N_17827);
xnor UO_2018 (O_2018,N_17244,N_15469);
nand UO_2019 (O_2019,N_15271,N_17498);
or UO_2020 (O_2020,N_17526,N_18825);
nand UO_2021 (O_2021,N_18022,N_16381);
xnor UO_2022 (O_2022,N_17208,N_17774);
or UO_2023 (O_2023,N_18108,N_15444);
nor UO_2024 (O_2024,N_19396,N_15901);
nor UO_2025 (O_2025,N_15499,N_16449);
and UO_2026 (O_2026,N_16646,N_19993);
nand UO_2027 (O_2027,N_18184,N_17948);
and UO_2028 (O_2028,N_15237,N_17075);
nor UO_2029 (O_2029,N_15285,N_15230);
and UO_2030 (O_2030,N_16965,N_15507);
xor UO_2031 (O_2031,N_16837,N_17369);
and UO_2032 (O_2032,N_17507,N_16658);
nor UO_2033 (O_2033,N_19445,N_15552);
nand UO_2034 (O_2034,N_19249,N_15697);
and UO_2035 (O_2035,N_17850,N_19692);
nor UO_2036 (O_2036,N_15702,N_19214);
or UO_2037 (O_2037,N_18050,N_15406);
or UO_2038 (O_2038,N_17243,N_17175);
nor UO_2039 (O_2039,N_18303,N_15049);
nand UO_2040 (O_2040,N_16610,N_19217);
xnor UO_2041 (O_2041,N_19705,N_16523);
nand UO_2042 (O_2042,N_16302,N_15144);
nor UO_2043 (O_2043,N_19056,N_15264);
nor UO_2044 (O_2044,N_17897,N_17543);
nand UO_2045 (O_2045,N_16462,N_15795);
xnor UO_2046 (O_2046,N_19771,N_15253);
and UO_2047 (O_2047,N_19720,N_19612);
or UO_2048 (O_2048,N_19531,N_19055);
nand UO_2049 (O_2049,N_17861,N_17819);
nand UO_2050 (O_2050,N_15154,N_15520);
nor UO_2051 (O_2051,N_16429,N_18668);
nor UO_2052 (O_2052,N_18757,N_17246);
and UO_2053 (O_2053,N_19433,N_17980);
and UO_2054 (O_2054,N_17495,N_19484);
or UO_2055 (O_2055,N_18420,N_15104);
or UO_2056 (O_2056,N_19768,N_17858);
nor UO_2057 (O_2057,N_19753,N_15644);
or UO_2058 (O_2058,N_16963,N_15547);
or UO_2059 (O_2059,N_15338,N_15251);
nand UO_2060 (O_2060,N_18804,N_16066);
and UO_2061 (O_2061,N_15257,N_16109);
nand UO_2062 (O_2062,N_18275,N_18813);
and UO_2063 (O_2063,N_18494,N_18442);
or UO_2064 (O_2064,N_18597,N_16376);
or UO_2065 (O_2065,N_19423,N_17638);
or UO_2066 (O_2066,N_16250,N_15211);
and UO_2067 (O_2067,N_15804,N_18224);
or UO_2068 (O_2068,N_18374,N_16165);
or UO_2069 (O_2069,N_17161,N_16308);
or UO_2070 (O_2070,N_17347,N_17996);
nor UO_2071 (O_2071,N_17389,N_16953);
and UO_2072 (O_2072,N_19546,N_19654);
or UO_2073 (O_2073,N_19712,N_16036);
and UO_2074 (O_2074,N_19783,N_19431);
nor UO_2075 (O_2075,N_19969,N_17064);
and UO_2076 (O_2076,N_16175,N_15821);
nor UO_2077 (O_2077,N_17003,N_17407);
or UO_2078 (O_2078,N_16621,N_15707);
and UO_2079 (O_2079,N_15079,N_15170);
and UO_2080 (O_2080,N_15527,N_16217);
nand UO_2081 (O_2081,N_19250,N_19494);
and UO_2082 (O_2082,N_16644,N_17106);
xnor UO_2083 (O_2083,N_16316,N_16237);
nand UO_2084 (O_2084,N_15871,N_19281);
or UO_2085 (O_2085,N_16350,N_18065);
or UO_2086 (O_2086,N_16275,N_17023);
xor UO_2087 (O_2087,N_16582,N_16488);
or UO_2088 (O_2088,N_16254,N_15309);
or UO_2089 (O_2089,N_17552,N_15024);
or UO_2090 (O_2090,N_18568,N_19758);
nand UO_2091 (O_2091,N_17298,N_15161);
nor UO_2092 (O_2092,N_15156,N_16721);
or UO_2093 (O_2093,N_18591,N_16476);
and UO_2094 (O_2094,N_17034,N_18575);
nand UO_2095 (O_2095,N_16830,N_19609);
or UO_2096 (O_2096,N_19289,N_18246);
nor UO_2097 (O_2097,N_15549,N_17615);
nor UO_2098 (O_2098,N_16077,N_16768);
nor UO_2099 (O_2099,N_19234,N_19958);
or UO_2100 (O_2100,N_18870,N_19317);
xor UO_2101 (O_2101,N_19370,N_19873);
and UO_2102 (O_2102,N_19680,N_17044);
nor UO_2103 (O_2103,N_18549,N_18933);
nor UO_2104 (O_2104,N_19558,N_18622);
nand UO_2105 (O_2105,N_15882,N_19957);
or UO_2106 (O_2106,N_17141,N_18950);
nor UO_2107 (O_2107,N_15212,N_15595);
and UO_2108 (O_2108,N_15019,N_19880);
or UO_2109 (O_2109,N_18767,N_18690);
nor UO_2110 (O_2110,N_15999,N_15891);
nor UO_2111 (O_2111,N_18789,N_16781);
xnor UO_2112 (O_2112,N_16944,N_17433);
xor UO_2113 (O_2113,N_15627,N_15905);
nand UO_2114 (O_2114,N_18042,N_15592);
nand UO_2115 (O_2115,N_17469,N_18382);
nand UO_2116 (O_2116,N_19316,N_17812);
nor UO_2117 (O_2117,N_18161,N_19220);
nor UO_2118 (O_2118,N_15852,N_18910);
xor UO_2119 (O_2119,N_15242,N_15333);
and UO_2120 (O_2120,N_19095,N_16820);
nand UO_2121 (O_2121,N_16408,N_15767);
nand UO_2122 (O_2122,N_15249,N_17300);
or UO_2123 (O_2123,N_15442,N_18773);
nand UO_2124 (O_2124,N_15982,N_18031);
nand UO_2125 (O_2125,N_16723,N_19823);
or UO_2126 (O_2126,N_15738,N_16777);
xnor UO_2127 (O_2127,N_17007,N_15730);
and UO_2128 (O_2128,N_16354,N_19700);
nand UO_2129 (O_2129,N_15737,N_16724);
or UO_2130 (O_2130,N_19662,N_19184);
or UO_2131 (O_2131,N_16485,N_18248);
or UO_2132 (O_2132,N_19106,N_19881);
or UO_2133 (O_2133,N_18626,N_16490);
nand UO_2134 (O_2134,N_16915,N_17694);
nand UO_2135 (O_2135,N_15825,N_19850);
nand UO_2136 (O_2136,N_18019,N_19919);
xnor UO_2137 (O_2137,N_16722,N_17825);
nand UO_2138 (O_2138,N_18763,N_18816);
and UO_2139 (O_2139,N_16464,N_18711);
nand UO_2140 (O_2140,N_19022,N_15025);
xor UO_2141 (O_2141,N_19432,N_19357);
or UO_2142 (O_2142,N_15379,N_19098);
or UO_2143 (O_2143,N_16278,N_16168);
or UO_2144 (O_2144,N_16720,N_17086);
or UO_2145 (O_2145,N_16149,N_19610);
and UO_2146 (O_2146,N_15898,N_18567);
or UO_2147 (O_2147,N_15004,N_15267);
or UO_2148 (O_2148,N_19626,N_15345);
or UO_2149 (O_2149,N_19591,N_18641);
nand UO_2150 (O_2150,N_19050,N_16801);
or UO_2151 (O_2151,N_17073,N_17678);
nand UO_2152 (O_2152,N_15295,N_15798);
nor UO_2153 (O_2153,N_15146,N_18977);
and UO_2154 (O_2154,N_17505,N_15766);
nand UO_2155 (O_2155,N_16627,N_16294);
or UO_2156 (O_2156,N_15820,N_15681);
nor UO_2157 (O_2157,N_18426,N_17305);
nor UO_2158 (O_2158,N_18168,N_15280);
and UO_2159 (O_2159,N_16650,N_19632);
and UO_2160 (O_2160,N_16398,N_17908);
or UO_2161 (O_2161,N_15892,N_18386);
xor UO_2162 (O_2162,N_19389,N_16122);
nor UO_2163 (O_2163,N_19160,N_15141);
nor UO_2164 (O_2164,N_15364,N_15409);
nand UO_2165 (O_2165,N_19185,N_15408);
or UO_2166 (O_2166,N_19387,N_15529);
nor UO_2167 (O_2167,N_18645,N_18724);
and UO_2168 (O_2168,N_15765,N_17637);
xor UO_2169 (O_2169,N_19061,N_18377);
xnor UO_2170 (O_2170,N_19161,N_16751);
nand UO_2171 (O_2171,N_18485,N_19960);
nand UO_2172 (O_2172,N_19847,N_15818);
nand UO_2173 (O_2173,N_17422,N_16063);
nor UO_2174 (O_2174,N_15065,N_19678);
nor UO_2175 (O_2175,N_19090,N_19426);
and UO_2176 (O_2176,N_19151,N_19622);
nor UO_2177 (O_2177,N_17272,N_18852);
or UO_2178 (O_2178,N_15628,N_15654);
nand UO_2179 (O_2179,N_19904,N_17791);
nand UO_2180 (O_2180,N_15116,N_19563);
and UO_2181 (O_2181,N_16555,N_18845);
nand UO_2182 (O_2182,N_19043,N_16932);
or UO_2183 (O_2183,N_18453,N_16689);
and UO_2184 (O_2184,N_17459,N_18609);
nand UO_2185 (O_2185,N_19024,N_17132);
nand UO_2186 (O_2186,N_18366,N_18281);
nand UO_2187 (O_2187,N_17737,N_18389);
or UO_2188 (O_2188,N_18906,N_19755);
or UO_2189 (O_2189,N_15220,N_19814);
or UO_2190 (O_2190,N_15736,N_18847);
nor UO_2191 (O_2191,N_18466,N_15932);
nor UO_2192 (O_2192,N_19458,N_18868);
xnor UO_2193 (O_2193,N_15731,N_18140);
or UO_2194 (O_2194,N_15000,N_16019);
or UO_2195 (O_2195,N_17950,N_18416);
and UO_2196 (O_2196,N_17125,N_17998);
or UO_2197 (O_2197,N_19997,N_19241);
xnor UO_2198 (O_2198,N_16579,N_16193);
nor UO_2199 (O_2199,N_18274,N_17641);
nor UO_2200 (O_2200,N_15700,N_16375);
and UO_2201 (O_2201,N_18987,N_18298);
xor UO_2202 (O_2202,N_18543,N_18086);
and UO_2203 (O_2203,N_17341,N_19155);
and UO_2204 (O_2204,N_15861,N_17562);
nand UO_2205 (O_2205,N_18624,N_18943);
nor UO_2206 (O_2206,N_15667,N_15415);
nor UO_2207 (O_2207,N_15847,N_18073);
and UO_2208 (O_2208,N_17464,N_18265);
nand UO_2209 (O_2209,N_15386,N_17216);
or UO_2210 (O_2210,N_16612,N_19968);
nand UO_2211 (O_2211,N_19425,N_16732);
and UO_2212 (O_2212,N_18559,N_17763);
nand UO_2213 (O_2213,N_19836,N_19573);
nand UO_2214 (O_2214,N_17978,N_17015);
nor UO_2215 (O_2215,N_18921,N_19307);
or UO_2216 (O_2216,N_15729,N_16183);
or UO_2217 (O_2217,N_19364,N_16826);
nand UO_2218 (O_2218,N_19089,N_17205);
nor UO_2219 (O_2219,N_16608,N_15866);
nor UO_2220 (O_2220,N_16204,N_16694);
nand UO_2221 (O_2221,N_17849,N_16853);
and UO_2222 (O_2222,N_18380,N_16009);
nor UO_2223 (O_2223,N_17428,N_15705);
and UO_2224 (O_2224,N_19393,N_16151);
or UO_2225 (O_2225,N_15142,N_17333);
and UO_2226 (O_2226,N_15519,N_15894);
or UO_2227 (O_2227,N_16946,N_15373);
or UO_2228 (O_2228,N_16027,N_19144);
or UO_2229 (O_2229,N_16410,N_18701);
nor UO_2230 (O_2230,N_15010,N_17680);
or UO_2231 (O_2231,N_15178,N_15817);
nor UO_2232 (O_2232,N_18721,N_18052);
and UO_2233 (O_2233,N_16343,N_17067);
nor UO_2234 (O_2234,N_17831,N_16420);
nand UO_2235 (O_2235,N_19731,N_16486);
and UO_2236 (O_2236,N_17884,N_15077);
xor UO_2237 (O_2237,N_15703,N_19834);
and UO_2238 (O_2238,N_18907,N_17189);
and UO_2239 (O_2239,N_18365,N_17232);
or UO_2240 (O_2240,N_16635,N_16970);
and UO_2241 (O_2241,N_19821,N_19991);
nand UO_2242 (O_2242,N_17720,N_18202);
nor UO_2243 (O_2243,N_16955,N_16017);
and UO_2244 (O_2244,N_19288,N_18429);
xor UO_2245 (O_2245,N_15180,N_19274);
nand UO_2246 (O_2246,N_19659,N_19018);
nor UO_2247 (O_2247,N_18738,N_17022);
nor UO_2248 (O_2248,N_18634,N_16883);
or UO_2249 (O_2249,N_17412,N_15419);
nand UO_2250 (O_2250,N_17623,N_18436);
and UO_2251 (O_2251,N_18110,N_18390);
and UO_2252 (O_2252,N_18063,N_19746);
and UO_2253 (O_2253,N_17860,N_15291);
or UO_2254 (O_2254,N_16918,N_15807);
or UO_2255 (O_2255,N_17558,N_16958);
xor UO_2256 (O_2256,N_17862,N_16606);
nand UO_2257 (O_2257,N_16735,N_17739);
and UO_2258 (O_2258,N_19939,N_19751);
and UO_2259 (O_2259,N_15363,N_17194);
nor UO_2260 (O_2260,N_16632,N_18875);
nand UO_2261 (O_2261,N_17129,N_18951);
xnor UO_2262 (O_2262,N_17301,N_19959);
nand UO_2263 (O_2263,N_17318,N_17173);
nand UO_2264 (O_2264,N_17276,N_15503);
nor UO_2265 (O_2265,N_16990,N_19035);
nor UO_2266 (O_2266,N_15917,N_19483);
xor UO_2267 (O_2267,N_15110,N_17966);
xnor UO_2268 (O_2268,N_17217,N_17118);
xnor UO_2269 (O_2269,N_17914,N_18623);
and UO_2270 (O_2270,N_16040,N_16638);
xnor UO_2271 (O_2271,N_16824,N_16676);
nand UO_2272 (O_2272,N_16769,N_15564);
or UO_2273 (O_2273,N_15919,N_17271);
xor UO_2274 (O_2274,N_18554,N_18889);
nand UO_2275 (O_2275,N_15140,N_15713);
xnor UO_2276 (O_2276,N_15354,N_15727);
nand UO_2277 (O_2277,N_15411,N_16776);
nand UO_2278 (O_2278,N_15735,N_15268);
and UO_2279 (O_2279,N_16805,N_15749);
or UO_2280 (O_2280,N_18099,N_15027);
or UO_2281 (O_2281,N_15877,N_18199);
or UO_2282 (O_2282,N_15836,N_18694);
nor UO_2283 (O_2283,N_15728,N_19008);
nor UO_2284 (O_2284,N_18333,N_19508);
or UO_2285 (O_2285,N_15189,N_18006);
nand UO_2286 (O_2286,N_15696,N_15197);
nor UO_2287 (O_2287,N_16549,N_15954);
nor UO_2288 (O_2288,N_17692,N_16328);
and UO_2289 (O_2289,N_15909,N_19675);
nand UO_2290 (O_2290,N_19690,N_16229);
nor UO_2291 (O_2291,N_16466,N_15355);
nand UO_2292 (O_2292,N_15417,N_17541);
xnor UO_2293 (O_2293,N_16224,N_18422);
xor UO_2294 (O_2294,N_17493,N_17659);
xor UO_2295 (O_2295,N_19529,N_19828);
xnor UO_2296 (O_2296,N_19292,N_18698);
nor UO_2297 (O_2297,N_19309,N_16878);
nor UO_2298 (O_2298,N_16974,N_17814);
and UO_2299 (O_2299,N_17384,N_18571);
and UO_2300 (O_2300,N_15446,N_19729);
nand UO_2301 (O_2301,N_19848,N_18109);
nor UO_2302 (O_2302,N_19369,N_15585);
and UO_2303 (O_2303,N_17165,N_19004);
nand UO_2304 (O_2304,N_18515,N_19974);
and UO_2305 (O_2305,N_18796,N_15684);
or UO_2306 (O_2306,N_15402,N_15112);
nor UO_2307 (O_2307,N_18129,N_16617);
or UO_2308 (O_2308,N_15997,N_17833);
nor UO_2309 (O_2309,N_15017,N_17569);
or UO_2310 (O_2310,N_15559,N_16322);
or UO_2311 (O_2311,N_18125,N_16365);
and UO_2312 (O_2312,N_16245,N_17855);
nand UO_2313 (O_2313,N_17080,N_17759);
or UO_2314 (O_2314,N_19988,N_16609);
xor UO_2315 (O_2315,N_17502,N_17116);
or UO_2316 (O_2316,N_17240,N_16502);
nor UO_2317 (O_2317,N_19740,N_19616);
and UO_2318 (O_2318,N_17920,N_19552);
nor UO_2319 (O_2319,N_19039,N_15523);
nor UO_2320 (O_2320,N_19077,N_15981);
nor UO_2321 (O_2321,N_17754,N_19402);
and UO_2322 (O_2322,N_18372,N_15838);
or UO_2323 (O_2323,N_15930,N_18430);
nor UO_2324 (O_2324,N_19806,N_18283);
or UO_2325 (O_2325,N_15462,N_15286);
nor UO_2326 (O_2326,N_15790,N_19647);
and UO_2327 (O_2327,N_15174,N_17647);
nor UO_2328 (O_2328,N_16239,N_19981);
or UO_2329 (O_2329,N_19013,N_17824);
and UO_2330 (O_2330,N_18093,N_16756);
and UO_2331 (O_2331,N_15420,N_16301);
nor UO_2332 (O_2332,N_18604,N_16925);
and UO_2333 (O_2333,N_19042,N_17793);
or UO_2334 (O_2334,N_16384,N_17202);
nand UO_2335 (O_2335,N_18320,N_15346);
xnor UO_2336 (O_2336,N_19554,N_19041);
and UO_2337 (O_2337,N_19518,N_15509);
or UO_2338 (O_2338,N_16256,N_15193);
xor UO_2339 (O_2339,N_15983,N_18177);
nor UO_2340 (O_2340,N_16164,N_16637);
nand UO_2341 (O_2341,N_17755,N_15688);
xnor UO_2342 (O_2342,N_18096,N_17917);
or UO_2343 (O_2343,N_17017,N_19383);
and UO_2344 (O_2344,N_18316,N_19944);
or UO_2345 (O_2345,N_19864,N_18835);
nand UO_2346 (O_2346,N_17144,N_15283);
and UO_2347 (O_2347,N_15375,N_17581);
and UO_2348 (O_2348,N_17788,N_18803);
or UO_2349 (O_2349,N_18560,N_18152);
nor UO_2350 (O_2350,N_16018,N_15085);
and UO_2351 (O_2351,N_17455,N_15947);
xor UO_2352 (O_2352,N_15780,N_18732);
xor UO_2353 (O_2353,N_17504,N_15637);
nand UO_2354 (O_2354,N_18896,N_16839);
or UO_2355 (O_2355,N_17904,N_18163);
and UO_2356 (O_2356,N_16182,N_15279);
and UO_2357 (O_2357,N_15613,N_15504);
or UO_2358 (O_2358,N_15953,N_16267);
and UO_2359 (O_2359,N_18706,N_17191);
xnor UO_2360 (O_2360,N_19673,N_17002);
nor UO_2361 (O_2361,N_18684,N_16940);
or UO_2362 (O_2362,N_16645,N_15612);
nor UO_2363 (O_2363,N_18413,N_19054);
or UO_2364 (O_2364,N_15812,N_18646);
or UO_2365 (O_2365,N_15908,N_19767);
nand UO_2366 (O_2366,N_18425,N_18811);
or UO_2367 (O_2367,N_17404,N_15433);
and UO_2368 (O_2368,N_15208,N_16696);
xor UO_2369 (O_2369,N_16713,N_19764);
and UO_2370 (O_2370,N_19689,N_17875);
or UO_2371 (O_2371,N_15007,N_19769);
or UO_2372 (O_2372,N_18087,N_18499);
nand UO_2373 (O_2373,N_18760,N_17215);
nand UO_2374 (O_2374,N_19100,N_18107);
and UO_2375 (O_2375,N_19787,N_16352);
xor UO_2376 (O_2376,N_19105,N_18288);
and UO_2377 (O_2377,N_17351,N_18251);
or UO_2378 (O_2378,N_18434,N_18139);
or UO_2379 (O_2379,N_16573,N_17229);
nand UO_2380 (O_2380,N_16083,N_17079);
and UO_2381 (O_2381,N_18526,N_15191);
or UO_2382 (O_2382,N_18359,N_18747);
or UO_2383 (O_2383,N_16059,N_16058);
or UO_2384 (O_2384,N_19813,N_18433);
xnor UO_2385 (O_2385,N_17836,N_17962);
nor UO_2386 (O_2386,N_19799,N_15927);
nand UO_2387 (O_2387,N_15452,N_15312);
and UO_2388 (O_2388,N_15209,N_15425);
nand UO_2389 (O_2389,N_15488,N_17854);
and UO_2390 (O_2390,N_17188,N_17514);
or UO_2391 (O_2391,N_19080,N_18547);
and UO_2392 (O_2392,N_19163,N_16454);
or UO_2393 (O_2393,N_18344,N_16284);
and UO_2394 (O_2394,N_18778,N_16088);
nor UO_2395 (O_2395,N_16559,N_16140);
nor UO_2396 (O_2396,N_17284,N_17586);
or UO_2397 (O_2397,N_16422,N_18400);
and UO_2398 (O_2398,N_19148,N_19313);
or UO_2399 (O_2399,N_16512,N_18186);
nand UO_2400 (O_2400,N_18402,N_19520);
nor UO_2401 (O_2401,N_15172,N_18996);
nor UO_2402 (O_2402,N_15316,N_15250);
xor UO_2403 (O_2403,N_17374,N_18257);
nor UO_2404 (O_2404,N_15044,N_18744);
nor UO_2405 (O_2405,N_18409,N_16903);
or UO_2406 (O_2406,N_16520,N_17051);
and UO_2407 (O_2407,N_15636,N_16943);
xnor UO_2408 (O_2408,N_15535,N_19046);
xor UO_2409 (O_2409,N_18067,N_15936);
nand UO_2410 (O_2410,N_16081,N_19462);
or UO_2411 (O_2411,N_19619,N_16541);
or UO_2412 (O_2412,N_17294,N_18254);
nand UO_2413 (O_2413,N_19636,N_19231);
and UO_2414 (O_2414,N_18975,N_16115);
nand UO_2415 (O_2415,N_17396,N_17636);
and UO_2416 (O_2416,N_15261,N_19854);
and UO_2417 (O_2417,N_17682,N_15819);
nor UO_2418 (O_2418,N_19596,N_16730);
nand UO_2419 (O_2419,N_15665,N_18533);
and UO_2420 (O_2420,N_15458,N_18959);
or UO_2421 (O_2421,N_16684,N_16086);
nor UO_2422 (O_2422,N_19668,N_19615);
xnor UO_2423 (O_2423,N_17314,N_15540);
nand UO_2424 (O_2424,N_15365,N_19942);
nor UO_2425 (O_2425,N_17453,N_19186);
nand UO_2426 (O_2426,N_17844,N_19112);
and UO_2427 (O_2427,N_16594,N_15546);
nand UO_2428 (O_2428,N_19223,N_19789);
or UO_2429 (O_2429,N_16252,N_16251);
or UO_2430 (O_2430,N_18054,N_17425);
nand UO_2431 (O_2431,N_19849,N_17001);
or UO_2432 (O_2432,N_19743,N_18451);
nor UO_2433 (O_2433,N_16910,N_16761);
nor UO_2434 (O_2434,N_16055,N_19717);
nor UO_2435 (O_2435,N_15490,N_17104);
and UO_2436 (O_2436,N_16481,N_19358);
nand UO_2437 (O_2437,N_18361,N_15635);
nand UO_2438 (O_2438,N_19339,N_19592);
and UO_2439 (O_2439,N_16282,N_15472);
and UO_2440 (O_2440,N_17778,N_19815);
or UO_2441 (O_2441,N_19427,N_18391);
and UO_2442 (O_2442,N_16344,N_17488);
xnor UO_2443 (O_2443,N_17186,N_18472);
xor UO_2444 (O_2444,N_18260,N_16679);
nand UO_2445 (O_2445,N_17671,N_16248);
nand UO_2446 (O_2446,N_18493,N_19139);
and UO_2447 (O_2447,N_16570,N_18866);
and UO_2448 (O_2448,N_17684,N_16056);
or UO_2449 (O_2449,N_19489,N_15443);
nor UO_2450 (O_2450,N_18302,N_19952);
nor UO_2451 (O_2451,N_15974,N_19954);
xnor UO_2452 (O_2452,N_15858,N_16123);
or UO_2453 (O_2453,N_15199,N_16074);
nand UO_2454 (O_2454,N_17525,N_19869);
xnor UO_2455 (O_2455,N_17771,N_17524);
nor UO_2456 (O_2456,N_19017,N_17181);
nand UO_2457 (O_2457,N_16507,N_18957);
and UO_2458 (O_2458,N_16984,N_16324);
and UO_2459 (O_2459,N_18503,N_17446);
nand UO_2460 (O_2460,N_19504,N_18203);
nor UO_2461 (O_2461,N_15814,N_19490);
nor UO_2462 (O_2462,N_16531,N_16315);
and UO_2463 (O_2463,N_17124,N_17005);
nor UO_2464 (O_2464,N_18980,N_19670);
xnor UO_2465 (O_2465,N_19002,N_16395);
nand UO_2466 (O_2466,N_16062,N_19455);
nor UO_2467 (O_2467,N_15687,N_19373);
xnor UO_2468 (O_2468,N_19543,N_19578);
nand UO_2469 (O_2469,N_18590,N_19142);
nor UO_2470 (O_2470,N_15218,N_16596);
nor UO_2471 (O_2471,N_19601,N_15058);
nand UO_2472 (O_2472,N_18858,N_15875);
nand UO_2473 (O_2473,N_18642,N_18705);
and UO_2474 (O_2474,N_15491,N_17987);
xor UO_2475 (O_2475,N_19866,N_18345);
nand UO_2476 (O_2476,N_19096,N_17580);
xnor UO_2477 (O_2477,N_15012,N_15768);
nand UO_2478 (O_2478,N_16125,N_18940);
nand UO_2479 (O_2479,N_19865,N_17942);
nor UO_2480 (O_2480,N_19963,N_18536);
xnor UO_2481 (O_2481,N_16438,N_15374);
or UO_2482 (O_2482,N_17745,N_19916);
or UO_2483 (O_2483,N_19841,N_17376);
or UO_2484 (O_2484,N_16035,N_19014);
nand UO_2485 (O_2485,N_16178,N_17450);
nand UO_2486 (O_2486,N_16461,N_15888);
nand UO_2487 (O_2487,N_16551,N_17107);
and UO_2488 (O_2488,N_18640,N_19343);
nand UO_2489 (O_2489,N_17383,N_16285);
or UO_2490 (O_2490,N_17419,N_15245);
and UO_2491 (O_2491,N_17295,N_16894);
nand UO_2492 (O_2492,N_18631,N_16257);
and UO_2493 (O_2493,N_17214,N_18941);
and UO_2494 (O_2494,N_18755,N_15889);
or UO_2495 (O_2495,N_18363,N_18440);
xnor UO_2496 (O_2496,N_19693,N_15416);
or UO_2497 (O_2497,N_17714,N_16455);
xnor UO_2498 (O_2498,N_15762,N_19571);
or UO_2499 (O_2499,N_18614,N_17515);
endmodule