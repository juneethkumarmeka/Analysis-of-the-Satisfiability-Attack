module basic_1500_15000_2000_20_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_1240,In_532);
or U1 (N_1,In_738,In_197);
or U2 (N_2,In_817,In_880);
and U3 (N_3,In_1044,In_1392);
or U4 (N_4,In_494,In_29);
nor U5 (N_5,In_581,In_1223);
or U6 (N_6,In_316,In_1219);
xor U7 (N_7,In_806,In_641);
nor U8 (N_8,In_527,In_1257);
xor U9 (N_9,In_763,In_1262);
and U10 (N_10,In_1290,In_209);
xnor U11 (N_11,In_1425,In_673);
or U12 (N_12,In_666,In_377);
nand U13 (N_13,In_1135,In_477);
xnor U14 (N_14,In_597,In_905);
and U15 (N_15,In_337,In_621);
nor U16 (N_16,In_204,In_678);
or U17 (N_17,In_616,In_350);
nor U18 (N_18,In_155,In_1294);
nand U19 (N_19,In_1118,In_784);
and U20 (N_20,In_555,In_694);
xnor U21 (N_21,In_891,In_145);
or U22 (N_22,In_577,In_130);
and U23 (N_23,In_733,In_269);
nand U24 (N_24,In_542,In_1170);
or U25 (N_25,In_643,In_681);
or U26 (N_26,In_361,In_1353);
or U27 (N_27,In_1145,In_381);
or U28 (N_28,In_998,In_1228);
and U29 (N_29,In_1277,In_240);
xnor U30 (N_30,In_167,In_900);
xor U31 (N_31,In_19,In_1097);
nand U32 (N_32,In_811,In_1098);
nor U33 (N_33,In_973,In_1288);
xnor U34 (N_34,In_97,In_1008);
nand U35 (N_35,In_728,In_1115);
and U36 (N_36,In_725,In_987);
nor U37 (N_37,In_1347,In_523);
nor U38 (N_38,In_576,In_967);
nor U39 (N_39,In_70,In_10);
xor U40 (N_40,In_612,In_910);
xor U41 (N_41,In_338,In_774);
xor U42 (N_42,In_283,In_384);
or U43 (N_43,In_76,In_290);
or U44 (N_44,In_849,In_399);
and U45 (N_45,In_1226,In_75);
xor U46 (N_46,In_1176,In_1171);
nand U47 (N_47,In_1004,In_1409);
xor U48 (N_48,In_408,In_132);
xor U49 (N_49,In_321,In_1218);
nand U50 (N_50,In_1087,In_1427);
nor U51 (N_51,In_847,In_1352);
and U52 (N_52,In_1393,In_509);
nand U53 (N_53,In_92,In_633);
and U54 (N_54,In_263,In_1143);
nor U55 (N_55,In_918,In_100);
nor U56 (N_56,In_185,In_933);
xor U57 (N_57,In_1108,In_1447);
or U58 (N_58,In_789,In_552);
or U59 (N_59,In_1448,In_833);
and U60 (N_60,In_504,In_1330);
nor U61 (N_61,In_1010,In_574);
or U62 (N_62,In_49,In_1040);
nand U63 (N_63,In_721,In_432);
nor U64 (N_64,In_637,In_1178);
nand U65 (N_65,In_1112,In_88);
xor U66 (N_66,In_859,In_654);
nand U67 (N_67,In_618,In_915);
or U68 (N_68,In_1064,In_1291);
nand U69 (N_69,In_1187,In_688);
nor U70 (N_70,In_447,In_729);
nor U71 (N_71,In_151,In_841);
nand U72 (N_72,In_761,In_1305);
or U73 (N_73,In_1092,In_780);
and U74 (N_74,In_246,In_117);
nand U75 (N_75,In_352,In_1263);
xnor U76 (N_76,In_333,In_383);
nor U77 (N_77,In_1095,In_496);
or U78 (N_78,In_1342,In_1308);
nand U79 (N_79,In_1276,In_230);
xor U80 (N_80,In_411,In_1488);
and U81 (N_81,In_1315,In_547);
or U82 (N_82,In_309,In_187);
nor U83 (N_83,In_726,In_439);
or U84 (N_84,In_273,In_1314);
and U85 (N_85,In_1244,In_687);
nor U86 (N_86,In_964,In_975);
and U87 (N_87,In_1150,In_242);
nand U88 (N_88,In_1039,In_205);
nand U89 (N_89,In_6,In_247);
xnor U90 (N_90,In_1116,In_1117);
nor U91 (N_91,In_1439,In_77);
and U92 (N_92,In_356,In_739);
xor U93 (N_93,In_1364,In_1198);
nor U94 (N_94,In_512,In_1164);
and U95 (N_95,In_1378,In_808);
xnor U96 (N_96,In_434,In_219);
and U97 (N_97,In_645,In_1453);
nand U98 (N_98,In_1367,In_1355);
or U99 (N_99,In_1042,In_138);
nand U100 (N_100,In_773,In_691);
xnor U101 (N_101,In_546,In_1062);
nor U102 (N_102,In_732,In_85);
nor U103 (N_103,In_1402,In_116);
nor U104 (N_104,In_1272,In_1376);
xnor U105 (N_105,In_602,In_161);
and U106 (N_106,In_909,In_259);
and U107 (N_107,In_793,In_851);
xor U108 (N_108,In_96,In_751);
nand U109 (N_109,In_30,In_353);
nand U110 (N_110,In_1398,In_697);
nand U111 (N_111,In_1451,In_1438);
nand U112 (N_112,In_340,In_270);
and U113 (N_113,In_924,In_680);
xnor U114 (N_114,In_951,In_169);
nor U115 (N_115,In_565,In_332);
nand U116 (N_116,In_1254,In_329);
or U117 (N_117,In_1450,In_1387);
xor U118 (N_118,In_20,In_314);
or U119 (N_119,In_1014,In_1437);
or U120 (N_120,In_939,In_336);
and U121 (N_121,In_87,In_813);
nor U122 (N_122,In_221,In_1137);
xnor U123 (N_123,In_1020,In_456);
xor U124 (N_124,In_727,In_364);
or U125 (N_125,In_184,In_443);
and U126 (N_126,In_896,In_1496);
and U127 (N_127,In_1124,In_233);
or U128 (N_128,In_1283,In_143);
or U129 (N_129,In_1037,In_716);
nand U130 (N_130,In_125,In_380);
nor U131 (N_131,In_1078,In_82);
nand U132 (N_132,In_579,In_1468);
nand U133 (N_133,In_535,In_220);
or U134 (N_134,In_959,In_163);
or U135 (N_135,In_611,In_315);
and U136 (N_136,In_674,In_531);
or U137 (N_137,In_128,In_809);
or U138 (N_138,In_825,In_1027);
xor U139 (N_139,In_279,In_1180);
nor U140 (N_140,In_1173,In_1);
nand U141 (N_141,In_928,In_1227);
xnor U142 (N_142,In_892,In_72);
and U143 (N_143,In_79,In_559);
or U144 (N_144,In_1071,In_649);
nor U145 (N_145,In_414,In_965);
or U146 (N_146,In_797,In_278);
nand U147 (N_147,In_908,In_341);
or U148 (N_148,In_904,In_196);
and U149 (N_149,In_706,In_1024);
nor U150 (N_150,In_249,In_1298);
xor U151 (N_151,In_113,In_207);
and U152 (N_152,In_55,In_174);
nor U153 (N_153,In_1432,In_717);
nand U154 (N_154,In_1499,In_107);
and U155 (N_155,In_563,In_1375);
nor U156 (N_156,In_1192,In_1394);
nand U157 (N_157,In_917,In_391);
xnor U158 (N_158,In_460,In_1300);
nand U159 (N_159,In_1172,In_888);
and U160 (N_160,In_1079,In_1083);
nand U161 (N_161,In_1316,In_650);
xor U162 (N_162,In_1275,In_295);
nand U163 (N_163,In_451,In_265);
or U164 (N_164,In_418,In_506);
xor U165 (N_165,In_348,In_93);
nand U166 (N_166,In_179,In_1031);
and U167 (N_167,In_713,In_1446);
or U168 (N_168,In_1434,In_254);
nand U169 (N_169,In_1128,In_598);
and U170 (N_170,In_567,In_54);
nor U171 (N_171,In_371,In_1224);
and U172 (N_172,In_44,In_960);
xor U173 (N_173,In_1174,In_1109);
and U174 (N_174,In_108,In_359);
xor U175 (N_175,In_1038,In_448);
nand U176 (N_176,In_1400,In_1047);
and U177 (N_177,In_991,In_16);
nand U178 (N_178,In_213,In_1114);
nand U179 (N_179,In_66,In_684);
xor U180 (N_180,In_1041,In_166);
and U181 (N_181,In_1374,In_421);
xnor U182 (N_182,In_306,In_989);
nand U183 (N_183,In_764,In_1075);
and U184 (N_184,In_877,In_976);
nor U185 (N_185,In_1362,In_172);
nor U186 (N_186,In_566,In_1296);
and U187 (N_187,In_1259,In_354);
nor U188 (N_188,In_189,In_475);
xor U189 (N_189,In_935,In_214);
xor U190 (N_190,In_529,In_689);
and U191 (N_191,In_1233,In_50);
and U192 (N_192,In_1230,In_995);
and U193 (N_193,In_902,In_483);
and U194 (N_194,In_497,In_1269);
and U195 (N_195,In_394,In_554);
or U196 (N_196,In_1026,In_1054);
and U197 (N_197,In_368,In_236);
or U198 (N_198,In_1306,In_1472);
xnor U199 (N_199,In_1335,In_626);
xnor U200 (N_200,In_94,In_1013);
or U201 (N_201,In_26,In_1181);
or U202 (N_202,In_826,In_150);
and U203 (N_203,In_842,In_1481);
nand U204 (N_204,In_1410,In_832);
xnor U205 (N_205,In_517,In_946);
nand U206 (N_206,In_24,In_575);
and U207 (N_207,In_17,In_1297);
and U208 (N_208,In_570,In_328);
and U209 (N_209,In_792,In_744);
xnor U210 (N_210,In_1415,In_1274);
xor U211 (N_211,In_0,In_203);
or U212 (N_212,In_1161,In_1282);
nor U213 (N_213,In_258,In_790);
xnor U214 (N_214,In_63,In_1215);
and U215 (N_215,In_1480,In_1035);
and U216 (N_216,In_662,In_735);
nand U217 (N_217,In_747,In_667);
or U218 (N_218,In_1323,In_420);
nand U219 (N_219,In_105,In_927);
nor U220 (N_220,In_796,In_1067);
and U221 (N_221,In_635,In_302);
nor U222 (N_222,In_1455,In_1431);
xor U223 (N_223,In_1489,In_1310);
nor U224 (N_224,In_1221,In_589);
or U225 (N_225,In_64,In_1319);
and U226 (N_226,In_776,In_1264);
or U227 (N_227,In_1383,In_1159);
or U228 (N_228,In_1255,In_818);
nor U229 (N_229,In_1491,In_966);
nand U230 (N_230,In_1204,In_1022);
nand U231 (N_231,In_536,In_1140);
or U232 (N_232,In_365,In_968);
or U233 (N_233,In_86,In_415);
xor U234 (N_234,In_1278,In_62);
or U235 (N_235,In_801,In_264);
and U236 (N_236,In_1080,In_1162);
nor U237 (N_237,In_370,In_1424);
or U238 (N_238,In_834,In_1336);
nand U239 (N_239,In_953,In_1327);
nand U240 (N_240,In_608,In_934);
xor U241 (N_241,In_664,In_1470);
xnor U242 (N_242,In_768,In_461);
xnor U243 (N_243,In_1273,In_955);
xnor U244 (N_244,In_390,In_190);
or U245 (N_245,In_164,In_1068);
xor U246 (N_246,In_1185,In_115);
xor U247 (N_247,In_1048,In_1261);
xnor U248 (N_248,In_136,In_299);
and U249 (N_249,In_1399,In_837);
and U250 (N_250,In_525,In_863);
and U251 (N_251,In_986,In_941);
nand U252 (N_252,In_1236,In_395);
xnor U253 (N_253,In_25,In_1129);
and U254 (N_254,In_875,In_585);
nand U255 (N_255,In_515,In_7);
nand U256 (N_256,In_60,In_1443);
nand U257 (N_257,In_1205,In_510);
or U258 (N_258,In_514,In_1006);
nor U259 (N_259,In_972,In_393);
or U260 (N_260,In_1459,In_835);
xnor U261 (N_261,In_1485,In_1193);
xor U262 (N_262,In_709,In_1390);
xnor U263 (N_263,In_1477,In_405);
nor U264 (N_264,In_556,In_590);
or U265 (N_265,In_921,In_994);
nor U266 (N_266,In_596,In_317);
or U267 (N_267,In_1131,In_1211);
xor U268 (N_268,In_656,In_137);
xnor U269 (N_269,In_1321,In_1304);
and U270 (N_270,In_519,In_839);
xor U271 (N_271,In_152,In_1133);
nor U272 (N_272,In_550,In_992);
nor U273 (N_273,In_631,In_846);
xor U274 (N_274,In_472,In_84);
xor U275 (N_275,In_1414,In_471);
or U276 (N_276,In_226,In_1452);
or U277 (N_277,In_1000,In_58);
xnor U278 (N_278,In_199,In_42);
nand U279 (N_279,In_28,In_1464);
and U280 (N_280,In_245,In_490);
xor U281 (N_281,In_1260,In_442);
and U282 (N_282,In_996,In_1358);
nand U283 (N_283,In_677,In_281);
and U284 (N_284,In_925,In_1169);
or U285 (N_285,In_874,In_293);
or U286 (N_286,In_518,In_1146);
or U287 (N_287,In_224,In_215);
nor U288 (N_288,In_268,In_285);
nand U289 (N_289,In_47,In_1476);
and U290 (N_290,In_294,In_144);
and U291 (N_291,In_718,In_816);
and U292 (N_292,In_1337,In_1359);
or U293 (N_293,In_1365,In_173);
nor U294 (N_294,In_256,In_671);
and U295 (N_295,In_700,In_69);
nor U296 (N_296,In_1081,In_1416);
and U297 (N_297,In_1265,In_828);
nand U298 (N_298,In_736,In_398);
nor U299 (N_299,In_931,In_454);
nor U300 (N_300,In_441,In_305);
and U301 (N_301,In_889,In_600);
and U302 (N_302,In_1465,In_267);
and U303 (N_303,In_1235,In_118);
xnor U304 (N_304,In_1188,In_508);
and U305 (N_305,In_252,In_819);
and U306 (N_306,In_881,In_831);
nand U307 (N_307,In_952,In_1163);
or U308 (N_308,In_1053,In_404);
and U309 (N_309,In_1307,In_119);
and U310 (N_310,In_38,In_771);
or U311 (N_311,In_274,In_158);
and U312 (N_312,In_1134,In_344);
or U313 (N_313,In_111,In_482);
nand U314 (N_314,In_1203,In_110);
nor U315 (N_315,In_1096,In_244);
and U316 (N_316,In_607,In_466);
xor U317 (N_317,In_1104,In_544);
xnor U318 (N_318,In_153,In_286);
nor U319 (N_319,In_1326,In_628);
or U320 (N_320,In_90,In_410);
or U321 (N_321,In_1072,In_1046);
and U322 (N_322,In_804,In_375);
xnor U323 (N_323,In_630,In_1350);
xor U324 (N_324,In_533,In_812);
or U325 (N_325,In_593,In_1429);
or U326 (N_326,In_192,In_1066);
and U327 (N_327,In_502,In_1011);
and U328 (N_328,In_1475,In_201);
nor U329 (N_329,In_131,In_873);
nand U330 (N_330,In_346,In_791);
xnor U331 (N_331,In_438,In_1312);
xnor U332 (N_332,In_369,In_1132);
xor U333 (N_333,In_15,In_724);
nor U334 (N_334,In_343,In_433);
or U335 (N_335,In_919,In_1421);
nor U336 (N_336,In_1340,In_1206);
nor U337 (N_337,In_1442,In_853);
xnor U338 (N_338,In_289,In_363);
nand U339 (N_339,In_342,In_308);
nor U340 (N_340,In_1152,In_385);
or U341 (N_341,In_1060,In_313);
or U342 (N_342,In_379,In_1397);
nor U343 (N_343,In_657,In_14);
xor U344 (N_344,In_1052,In_1498);
nor U345 (N_345,In_133,In_1103);
or U346 (N_346,In_248,In_1287);
and U347 (N_347,In_1248,In_795);
and U348 (N_348,In_355,In_558);
xor U349 (N_349,In_291,In_1369);
and U350 (N_350,In_34,In_492);
nor U351 (N_351,In_489,In_1076);
or U352 (N_352,In_668,In_401);
or U353 (N_353,In_1320,In_445);
xor U354 (N_354,In_1231,In_5);
or U355 (N_355,In_759,In_13);
xor U356 (N_356,In_652,In_1368);
or U357 (N_357,In_1030,In_683);
xor U358 (N_358,In_663,In_288);
nor U359 (N_359,In_182,In_104);
nor U360 (N_360,In_945,In_1085);
xnor U361 (N_361,In_1395,In_943);
nor U362 (N_362,In_1253,In_1002);
nand U363 (N_363,In_893,In_1411);
nand U364 (N_364,In_580,In_194);
nor U365 (N_365,In_1474,In_1418);
or U366 (N_366,In_1045,In_753);
and U367 (N_367,In_323,In_926);
or U368 (N_368,In_869,In_993);
or U369 (N_369,In_500,In_389);
and U370 (N_370,In_982,In_798);
xor U371 (N_371,In_53,In_1413);
or U372 (N_372,In_11,In_412);
nand U373 (N_373,In_127,In_1458);
xnor U374 (N_374,In_659,In_1050);
xor U375 (N_375,In_498,In_990);
xnor U376 (N_376,In_123,In_857);
or U377 (N_377,In_1217,In_266);
or U378 (N_378,In_1069,In_862);
xnor U379 (N_379,In_175,In_178);
nand U380 (N_380,In_1461,In_815);
xor U381 (N_381,In_1302,In_534);
xor U382 (N_382,In_303,In_690);
nand U383 (N_383,In_962,In_80);
or U384 (N_384,In_397,In_914);
and U385 (N_385,In_83,In_446);
and U386 (N_386,In_682,In_146);
or U387 (N_387,In_465,In_1061);
nand U388 (N_388,In_954,In_894);
nand U389 (N_389,In_624,In_1322);
nand U390 (N_390,In_1216,In_387);
nor U391 (N_391,In_1249,In_1423);
nor U392 (N_392,In_604,In_619);
nand U393 (N_393,In_564,In_311);
or U394 (N_394,In_553,In_1331);
xor U395 (N_395,In_310,In_416);
xnor U396 (N_396,In_177,In_1207);
and U397 (N_397,In_805,In_750);
nor U398 (N_398,In_1293,In_1126);
or U399 (N_399,In_217,In_2);
nor U400 (N_400,In_35,In_231);
nand U401 (N_401,In_513,In_1239);
nand U402 (N_402,In_463,In_1184);
and U403 (N_403,In_899,In_913);
and U404 (N_404,In_594,In_436);
nor U405 (N_405,In_124,In_605);
nor U406 (N_406,In_686,In_571);
xor U407 (N_407,In_1292,In_757);
and U408 (N_408,In_239,In_947);
or U409 (N_409,In_1033,In_1333);
nand U410 (N_410,In_836,In_560);
and U411 (N_411,In_658,In_984);
and U412 (N_412,In_480,In_614);
or U413 (N_413,In_501,In_1089);
nor U414 (N_414,In_1311,In_425);
nor U415 (N_415,In_661,In_710);
or U416 (N_416,In_271,In_625);
xnor U417 (N_417,In_1229,In_1436);
nor U418 (N_418,In_481,In_1165);
and U419 (N_419,In_413,In_978);
nand U420 (N_420,In_1256,In_821);
nor U421 (N_421,In_1247,In_388);
nor U422 (N_422,In_582,In_511);
nand U423 (N_423,In_890,In_71);
and U424 (N_424,In_165,In_1242);
nand U425 (N_425,In_872,In_1271);
xor U426 (N_426,In_435,In_1377);
nor U427 (N_427,In_866,In_51);
nor U428 (N_428,In_699,In_296);
nor U429 (N_429,In_923,In_591);
nand U430 (N_430,In_40,In_21);
xnor U431 (N_431,In_1210,In_495);
nand U432 (N_432,In_1058,In_723);
or U433 (N_433,In_646,In_1074);
or U434 (N_434,In_1258,In_424);
nor U435 (N_435,In_1467,In_695);
or U436 (N_436,In_1268,In_339);
nor U437 (N_437,In_609,In_1049);
or U438 (N_438,In_1160,In_644);
and U439 (N_439,In_1325,In_1125);
nor U440 (N_440,In_606,In_772);
nand U441 (N_441,In_999,In_882);
nor U442 (N_442,In_1366,In_755);
and U443 (N_443,In_1107,In_134);
xnor U444 (N_444,In_1101,In_1445);
or U445 (N_445,In_1401,In_1281);
and U446 (N_446,In_176,In_255);
and U447 (N_447,In_1497,In_722);
and U448 (N_448,In_330,In_1435);
nor U449 (N_449,In_852,In_940);
and U450 (N_450,In_491,In_1286);
or U451 (N_451,In_911,In_431);
nor U452 (N_452,In_423,In_760);
or U453 (N_453,In_814,In_997);
nand U454 (N_454,In_1005,In_1252);
or U455 (N_455,In_357,In_861);
or U456 (N_456,In_1245,In_140);
or U457 (N_457,In_36,In_767);
nand U458 (N_458,In_1121,In_366);
nor U459 (N_459,In_1403,In_487);
xnor U460 (N_460,In_334,In_854);
xor U461 (N_461,In_467,In_180);
nand U462 (N_462,In_1384,In_298);
and U463 (N_463,In_301,In_592);
xor U464 (N_464,In_406,In_1404);
or U465 (N_465,In_1212,In_1009);
nand U466 (N_466,In_429,In_783);
and U467 (N_467,In_670,In_208);
and U468 (N_468,In_1151,In_551);
nor U469 (N_469,In_89,In_1482);
nand U470 (N_470,In_901,In_122);
or U471 (N_471,In_1479,In_1139);
nand U472 (N_472,In_374,In_613);
or U473 (N_473,In_610,In_195);
xor U474 (N_474,In_855,In_787);
xnor U475 (N_475,In_452,In_37);
nor U476 (N_476,In_586,In_503);
nor U477 (N_477,In_32,In_1130);
or U478 (N_478,In_1088,In_1332);
and U479 (N_479,In_932,In_1357);
nand U480 (N_480,In_1483,In_845);
nand U481 (N_481,In_1370,In_1199);
and U482 (N_482,In_1186,In_400);
and U483 (N_483,In_257,In_745);
nor U484 (N_484,In_632,In_1462);
nand U485 (N_485,In_78,In_135);
or U486 (N_486,In_52,In_101);
xnor U487 (N_487,In_693,In_428);
nor U488 (N_488,In_73,In_227);
or U489 (N_489,In_1241,In_162);
nor U490 (N_490,In_358,In_1086);
nand U491 (N_491,In_1486,In_944);
xnor U492 (N_492,In_1487,In_1454);
xnor U493 (N_493,In_1191,In_322);
nor U494 (N_494,In_521,In_648);
nor U495 (N_495,In_974,In_1407);
and U496 (N_496,In_198,In_449);
xnor U497 (N_497,In_427,In_1141);
or U498 (N_498,In_543,In_121);
and U499 (N_499,In_129,In_27);
nor U500 (N_500,In_1484,In_1351);
nand U501 (N_501,In_620,In_1120);
and U502 (N_502,In_468,In_1243);
xnor U503 (N_503,In_782,In_827);
xnor U504 (N_504,In_737,In_584);
nand U505 (N_505,In_170,In_1019);
or U506 (N_506,In_765,In_985);
nor U507 (N_507,In_23,In_640);
nand U508 (N_508,In_1457,In_484);
or U509 (N_509,In_106,In_803);
xnor U510 (N_510,In_743,In_1070);
and U511 (N_511,In_1090,In_1209);
or U512 (N_512,In_473,In_280);
nand U513 (N_513,In_486,In_1280);
nand U514 (N_514,In_1102,In_820);
and U515 (N_515,In_1166,In_95);
nand U516 (N_516,In_1084,In_898);
nand U517 (N_517,In_588,In_1222);
nor U518 (N_518,In_1168,In_884);
xnor U519 (N_519,In_458,In_1189);
and U520 (N_520,In_698,In_1412);
or U521 (N_521,In_858,In_1167);
xnor U522 (N_522,In_950,In_300);
nand U523 (N_523,In_599,In_868);
and U524 (N_524,In_98,In_1380);
xnor U525 (N_525,In_1344,In_887);
nor U526 (N_526,In_277,In_250);
nand U527 (N_527,In_488,In_524);
or U528 (N_528,In_45,In_212);
or U529 (N_529,In_856,In_638);
nand U530 (N_530,In_43,In_91);
or U531 (N_531,In_1341,In_1386);
nor U532 (N_532,In_879,In_41);
nor U533 (N_533,In_634,In_778);
xnor U534 (N_534,In_867,In_838);
nand U535 (N_535,In_655,In_669);
or U536 (N_536,In_292,In_1303);
or U537 (N_537,In_516,In_1153);
xor U538 (N_538,In_642,In_886);
xnor U539 (N_539,In_1111,In_1284);
or U540 (N_540,In_963,In_1059);
and U541 (N_541,In_865,In_362);
nand U542 (N_542,In_1001,In_1346);
nor U543 (N_543,In_1177,In_1148);
or U544 (N_544,In_748,In_287);
xnor U545 (N_545,In_741,In_720);
or U546 (N_546,In_777,In_1182);
nand U547 (N_547,In_1036,In_469);
nand U548 (N_548,In_272,In_1238);
and U549 (N_549,In_708,In_758);
or U550 (N_550,In_1220,In_440);
nand U551 (N_551,In_112,In_1029);
and U552 (N_552,In_1099,In_148);
or U553 (N_553,In_526,In_22);
nor U554 (N_554,In_949,In_528);
xnor U555 (N_555,In_561,In_282);
xnor U556 (N_556,In_1328,In_253);
nand U557 (N_557,In_1025,In_1419);
and U558 (N_558,In_304,In_977);
xor U559 (N_559,In_1441,In_331);
nor U560 (N_560,In_746,In_1373);
nor U561 (N_561,In_623,In_1417);
nor U562 (N_562,In_403,In_1356);
or U563 (N_563,In_360,In_829);
or U564 (N_564,In_324,In_1430);
nand U565 (N_565,In_734,In_1385);
nor U566 (N_566,In_961,In_1433);
and U567 (N_567,In_540,In_378);
and U568 (N_568,In_830,In_462);
nand U569 (N_569,In_731,In_275);
xnor U570 (N_570,In_1471,In_225);
nand U571 (N_571,In_126,In_1100);
or U572 (N_572,In_48,In_1043);
xnor U573 (N_573,In_1301,In_636);
nand U574 (N_574,In_1440,In_1237);
nor U575 (N_575,In_948,In_844);
or U576 (N_576,In_68,In_864);
nor U577 (N_577,In_679,In_979);
or U578 (N_578,In_522,In_318);
or U579 (N_579,In_312,In_1382);
and U580 (N_580,In_1214,In_33);
nand U581 (N_581,In_1196,In_1391);
and U582 (N_582,In_929,In_568);
nor U583 (N_583,In_74,In_186);
and U584 (N_584,In_794,In_883);
nand U585 (N_585,In_1156,In_450);
and U586 (N_586,In_8,In_920);
nand U587 (N_587,In_216,In_770);
or U588 (N_588,In_1361,In_702);
or U589 (N_589,In_860,In_479);
nand U590 (N_590,In_1408,In_56);
or U591 (N_591,In_807,In_261);
nor U592 (N_592,In_980,In_1015);
and U593 (N_593,In_31,In_505);
or U594 (N_594,In_1077,In_326);
xor U595 (N_595,In_703,In_1113);
nor U596 (N_596,In_823,In_234);
nand U597 (N_597,In_1144,In_499);
xnor U598 (N_598,In_1456,In_297);
and U599 (N_599,In_9,In_61);
xnor U600 (N_600,In_1091,In_1478);
and U601 (N_601,In_1279,In_969);
nor U602 (N_602,In_1213,In_749);
xnor U603 (N_603,In_1028,In_1021);
nor U604 (N_604,In_587,In_870);
and U605 (N_605,In_478,In_956);
or U606 (N_606,In_895,In_1317);
nand U607 (N_607,In_276,In_1406);
nand U608 (N_608,In_417,In_453);
or U609 (N_609,In_701,In_154);
or U610 (N_610,In_210,In_622);
or U611 (N_611,In_444,In_211);
nor U612 (N_612,In_1285,In_485);
nand U613 (N_613,In_1208,In_1057);
or U614 (N_614,In_983,In_583);
and U615 (N_615,In_1007,In_1179);
and U616 (N_616,In_262,In_1363);
and U617 (N_617,In_719,In_367);
xor U618 (N_618,In_1197,In_897);
or U619 (N_619,In_1372,In_325);
xor U620 (N_620,In_756,In_676);
xnor U621 (N_621,In_1138,In_549);
nand U622 (N_622,In_840,In_426);
nand U623 (N_623,In_1094,In_206);
nor U624 (N_624,In_1460,In_181);
xor U625 (N_625,In_422,In_685);
or U626 (N_626,In_675,In_1201);
nor U627 (N_627,In_1267,In_12);
xnor U628 (N_628,In_139,In_1119);
xnor U629 (N_629,In_730,In_541);
nor U630 (N_630,In_1324,In_711);
nand U631 (N_631,In_243,In_754);
nor U632 (N_632,In_57,In_1270);
or U633 (N_633,In_930,In_1313);
xor U634 (N_634,In_1110,In_1338);
xnor U635 (N_635,In_1034,In_419);
and U636 (N_636,In_573,In_988);
and U637 (N_637,In_712,In_59);
or U638 (N_638,In_1494,In_1339);
or U639 (N_639,In_156,In_742);
nor U640 (N_640,In_171,In_1055);
and U641 (N_641,In_871,In_141);
or U642 (N_642,In_848,In_627);
nor U643 (N_643,In_1492,In_707);
or U644 (N_644,In_810,In_319);
or U645 (N_645,In_103,In_1426);
nor U646 (N_646,In_1093,In_1202);
nand U647 (N_647,In_692,In_672);
nor U648 (N_648,In_335,In_1122);
nor U649 (N_649,In_1142,In_1354);
xnor U650 (N_650,In_228,In_1422);
or U651 (N_651,In_906,In_1136);
nor U652 (N_652,In_766,In_545);
and U653 (N_653,In_222,In_1017);
and U654 (N_654,In_572,In_665);
xor U655 (N_655,In_1194,In_878);
or U656 (N_656,In_537,In_1379);
nand U657 (N_657,In_1428,In_1490);
xnor U658 (N_658,In_1023,In_251);
nand U659 (N_659,In_168,In_907);
xor U660 (N_660,In_351,In_147);
nor U661 (N_661,In_238,In_971);
and U662 (N_662,In_769,In_1149);
nor U663 (N_663,In_651,In_824);
xor U664 (N_664,In_639,In_1016);
nor U665 (N_665,In_386,In_1032);
nor U666 (N_666,In_99,In_885);
xnor U667 (N_667,In_660,In_493);
xor U668 (N_668,In_970,In_781);
or U669 (N_669,In_1250,In_1329);
nor U670 (N_670,In_1469,In_218);
nor U671 (N_671,In_1157,In_705);
nand U672 (N_672,In_1018,In_538);
or U673 (N_673,In_1345,In_373);
nor U674 (N_674,In_530,In_507);
xnor U675 (N_675,In_1493,In_1334);
and U676 (N_676,In_539,In_942);
nand U677 (N_677,In_1463,In_938);
nor U678 (N_678,In_1246,In_1147);
or U679 (N_679,In_936,In_601);
and U680 (N_680,In_3,In_916);
nor U681 (N_681,In_843,In_775);
and U682 (N_682,In_320,In_740);
nor U683 (N_683,In_1495,In_160);
xnor U684 (N_684,In_392,In_595);
and U685 (N_685,In_696,In_376);
and U686 (N_686,In_67,In_1106);
or U687 (N_687,In_903,In_200);
nor U688 (N_688,In_81,In_191);
nand U689 (N_689,In_1289,In_188);
or U690 (N_690,In_109,In_957);
nand U691 (N_691,In_1371,In_548);
xor U692 (N_692,In_876,In_1444);
nor U693 (N_693,In_1299,In_142);
xnor U694 (N_694,In_46,In_396);
nor U695 (N_695,In_1309,In_232);
xor U696 (N_696,In_284,In_1073);
and U697 (N_697,In_4,In_159);
nor U698 (N_698,In_617,In_1389);
nand U699 (N_699,In_786,In_223);
and U700 (N_700,In_402,In_345);
nor U701 (N_701,In_464,In_785);
or U702 (N_702,In_407,In_1105);
or U703 (N_703,In_459,In_520);
xor U704 (N_704,In_850,In_788);
or U705 (N_705,In_752,In_1405);
xnor U706 (N_706,In_1082,In_1318);
or U707 (N_707,In_1396,In_1195);
xnor U708 (N_708,In_1183,In_799);
and U709 (N_709,In_120,In_1232);
xor U710 (N_710,In_1266,In_476);
and U711 (N_711,In_1295,In_1155);
or U712 (N_712,In_382,In_704);
xnor U713 (N_713,In_1003,In_779);
nand U714 (N_714,In_455,In_562);
xnor U715 (N_715,In_1420,In_1154);
nor U716 (N_716,In_569,In_241);
xnor U717 (N_717,In_457,In_114);
xnor U718 (N_718,In_65,In_557);
nor U719 (N_719,In_229,In_714);
xnor U720 (N_720,In_922,In_1473);
and U721 (N_721,In_149,In_1051);
nand U722 (N_722,In_1449,In_1063);
xnor U723 (N_723,In_822,In_1349);
or U724 (N_724,In_202,In_762);
and U725 (N_725,In_102,In_430);
or U726 (N_726,In_958,In_715);
xnor U727 (N_727,In_937,In_1360);
xnor U728 (N_728,In_1348,In_1012);
and U729 (N_729,In_18,In_1381);
nor U730 (N_730,In_183,In_1190);
nand U731 (N_731,In_193,In_615);
and U732 (N_732,In_409,In_1251);
and U733 (N_733,In_39,In_981);
nor U734 (N_734,In_237,In_1234);
nand U735 (N_735,In_1056,In_1225);
xnor U736 (N_736,In_578,In_307);
nor U737 (N_737,In_474,In_1158);
nand U738 (N_738,In_327,In_802);
and U739 (N_739,In_1388,In_912);
nor U740 (N_740,In_470,In_349);
and U741 (N_741,In_629,In_800);
xnor U742 (N_742,In_1466,In_1175);
nand U743 (N_743,In_1065,In_1123);
and U744 (N_744,In_157,In_1127);
or U745 (N_745,In_647,In_260);
nand U746 (N_746,In_1200,In_653);
xor U747 (N_747,In_603,In_1343);
nor U748 (N_748,In_437,In_347);
and U749 (N_749,In_372,In_235);
or U750 (N_750,N_647,N_420);
nor U751 (N_751,N_626,N_72);
nor U752 (N_752,N_443,N_23);
and U753 (N_753,N_291,N_357);
nand U754 (N_754,N_161,N_704);
nand U755 (N_755,N_606,N_731);
xor U756 (N_756,N_693,N_63);
and U757 (N_757,N_471,N_352);
xnor U758 (N_758,N_502,N_143);
xor U759 (N_759,N_610,N_430);
nand U760 (N_760,N_301,N_111);
nor U761 (N_761,N_87,N_677);
nor U762 (N_762,N_282,N_485);
and U763 (N_763,N_36,N_317);
xor U764 (N_764,N_455,N_312);
nor U765 (N_765,N_32,N_271);
and U766 (N_766,N_456,N_712);
or U767 (N_767,N_354,N_460);
nand U768 (N_768,N_434,N_5);
nand U769 (N_769,N_165,N_686);
and U770 (N_770,N_179,N_692);
nor U771 (N_771,N_322,N_432);
and U772 (N_772,N_164,N_40);
nand U773 (N_773,N_260,N_578);
nor U774 (N_774,N_453,N_721);
xnor U775 (N_775,N_487,N_214);
nand U776 (N_776,N_550,N_113);
or U777 (N_777,N_611,N_575);
nand U778 (N_778,N_457,N_679);
or U779 (N_779,N_139,N_172);
nand U780 (N_780,N_366,N_296);
xnor U781 (N_781,N_532,N_86);
nand U782 (N_782,N_309,N_645);
nand U783 (N_783,N_374,N_600);
nor U784 (N_784,N_559,N_137);
or U785 (N_785,N_701,N_427);
and U786 (N_786,N_153,N_173);
nor U787 (N_787,N_13,N_325);
or U788 (N_788,N_725,N_269);
and U789 (N_789,N_740,N_705);
or U790 (N_790,N_431,N_233);
nand U791 (N_791,N_551,N_724);
or U792 (N_792,N_386,N_560);
nor U793 (N_793,N_359,N_496);
nand U794 (N_794,N_574,N_425);
xor U795 (N_795,N_672,N_320);
and U796 (N_796,N_255,N_470);
xor U797 (N_797,N_394,N_397);
xor U798 (N_798,N_58,N_120);
xor U799 (N_799,N_492,N_642);
and U800 (N_800,N_47,N_666);
or U801 (N_801,N_11,N_150);
xnor U802 (N_802,N_186,N_228);
and U803 (N_803,N_45,N_416);
nand U804 (N_804,N_71,N_553);
and U805 (N_805,N_115,N_155);
nor U806 (N_806,N_580,N_700);
nand U807 (N_807,N_730,N_225);
and U808 (N_808,N_229,N_627);
xor U809 (N_809,N_702,N_512);
or U810 (N_810,N_177,N_259);
nor U811 (N_811,N_449,N_567);
and U812 (N_812,N_735,N_646);
nor U813 (N_813,N_404,N_500);
or U814 (N_814,N_276,N_9);
and U815 (N_815,N_60,N_44);
or U816 (N_816,N_495,N_507);
and U817 (N_817,N_643,N_510);
or U818 (N_818,N_289,N_729);
nand U819 (N_819,N_438,N_586);
nor U820 (N_820,N_236,N_401);
or U821 (N_821,N_387,N_257);
nor U822 (N_822,N_323,N_622);
nor U823 (N_823,N_605,N_246);
xnor U824 (N_824,N_98,N_618);
and U825 (N_825,N_612,N_499);
nand U826 (N_826,N_659,N_253);
xnor U827 (N_827,N_213,N_201);
nor U828 (N_828,N_292,N_70);
or U829 (N_829,N_743,N_717);
or U830 (N_830,N_441,N_601);
xor U831 (N_831,N_189,N_744);
and U832 (N_832,N_587,N_445);
nor U833 (N_833,N_12,N_719);
nand U834 (N_834,N_442,N_100);
nand U835 (N_835,N_625,N_73);
xnor U836 (N_836,N_34,N_486);
and U837 (N_837,N_33,N_131);
nor U838 (N_838,N_262,N_699);
nand U839 (N_839,N_467,N_341);
nand U840 (N_840,N_261,N_344);
nor U841 (N_841,N_695,N_35);
or U842 (N_842,N_22,N_564);
or U843 (N_843,N_676,N_148);
nand U844 (N_844,N_110,N_336);
nand U845 (N_845,N_707,N_18);
nand U846 (N_846,N_294,N_392);
or U847 (N_847,N_267,N_716);
xor U848 (N_848,N_504,N_415);
nor U849 (N_849,N_285,N_491);
and U850 (N_850,N_603,N_193);
and U851 (N_851,N_440,N_175);
xnor U852 (N_852,N_210,N_351);
nand U853 (N_853,N_247,N_493);
or U854 (N_854,N_151,N_613);
nand U855 (N_855,N_408,N_377);
xnor U856 (N_856,N_304,N_51);
and U857 (N_857,N_656,N_452);
xnor U858 (N_858,N_321,N_745);
nand U859 (N_859,N_544,N_589);
xor U860 (N_860,N_683,N_0);
or U861 (N_861,N_212,N_117);
nand U862 (N_862,N_8,N_90);
nor U863 (N_863,N_383,N_414);
and U864 (N_864,N_615,N_142);
xor U865 (N_865,N_451,N_483);
or U866 (N_866,N_579,N_249);
nand U867 (N_867,N_160,N_526);
and U868 (N_868,N_118,N_385);
or U869 (N_869,N_494,N_81);
nor U870 (N_870,N_328,N_522);
nor U871 (N_871,N_97,N_3);
nand U872 (N_872,N_61,N_474);
and U873 (N_873,N_475,N_447);
and U874 (N_874,N_583,N_211);
nor U875 (N_875,N_537,N_690);
xnor U876 (N_876,N_528,N_251);
or U877 (N_877,N_250,N_67);
xnor U878 (N_878,N_450,N_382);
nor U879 (N_879,N_57,N_114);
or U880 (N_880,N_62,N_435);
nor U881 (N_881,N_402,N_169);
nand U882 (N_882,N_480,N_266);
nand U883 (N_883,N_335,N_88);
xnor U884 (N_884,N_314,N_190);
nand U885 (N_885,N_548,N_347);
xnor U886 (N_886,N_617,N_591);
and U887 (N_887,N_566,N_94);
or U888 (N_888,N_543,N_29);
and U889 (N_889,N_674,N_217);
nor U890 (N_890,N_644,N_123);
or U891 (N_891,N_222,N_597);
and U892 (N_892,N_562,N_28);
nand U893 (N_893,N_358,N_747);
or U894 (N_894,N_698,N_513);
and U895 (N_895,N_585,N_109);
or U896 (N_896,N_65,N_307);
nor U897 (N_897,N_555,N_516);
xor U898 (N_898,N_330,N_412);
and U899 (N_899,N_19,N_205);
xor U900 (N_900,N_302,N_78);
and U901 (N_901,N_519,N_466);
or U902 (N_902,N_552,N_657);
or U903 (N_903,N_422,N_157);
and U904 (N_904,N_207,N_390);
xor U905 (N_905,N_518,N_231);
nor U906 (N_906,N_168,N_662);
xor U907 (N_907,N_84,N_361);
xnor U908 (N_908,N_632,N_459);
nand U909 (N_909,N_636,N_80);
or U910 (N_910,N_623,N_732);
or U911 (N_911,N_506,N_396);
nand U912 (N_912,N_595,N_203);
nand U913 (N_913,N_718,N_264);
and U914 (N_914,N_16,N_50);
and U915 (N_915,N_99,N_194);
and U916 (N_916,N_215,N_378);
xnor U917 (N_917,N_85,N_140);
xor U918 (N_918,N_75,N_572);
nand U919 (N_919,N_428,N_30);
and U920 (N_920,N_180,N_181);
nand U921 (N_921,N_68,N_235);
nor U922 (N_922,N_239,N_192);
nor U923 (N_923,N_391,N_184);
or U924 (N_924,N_542,N_631);
nand U925 (N_925,N_316,N_748);
and U926 (N_926,N_82,N_220);
or U927 (N_927,N_688,N_310);
and U928 (N_928,N_568,N_54);
nor U929 (N_929,N_122,N_241);
nor U930 (N_930,N_458,N_399);
xor U931 (N_931,N_403,N_514);
or U932 (N_932,N_334,N_227);
or U933 (N_933,N_216,N_281);
and U934 (N_934,N_736,N_691);
and U935 (N_935,N_126,N_706);
nand U936 (N_936,N_405,N_167);
or U937 (N_937,N_571,N_288);
or U938 (N_938,N_533,N_746);
nor U939 (N_939,N_709,N_363);
nand U940 (N_940,N_678,N_268);
and U941 (N_941,N_664,N_365);
nor U942 (N_942,N_91,N_293);
or U943 (N_943,N_556,N_202);
and U944 (N_944,N_209,N_178);
and U945 (N_945,N_195,N_197);
nand U946 (N_946,N_448,N_703);
nand U947 (N_947,N_406,N_569);
or U948 (N_948,N_10,N_593);
or U949 (N_949,N_342,N_333);
and U950 (N_950,N_461,N_92);
or U951 (N_951,N_614,N_654);
or U952 (N_952,N_708,N_380);
or U953 (N_953,N_232,N_738);
nor U954 (N_954,N_125,N_208);
and U955 (N_955,N_713,N_633);
xor U956 (N_956,N_287,N_132);
and U957 (N_957,N_530,N_665);
and U958 (N_958,N_185,N_355);
or U959 (N_959,N_4,N_711);
nand U960 (N_960,N_558,N_462);
nand U961 (N_961,N_668,N_478);
and U962 (N_962,N_102,N_93);
nor U963 (N_963,N_609,N_174);
xnor U964 (N_964,N_147,N_444);
nand U965 (N_965,N_364,N_162);
xnor U966 (N_966,N_101,N_411);
nor U967 (N_967,N_539,N_655);
xnor U968 (N_968,N_594,N_608);
nand U969 (N_969,N_669,N_136);
and U970 (N_970,N_219,N_588);
or U971 (N_971,N_557,N_521);
nor U972 (N_972,N_598,N_25);
nor U973 (N_973,N_53,N_728);
or U974 (N_974,N_697,N_529);
nor U975 (N_975,N_682,N_371);
or U976 (N_976,N_436,N_469);
xor U977 (N_977,N_410,N_224);
nor U978 (N_978,N_508,N_515);
and U979 (N_979,N_472,N_327);
or U980 (N_980,N_742,N_69);
nor U981 (N_981,N_297,N_226);
and U982 (N_982,N_400,N_339);
nand U983 (N_983,N_733,N_258);
xor U984 (N_984,N_89,N_254);
nand U985 (N_985,N_437,N_577);
nor U986 (N_986,N_104,N_21);
nand U987 (N_987,N_734,N_630);
or U988 (N_988,N_720,N_554);
or U989 (N_989,N_372,N_134);
and U990 (N_990,N_503,N_103);
nand U991 (N_991,N_26,N_221);
nor U992 (N_992,N_663,N_311);
nand U993 (N_993,N_124,N_581);
or U994 (N_994,N_350,N_576);
nand U995 (N_995,N_680,N_135);
nand U996 (N_996,N_64,N_183);
nor U997 (N_997,N_619,N_129);
and U998 (N_998,N_74,N_607);
xor U999 (N_999,N_163,N_17);
nor U1000 (N_1000,N_628,N_156);
and U1001 (N_1001,N_7,N_353);
or U1002 (N_1002,N_737,N_433);
or U1003 (N_1003,N_38,N_272);
nand U1004 (N_1004,N_421,N_170);
xnor U1005 (N_1005,N_468,N_545);
or U1006 (N_1006,N_592,N_710);
or U1007 (N_1007,N_127,N_395);
xor U1008 (N_1008,N_685,N_138);
or U1009 (N_1009,N_429,N_83);
and U1010 (N_1010,N_270,N_343);
xor U1011 (N_1011,N_349,N_240);
or U1012 (N_1012,N_237,N_324);
nand U1013 (N_1013,N_423,N_417);
and U1014 (N_1014,N_546,N_234);
or U1015 (N_1015,N_375,N_370);
and U1016 (N_1016,N_20,N_24);
xor U1017 (N_1017,N_749,N_439);
nor U1018 (N_1018,N_723,N_348);
and U1019 (N_1019,N_463,N_96);
nand U1020 (N_1020,N_200,N_306);
nor U1021 (N_1021,N_223,N_536);
xor U1022 (N_1022,N_384,N_121);
or U1023 (N_1023,N_256,N_55);
nor U1024 (N_1024,N_482,N_540);
and U1025 (N_1025,N_315,N_652);
nor U1026 (N_1026,N_182,N_641);
xnor U1027 (N_1027,N_473,N_604);
xnor U1028 (N_1028,N_105,N_230);
or U1029 (N_1029,N_204,N_727);
or U1030 (N_1030,N_191,N_649);
and U1031 (N_1031,N_141,N_484);
nor U1032 (N_1032,N_218,N_629);
nor U1033 (N_1033,N_95,N_245);
xnor U1034 (N_1034,N_393,N_76);
nand U1035 (N_1035,N_599,N_318);
xnor U1036 (N_1036,N_582,N_43);
or U1037 (N_1037,N_52,N_283);
or U1038 (N_1038,N_525,N_284);
nor U1039 (N_1039,N_345,N_419);
nand U1040 (N_1040,N_639,N_37);
nand U1041 (N_1041,N_476,N_653);
xnor U1042 (N_1042,N_108,N_166);
or U1043 (N_1043,N_242,N_517);
or U1044 (N_1044,N_244,N_549);
and U1045 (N_1045,N_689,N_501);
or U1046 (N_1046,N_278,N_671);
xor U1047 (N_1047,N_389,N_332);
or U1048 (N_1048,N_726,N_319);
nor U1049 (N_1049,N_326,N_409);
nor U1050 (N_1050,N_159,N_128);
nor U1051 (N_1051,N_238,N_722);
nand U1052 (N_1052,N_398,N_15);
xnor U1053 (N_1053,N_154,N_481);
and U1054 (N_1054,N_534,N_684);
nand U1055 (N_1055,N_369,N_424);
nand U1056 (N_1056,N_56,N_477);
and U1057 (N_1057,N_313,N_621);
nor U1058 (N_1058,N_305,N_446);
xnor U1059 (N_1059,N_658,N_547);
xnor U1060 (N_1060,N_407,N_651);
and U1061 (N_1061,N_171,N_464);
nor U1062 (N_1062,N_6,N_290);
xor U1063 (N_1063,N_252,N_498);
xor U1064 (N_1064,N_41,N_300);
nand U1065 (N_1065,N_14,N_48);
and U1066 (N_1066,N_362,N_381);
xor U1067 (N_1067,N_158,N_176);
nor U1068 (N_1068,N_146,N_338);
nor U1069 (N_1069,N_596,N_295);
and U1070 (N_1070,N_133,N_673);
or U1071 (N_1071,N_714,N_303);
or U1072 (N_1072,N_561,N_79);
and U1073 (N_1073,N_340,N_199);
nor U1074 (N_1074,N_505,N_1);
nand U1075 (N_1075,N_681,N_488);
nor U1076 (N_1076,N_538,N_275);
nand U1077 (N_1077,N_520,N_624);
and U1078 (N_1078,N_661,N_274);
xnor U1079 (N_1079,N_59,N_308);
xor U1080 (N_1080,N_489,N_379);
and U1081 (N_1081,N_635,N_198);
and U1082 (N_1082,N_187,N_145);
nor U1083 (N_1083,N_511,N_31);
xor U1084 (N_1084,N_616,N_565);
xnor U1085 (N_1085,N_106,N_265);
and U1086 (N_1086,N_367,N_49);
and U1087 (N_1087,N_675,N_280);
and U1088 (N_1088,N_413,N_524);
or U1089 (N_1089,N_715,N_42);
nor U1090 (N_1090,N_454,N_523);
or U1091 (N_1091,N_490,N_66);
and U1092 (N_1092,N_563,N_527);
nand U1093 (N_1093,N_741,N_648);
nor U1094 (N_1094,N_650,N_573);
nor U1095 (N_1095,N_243,N_509);
nor U1096 (N_1096,N_77,N_634);
and U1097 (N_1097,N_196,N_152);
nand U1098 (N_1098,N_27,N_667);
xnor U1099 (N_1099,N_356,N_368);
xor U1100 (N_1100,N_376,N_112);
or U1101 (N_1101,N_479,N_144);
and U1102 (N_1102,N_277,N_286);
or U1103 (N_1103,N_188,N_418);
nand U1104 (N_1104,N_329,N_46);
nand U1105 (N_1105,N_620,N_263);
nand U1106 (N_1106,N_426,N_116);
or U1107 (N_1107,N_590,N_248);
xor U1108 (N_1108,N_531,N_331);
nand U1109 (N_1109,N_638,N_694);
nor U1110 (N_1110,N_298,N_299);
xor U1111 (N_1111,N_346,N_39);
nor U1112 (N_1112,N_388,N_670);
and U1113 (N_1113,N_107,N_2);
nand U1114 (N_1114,N_739,N_584);
and U1115 (N_1115,N_149,N_535);
nor U1116 (N_1116,N_273,N_119);
or U1117 (N_1117,N_130,N_696);
and U1118 (N_1118,N_337,N_602);
or U1119 (N_1119,N_637,N_687);
xnor U1120 (N_1120,N_640,N_360);
nand U1121 (N_1121,N_541,N_570);
xor U1122 (N_1122,N_497,N_206);
nand U1123 (N_1123,N_660,N_465);
xnor U1124 (N_1124,N_373,N_279);
nand U1125 (N_1125,N_119,N_478);
nor U1126 (N_1126,N_749,N_685);
or U1127 (N_1127,N_408,N_636);
nand U1128 (N_1128,N_642,N_341);
or U1129 (N_1129,N_82,N_166);
or U1130 (N_1130,N_121,N_632);
or U1131 (N_1131,N_56,N_505);
xor U1132 (N_1132,N_671,N_183);
nor U1133 (N_1133,N_601,N_312);
and U1134 (N_1134,N_215,N_628);
or U1135 (N_1135,N_115,N_710);
or U1136 (N_1136,N_248,N_682);
xnor U1137 (N_1137,N_537,N_44);
and U1138 (N_1138,N_66,N_436);
or U1139 (N_1139,N_677,N_744);
nand U1140 (N_1140,N_215,N_487);
xnor U1141 (N_1141,N_458,N_267);
nand U1142 (N_1142,N_283,N_135);
xnor U1143 (N_1143,N_261,N_424);
xnor U1144 (N_1144,N_77,N_362);
and U1145 (N_1145,N_284,N_586);
and U1146 (N_1146,N_302,N_723);
nor U1147 (N_1147,N_250,N_416);
nand U1148 (N_1148,N_420,N_687);
and U1149 (N_1149,N_625,N_319);
xor U1150 (N_1150,N_503,N_39);
or U1151 (N_1151,N_435,N_85);
nand U1152 (N_1152,N_48,N_28);
and U1153 (N_1153,N_666,N_730);
xnor U1154 (N_1154,N_377,N_561);
nand U1155 (N_1155,N_568,N_319);
or U1156 (N_1156,N_38,N_538);
xor U1157 (N_1157,N_41,N_335);
nor U1158 (N_1158,N_58,N_704);
xnor U1159 (N_1159,N_305,N_511);
or U1160 (N_1160,N_451,N_608);
and U1161 (N_1161,N_94,N_541);
nand U1162 (N_1162,N_347,N_209);
or U1163 (N_1163,N_697,N_51);
and U1164 (N_1164,N_663,N_131);
xnor U1165 (N_1165,N_326,N_94);
xnor U1166 (N_1166,N_637,N_702);
nor U1167 (N_1167,N_736,N_418);
xor U1168 (N_1168,N_39,N_656);
or U1169 (N_1169,N_694,N_196);
or U1170 (N_1170,N_594,N_491);
nand U1171 (N_1171,N_418,N_227);
or U1172 (N_1172,N_690,N_518);
nor U1173 (N_1173,N_258,N_358);
nand U1174 (N_1174,N_123,N_500);
nor U1175 (N_1175,N_508,N_387);
and U1176 (N_1176,N_652,N_266);
nand U1177 (N_1177,N_420,N_677);
or U1178 (N_1178,N_586,N_616);
and U1179 (N_1179,N_624,N_505);
and U1180 (N_1180,N_300,N_715);
or U1181 (N_1181,N_412,N_88);
and U1182 (N_1182,N_472,N_20);
and U1183 (N_1183,N_174,N_477);
or U1184 (N_1184,N_572,N_59);
xnor U1185 (N_1185,N_270,N_125);
and U1186 (N_1186,N_173,N_322);
nand U1187 (N_1187,N_117,N_249);
nor U1188 (N_1188,N_678,N_392);
nor U1189 (N_1189,N_565,N_406);
nor U1190 (N_1190,N_432,N_204);
or U1191 (N_1191,N_432,N_460);
or U1192 (N_1192,N_600,N_496);
or U1193 (N_1193,N_466,N_568);
xnor U1194 (N_1194,N_677,N_570);
nand U1195 (N_1195,N_480,N_119);
nand U1196 (N_1196,N_423,N_340);
or U1197 (N_1197,N_360,N_307);
nor U1198 (N_1198,N_320,N_415);
xnor U1199 (N_1199,N_573,N_379);
xor U1200 (N_1200,N_87,N_443);
nor U1201 (N_1201,N_330,N_319);
nand U1202 (N_1202,N_663,N_586);
and U1203 (N_1203,N_740,N_412);
or U1204 (N_1204,N_525,N_141);
or U1205 (N_1205,N_292,N_161);
or U1206 (N_1206,N_203,N_570);
and U1207 (N_1207,N_178,N_289);
nor U1208 (N_1208,N_216,N_24);
nor U1209 (N_1209,N_311,N_211);
or U1210 (N_1210,N_376,N_561);
or U1211 (N_1211,N_140,N_694);
or U1212 (N_1212,N_100,N_10);
or U1213 (N_1213,N_683,N_464);
xnor U1214 (N_1214,N_179,N_217);
nor U1215 (N_1215,N_202,N_284);
nor U1216 (N_1216,N_216,N_441);
or U1217 (N_1217,N_230,N_90);
or U1218 (N_1218,N_724,N_432);
nand U1219 (N_1219,N_475,N_155);
xor U1220 (N_1220,N_583,N_625);
nand U1221 (N_1221,N_637,N_507);
and U1222 (N_1222,N_656,N_201);
nand U1223 (N_1223,N_0,N_409);
xor U1224 (N_1224,N_34,N_573);
nor U1225 (N_1225,N_470,N_644);
nand U1226 (N_1226,N_95,N_141);
or U1227 (N_1227,N_211,N_444);
xnor U1228 (N_1228,N_228,N_307);
nor U1229 (N_1229,N_94,N_495);
and U1230 (N_1230,N_596,N_503);
xnor U1231 (N_1231,N_364,N_340);
nor U1232 (N_1232,N_516,N_417);
nand U1233 (N_1233,N_212,N_78);
or U1234 (N_1234,N_34,N_173);
nand U1235 (N_1235,N_693,N_736);
nand U1236 (N_1236,N_483,N_121);
and U1237 (N_1237,N_134,N_47);
xnor U1238 (N_1238,N_704,N_559);
and U1239 (N_1239,N_17,N_738);
nor U1240 (N_1240,N_393,N_592);
nand U1241 (N_1241,N_691,N_706);
nor U1242 (N_1242,N_309,N_54);
xor U1243 (N_1243,N_486,N_455);
nor U1244 (N_1244,N_568,N_152);
nor U1245 (N_1245,N_747,N_258);
nor U1246 (N_1246,N_617,N_284);
nand U1247 (N_1247,N_51,N_738);
and U1248 (N_1248,N_106,N_316);
and U1249 (N_1249,N_16,N_342);
and U1250 (N_1250,N_419,N_431);
xnor U1251 (N_1251,N_442,N_513);
nor U1252 (N_1252,N_104,N_594);
xnor U1253 (N_1253,N_655,N_4);
nor U1254 (N_1254,N_466,N_675);
or U1255 (N_1255,N_137,N_140);
xnor U1256 (N_1256,N_414,N_125);
nand U1257 (N_1257,N_252,N_132);
or U1258 (N_1258,N_682,N_59);
or U1259 (N_1259,N_461,N_344);
or U1260 (N_1260,N_582,N_252);
and U1261 (N_1261,N_234,N_94);
xnor U1262 (N_1262,N_365,N_178);
nand U1263 (N_1263,N_432,N_709);
and U1264 (N_1264,N_11,N_466);
nor U1265 (N_1265,N_371,N_320);
or U1266 (N_1266,N_312,N_488);
nor U1267 (N_1267,N_79,N_504);
nor U1268 (N_1268,N_612,N_287);
xnor U1269 (N_1269,N_408,N_238);
or U1270 (N_1270,N_616,N_27);
xnor U1271 (N_1271,N_623,N_7);
nand U1272 (N_1272,N_412,N_696);
nor U1273 (N_1273,N_545,N_341);
xor U1274 (N_1274,N_152,N_11);
and U1275 (N_1275,N_425,N_457);
xor U1276 (N_1276,N_599,N_628);
xor U1277 (N_1277,N_667,N_57);
nor U1278 (N_1278,N_187,N_157);
nor U1279 (N_1279,N_455,N_108);
xor U1280 (N_1280,N_198,N_144);
nand U1281 (N_1281,N_677,N_323);
or U1282 (N_1282,N_590,N_656);
nand U1283 (N_1283,N_46,N_599);
nor U1284 (N_1284,N_725,N_40);
nor U1285 (N_1285,N_270,N_292);
nor U1286 (N_1286,N_568,N_455);
or U1287 (N_1287,N_506,N_319);
xnor U1288 (N_1288,N_632,N_495);
xnor U1289 (N_1289,N_533,N_701);
nor U1290 (N_1290,N_315,N_236);
nand U1291 (N_1291,N_114,N_412);
and U1292 (N_1292,N_506,N_394);
nand U1293 (N_1293,N_294,N_187);
or U1294 (N_1294,N_211,N_356);
and U1295 (N_1295,N_694,N_213);
and U1296 (N_1296,N_55,N_667);
and U1297 (N_1297,N_176,N_505);
xor U1298 (N_1298,N_154,N_31);
nor U1299 (N_1299,N_2,N_709);
nor U1300 (N_1300,N_697,N_473);
nor U1301 (N_1301,N_383,N_69);
xor U1302 (N_1302,N_372,N_421);
nand U1303 (N_1303,N_523,N_510);
or U1304 (N_1304,N_308,N_271);
or U1305 (N_1305,N_403,N_367);
and U1306 (N_1306,N_74,N_475);
and U1307 (N_1307,N_539,N_624);
and U1308 (N_1308,N_354,N_212);
xnor U1309 (N_1309,N_473,N_587);
and U1310 (N_1310,N_746,N_241);
nand U1311 (N_1311,N_317,N_349);
or U1312 (N_1312,N_442,N_53);
nand U1313 (N_1313,N_257,N_652);
nand U1314 (N_1314,N_396,N_478);
or U1315 (N_1315,N_466,N_590);
xnor U1316 (N_1316,N_588,N_638);
nand U1317 (N_1317,N_515,N_243);
or U1318 (N_1318,N_160,N_331);
xnor U1319 (N_1319,N_610,N_378);
nor U1320 (N_1320,N_345,N_446);
and U1321 (N_1321,N_485,N_301);
xor U1322 (N_1322,N_655,N_88);
and U1323 (N_1323,N_722,N_394);
or U1324 (N_1324,N_308,N_435);
xnor U1325 (N_1325,N_453,N_45);
nand U1326 (N_1326,N_536,N_361);
nand U1327 (N_1327,N_327,N_412);
xnor U1328 (N_1328,N_345,N_44);
nand U1329 (N_1329,N_278,N_376);
and U1330 (N_1330,N_656,N_355);
nand U1331 (N_1331,N_407,N_733);
or U1332 (N_1332,N_743,N_273);
nor U1333 (N_1333,N_161,N_135);
and U1334 (N_1334,N_252,N_435);
nor U1335 (N_1335,N_707,N_466);
xor U1336 (N_1336,N_536,N_6);
or U1337 (N_1337,N_168,N_581);
xnor U1338 (N_1338,N_701,N_712);
nor U1339 (N_1339,N_135,N_206);
and U1340 (N_1340,N_421,N_615);
nand U1341 (N_1341,N_255,N_416);
nor U1342 (N_1342,N_219,N_717);
nor U1343 (N_1343,N_432,N_311);
xnor U1344 (N_1344,N_202,N_250);
nor U1345 (N_1345,N_138,N_410);
xnor U1346 (N_1346,N_513,N_100);
and U1347 (N_1347,N_254,N_630);
nand U1348 (N_1348,N_462,N_151);
nand U1349 (N_1349,N_450,N_384);
nand U1350 (N_1350,N_495,N_235);
or U1351 (N_1351,N_290,N_581);
or U1352 (N_1352,N_489,N_87);
nor U1353 (N_1353,N_661,N_666);
nor U1354 (N_1354,N_420,N_603);
nand U1355 (N_1355,N_480,N_377);
nor U1356 (N_1356,N_490,N_296);
nand U1357 (N_1357,N_360,N_555);
or U1358 (N_1358,N_340,N_216);
nor U1359 (N_1359,N_445,N_569);
nand U1360 (N_1360,N_252,N_547);
nor U1361 (N_1361,N_502,N_417);
nor U1362 (N_1362,N_334,N_608);
and U1363 (N_1363,N_669,N_162);
and U1364 (N_1364,N_673,N_423);
or U1365 (N_1365,N_322,N_712);
xnor U1366 (N_1366,N_534,N_446);
and U1367 (N_1367,N_601,N_334);
or U1368 (N_1368,N_68,N_745);
and U1369 (N_1369,N_589,N_258);
xnor U1370 (N_1370,N_69,N_609);
nand U1371 (N_1371,N_303,N_82);
nand U1372 (N_1372,N_105,N_178);
nand U1373 (N_1373,N_35,N_221);
or U1374 (N_1374,N_15,N_6);
or U1375 (N_1375,N_314,N_84);
xor U1376 (N_1376,N_66,N_714);
nand U1377 (N_1377,N_557,N_113);
nor U1378 (N_1378,N_517,N_396);
nand U1379 (N_1379,N_524,N_358);
xnor U1380 (N_1380,N_570,N_473);
or U1381 (N_1381,N_122,N_303);
nand U1382 (N_1382,N_389,N_488);
and U1383 (N_1383,N_546,N_592);
or U1384 (N_1384,N_20,N_360);
xor U1385 (N_1385,N_675,N_43);
xnor U1386 (N_1386,N_329,N_416);
nand U1387 (N_1387,N_280,N_721);
or U1388 (N_1388,N_378,N_516);
or U1389 (N_1389,N_701,N_417);
xor U1390 (N_1390,N_518,N_572);
nand U1391 (N_1391,N_281,N_363);
and U1392 (N_1392,N_528,N_71);
xor U1393 (N_1393,N_40,N_559);
and U1394 (N_1394,N_381,N_198);
nor U1395 (N_1395,N_141,N_602);
or U1396 (N_1396,N_720,N_569);
xnor U1397 (N_1397,N_532,N_330);
nor U1398 (N_1398,N_445,N_245);
nand U1399 (N_1399,N_657,N_539);
nand U1400 (N_1400,N_730,N_669);
or U1401 (N_1401,N_327,N_28);
or U1402 (N_1402,N_275,N_78);
or U1403 (N_1403,N_543,N_136);
nand U1404 (N_1404,N_315,N_566);
and U1405 (N_1405,N_416,N_210);
or U1406 (N_1406,N_535,N_714);
or U1407 (N_1407,N_281,N_95);
xnor U1408 (N_1408,N_132,N_517);
or U1409 (N_1409,N_489,N_460);
and U1410 (N_1410,N_669,N_15);
xor U1411 (N_1411,N_187,N_673);
or U1412 (N_1412,N_383,N_128);
nand U1413 (N_1413,N_450,N_581);
nor U1414 (N_1414,N_562,N_329);
xor U1415 (N_1415,N_529,N_498);
nor U1416 (N_1416,N_658,N_363);
or U1417 (N_1417,N_570,N_173);
and U1418 (N_1418,N_448,N_267);
xnor U1419 (N_1419,N_219,N_708);
nand U1420 (N_1420,N_174,N_542);
xor U1421 (N_1421,N_455,N_693);
xnor U1422 (N_1422,N_407,N_195);
nand U1423 (N_1423,N_295,N_450);
xnor U1424 (N_1424,N_543,N_189);
nand U1425 (N_1425,N_488,N_155);
or U1426 (N_1426,N_256,N_278);
xor U1427 (N_1427,N_40,N_121);
xnor U1428 (N_1428,N_716,N_408);
or U1429 (N_1429,N_641,N_247);
xor U1430 (N_1430,N_435,N_610);
or U1431 (N_1431,N_79,N_338);
nand U1432 (N_1432,N_639,N_678);
or U1433 (N_1433,N_199,N_727);
nand U1434 (N_1434,N_456,N_23);
or U1435 (N_1435,N_35,N_426);
nand U1436 (N_1436,N_186,N_102);
nand U1437 (N_1437,N_664,N_351);
nor U1438 (N_1438,N_95,N_426);
nor U1439 (N_1439,N_349,N_552);
nor U1440 (N_1440,N_673,N_249);
or U1441 (N_1441,N_320,N_450);
nand U1442 (N_1442,N_629,N_467);
or U1443 (N_1443,N_619,N_433);
and U1444 (N_1444,N_744,N_224);
or U1445 (N_1445,N_470,N_194);
xnor U1446 (N_1446,N_591,N_351);
nor U1447 (N_1447,N_425,N_163);
xor U1448 (N_1448,N_365,N_687);
or U1449 (N_1449,N_399,N_124);
or U1450 (N_1450,N_675,N_236);
nand U1451 (N_1451,N_375,N_42);
nand U1452 (N_1452,N_489,N_60);
and U1453 (N_1453,N_240,N_681);
xor U1454 (N_1454,N_292,N_697);
or U1455 (N_1455,N_106,N_359);
nor U1456 (N_1456,N_511,N_693);
and U1457 (N_1457,N_149,N_0);
and U1458 (N_1458,N_10,N_72);
and U1459 (N_1459,N_251,N_694);
or U1460 (N_1460,N_361,N_393);
xnor U1461 (N_1461,N_223,N_207);
nor U1462 (N_1462,N_434,N_199);
nand U1463 (N_1463,N_199,N_119);
and U1464 (N_1464,N_614,N_485);
and U1465 (N_1465,N_437,N_216);
xnor U1466 (N_1466,N_138,N_429);
xor U1467 (N_1467,N_77,N_435);
nor U1468 (N_1468,N_744,N_325);
xnor U1469 (N_1469,N_344,N_123);
and U1470 (N_1470,N_635,N_663);
or U1471 (N_1471,N_720,N_659);
nand U1472 (N_1472,N_364,N_30);
and U1473 (N_1473,N_235,N_360);
xnor U1474 (N_1474,N_94,N_267);
and U1475 (N_1475,N_167,N_646);
or U1476 (N_1476,N_228,N_451);
nand U1477 (N_1477,N_472,N_143);
xnor U1478 (N_1478,N_52,N_329);
nand U1479 (N_1479,N_744,N_699);
or U1480 (N_1480,N_96,N_158);
and U1481 (N_1481,N_320,N_610);
or U1482 (N_1482,N_543,N_509);
nor U1483 (N_1483,N_284,N_700);
xor U1484 (N_1484,N_35,N_55);
and U1485 (N_1485,N_179,N_594);
and U1486 (N_1486,N_374,N_673);
nand U1487 (N_1487,N_103,N_557);
xnor U1488 (N_1488,N_475,N_643);
nand U1489 (N_1489,N_148,N_48);
and U1490 (N_1490,N_731,N_318);
and U1491 (N_1491,N_309,N_99);
or U1492 (N_1492,N_50,N_416);
nand U1493 (N_1493,N_129,N_136);
and U1494 (N_1494,N_266,N_572);
xnor U1495 (N_1495,N_89,N_511);
nor U1496 (N_1496,N_107,N_435);
or U1497 (N_1497,N_415,N_428);
or U1498 (N_1498,N_658,N_180);
xor U1499 (N_1499,N_591,N_369);
xor U1500 (N_1500,N_1256,N_1401);
nor U1501 (N_1501,N_920,N_818);
nor U1502 (N_1502,N_1064,N_1228);
and U1503 (N_1503,N_1035,N_1049);
or U1504 (N_1504,N_1272,N_1428);
nor U1505 (N_1505,N_1004,N_803);
or U1506 (N_1506,N_884,N_1381);
xor U1507 (N_1507,N_1138,N_1226);
and U1508 (N_1508,N_1386,N_915);
nand U1509 (N_1509,N_1392,N_1061);
nand U1510 (N_1510,N_1133,N_758);
or U1511 (N_1511,N_913,N_1063);
or U1512 (N_1512,N_1053,N_1185);
xnor U1513 (N_1513,N_1165,N_759);
or U1514 (N_1514,N_909,N_1253);
nor U1515 (N_1515,N_788,N_1070);
or U1516 (N_1516,N_1172,N_1105);
xnor U1517 (N_1517,N_1097,N_1075);
nor U1518 (N_1518,N_1385,N_1332);
and U1519 (N_1519,N_1407,N_1171);
xor U1520 (N_1520,N_1236,N_1176);
and U1521 (N_1521,N_1391,N_1052);
and U1522 (N_1522,N_1247,N_937);
and U1523 (N_1523,N_1473,N_1451);
and U1524 (N_1524,N_1340,N_959);
nand U1525 (N_1525,N_916,N_1325);
nor U1526 (N_1526,N_1085,N_1042);
and U1527 (N_1527,N_875,N_1060);
nor U1528 (N_1528,N_771,N_857);
or U1529 (N_1529,N_1214,N_756);
xnor U1530 (N_1530,N_1131,N_1187);
nor U1531 (N_1531,N_1020,N_876);
nor U1532 (N_1532,N_1339,N_1455);
nand U1533 (N_1533,N_750,N_873);
and U1534 (N_1534,N_940,N_1076);
or U1535 (N_1535,N_800,N_1229);
or U1536 (N_1536,N_903,N_1371);
and U1537 (N_1537,N_1373,N_1241);
nor U1538 (N_1538,N_802,N_789);
xor U1539 (N_1539,N_1243,N_1478);
nor U1540 (N_1540,N_1426,N_1352);
nand U1541 (N_1541,N_1300,N_1013);
xnor U1542 (N_1542,N_1047,N_919);
and U1543 (N_1543,N_848,N_1203);
and U1544 (N_1544,N_1080,N_1231);
and U1545 (N_1545,N_1009,N_964);
xnor U1546 (N_1546,N_1434,N_1152);
nand U1547 (N_1547,N_1424,N_1178);
nand U1548 (N_1548,N_825,N_877);
xnor U1549 (N_1549,N_1462,N_1184);
nor U1550 (N_1550,N_1397,N_1018);
nand U1551 (N_1551,N_1314,N_1412);
or U1552 (N_1552,N_1452,N_979);
xnor U1553 (N_1553,N_1069,N_1395);
xor U1554 (N_1554,N_1007,N_1414);
or U1555 (N_1555,N_1273,N_1123);
nor U1556 (N_1556,N_1374,N_863);
or U1557 (N_1557,N_1248,N_1202);
xnor U1558 (N_1558,N_1393,N_1269);
and U1559 (N_1559,N_1274,N_838);
or U1560 (N_1560,N_1121,N_924);
xnor U1561 (N_1561,N_1162,N_1227);
nor U1562 (N_1562,N_1302,N_1305);
and U1563 (N_1563,N_1427,N_858);
nand U1564 (N_1564,N_1217,N_994);
or U1565 (N_1565,N_815,N_932);
nand U1566 (N_1566,N_1458,N_1006);
or U1567 (N_1567,N_1118,N_1206);
nand U1568 (N_1568,N_1086,N_898);
nor U1569 (N_1569,N_1139,N_1117);
nand U1570 (N_1570,N_1014,N_1278);
or U1571 (N_1571,N_816,N_1435);
or U1572 (N_1572,N_939,N_1467);
or U1573 (N_1573,N_1448,N_1192);
xnor U1574 (N_1574,N_904,N_753);
xnor U1575 (N_1575,N_1491,N_912);
nor U1576 (N_1576,N_1372,N_882);
nor U1577 (N_1577,N_930,N_1023);
nor U1578 (N_1578,N_767,N_963);
nor U1579 (N_1579,N_972,N_837);
or U1580 (N_1580,N_1328,N_755);
or U1581 (N_1581,N_1005,N_1250);
and U1582 (N_1582,N_1144,N_1183);
nor U1583 (N_1583,N_1111,N_1084);
and U1584 (N_1584,N_1000,N_1148);
or U1585 (N_1585,N_1220,N_861);
xor U1586 (N_1586,N_1350,N_859);
nand U1587 (N_1587,N_1147,N_1358);
nor U1588 (N_1588,N_809,N_929);
or U1589 (N_1589,N_1038,N_1254);
or U1590 (N_1590,N_1057,N_948);
nand U1591 (N_1591,N_1215,N_1021);
or U1592 (N_1592,N_1164,N_1223);
or U1593 (N_1593,N_1208,N_1001);
or U1594 (N_1594,N_1488,N_869);
or U1595 (N_1595,N_1126,N_786);
nand U1596 (N_1596,N_834,N_1091);
nand U1597 (N_1597,N_1177,N_1234);
or U1598 (N_1598,N_1485,N_1324);
nor U1599 (N_1599,N_1489,N_1114);
nand U1600 (N_1600,N_1341,N_1211);
or U1601 (N_1601,N_1298,N_949);
and U1602 (N_1602,N_1096,N_1045);
nor U1603 (N_1603,N_1481,N_1389);
or U1604 (N_1604,N_1443,N_791);
and U1605 (N_1605,N_852,N_887);
nand U1606 (N_1606,N_1166,N_1263);
or U1607 (N_1607,N_796,N_1150);
nand U1608 (N_1608,N_1050,N_1257);
and U1609 (N_1609,N_1167,N_1470);
nand U1610 (N_1610,N_926,N_1191);
nand U1611 (N_1611,N_787,N_813);
and U1612 (N_1612,N_1471,N_1225);
or U1613 (N_1613,N_1319,N_1040);
or U1614 (N_1614,N_969,N_1270);
nor U1615 (N_1615,N_1317,N_778);
xnor U1616 (N_1616,N_1079,N_1318);
nor U1617 (N_1617,N_1051,N_1090);
and U1618 (N_1618,N_901,N_907);
nand U1619 (N_1619,N_1265,N_989);
xnor U1620 (N_1620,N_1495,N_1286);
or U1621 (N_1621,N_1357,N_981);
or U1622 (N_1622,N_1017,N_761);
nand U1623 (N_1623,N_1204,N_1116);
nor U1624 (N_1624,N_1292,N_936);
nand U1625 (N_1625,N_954,N_974);
or U1626 (N_1626,N_1043,N_1271);
and U1627 (N_1627,N_997,N_1010);
nor U1628 (N_1628,N_911,N_1440);
and U1629 (N_1629,N_1266,N_812);
nand U1630 (N_1630,N_1333,N_878);
nand U1631 (N_1631,N_950,N_794);
xnor U1632 (N_1632,N_1343,N_1024);
xnor U1633 (N_1633,N_1125,N_1375);
and U1634 (N_1634,N_941,N_1337);
and U1635 (N_1635,N_953,N_1313);
xor U1636 (N_1636,N_1346,N_895);
nor U1637 (N_1637,N_1033,N_1342);
and U1638 (N_1638,N_811,N_1246);
and U1639 (N_1639,N_1255,N_764);
nor U1640 (N_1640,N_1486,N_1413);
nand U1641 (N_1641,N_1493,N_1264);
xor U1642 (N_1642,N_1367,N_872);
or U1643 (N_1643,N_831,N_1406);
nand U1644 (N_1644,N_770,N_850);
xor U1645 (N_1645,N_938,N_1044);
nor U1646 (N_1646,N_917,N_1262);
xor U1647 (N_1647,N_1088,N_1380);
nand U1648 (N_1648,N_792,N_1410);
nand U1649 (N_1649,N_933,N_1019);
and U1650 (N_1650,N_996,N_1170);
xnor U1651 (N_1651,N_1487,N_1334);
nand U1652 (N_1652,N_1276,N_1331);
and U1653 (N_1653,N_1194,N_1260);
nand U1654 (N_1654,N_1107,N_993);
nand U1655 (N_1655,N_958,N_1160);
nor U1656 (N_1656,N_1074,N_1354);
and U1657 (N_1657,N_752,N_1041);
and U1658 (N_1658,N_1415,N_1450);
and U1659 (N_1659,N_890,N_1089);
nand U1660 (N_1660,N_868,N_923);
nand U1661 (N_1661,N_1154,N_1388);
and U1662 (N_1662,N_1128,N_1062);
xnor U1663 (N_1663,N_760,N_1281);
and U1664 (N_1664,N_982,N_1320);
nand U1665 (N_1665,N_1425,N_1499);
and U1666 (N_1666,N_1015,N_1046);
nand U1667 (N_1667,N_1098,N_1219);
and U1668 (N_1668,N_851,N_1296);
and U1669 (N_1669,N_1078,N_1408);
and U1670 (N_1670,N_1011,N_888);
xor U1671 (N_1671,N_1457,N_1390);
and U1672 (N_1672,N_1136,N_1418);
nor U1673 (N_1673,N_801,N_1028);
or U1674 (N_1674,N_1149,N_1259);
xnor U1675 (N_1675,N_1119,N_1484);
nor U1676 (N_1676,N_1315,N_976);
or U1677 (N_1677,N_992,N_1093);
and U1678 (N_1678,N_807,N_1200);
nand U1679 (N_1679,N_1222,N_1411);
or U1680 (N_1680,N_1309,N_1399);
and U1681 (N_1681,N_862,N_1235);
or U1682 (N_1682,N_1291,N_952);
or U1683 (N_1683,N_847,N_1277);
nand U1684 (N_1684,N_998,N_1453);
nor U1685 (N_1685,N_1361,N_1109);
nand U1686 (N_1686,N_1081,N_1433);
nor U1687 (N_1687,N_980,N_1168);
xor U1688 (N_1688,N_769,N_1447);
xnor U1689 (N_1689,N_1135,N_1245);
xor U1690 (N_1690,N_846,N_880);
xor U1691 (N_1691,N_1446,N_1155);
and U1692 (N_1692,N_1476,N_1032);
nor U1693 (N_1693,N_957,N_1179);
nor U1694 (N_1694,N_819,N_1025);
or U1695 (N_1695,N_1303,N_1110);
xor U1696 (N_1696,N_1363,N_751);
nand U1697 (N_1697,N_871,N_1238);
nand U1698 (N_1698,N_922,N_1330);
nor U1699 (N_1699,N_855,N_779);
nor U1700 (N_1700,N_1294,N_1301);
or U1701 (N_1701,N_1356,N_1244);
nor U1702 (N_1702,N_1327,N_1345);
and U1703 (N_1703,N_1360,N_983);
nor U1704 (N_1704,N_891,N_1233);
nand U1705 (N_1705,N_1077,N_1376);
and U1706 (N_1706,N_1113,N_991);
or U1707 (N_1707,N_1437,N_765);
nand U1708 (N_1708,N_1251,N_925);
or U1709 (N_1709,N_827,N_808);
or U1710 (N_1710,N_1095,N_828);
nor U1711 (N_1711,N_1326,N_951);
xor U1712 (N_1712,N_845,N_1420);
xor U1713 (N_1713,N_910,N_1163);
nor U1714 (N_1714,N_935,N_804);
nand U1715 (N_1715,N_879,N_1379);
or U1716 (N_1716,N_1029,N_1188);
and U1717 (N_1717,N_1349,N_970);
or U1718 (N_1718,N_1221,N_943);
nand U1719 (N_1719,N_885,N_1087);
nand U1720 (N_1720,N_1218,N_843);
nor U1721 (N_1721,N_1384,N_896);
nand U1722 (N_1722,N_1196,N_1338);
nor U1723 (N_1723,N_965,N_1102);
xor U1724 (N_1724,N_1285,N_962);
or U1725 (N_1725,N_1132,N_1056);
nor U1726 (N_1726,N_1100,N_1182);
or U1727 (N_1727,N_1068,N_1477);
and U1728 (N_1728,N_975,N_1103);
and U1729 (N_1729,N_984,N_854);
and U1730 (N_1730,N_775,N_782);
or U1731 (N_1731,N_1366,N_1175);
xor U1732 (N_1732,N_900,N_1293);
nand U1733 (N_1733,N_1383,N_781);
nor U1734 (N_1734,N_1072,N_1468);
or U1735 (N_1735,N_1387,N_1423);
nand U1736 (N_1736,N_1490,N_1459);
and U1737 (N_1737,N_866,N_1210);
xor U1738 (N_1738,N_844,N_773);
nor U1739 (N_1739,N_955,N_1304);
and U1740 (N_1740,N_1134,N_931);
and U1741 (N_1741,N_1067,N_823);
and U1742 (N_1742,N_1288,N_892);
nand U1743 (N_1743,N_1321,N_927);
or U1744 (N_1744,N_894,N_1082);
nor U1745 (N_1745,N_1066,N_840);
nor U1746 (N_1746,N_1012,N_1279);
nor U1747 (N_1747,N_1055,N_960);
or U1748 (N_1748,N_966,N_1430);
nor U1749 (N_1749,N_1353,N_1027);
nor U1750 (N_1750,N_867,N_914);
or U1751 (N_1751,N_1444,N_987);
or U1752 (N_1752,N_1496,N_1394);
and U1753 (N_1753,N_1416,N_1365);
nor U1754 (N_1754,N_777,N_1369);
xor U1755 (N_1755,N_1198,N_1120);
and U1756 (N_1756,N_841,N_1159);
and U1757 (N_1757,N_1405,N_1466);
nand U1758 (N_1758,N_973,N_1022);
nand U1759 (N_1759,N_1438,N_799);
or U1760 (N_1760,N_1094,N_820);
nand U1761 (N_1761,N_1130,N_1335);
and U1762 (N_1762,N_1355,N_1242);
or U1763 (N_1763,N_1382,N_978);
and U1764 (N_1764,N_797,N_1181);
and U1765 (N_1765,N_988,N_1216);
nor U1766 (N_1766,N_1480,N_886);
or U1767 (N_1767,N_1195,N_1475);
xor U1768 (N_1768,N_1143,N_1449);
xnor U1769 (N_1769,N_1429,N_1421);
nor U1770 (N_1770,N_824,N_906);
or U1771 (N_1771,N_1403,N_1445);
xnor U1772 (N_1772,N_1460,N_1140);
xor U1773 (N_1773,N_817,N_1173);
and U1774 (N_1774,N_1290,N_1065);
xor U1775 (N_1775,N_956,N_934);
or U1776 (N_1776,N_1039,N_1432);
xor U1777 (N_1777,N_1205,N_1261);
nand U1778 (N_1778,N_798,N_1058);
xnor U1779 (N_1779,N_1400,N_1402);
xor U1780 (N_1780,N_1240,N_1295);
nand U1781 (N_1781,N_961,N_1311);
and U1782 (N_1782,N_1212,N_839);
nand U1783 (N_1783,N_1036,N_842);
xnor U1784 (N_1784,N_860,N_1479);
xor U1785 (N_1785,N_1157,N_968);
or U1786 (N_1786,N_1054,N_1283);
and U1787 (N_1787,N_1336,N_1071);
or U1788 (N_1788,N_944,N_1031);
nor U1789 (N_1789,N_1141,N_1268);
and U1790 (N_1790,N_1362,N_822);
nand U1791 (N_1791,N_995,N_826);
and U1792 (N_1792,N_793,N_874);
and U1793 (N_1793,N_790,N_1454);
or U1794 (N_1794,N_1316,N_830);
xnor U1795 (N_1795,N_1378,N_1282);
nor U1796 (N_1796,N_849,N_1092);
nor U1797 (N_1797,N_1127,N_1230);
and U1798 (N_1798,N_1441,N_774);
xnor U1799 (N_1799,N_1197,N_1101);
nand U1800 (N_1800,N_1104,N_918);
xor U1801 (N_1801,N_1142,N_1124);
xnor U1802 (N_1802,N_1370,N_1156);
and U1803 (N_1803,N_1280,N_1189);
and U1804 (N_1804,N_836,N_853);
and U1805 (N_1805,N_942,N_1310);
xor U1806 (N_1806,N_1494,N_1151);
nand U1807 (N_1807,N_985,N_1258);
xnor U1808 (N_1808,N_1348,N_1483);
xor U1809 (N_1809,N_1289,N_1364);
and U1810 (N_1810,N_757,N_829);
and U1811 (N_1811,N_763,N_870);
nand U1812 (N_1812,N_1115,N_1465);
and U1813 (N_1813,N_1213,N_1431);
nor U1814 (N_1814,N_1396,N_1193);
nor U1815 (N_1815,N_1249,N_893);
or U1816 (N_1816,N_1186,N_1497);
or U1817 (N_1817,N_897,N_977);
xor U1818 (N_1818,N_1073,N_1112);
nor U1819 (N_1819,N_1275,N_806);
and U1820 (N_1820,N_1442,N_1083);
xnor U1821 (N_1821,N_1422,N_1003);
nand U1822 (N_1822,N_947,N_1474);
and U1823 (N_1823,N_905,N_1207);
nand U1824 (N_1824,N_864,N_1158);
nor U1825 (N_1825,N_1347,N_1224);
xor U1826 (N_1826,N_971,N_1030);
or U1827 (N_1827,N_881,N_1034);
and U1828 (N_1828,N_1329,N_1232);
and U1829 (N_1829,N_1169,N_1201);
xor U1830 (N_1830,N_1306,N_1498);
nor U1831 (N_1831,N_776,N_1190);
nand U1832 (N_1832,N_1308,N_1322);
nor U1833 (N_1833,N_1237,N_1439);
xor U1834 (N_1834,N_821,N_1059);
nor U1835 (N_1835,N_946,N_1267);
and U1836 (N_1836,N_1026,N_784);
nand U1837 (N_1837,N_1209,N_1492);
nor U1838 (N_1838,N_990,N_1299);
or U1839 (N_1839,N_1048,N_810);
xnor U1840 (N_1840,N_1368,N_783);
xnor U1841 (N_1841,N_1464,N_1284);
nor U1842 (N_1842,N_1037,N_928);
xnor U1843 (N_1843,N_999,N_1463);
and U1844 (N_1844,N_1174,N_902);
and U1845 (N_1845,N_762,N_1122);
xnor U1846 (N_1846,N_1106,N_814);
and U1847 (N_1847,N_833,N_883);
xor U1848 (N_1848,N_1180,N_832);
or U1849 (N_1849,N_1129,N_1099);
nand U1850 (N_1850,N_1461,N_1199);
nand U1851 (N_1851,N_1377,N_1297);
nand U1852 (N_1852,N_945,N_1472);
nand U1853 (N_1853,N_835,N_1398);
xnor U1854 (N_1854,N_1419,N_1351);
nor U1855 (N_1855,N_780,N_986);
nor U1856 (N_1856,N_1344,N_899);
or U1857 (N_1857,N_772,N_1409);
nand U1858 (N_1858,N_1307,N_967);
and U1859 (N_1859,N_865,N_1161);
and U1860 (N_1860,N_754,N_1482);
and U1861 (N_1861,N_1456,N_768);
nor U1862 (N_1862,N_1252,N_908);
and U1863 (N_1863,N_1359,N_1404);
xor U1864 (N_1864,N_889,N_1108);
xor U1865 (N_1865,N_1436,N_856);
or U1866 (N_1866,N_921,N_1312);
or U1867 (N_1867,N_795,N_1287);
xor U1868 (N_1868,N_1145,N_766);
nor U1869 (N_1869,N_1016,N_805);
and U1870 (N_1870,N_1137,N_1146);
or U1871 (N_1871,N_1002,N_1239);
and U1872 (N_1872,N_1469,N_1008);
and U1873 (N_1873,N_1153,N_785);
xnor U1874 (N_1874,N_1323,N_1417);
xnor U1875 (N_1875,N_965,N_989);
and U1876 (N_1876,N_1329,N_896);
nor U1877 (N_1877,N_1090,N_1077);
xnor U1878 (N_1878,N_825,N_1316);
and U1879 (N_1879,N_968,N_1124);
or U1880 (N_1880,N_871,N_1457);
nand U1881 (N_1881,N_1415,N_909);
xor U1882 (N_1882,N_966,N_1433);
xnor U1883 (N_1883,N_1449,N_1036);
and U1884 (N_1884,N_785,N_802);
xnor U1885 (N_1885,N_937,N_1404);
nand U1886 (N_1886,N_1115,N_1253);
nand U1887 (N_1887,N_1390,N_1375);
and U1888 (N_1888,N_1342,N_778);
nand U1889 (N_1889,N_955,N_1224);
nor U1890 (N_1890,N_971,N_1157);
xnor U1891 (N_1891,N_1064,N_1326);
nor U1892 (N_1892,N_1464,N_1169);
xor U1893 (N_1893,N_1148,N_965);
nand U1894 (N_1894,N_861,N_1269);
xor U1895 (N_1895,N_1437,N_876);
nand U1896 (N_1896,N_891,N_1380);
or U1897 (N_1897,N_1478,N_1022);
or U1898 (N_1898,N_1086,N_890);
nor U1899 (N_1899,N_1277,N_1439);
nor U1900 (N_1900,N_1007,N_1028);
or U1901 (N_1901,N_908,N_920);
nor U1902 (N_1902,N_895,N_1105);
nor U1903 (N_1903,N_974,N_894);
xnor U1904 (N_1904,N_1245,N_886);
or U1905 (N_1905,N_789,N_1131);
xnor U1906 (N_1906,N_917,N_798);
nand U1907 (N_1907,N_1215,N_775);
or U1908 (N_1908,N_970,N_756);
and U1909 (N_1909,N_755,N_1156);
nor U1910 (N_1910,N_1061,N_757);
nor U1911 (N_1911,N_1265,N_1328);
xnor U1912 (N_1912,N_1121,N_793);
or U1913 (N_1913,N_1388,N_1009);
or U1914 (N_1914,N_814,N_933);
nand U1915 (N_1915,N_1208,N_851);
xor U1916 (N_1916,N_1415,N_1088);
xor U1917 (N_1917,N_832,N_1188);
xnor U1918 (N_1918,N_1355,N_1162);
nor U1919 (N_1919,N_872,N_905);
nor U1920 (N_1920,N_1126,N_1407);
xnor U1921 (N_1921,N_1266,N_1271);
nor U1922 (N_1922,N_942,N_1158);
nand U1923 (N_1923,N_1178,N_1123);
xor U1924 (N_1924,N_925,N_1221);
nor U1925 (N_1925,N_1312,N_1141);
or U1926 (N_1926,N_1102,N_1249);
xor U1927 (N_1927,N_907,N_895);
xnor U1928 (N_1928,N_1434,N_1334);
or U1929 (N_1929,N_996,N_1495);
nand U1930 (N_1930,N_1378,N_804);
nor U1931 (N_1931,N_867,N_823);
xnor U1932 (N_1932,N_1045,N_1129);
nand U1933 (N_1933,N_1099,N_1013);
and U1934 (N_1934,N_871,N_1264);
nor U1935 (N_1935,N_962,N_1336);
nand U1936 (N_1936,N_872,N_1473);
nor U1937 (N_1937,N_1389,N_777);
or U1938 (N_1938,N_1361,N_1070);
nor U1939 (N_1939,N_1176,N_775);
nand U1940 (N_1940,N_1078,N_1112);
or U1941 (N_1941,N_1169,N_1034);
or U1942 (N_1942,N_1048,N_953);
and U1943 (N_1943,N_1413,N_1330);
xnor U1944 (N_1944,N_1451,N_1444);
and U1945 (N_1945,N_1165,N_753);
nor U1946 (N_1946,N_1176,N_1386);
nand U1947 (N_1947,N_1008,N_1199);
xnor U1948 (N_1948,N_1109,N_1055);
and U1949 (N_1949,N_1299,N_1213);
and U1950 (N_1950,N_1146,N_1075);
and U1951 (N_1951,N_755,N_1432);
xnor U1952 (N_1952,N_1098,N_1379);
and U1953 (N_1953,N_1406,N_1186);
or U1954 (N_1954,N_1296,N_880);
or U1955 (N_1955,N_1269,N_953);
nor U1956 (N_1956,N_1351,N_1402);
nor U1957 (N_1957,N_1430,N_1086);
xor U1958 (N_1958,N_1276,N_760);
and U1959 (N_1959,N_1059,N_931);
and U1960 (N_1960,N_1065,N_1254);
nor U1961 (N_1961,N_970,N_1444);
or U1962 (N_1962,N_1014,N_841);
xor U1963 (N_1963,N_1296,N_1077);
nand U1964 (N_1964,N_984,N_1164);
or U1965 (N_1965,N_937,N_812);
or U1966 (N_1966,N_1375,N_978);
xnor U1967 (N_1967,N_1295,N_989);
and U1968 (N_1968,N_974,N_1230);
xor U1969 (N_1969,N_997,N_1217);
xnor U1970 (N_1970,N_986,N_1307);
xor U1971 (N_1971,N_1125,N_939);
or U1972 (N_1972,N_811,N_1316);
nor U1973 (N_1973,N_1004,N_849);
nor U1974 (N_1974,N_1369,N_1496);
nand U1975 (N_1975,N_881,N_1126);
nand U1976 (N_1976,N_874,N_1269);
xnor U1977 (N_1977,N_1408,N_1250);
xor U1978 (N_1978,N_961,N_956);
nor U1979 (N_1979,N_924,N_1200);
xor U1980 (N_1980,N_1264,N_818);
nor U1981 (N_1981,N_1152,N_1096);
nor U1982 (N_1982,N_1432,N_1368);
nor U1983 (N_1983,N_920,N_1008);
or U1984 (N_1984,N_1433,N_1400);
nor U1985 (N_1985,N_785,N_912);
and U1986 (N_1986,N_815,N_1080);
and U1987 (N_1987,N_1128,N_1377);
or U1988 (N_1988,N_761,N_1279);
or U1989 (N_1989,N_1309,N_803);
and U1990 (N_1990,N_1325,N_1375);
or U1991 (N_1991,N_776,N_1000);
nand U1992 (N_1992,N_1347,N_1354);
xnor U1993 (N_1993,N_1286,N_1417);
or U1994 (N_1994,N_1304,N_1173);
xor U1995 (N_1995,N_1101,N_1462);
or U1996 (N_1996,N_872,N_1229);
or U1997 (N_1997,N_866,N_1025);
or U1998 (N_1998,N_1405,N_768);
nand U1999 (N_1999,N_1022,N_1144);
or U2000 (N_2000,N_1264,N_1459);
or U2001 (N_2001,N_1249,N_861);
nand U2002 (N_2002,N_944,N_1075);
nor U2003 (N_2003,N_1081,N_1058);
xnor U2004 (N_2004,N_1145,N_1274);
xnor U2005 (N_2005,N_834,N_1026);
and U2006 (N_2006,N_1097,N_1007);
nor U2007 (N_2007,N_1351,N_1137);
nor U2008 (N_2008,N_929,N_1090);
or U2009 (N_2009,N_1472,N_906);
nand U2010 (N_2010,N_1350,N_808);
or U2011 (N_2011,N_788,N_1440);
and U2012 (N_2012,N_1336,N_1408);
and U2013 (N_2013,N_1347,N_1455);
nand U2014 (N_2014,N_980,N_882);
or U2015 (N_2015,N_1104,N_1482);
xnor U2016 (N_2016,N_1354,N_1239);
xor U2017 (N_2017,N_1029,N_1065);
nor U2018 (N_2018,N_844,N_1470);
and U2019 (N_2019,N_1127,N_1015);
and U2020 (N_2020,N_1309,N_984);
or U2021 (N_2021,N_1112,N_1139);
nand U2022 (N_2022,N_762,N_1376);
or U2023 (N_2023,N_864,N_1450);
nand U2024 (N_2024,N_794,N_1126);
nand U2025 (N_2025,N_1017,N_1191);
xnor U2026 (N_2026,N_844,N_1194);
xnor U2027 (N_2027,N_1255,N_781);
or U2028 (N_2028,N_901,N_1001);
nand U2029 (N_2029,N_842,N_1317);
nor U2030 (N_2030,N_916,N_1245);
and U2031 (N_2031,N_922,N_1288);
nand U2032 (N_2032,N_799,N_1337);
and U2033 (N_2033,N_1212,N_1244);
and U2034 (N_2034,N_1028,N_850);
nand U2035 (N_2035,N_776,N_1060);
nor U2036 (N_2036,N_1313,N_1449);
and U2037 (N_2037,N_930,N_853);
or U2038 (N_2038,N_1222,N_795);
xnor U2039 (N_2039,N_770,N_869);
nor U2040 (N_2040,N_1074,N_1374);
xor U2041 (N_2041,N_790,N_1064);
or U2042 (N_2042,N_990,N_1168);
nor U2043 (N_2043,N_1332,N_1477);
nor U2044 (N_2044,N_870,N_1081);
nand U2045 (N_2045,N_1032,N_976);
xnor U2046 (N_2046,N_965,N_1042);
nand U2047 (N_2047,N_1433,N_1468);
nand U2048 (N_2048,N_1315,N_1471);
xor U2049 (N_2049,N_779,N_757);
or U2050 (N_2050,N_781,N_1345);
nand U2051 (N_2051,N_1020,N_963);
nand U2052 (N_2052,N_961,N_872);
nand U2053 (N_2053,N_759,N_1195);
and U2054 (N_2054,N_1414,N_880);
nor U2055 (N_2055,N_1278,N_750);
or U2056 (N_2056,N_1363,N_1435);
and U2057 (N_2057,N_1422,N_1163);
nand U2058 (N_2058,N_764,N_877);
xnor U2059 (N_2059,N_1082,N_1412);
and U2060 (N_2060,N_955,N_1050);
nand U2061 (N_2061,N_988,N_1117);
and U2062 (N_2062,N_984,N_899);
nor U2063 (N_2063,N_1411,N_854);
xor U2064 (N_2064,N_936,N_1365);
and U2065 (N_2065,N_1467,N_1214);
xnor U2066 (N_2066,N_1444,N_1279);
nor U2067 (N_2067,N_1075,N_970);
and U2068 (N_2068,N_1020,N_1101);
or U2069 (N_2069,N_1403,N_1241);
xnor U2070 (N_2070,N_1439,N_1344);
nor U2071 (N_2071,N_834,N_826);
or U2072 (N_2072,N_806,N_767);
nand U2073 (N_2073,N_984,N_786);
or U2074 (N_2074,N_1241,N_1006);
nor U2075 (N_2075,N_917,N_1286);
and U2076 (N_2076,N_822,N_1125);
and U2077 (N_2077,N_1183,N_1444);
nor U2078 (N_2078,N_896,N_957);
nand U2079 (N_2079,N_1241,N_1144);
nor U2080 (N_2080,N_914,N_1015);
and U2081 (N_2081,N_1232,N_1150);
nand U2082 (N_2082,N_1388,N_753);
and U2083 (N_2083,N_1000,N_1209);
nor U2084 (N_2084,N_992,N_790);
and U2085 (N_2085,N_1037,N_1268);
nand U2086 (N_2086,N_1185,N_1099);
nor U2087 (N_2087,N_941,N_1112);
nor U2088 (N_2088,N_1474,N_921);
nand U2089 (N_2089,N_857,N_986);
nand U2090 (N_2090,N_852,N_1384);
nand U2091 (N_2091,N_1322,N_1428);
nor U2092 (N_2092,N_1014,N_792);
and U2093 (N_2093,N_1488,N_812);
and U2094 (N_2094,N_1193,N_1149);
nor U2095 (N_2095,N_1482,N_1322);
or U2096 (N_2096,N_872,N_1345);
or U2097 (N_2097,N_989,N_1089);
or U2098 (N_2098,N_1160,N_1394);
nor U2099 (N_2099,N_1353,N_1159);
nand U2100 (N_2100,N_1063,N_939);
and U2101 (N_2101,N_1322,N_1248);
nor U2102 (N_2102,N_872,N_1090);
nand U2103 (N_2103,N_1320,N_1360);
nand U2104 (N_2104,N_1265,N_827);
or U2105 (N_2105,N_922,N_1215);
xnor U2106 (N_2106,N_1027,N_1163);
nand U2107 (N_2107,N_1418,N_966);
nand U2108 (N_2108,N_1033,N_1090);
nand U2109 (N_2109,N_1372,N_1274);
nor U2110 (N_2110,N_814,N_859);
nand U2111 (N_2111,N_938,N_1436);
or U2112 (N_2112,N_1495,N_915);
xnor U2113 (N_2113,N_1310,N_1409);
or U2114 (N_2114,N_878,N_1179);
and U2115 (N_2115,N_1142,N_1398);
nor U2116 (N_2116,N_811,N_1432);
nand U2117 (N_2117,N_779,N_1066);
xnor U2118 (N_2118,N_1409,N_1171);
nor U2119 (N_2119,N_1250,N_836);
nor U2120 (N_2120,N_1380,N_1208);
or U2121 (N_2121,N_1159,N_1263);
nand U2122 (N_2122,N_1249,N_977);
xor U2123 (N_2123,N_1277,N_1319);
nor U2124 (N_2124,N_1007,N_1148);
nand U2125 (N_2125,N_896,N_1215);
or U2126 (N_2126,N_1491,N_1121);
xor U2127 (N_2127,N_1072,N_1235);
nand U2128 (N_2128,N_828,N_1078);
or U2129 (N_2129,N_1186,N_980);
nor U2130 (N_2130,N_763,N_1330);
and U2131 (N_2131,N_1342,N_965);
nand U2132 (N_2132,N_971,N_863);
and U2133 (N_2133,N_760,N_1457);
xnor U2134 (N_2134,N_1498,N_1285);
nand U2135 (N_2135,N_1352,N_1475);
nor U2136 (N_2136,N_1018,N_859);
nand U2137 (N_2137,N_1456,N_1470);
xnor U2138 (N_2138,N_1232,N_787);
nor U2139 (N_2139,N_1379,N_1384);
nor U2140 (N_2140,N_1492,N_915);
and U2141 (N_2141,N_1025,N_845);
nor U2142 (N_2142,N_959,N_1183);
nand U2143 (N_2143,N_1481,N_1353);
and U2144 (N_2144,N_1385,N_1108);
and U2145 (N_2145,N_936,N_1485);
nand U2146 (N_2146,N_1337,N_1105);
or U2147 (N_2147,N_1499,N_828);
or U2148 (N_2148,N_1369,N_1245);
xnor U2149 (N_2149,N_1433,N_1052);
nand U2150 (N_2150,N_1207,N_1281);
nor U2151 (N_2151,N_1004,N_784);
or U2152 (N_2152,N_1236,N_1115);
and U2153 (N_2153,N_904,N_1009);
and U2154 (N_2154,N_1182,N_803);
or U2155 (N_2155,N_1459,N_1329);
xor U2156 (N_2156,N_914,N_1411);
and U2157 (N_2157,N_859,N_984);
or U2158 (N_2158,N_890,N_838);
xor U2159 (N_2159,N_1274,N_1068);
xnor U2160 (N_2160,N_1299,N_1410);
nand U2161 (N_2161,N_1235,N_918);
and U2162 (N_2162,N_1066,N_1406);
nor U2163 (N_2163,N_1081,N_978);
and U2164 (N_2164,N_1142,N_1081);
nand U2165 (N_2165,N_1088,N_1313);
or U2166 (N_2166,N_882,N_1480);
or U2167 (N_2167,N_1343,N_1279);
nand U2168 (N_2168,N_1358,N_1019);
or U2169 (N_2169,N_934,N_988);
xor U2170 (N_2170,N_1264,N_1096);
and U2171 (N_2171,N_1234,N_1056);
nor U2172 (N_2172,N_1488,N_1141);
xnor U2173 (N_2173,N_960,N_847);
nand U2174 (N_2174,N_1019,N_872);
and U2175 (N_2175,N_1099,N_761);
or U2176 (N_2176,N_1197,N_1276);
xnor U2177 (N_2177,N_985,N_814);
xor U2178 (N_2178,N_1374,N_1197);
nor U2179 (N_2179,N_1352,N_1183);
nand U2180 (N_2180,N_1239,N_1496);
nor U2181 (N_2181,N_835,N_1272);
xnor U2182 (N_2182,N_1028,N_793);
xor U2183 (N_2183,N_1317,N_985);
xor U2184 (N_2184,N_1296,N_875);
xor U2185 (N_2185,N_1178,N_1101);
or U2186 (N_2186,N_781,N_1027);
or U2187 (N_2187,N_962,N_1447);
nor U2188 (N_2188,N_1321,N_1476);
or U2189 (N_2189,N_755,N_1229);
nor U2190 (N_2190,N_799,N_1233);
xor U2191 (N_2191,N_1116,N_1211);
nand U2192 (N_2192,N_1050,N_1182);
xnor U2193 (N_2193,N_779,N_1381);
or U2194 (N_2194,N_1082,N_999);
nand U2195 (N_2195,N_1289,N_1476);
nand U2196 (N_2196,N_854,N_994);
or U2197 (N_2197,N_966,N_1151);
nor U2198 (N_2198,N_1129,N_1325);
nor U2199 (N_2199,N_805,N_798);
nand U2200 (N_2200,N_834,N_1328);
nor U2201 (N_2201,N_1083,N_849);
xnor U2202 (N_2202,N_1066,N_1378);
xnor U2203 (N_2203,N_1041,N_995);
xor U2204 (N_2204,N_1416,N_1113);
nand U2205 (N_2205,N_1277,N_910);
nand U2206 (N_2206,N_1004,N_1029);
or U2207 (N_2207,N_855,N_798);
or U2208 (N_2208,N_1404,N_1119);
xor U2209 (N_2209,N_1433,N_782);
or U2210 (N_2210,N_897,N_1256);
nor U2211 (N_2211,N_1162,N_872);
nand U2212 (N_2212,N_1171,N_1100);
nor U2213 (N_2213,N_1130,N_1208);
nor U2214 (N_2214,N_1029,N_1025);
nor U2215 (N_2215,N_1453,N_919);
or U2216 (N_2216,N_1155,N_1243);
nand U2217 (N_2217,N_1308,N_1218);
nand U2218 (N_2218,N_1386,N_1283);
nand U2219 (N_2219,N_1304,N_1332);
and U2220 (N_2220,N_1138,N_1418);
or U2221 (N_2221,N_1369,N_1044);
or U2222 (N_2222,N_1058,N_1424);
nor U2223 (N_2223,N_1023,N_1084);
nand U2224 (N_2224,N_1209,N_1272);
nor U2225 (N_2225,N_1039,N_935);
nand U2226 (N_2226,N_1052,N_1303);
nor U2227 (N_2227,N_1259,N_1424);
and U2228 (N_2228,N_1258,N_806);
or U2229 (N_2229,N_1137,N_1008);
nor U2230 (N_2230,N_897,N_1412);
or U2231 (N_2231,N_933,N_1028);
and U2232 (N_2232,N_1261,N_849);
nand U2233 (N_2233,N_1236,N_1099);
xnor U2234 (N_2234,N_1345,N_1309);
and U2235 (N_2235,N_1304,N_1426);
and U2236 (N_2236,N_898,N_1422);
xor U2237 (N_2237,N_1018,N_1269);
and U2238 (N_2238,N_803,N_1026);
nand U2239 (N_2239,N_1278,N_1327);
xnor U2240 (N_2240,N_1253,N_756);
xnor U2241 (N_2241,N_1447,N_1086);
or U2242 (N_2242,N_833,N_1277);
xor U2243 (N_2243,N_1055,N_1310);
nand U2244 (N_2244,N_1188,N_824);
xnor U2245 (N_2245,N_1401,N_1212);
xor U2246 (N_2246,N_952,N_1145);
nor U2247 (N_2247,N_978,N_1150);
xor U2248 (N_2248,N_1342,N_1431);
or U2249 (N_2249,N_755,N_1297);
and U2250 (N_2250,N_2193,N_1630);
and U2251 (N_2251,N_1980,N_2244);
or U2252 (N_2252,N_1807,N_1584);
or U2253 (N_2253,N_1733,N_1548);
or U2254 (N_2254,N_2038,N_1923);
nand U2255 (N_2255,N_2198,N_1776);
or U2256 (N_2256,N_2080,N_1782);
nand U2257 (N_2257,N_1576,N_1975);
nor U2258 (N_2258,N_1617,N_2046);
or U2259 (N_2259,N_2060,N_1608);
nor U2260 (N_2260,N_1528,N_1639);
and U2261 (N_2261,N_2133,N_2052);
xor U2262 (N_2262,N_2197,N_2100);
xnor U2263 (N_2263,N_2238,N_2073);
and U2264 (N_2264,N_1708,N_2087);
nor U2265 (N_2265,N_1764,N_2158);
xnor U2266 (N_2266,N_2191,N_2109);
and U2267 (N_2267,N_2248,N_2173);
nor U2268 (N_2268,N_1737,N_1832);
xor U2269 (N_2269,N_1623,N_1973);
and U2270 (N_2270,N_1751,N_1594);
and U2271 (N_2271,N_1819,N_1982);
or U2272 (N_2272,N_1673,N_2170);
xnor U2273 (N_2273,N_2008,N_2129);
nor U2274 (N_2274,N_1948,N_1785);
xor U2275 (N_2275,N_2218,N_1526);
or U2276 (N_2276,N_1981,N_1892);
and U2277 (N_2277,N_2010,N_2005);
and U2278 (N_2278,N_2171,N_1521);
xor U2279 (N_2279,N_1820,N_2051);
nand U2280 (N_2280,N_1582,N_1652);
nor U2281 (N_2281,N_2110,N_1882);
and U2282 (N_2282,N_1878,N_1543);
nand U2283 (N_2283,N_2172,N_1739);
or U2284 (N_2284,N_2131,N_2246);
xor U2285 (N_2285,N_1836,N_1653);
nand U2286 (N_2286,N_1924,N_2032);
nand U2287 (N_2287,N_1587,N_1602);
and U2288 (N_2288,N_2077,N_1760);
xor U2289 (N_2289,N_2071,N_2203);
nand U2290 (N_2290,N_1796,N_1884);
nor U2291 (N_2291,N_1964,N_1801);
and U2292 (N_2292,N_1599,N_2162);
nor U2293 (N_2293,N_1757,N_1985);
or U2294 (N_2294,N_2020,N_2088);
nand U2295 (N_2295,N_1978,N_2013);
and U2296 (N_2296,N_2009,N_1971);
or U2297 (N_2297,N_1694,N_1512);
xnor U2298 (N_2298,N_1937,N_1687);
and U2299 (N_2299,N_1644,N_2164);
xnor U2300 (N_2300,N_1508,N_1569);
nand U2301 (N_2301,N_2030,N_2095);
nand U2302 (N_2302,N_2112,N_2204);
and U2303 (N_2303,N_2002,N_2167);
xnor U2304 (N_2304,N_1645,N_2019);
and U2305 (N_2305,N_2120,N_1952);
or U2306 (N_2306,N_1936,N_2169);
nand U2307 (N_2307,N_1646,N_1993);
and U2308 (N_2308,N_1795,N_1724);
and U2309 (N_2309,N_2111,N_2039);
and U2310 (N_2310,N_1697,N_1792);
nand U2311 (N_2311,N_1956,N_2006);
or U2312 (N_2312,N_2083,N_1943);
or U2313 (N_2313,N_1953,N_1744);
or U2314 (N_2314,N_1632,N_1814);
or U2315 (N_2315,N_1949,N_1596);
or U2316 (N_2316,N_1709,N_1794);
and U2317 (N_2317,N_1773,N_1590);
or U2318 (N_2318,N_1509,N_1960);
nand U2319 (N_2319,N_1604,N_2078);
nor U2320 (N_2320,N_1929,N_1869);
and U2321 (N_2321,N_2176,N_1791);
and U2322 (N_2322,N_1532,N_1655);
nand U2323 (N_2323,N_2225,N_1585);
nor U2324 (N_2324,N_1809,N_2143);
nand U2325 (N_2325,N_2177,N_2175);
nand U2326 (N_2326,N_1925,N_1752);
nor U2327 (N_2327,N_1665,N_2042);
nor U2328 (N_2328,N_1805,N_2242);
nand U2329 (N_2329,N_1502,N_1988);
and U2330 (N_2330,N_1547,N_1802);
or U2331 (N_2331,N_2097,N_1777);
xnor U2332 (N_2332,N_1759,N_1771);
and U2333 (N_2333,N_1559,N_2145);
nand U2334 (N_2334,N_2174,N_1598);
or U2335 (N_2335,N_1831,N_1525);
nand U2336 (N_2336,N_2065,N_1911);
nor U2337 (N_2337,N_1810,N_2183);
or U2338 (N_2338,N_2163,N_1686);
xnor U2339 (N_2339,N_2081,N_2036);
and U2340 (N_2340,N_1550,N_2063);
nor U2341 (N_2341,N_1628,N_1983);
or U2342 (N_2342,N_1513,N_1866);
nand U2343 (N_2343,N_1511,N_2205);
xnor U2344 (N_2344,N_1835,N_1690);
xnor U2345 (N_2345,N_1530,N_1905);
nand U2346 (N_2346,N_2107,N_1830);
xnor U2347 (N_2347,N_1698,N_1660);
or U2348 (N_2348,N_2014,N_1664);
xnor U2349 (N_2349,N_1689,N_2138);
nand U2350 (N_2350,N_1638,N_1816);
xnor U2351 (N_2351,N_2223,N_1731);
nand U2352 (N_2352,N_1876,N_1597);
and U2353 (N_2353,N_1768,N_2216);
nor U2354 (N_2354,N_1755,N_1703);
and U2355 (N_2355,N_2072,N_1727);
xnor U2356 (N_2356,N_1877,N_1867);
xnor U2357 (N_2357,N_2058,N_1849);
xnor U2358 (N_2358,N_1812,N_1615);
nor U2359 (N_2359,N_1786,N_1568);
xnor U2360 (N_2360,N_2021,N_1620);
xnor U2361 (N_2361,N_1670,N_1987);
or U2362 (N_2362,N_1961,N_1804);
nor U2363 (N_2363,N_1691,N_1842);
or U2364 (N_2364,N_2245,N_1811);
nand U2365 (N_2365,N_1894,N_2214);
and U2366 (N_2366,N_2153,N_1790);
and U2367 (N_2367,N_2027,N_1534);
nand U2368 (N_2368,N_1838,N_2209);
nand U2369 (N_2369,N_2134,N_1589);
nor U2370 (N_2370,N_1552,N_1839);
nor U2371 (N_2371,N_1843,N_1900);
nand U2372 (N_2372,N_1588,N_1591);
and U2373 (N_2373,N_2229,N_2118);
nand U2374 (N_2374,N_1554,N_2055);
xor U2375 (N_2375,N_1780,N_1735);
nand U2376 (N_2376,N_2043,N_1827);
and U2377 (N_2377,N_1614,N_1979);
and U2378 (N_2378,N_2127,N_1868);
or U2379 (N_2379,N_1793,N_1817);
xor U2380 (N_2380,N_1613,N_1969);
nor U2381 (N_2381,N_1619,N_2182);
xor U2382 (N_2382,N_1542,N_1667);
and U2383 (N_2383,N_2011,N_1713);
or U2384 (N_2384,N_2213,N_1815);
or U2385 (N_2385,N_2104,N_1719);
or U2386 (N_2386,N_1500,N_1762);
xor U2387 (N_2387,N_1730,N_1607);
or U2388 (N_2388,N_1856,N_1947);
xor U2389 (N_2389,N_1912,N_1662);
and U2390 (N_2390,N_1996,N_1605);
and U2391 (N_2391,N_2026,N_2166);
nand U2392 (N_2392,N_2146,N_1743);
xnor U2393 (N_2393,N_2029,N_2233);
and U2394 (N_2394,N_2017,N_1705);
and U2395 (N_2395,N_1563,N_1693);
or U2396 (N_2396,N_2232,N_1518);
xor U2397 (N_2397,N_1540,N_1700);
nor U2398 (N_2398,N_2015,N_1716);
nor U2399 (N_2399,N_1846,N_2033);
xor U2400 (N_2400,N_1659,N_2211);
nand U2401 (N_2401,N_1889,N_1663);
xor U2402 (N_2402,N_2236,N_1834);
nand U2403 (N_2403,N_1908,N_1684);
or U2404 (N_2404,N_1636,N_1712);
or U2405 (N_2405,N_1860,N_1934);
nor U2406 (N_2406,N_1609,N_2093);
xor U2407 (N_2407,N_2076,N_1679);
nand U2408 (N_2408,N_2230,N_1756);
and U2409 (N_2409,N_1688,N_1910);
xnor U2410 (N_2410,N_1519,N_1968);
nand U2411 (N_2411,N_1896,N_1745);
nor U2412 (N_2412,N_1765,N_1580);
xor U2413 (N_2413,N_1682,N_1779);
nor U2414 (N_2414,N_2128,N_1573);
nor U2415 (N_2415,N_1618,N_1699);
or U2416 (N_2416,N_2240,N_1732);
nand U2417 (N_2417,N_1774,N_2160);
xor U2418 (N_2418,N_1875,N_1907);
nand U2419 (N_2419,N_1717,N_1649);
nand U2420 (N_2420,N_1959,N_1714);
and U2421 (N_2421,N_2003,N_2184);
and U2422 (N_2422,N_2125,N_1857);
xor U2423 (N_2423,N_1913,N_1909);
nand U2424 (N_2424,N_1593,N_2089);
nor U2425 (N_2425,N_1918,N_1977);
or U2426 (N_2426,N_1821,N_2059);
xnor U2427 (N_2427,N_1723,N_1854);
or U2428 (N_2428,N_1583,N_1904);
xnor U2429 (N_2429,N_2187,N_1886);
and U2430 (N_2430,N_2025,N_2220);
nand U2431 (N_2431,N_2147,N_1813);
and U2432 (N_2432,N_1772,N_1950);
nor U2433 (N_2433,N_2075,N_1631);
xnor U2434 (N_2434,N_1654,N_1972);
xor U2435 (N_2435,N_1763,N_1541);
and U2436 (N_2436,N_1888,N_1562);
and U2437 (N_2437,N_1668,N_2054);
or U2438 (N_2438,N_1635,N_1803);
xnor U2439 (N_2439,N_2168,N_2041);
nand U2440 (N_2440,N_2101,N_1874);
nor U2441 (N_2441,N_1845,N_1536);
or U2442 (N_2442,N_1951,N_1915);
nand U2443 (N_2443,N_2091,N_1938);
nand U2444 (N_2444,N_1800,N_2099);
or U2445 (N_2445,N_1880,N_1766);
xor U2446 (N_2446,N_2222,N_1883);
nor U2447 (N_2447,N_1529,N_1914);
nor U2448 (N_2448,N_2057,N_1676);
and U2449 (N_2449,N_1650,N_2108);
or U2450 (N_2450,N_1901,N_2066);
nand U2451 (N_2451,N_1930,N_1921);
nor U2452 (N_2452,N_1579,N_2115);
or U2453 (N_2453,N_1611,N_1505);
nand U2454 (N_2454,N_1558,N_2092);
and U2455 (N_2455,N_1787,N_1754);
or U2456 (N_2456,N_1577,N_2037);
or U2457 (N_2457,N_2188,N_1629);
or U2458 (N_2458,N_1967,N_1871);
nor U2459 (N_2459,N_1939,N_1781);
xor U2460 (N_2460,N_1535,N_2200);
xnor U2461 (N_2461,N_1678,N_2074);
or U2462 (N_2462,N_2207,N_2113);
and U2463 (N_2463,N_2035,N_1850);
or U2464 (N_2464,N_1958,N_1570);
or U2465 (N_2465,N_1680,N_2064);
xnor U2466 (N_2466,N_1507,N_1941);
nor U2467 (N_2467,N_1872,N_1643);
nor U2468 (N_2468,N_1704,N_1822);
xor U2469 (N_2469,N_2079,N_1851);
nand U2470 (N_2470,N_1966,N_1626);
and U2471 (N_2471,N_2045,N_2061);
xor U2472 (N_2472,N_1970,N_2106);
and U2473 (N_2473,N_2243,N_1954);
or U2474 (N_2474,N_1696,N_2228);
and U2475 (N_2475,N_1991,N_2049);
and U2476 (N_2476,N_1621,N_1571);
xor U2477 (N_2477,N_1504,N_1575);
nand U2478 (N_2478,N_1672,N_2028);
xor U2479 (N_2479,N_2050,N_1710);
or U2480 (N_2480,N_2227,N_1974);
and U2481 (N_2481,N_2149,N_1808);
nor U2482 (N_2482,N_1566,N_1533);
or U2483 (N_2483,N_2096,N_1788);
xnor U2484 (N_2484,N_1783,N_1879);
and U2485 (N_2485,N_1932,N_1840);
nand U2486 (N_2486,N_1557,N_2165);
xnor U2487 (N_2487,N_1610,N_1855);
or U2488 (N_2488,N_1612,N_1945);
xnor U2489 (N_2489,N_2192,N_2121);
nor U2490 (N_2490,N_2152,N_2070);
xnor U2491 (N_2491,N_2007,N_2085);
and U2492 (N_2492,N_2231,N_2126);
or U2493 (N_2493,N_1740,N_1863);
nand U2494 (N_2494,N_2024,N_2114);
and U2495 (N_2495,N_1778,N_1634);
xor U2496 (N_2496,N_2212,N_2040);
nand U2497 (N_2497,N_2151,N_2179);
nor U2498 (N_2498,N_2056,N_1720);
xor U2499 (N_2499,N_2084,N_1997);
nand U2500 (N_2500,N_1544,N_1707);
xnor U2501 (N_2501,N_1681,N_1881);
nor U2502 (N_2502,N_1858,N_1742);
or U2503 (N_2503,N_2181,N_1758);
xor U2504 (N_2504,N_1616,N_1935);
xnor U2505 (N_2505,N_1984,N_1677);
xor U2506 (N_2506,N_1514,N_1748);
nand U2507 (N_2507,N_2155,N_1728);
nand U2508 (N_2508,N_1606,N_2185);
and U2509 (N_2509,N_1887,N_2154);
or U2510 (N_2510,N_1722,N_1789);
nand U2511 (N_2511,N_1775,N_2103);
nor U2512 (N_2512,N_2217,N_2018);
xor U2513 (N_2513,N_1555,N_1920);
and U2514 (N_2514,N_1729,N_1675);
and U2515 (N_2515,N_2094,N_2234);
or U2516 (N_2516,N_1538,N_1873);
xor U2517 (N_2517,N_1671,N_1515);
xor U2518 (N_2518,N_1586,N_2122);
nand U2519 (N_2519,N_1683,N_1633);
nand U2520 (N_2520,N_2022,N_2241);
nor U2521 (N_2521,N_2067,N_2119);
nor U2522 (N_2522,N_2135,N_2137);
xor U2523 (N_2523,N_1556,N_1553);
nand U2524 (N_2524,N_1784,N_1761);
nor U2525 (N_2525,N_2102,N_1833);
nor U2526 (N_2526,N_1564,N_2062);
or U2527 (N_2527,N_1799,N_1940);
xnor U2528 (N_2528,N_1870,N_1647);
and U2529 (N_2529,N_1567,N_1899);
nand U2530 (N_2530,N_1825,N_1767);
or U2531 (N_2531,N_1847,N_1829);
nor U2532 (N_2532,N_1750,N_1641);
nand U2533 (N_2533,N_2224,N_1715);
nor U2534 (N_2534,N_1965,N_1844);
xnor U2535 (N_2535,N_1893,N_1551);
nor U2536 (N_2536,N_2156,N_1736);
xnor U2537 (N_2537,N_1746,N_1546);
nor U2538 (N_2538,N_2098,N_2086);
nor U2539 (N_2539,N_1510,N_1702);
and U2540 (N_2540,N_1990,N_1902);
nand U2541 (N_2541,N_1706,N_1642);
nand U2542 (N_2542,N_2196,N_1852);
or U2543 (N_2543,N_2124,N_1574);
and U2544 (N_2544,N_1865,N_1711);
or U2545 (N_2545,N_2117,N_1624);
and U2546 (N_2546,N_2178,N_2123);
or U2547 (N_2547,N_2148,N_1955);
xnor U2548 (N_2548,N_1640,N_1523);
and U2549 (N_2549,N_2249,N_2136);
and U2550 (N_2550,N_2201,N_2186);
and U2551 (N_2551,N_1818,N_1549);
and U2552 (N_2552,N_1581,N_2139);
and U2553 (N_2553,N_1917,N_2189);
xnor U2554 (N_2554,N_2157,N_1926);
nor U2555 (N_2555,N_1806,N_1595);
nor U2556 (N_2556,N_1753,N_1933);
nor U2557 (N_2557,N_1692,N_1992);
or U2558 (N_2558,N_2247,N_1995);
nor U2559 (N_2559,N_2053,N_2000);
nand U2560 (N_2560,N_2239,N_1749);
and U2561 (N_2561,N_1841,N_2190);
nand U2562 (N_2562,N_1962,N_1738);
xor U2563 (N_2563,N_1657,N_1592);
or U2564 (N_2564,N_1747,N_1837);
and U2565 (N_2565,N_2237,N_2069);
and U2566 (N_2566,N_1661,N_2202);
and U2567 (N_2567,N_1853,N_2044);
and U2568 (N_2568,N_2221,N_1897);
or U2569 (N_2569,N_2130,N_1798);
nor U2570 (N_2570,N_1545,N_1999);
nor U2571 (N_2571,N_1734,N_2144);
xor U2572 (N_2572,N_2208,N_1957);
and U2573 (N_2573,N_1862,N_1946);
nand U2574 (N_2574,N_1891,N_1674);
xor U2575 (N_2575,N_2034,N_2210);
nand U2576 (N_2576,N_2226,N_1928);
and U2577 (N_2577,N_1931,N_1578);
xor U2578 (N_2578,N_2194,N_1998);
and U2579 (N_2579,N_2180,N_1520);
nor U2580 (N_2580,N_2012,N_1637);
and U2581 (N_2581,N_2206,N_1517);
nor U2582 (N_2582,N_1826,N_1622);
nand U2583 (N_2583,N_2195,N_1848);
and U2584 (N_2584,N_2161,N_2001);
xnor U2585 (N_2585,N_2016,N_2090);
nand U2586 (N_2586,N_1501,N_1603);
or U2587 (N_2587,N_1539,N_2004);
nand U2588 (N_2588,N_1527,N_1741);
nor U2589 (N_2589,N_2048,N_1627);
xor U2590 (N_2590,N_1769,N_1895);
xnor U2591 (N_2591,N_2132,N_1890);
nand U2592 (N_2592,N_1828,N_2105);
or U2593 (N_2593,N_2023,N_1531);
nand U2594 (N_2594,N_2215,N_1725);
or U2595 (N_2595,N_1656,N_1721);
and U2596 (N_2596,N_1976,N_1522);
xnor U2597 (N_2597,N_1922,N_2082);
xnor U2598 (N_2598,N_1861,N_1824);
nor U2599 (N_2599,N_2159,N_1903);
or U2600 (N_2600,N_1859,N_1658);
and U2601 (N_2601,N_2219,N_1565);
or U2602 (N_2602,N_1516,N_1823);
and U2603 (N_2603,N_1601,N_1797);
or U2604 (N_2604,N_1701,N_1503);
and U2605 (N_2605,N_1669,N_1625);
or U2606 (N_2606,N_1718,N_1906);
and U2607 (N_2607,N_2047,N_2141);
nor U2608 (N_2608,N_1916,N_1560);
nand U2609 (N_2609,N_2199,N_1685);
or U2610 (N_2610,N_1695,N_1994);
or U2611 (N_2611,N_2116,N_1944);
xnor U2612 (N_2612,N_1986,N_1919);
xnor U2613 (N_2613,N_1651,N_2235);
xor U2614 (N_2614,N_1648,N_2031);
nor U2615 (N_2615,N_1989,N_1572);
nand U2616 (N_2616,N_1666,N_1963);
and U2617 (N_2617,N_1927,N_1524);
or U2618 (N_2618,N_1942,N_2142);
or U2619 (N_2619,N_1600,N_2150);
nor U2620 (N_2620,N_1885,N_1864);
or U2621 (N_2621,N_1537,N_2068);
xnor U2622 (N_2622,N_1561,N_2140);
xor U2623 (N_2623,N_1770,N_1726);
nand U2624 (N_2624,N_1898,N_1506);
and U2625 (N_2625,N_1837,N_1546);
nand U2626 (N_2626,N_2097,N_1732);
nor U2627 (N_2627,N_1873,N_1790);
and U2628 (N_2628,N_1788,N_1793);
xor U2629 (N_2629,N_1749,N_1606);
and U2630 (N_2630,N_1906,N_1526);
or U2631 (N_2631,N_2124,N_1558);
or U2632 (N_2632,N_1885,N_2030);
nor U2633 (N_2633,N_2249,N_1875);
nor U2634 (N_2634,N_2235,N_1825);
and U2635 (N_2635,N_1561,N_1799);
xnor U2636 (N_2636,N_1614,N_2086);
or U2637 (N_2637,N_2167,N_1644);
xnor U2638 (N_2638,N_1887,N_1734);
or U2639 (N_2639,N_1650,N_2183);
nor U2640 (N_2640,N_1841,N_2066);
nor U2641 (N_2641,N_1619,N_1572);
xnor U2642 (N_2642,N_2171,N_1822);
nor U2643 (N_2643,N_1607,N_1525);
or U2644 (N_2644,N_2218,N_2050);
xnor U2645 (N_2645,N_1943,N_2238);
or U2646 (N_2646,N_1961,N_2021);
and U2647 (N_2647,N_1796,N_1714);
nand U2648 (N_2648,N_1970,N_1866);
xnor U2649 (N_2649,N_1761,N_1999);
and U2650 (N_2650,N_2040,N_1641);
nor U2651 (N_2651,N_2117,N_1820);
and U2652 (N_2652,N_1846,N_1609);
nand U2653 (N_2653,N_2142,N_1509);
or U2654 (N_2654,N_2097,N_2133);
nor U2655 (N_2655,N_1844,N_1571);
and U2656 (N_2656,N_2008,N_1847);
nand U2657 (N_2657,N_1932,N_1868);
and U2658 (N_2658,N_2243,N_2208);
nor U2659 (N_2659,N_2193,N_1997);
nor U2660 (N_2660,N_1759,N_1743);
xor U2661 (N_2661,N_2172,N_1528);
nand U2662 (N_2662,N_1729,N_1578);
nor U2663 (N_2663,N_1951,N_2000);
or U2664 (N_2664,N_1981,N_1955);
xnor U2665 (N_2665,N_2007,N_1605);
nor U2666 (N_2666,N_2076,N_2082);
and U2667 (N_2667,N_2232,N_1621);
nor U2668 (N_2668,N_1965,N_1567);
and U2669 (N_2669,N_2035,N_1848);
xor U2670 (N_2670,N_1571,N_1977);
or U2671 (N_2671,N_1694,N_2116);
xor U2672 (N_2672,N_1762,N_1663);
or U2673 (N_2673,N_1641,N_2192);
or U2674 (N_2674,N_1825,N_2176);
nand U2675 (N_2675,N_1625,N_1972);
or U2676 (N_2676,N_1858,N_1611);
or U2677 (N_2677,N_1799,N_1676);
nand U2678 (N_2678,N_1916,N_2054);
and U2679 (N_2679,N_1882,N_1590);
xnor U2680 (N_2680,N_1610,N_1751);
and U2681 (N_2681,N_1878,N_1600);
nor U2682 (N_2682,N_1873,N_2245);
or U2683 (N_2683,N_2198,N_1527);
nor U2684 (N_2684,N_2181,N_2175);
or U2685 (N_2685,N_2008,N_1837);
and U2686 (N_2686,N_1586,N_1924);
or U2687 (N_2687,N_1895,N_2044);
and U2688 (N_2688,N_1657,N_1848);
and U2689 (N_2689,N_1745,N_2151);
and U2690 (N_2690,N_1930,N_1570);
nor U2691 (N_2691,N_1894,N_1645);
xor U2692 (N_2692,N_2194,N_1644);
or U2693 (N_2693,N_1997,N_1695);
xnor U2694 (N_2694,N_1752,N_1756);
xnor U2695 (N_2695,N_1768,N_1715);
and U2696 (N_2696,N_2196,N_1565);
xor U2697 (N_2697,N_1678,N_1629);
xnor U2698 (N_2698,N_1775,N_2185);
nor U2699 (N_2699,N_1738,N_1873);
and U2700 (N_2700,N_1667,N_2175);
nor U2701 (N_2701,N_1658,N_2155);
or U2702 (N_2702,N_1667,N_1775);
nor U2703 (N_2703,N_1714,N_2111);
or U2704 (N_2704,N_1985,N_2038);
xor U2705 (N_2705,N_1728,N_1770);
and U2706 (N_2706,N_2218,N_2076);
nor U2707 (N_2707,N_1797,N_1602);
nor U2708 (N_2708,N_2035,N_1747);
and U2709 (N_2709,N_2046,N_1876);
nand U2710 (N_2710,N_1890,N_2040);
and U2711 (N_2711,N_2202,N_1733);
or U2712 (N_2712,N_1524,N_1687);
xor U2713 (N_2713,N_2012,N_2175);
nand U2714 (N_2714,N_1651,N_1857);
or U2715 (N_2715,N_1748,N_1618);
xnor U2716 (N_2716,N_1689,N_1848);
nor U2717 (N_2717,N_2209,N_2009);
nand U2718 (N_2718,N_1809,N_2060);
nor U2719 (N_2719,N_1502,N_1729);
nor U2720 (N_2720,N_2036,N_2031);
nand U2721 (N_2721,N_1741,N_2126);
or U2722 (N_2722,N_1967,N_2097);
nor U2723 (N_2723,N_1823,N_1905);
nor U2724 (N_2724,N_1818,N_1569);
xnor U2725 (N_2725,N_1881,N_1850);
nand U2726 (N_2726,N_1992,N_1732);
and U2727 (N_2727,N_2224,N_1801);
xnor U2728 (N_2728,N_1959,N_1570);
nand U2729 (N_2729,N_1711,N_1912);
and U2730 (N_2730,N_1811,N_1663);
and U2731 (N_2731,N_1992,N_1904);
nor U2732 (N_2732,N_1915,N_2243);
or U2733 (N_2733,N_1607,N_1723);
or U2734 (N_2734,N_1666,N_1894);
xnor U2735 (N_2735,N_1698,N_1816);
xor U2736 (N_2736,N_1972,N_1505);
or U2737 (N_2737,N_2108,N_1605);
xnor U2738 (N_2738,N_1567,N_1856);
and U2739 (N_2739,N_2003,N_1674);
nor U2740 (N_2740,N_2228,N_1859);
or U2741 (N_2741,N_2105,N_2238);
xor U2742 (N_2742,N_1896,N_1767);
xor U2743 (N_2743,N_2224,N_1667);
nand U2744 (N_2744,N_1824,N_1699);
and U2745 (N_2745,N_1594,N_2178);
nand U2746 (N_2746,N_1984,N_1517);
nand U2747 (N_2747,N_1755,N_2222);
and U2748 (N_2748,N_2192,N_2076);
or U2749 (N_2749,N_1990,N_1631);
nand U2750 (N_2750,N_1992,N_1856);
nor U2751 (N_2751,N_1603,N_2122);
or U2752 (N_2752,N_1884,N_2136);
nand U2753 (N_2753,N_1559,N_1966);
nand U2754 (N_2754,N_1672,N_1817);
or U2755 (N_2755,N_1596,N_1978);
or U2756 (N_2756,N_1688,N_2225);
xor U2757 (N_2757,N_2220,N_2138);
or U2758 (N_2758,N_1636,N_1695);
or U2759 (N_2759,N_1967,N_1842);
nor U2760 (N_2760,N_2075,N_2161);
nand U2761 (N_2761,N_1782,N_1626);
nor U2762 (N_2762,N_1638,N_1937);
xnor U2763 (N_2763,N_2039,N_1896);
xor U2764 (N_2764,N_1679,N_1823);
xnor U2765 (N_2765,N_1728,N_2121);
or U2766 (N_2766,N_1509,N_1879);
or U2767 (N_2767,N_2042,N_1986);
xnor U2768 (N_2768,N_1884,N_2218);
or U2769 (N_2769,N_2215,N_1827);
or U2770 (N_2770,N_2199,N_1721);
nand U2771 (N_2771,N_2057,N_2215);
or U2772 (N_2772,N_2039,N_2248);
or U2773 (N_2773,N_1523,N_1934);
and U2774 (N_2774,N_1632,N_1855);
and U2775 (N_2775,N_1825,N_1501);
nand U2776 (N_2776,N_1911,N_1896);
xor U2777 (N_2777,N_2022,N_2017);
xnor U2778 (N_2778,N_1730,N_1905);
nand U2779 (N_2779,N_1688,N_2152);
and U2780 (N_2780,N_1912,N_1918);
nand U2781 (N_2781,N_1935,N_1533);
and U2782 (N_2782,N_2085,N_1778);
or U2783 (N_2783,N_1612,N_1884);
or U2784 (N_2784,N_1615,N_2047);
or U2785 (N_2785,N_2193,N_1864);
and U2786 (N_2786,N_1594,N_1869);
nor U2787 (N_2787,N_1907,N_2007);
and U2788 (N_2788,N_1698,N_1962);
or U2789 (N_2789,N_1972,N_1727);
xnor U2790 (N_2790,N_2144,N_1622);
nor U2791 (N_2791,N_1853,N_2030);
or U2792 (N_2792,N_1795,N_1919);
and U2793 (N_2793,N_2206,N_2093);
xor U2794 (N_2794,N_1571,N_2075);
nand U2795 (N_2795,N_1883,N_1513);
nor U2796 (N_2796,N_2063,N_2069);
nand U2797 (N_2797,N_1907,N_1656);
and U2798 (N_2798,N_2244,N_1911);
and U2799 (N_2799,N_1622,N_1920);
nor U2800 (N_2800,N_1843,N_1726);
nand U2801 (N_2801,N_1743,N_2163);
and U2802 (N_2802,N_1922,N_2044);
and U2803 (N_2803,N_1546,N_2030);
nor U2804 (N_2804,N_1844,N_2123);
or U2805 (N_2805,N_1646,N_2189);
xnor U2806 (N_2806,N_1927,N_2002);
and U2807 (N_2807,N_1696,N_2131);
or U2808 (N_2808,N_2152,N_1961);
or U2809 (N_2809,N_1905,N_2118);
xor U2810 (N_2810,N_1792,N_1534);
nand U2811 (N_2811,N_1677,N_1588);
nor U2812 (N_2812,N_2142,N_1988);
and U2813 (N_2813,N_2046,N_1936);
nor U2814 (N_2814,N_2013,N_2008);
xnor U2815 (N_2815,N_1868,N_2090);
nand U2816 (N_2816,N_1835,N_1575);
nor U2817 (N_2817,N_1828,N_2096);
or U2818 (N_2818,N_1863,N_1916);
nor U2819 (N_2819,N_1944,N_2167);
nor U2820 (N_2820,N_1602,N_1752);
nand U2821 (N_2821,N_1522,N_1782);
and U2822 (N_2822,N_1894,N_1973);
nor U2823 (N_2823,N_1912,N_1962);
xnor U2824 (N_2824,N_1629,N_2246);
or U2825 (N_2825,N_1787,N_1706);
and U2826 (N_2826,N_1816,N_2075);
or U2827 (N_2827,N_2150,N_2072);
nand U2828 (N_2828,N_2193,N_1819);
nor U2829 (N_2829,N_1747,N_2016);
xnor U2830 (N_2830,N_1856,N_2025);
and U2831 (N_2831,N_1890,N_1559);
xor U2832 (N_2832,N_1598,N_2012);
and U2833 (N_2833,N_1594,N_1880);
nand U2834 (N_2834,N_1950,N_2003);
or U2835 (N_2835,N_2081,N_1980);
or U2836 (N_2836,N_2019,N_1804);
nand U2837 (N_2837,N_2101,N_2070);
and U2838 (N_2838,N_2223,N_1918);
nor U2839 (N_2839,N_2052,N_1651);
xor U2840 (N_2840,N_1574,N_1619);
xor U2841 (N_2841,N_1602,N_1596);
nor U2842 (N_2842,N_1985,N_1831);
and U2843 (N_2843,N_1973,N_1736);
nor U2844 (N_2844,N_1768,N_1782);
nand U2845 (N_2845,N_2002,N_1825);
or U2846 (N_2846,N_2092,N_1952);
xnor U2847 (N_2847,N_1551,N_2193);
xor U2848 (N_2848,N_2092,N_1540);
nor U2849 (N_2849,N_2239,N_1726);
or U2850 (N_2850,N_1751,N_1721);
or U2851 (N_2851,N_1561,N_1997);
and U2852 (N_2852,N_1602,N_1871);
or U2853 (N_2853,N_1513,N_1803);
xor U2854 (N_2854,N_1935,N_1785);
nor U2855 (N_2855,N_1848,N_1959);
xor U2856 (N_2856,N_1650,N_2037);
and U2857 (N_2857,N_1856,N_2099);
or U2858 (N_2858,N_1590,N_1576);
nor U2859 (N_2859,N_1842,N_1738);
xor U2860 (N_2860,N_2026,N_1729);
or U2861 (N_2861,N_2220,N_1637);
xor U2862 (N_2862,N_2100,N_1867);
xnor U2863 (N_2863,N_2013,N_1685);
xor U2864 (N_2864,N_1626,N_1722);
nand U2865 (N_2865,N_1579,N_1782);
and U2866 (N_2866,N_2199,N_2192);
or U2867 (N_2867,N_2236,N_2136);
nand U2868 (N_2868,N_1632,N_1886);
or U2869 (N_2869,N_1802,N_2187);
nand U2870 (N_2870,N_1724,N_1950);
nor U2871 (N_2871,N_2211,N_1694);
nor U2872 (N_2872,N_2174,N_1834);
or U2873 (N_2873,N_1634,N_1525);
xnor U2874 (N_2874,N_1680,N_2103);
or U2875 (N_2875,N_1979,N_1870);
and U2876 (N_2876,N_1874,N_1539);
xor U2877 (N_2877,N_1947,N_1913);
xnor U2878 (N_2878,N_1696,N_1980);
and U2879 (N_2879,N_1852,N_2052);
and U2880 (N_2880,N_2201,N_1616);
xnor U2881 (N_2881,N_2125,N_1958);
nor U2882 (N_2882,N_1873,N_2249);
xor U2883 (N_2883,N_2046,N_1972);
or U2884 (N_2884,N_2243,N_1839);
nor U2885 (N_2885,N_2198,N_1944);
and U2886 (N_2886,N_1567,N_2015);
xor U2887 (N_2887,N_2016,N_1742);
or U2888 (N_2888,N_1930,N_2085);
and U2889 (N_2889,N_1769,N_1534);
and U2890 (N_2890,N_2222,N_1721);
nand U2891 (N_2891,N_1570,N_1836);
nor U2892 (N_2892,N_2058,N_2086);
xnor U2893 (N_2893,N_1814,N_1574);
or U2894 (N_2894,N_2237,N_2118);
nor U2895 (N_2895,N_1818,N_1766);
and U2896 (N_2896,N_1683,N_1687);
nand U2897 (N_2897,N_2154,N_1971);
nand U2898 (N_2898,N_1890,N_1961);
nor U2899 (N_2899,N_2118,N_1865);
xnor U2900 (N_2900,N_2245,N_1531);
nand U2901 (N_2901,N_2173,N_2069);
xnor U2902 (N_2902,N_1685,N_2155);
nand U2903 (N_2903,N_1873,N_2098);
or U2904 (N_2904,N_1672,N_2010);
nand U2905 (N_2905,N_1942,N_1606);
or U2906 (N_2906,N_1756,N_1873);
xor U2907 (N_2907,N_2049,N_1736);
nor U2908 (N_2908,N_1965,N_1565);
nor U2909 (N_2909,N_1624,N_1748);
and U2910 (N_2910,N_1920,N_1650);
xnor U2911 (N_2911,N_1581,N_1612);
and U2912 (N_2912,N_2134,N_2181);
nand U2913 (N_2913,N_1784,N_2054);
and U2914 (N_2914,N_1856,N_1597);
or U2915 (N_2915,N_1558,N_1792);
nand U2916 (N_2916,N_1605,N_2171);
or U2917 (N_2917,N_2088,N_1814);
xor U2918 (N_2918,N_2060,N_1574);
and U2919 (N_2919,N_2137,N_1828);
xnor U2920 (N_2920,N_2068,N_1722);
xor U2921 (N_2921,N_1624,N_1962);
nor U2922 (N_2922,N_1674,N_1515);
or U2923 (N_2923,N_1640,N_1691);
nor U2924 (N_2924,N_1560,N_2126);
or U2925 (N_2925,N_2131,N_1787);
nand U2926 (N_2926,N_2044,N_1675);
nor U2927 (N_2927,N_1813,N_2165);
nand U2928 (N_2928,N_1748,N_1553);
or U2929 (N_2929,N_1535,N_2223);
nor U2930 (N_2930,N_2201,N_1779);
or U2931 (N_2931,N_1663,N_2146);
or U2932 (N_2932,N_1540,N_1739);
nor U2933 (N_2933,N_1617,N_1886);
xnor U2934 (N_2934,N_2167,N_1725);
nand U2935 (N_2935,N_1686,N_1835);
nor U2936 (N_2936,N_1769,N_1923);
or U2937 (N_2937,N_2011,N_1537);
nor U2938 (N_2938,N_1980,N_1703);
or U2939 (N_2939,N_1638,N_1682);
or U2940 (N_2940,N_1856,N_1603);
or U2941 (N_2941,N_1678,N_1799);
and U2942 (N_2942,N_1603,N_1662);
and U2943 (N_2943,N_2006,N_1780);
and U2944 (N_2944,N_1533,N_1629);
nand U2945 (N_2945,N_1669,N_1685);
nand U2946 (N_2946,N_1961,N_1915);
and U2947 (N_2947,N_1732,N_2105);
xor U2948 (N_2948,N_1619,N_1976);
and U2949 (N_2949,N_1931,N_2190);
nor U2950 (N_2950,N_1757,N_1790);
nand U2951 (N_2951,N_2153,N_1954);
xor U2952 (N_2952,N_1670,N_1920);
nor U2953 (N_2953,N_1905,N_1623);
or U2954 (N_2954,N_1671,N_2126);
nand U2955 (N_2955,N_2070,N_1768);
nand U2956 (N_2956,N_2012,N_2232);
or U2957 (N_2957,N_1794,N_1957);
nor U2958 (N_2958,N_1731,N_1810);
nand U2959 (N_2959,N_1728,N_1741);
and U2960 (N_2960,N_1863,N_1959);
xnor U2961 (N_2961,N_1834,N_1761);
nor U2962 (N_2962,N_1524,N_1688);
nor U2963 (N_2963,N_1788,N_1762);
and U2964 (N_2964,N_1975,N_1567);
and U2965 (N_2965,N_1999,N_1882);
xnor U2966 (N_2966,N_1930,N_1540);
nor U2967 (N_2967,N_2097,N_2184);
nor U2968 (N_2968,N_2132,N_2092);
nor U2969 (N_2969,N_1650,N_2017);
or U2970 (N_2970,N_1942,N_1599);
xnor U2971 (N_2971,N_2210,N_1895);
and U2972 (N_2972,N_1680,N_1646);
nand U2973 (N_2973,N_1648,N_1879);
nand U2974 (N_2974,N_1597,N_1762);
nand U2975 (N_2975,N_1679,N_1582);
nor U2976 (N_2976,N_1549,N_1775);
nand U2977 (N_2977,N_1592,N_1724);
or U2978 (N_2978,N_1881,N_2109);
xnor U2979 (N_2979,N_2166,N_1515);
and U2980 (N_2980,N_1805,N_1815);
nor U2981 (N_2981,N_1594,N_1740);
xor U2982 (N_2982,N_2220,N_1683);
and U2983 (N_2983,N_2151,N_1706);
nor U2984 (N_2984,N_1876,N_2055);
nor U2985 (N_2985,N_2158,N_1609);
and U2986 (N_2986,N_1613,N_1546);
and U2987 (N_2987,N_1814,N_2008);
xor U2988 (N_2988,N_2020,N_1722);
or U2989 (N_2989,N_1567,N_1712);
nand U2990 (N_2990,N_1868,N_2130);
xnor U2991 (N_2991,N_1708,N_1662);
nand U2992 (N_2992,N_1621,N_1725);
or U2993 (N_2993,N_1976,N_1610);
nand U2994 (N_2994,N_2113,N_2059);
or U2995 (N_2995,N_1665,N_1610);
xor U2996 (N_2996,N_1515,N_1550);
nor U2997 (N_2997,N_1507,N_1650);
xor U2998 (N_2998,N_2200,N_1530);
nand U2999 (N_2999,N_1751,N_1656);
xor U3000 (N_3000,N_2605,N_2835);
nand U3001 (N_3001,N_2774,N_2617);
and U3002 (N_3002,N_2874,N_2913);
nand U3003 (N_3003,N_2902,N_2946);
nor U3004 (N_3004,N_2526,N_2776);
and U3005 (N_3005,N_2333,N_2330);
nand U3006 (N_3006,N_2788,N_2505);
and U3007 (N_3007,N_2613,N_2861);
nor U3008 (N_3008,N_2346,N_2479);
or U3009 (N_3009,N_2745,N_2489);
xor U3010 (N_3010,N_2881,N_2614);
or U3011 (N_3011,N_2537,N_2490);
or U3012 (N_3012,N_2910,N_2987);
and U3013 (N_3013,N_2596,N_2288);
xor U3014 (N_3014,N_2378,N_2264);
or U3015 (N_3015,N_2369,N_2901);
nor U3016 (N_3016,N_2293,N_2963);
nand U3017 (N_3017,N_2339,N_2252);
nand U3018 (N_3018,N_2680,N_2591);
nand U3019 (N_3019,N_2967,N_2522);
nor U3020 (N_3020,N_2924,N_2801);
nor U3021 (N_3021,N_2532,N_2803);
nor U3022 (N_3022,N_2312,N_2544);
and U3023 (N_3023,N_2748,N_2373);
nor U3024 (N_3024,N_2687,N_2736);
nand U3025 (N_3025,N_2494,N_2764);
nand U3026 (N_3026,N_2959,N_2599);
nor U3027 (N_3027,N_2447,N_2802);
xnor U3028 (N_3028,N_2253,N_2672);
xor U3029 (N_3029,N_2779,N_2506);
nand U3030 (N_3030,N_2844,N_2593);
xor U3031 (N_3031,N_2903,N_2527);
xnor U3032 (N_3032,N_2615,N_2649);
or U3033 (N_3033,N_2563,N_2931);
xor U3034 (N_3034,N_2568,N_2744);
xnor U3035 (N_3035,N_2360,N_2864);
and U3036 (N_3036,N_2463,N_2488);
or U3037 (N_3037,N_2289,N_2538);
and U3038 (N_3038,N_2906,N_2274);
nand U3039 (N_3039,N_2842,N_2768);
nand U3040 (N_3040,N_2318,N_2921);
xor U3041 (N_3041,N_2677,N_2493);
nand U3042 (N_3042,N_2958,N_2955);
nand U3043 (N_3043,N_2714,N_2944);
xor U3044 (N_3044,N_2763,N_2951);
nand U3045 (N_3045,N_2894,N_2860);
and U3046 (N_3046,N_2278,N_2357);
nand U3047 (N_3047,N_2974,N_2509);
and U3048 (N_3048,N_2303,N_2833);
nor U3049 (N_3049,N_2856,N_2740);
or U3050 (N_3050,N_2656,N_2707);
xnor U3051 (N_3051,N_2475,N_2790);
nand U3052 (N_3052,N_2683,N_2679);
or U3053 (N_3053,N_2941,N_2912);
nand U3054 (N_3054,N_2336,N_2923);
nor U3055 (N_3055,N_2272,N_2735);
and U3056 (N_3056,N_2807,N_2355);
xor U3057 (N_3057,N_2363,N_2420);
nand U3058 (N_3058,N_2328,N_2747);
xor U3059 (N_3059,N_2632,N_2811);
nor U3060 (N_3060,N_2405,N_2908);
xor U3061 (N_3061,N_2616,N_2705);
or U3062 (N_3062,N_2846,N_2364);
xor U3063 (N_3063,N_2478,N_2695);
or U3064 (N_3064,N_2928,N_2536);
xnor U3065 (N_3065,N_2503,N_2387);
and U3066 (N_3066,N_2316,N_2643);
nand U3067 (N_3067,N_2868,N_2356);
nor U3068 (N_3068,N_2467,N_2674);
xor U3069 (N_3069,N_2852,N_2650);
nand U3070 (N_3070,N_2323,N_2759);
and U3071 (N_3071,N_2853,N_2300);
nor U3072 (N_3072,N_2741,N_2935);
and U3073 (N_3073,N_2892,N_2354);
or U3074 (N_3074,N_2460,N_2628);
and U3075 (N_3075,N_2808,N_2480);
and U3076 (N_3076,N_2663,N_2399);
or U3077 (N_3077,N_2879,N_2326);
xor U3078 (N_3078,N_2895,N_2893);
nor U3079 (N_3079,N_2573,N_2444);
xnor U3080 (N_3080,N_2728,N_2971);
nor U3081 (N_3081,N_2546,N_2381);
or U3082 (N_3082,N_2507,N_2641);
and U3083 (N_3083,N_2584,N_2277);
nand U3084 (N_3084,N_2611,N_2535);
nand U3085 (N_3085,N_2800,N_2307);
nor U3086 (N_3086,N_2896,N_2849);
or U3087 (N_3087,N_2380,N_2256);
xnor U3088 (N_3088,N_2730,N_2750);
nand U3089 (N_3089,N_2789,N_2675);
or U3090 (N_3090,N_2766,N_2524);
xnor U3091 (N_3091,N_2290,N_2652);
nor U3092 (N_3092,N_2784,N_2697);
or U3093 (N_3093,N_2657,N_2442);
xnor U3094 (N_3094,N_2993,N_2285);
xor U3095 (N_3095,N_2454,N_2986);
nor U3096 (N_3096,N_2588,N_2783);
nor U3097 (N_3097,N_2309,N_2671);
and U3098 (N_3098,N_2753,N_2592);
nand U3099 (N_3099,N_2345,N_2712);
nor U3100 (N_3100,N_2491,N_2623);
nor U3101 (N_3101,N_2999,N_2761);
nor U3102 (N_3102,N_2638,N_2737);
xor U3103 (N_3103,N_2556,N_2976);
nor U3104 (N_3104,N_2580,N_2998);
nand U3105 (N_3105,N_2972,N_2438);
nor U3106 (N_3106,N_2443,N_2909);
nand U3107 (N_3107,N_2791,N_2820);
nand U3108 (N_3108,N_2283,N_2450);
nand U3109 (N_3109,N_2795,N_2659);
and U3110 (N_3110,N_2514,N_2678);
or U3111 (N_3111,N_2933,N_2839);
and U3112 (N_3112,N_2368,N_2934);
xnor U3113 (N_3113,N_2559,N_2587);
nor U3114 (N_3114,N_2704,N_2540);
and U3115 (N_3115,N_2973,N_2324);
and U3116 (N_3116,N_2406,N_2516);
xor U3117 (N_3117,N_2754,N_2732);
nand U3118 (N_3118,N_2694,N_2601);
xnor U3119 (N_3119,N_2942,N_2266);
nor U3120 (N_3120,N_2888,N_2670);
xnor U3121 (N_3121,N_2648,N_2301);
nor U3122 (N_3122,N_2334,N_2780);
or U3123 (N_3123,N_2470,N_2304);
xnor U3124 (N_3124,N_2622,N_2270);
nand U3125 (N_3125,N_2412,N_2669);
nor U3126 (N_3126,N_2257,N_2583);
and U3127 (N_3127,N_2499,N_2521);
or U3128 (N_3128,N_2558,N_2667);
nor U3129 (N_3129,N_2407,N_2726);
and U3130 (N_3130,N_2620,N_2402);
nand U3131 (N_3131,N_2448,N_2676);
or U3132 (N_3132,N_2701,N_2269);
and U3133 (N_3133,N_2459,N_2417);
nand U3134 (N_3134,N_2840,N_2518);
and U3135 (N_3135,N_2594,N_2729);
nor U3136 (N_3136,N_2792,N_2329);
xnor U3137 (N_3137,N_2566,N_2390);
nand U3138 (N_3138,N_2654,N_2557);
and U3139 (N_3139,N_2818,N_2922);
xor U3140 (N_3140,N_2477,N_2863);
and U3141 (N_3141,N_2651,N_2775);
nor U3142 (N_3142,N_2292,N_2600);
nor U3143 (N_3143,N_2569,N_2350);
nand U3144 (N_3144,N_2889,N_2688);
nand U3145 (N_3145,N_2857,N_2843);
and U3146 (N_3146,N_2372,N_2719);
and U3147 (N_3147,N_2919,N_2437);
nand U3148 (N_3148,N_2435,N_2481);
xor U3149 (N_3149,N_2658,N_2949);
or U3150 (N_3150,N_2286,N_2498);
nor U3151 (N_3151,N_2989,N_2630);
and U3152 (N_3152,N_2932,N_2692);
nand U3153 (N_3153,N_2547,N_2691);
and U3154 (N_3154,N_2310,N_2255);
xnor U3155 (N_3155,N_2751,N_2513);
xor U3156 (N_3156,N_2543,N_2890);
or U3157 (N_3157,N_2746,N_2867);
or U3158 (N_3158,N_2423,N_2383);
nand U3159 (N_3159,N_2268,N_2602);
xnor U3160 (N_3160,N_2830,N_2858);
xnor U3161 (N_3161,N_2436,N_2539);
and U3162 (N_3162,N_2351,N_2900);
and U3163 (N_3163,N_2512,N_2635);
nor U3164 (N_3164,N_2567,N_2552);
xor U3165 (N_3165,N_2782,N_2468);
nor U3166 (N_3166,N_2386,N_2296);
nand U3167 (N_3167,N_2608,N_2647);
nand U3168 (N_3168,N_2408,N_2709);
nand U3169 (N_3169,N_2353,N_2796);
xnor U3170 (N_3170,N_2703,N_2492);
xor U3171 (N_3171,N_2637,N_2664);
and U3172 (N_3172,N_2885,N_2957);
nor U3173 (N_3173,N_2717,N_2646);
or U3174 (N_3174,N_2434,N_2574);
nand U3175 (N_3175,N_2461,N_2545);
or U3176 (N_3176,N_2342,N_2331);
and U3177 (N_3177,N_2898,N_2904);
or U3178 (N_3178,N_2575,N_2716);
xor U3179 (N_3179,N_2873,N_2816);
or U3180 (N_3180,N_2361,N_2700);
nor U3181 (N_3181,N_2529,N_2422);
and U3182 (N_3182,N_2377,N_2362);
and U3183 (N_3183,N_2771,N_2549);
nor U3184 (N_3184,N_2590,N_2916);
nand U3185 (N_3185,N_2917,N_2606);
or U3186 (N_3186,N_2634,N_2837);
xor U3187 (N_3187,N_2721,N_2404);
nand U3188 (N_3188,N_2338,N_2483);
and U3189 (N_3189,N_2720,N_2562);
and U3190 (N_3190,N_2996,N_2340);
or U3191 (N_3191,N_2560,N_2668);
xor U3192 (N_3192,N_2317,N_2582);
nand U3193 (N_3193,N_2565,N_2884);
and U3194 (N_3194,N_2772,N_2409);
and U3195 (N_3195,N_2666,N_2827);
or U3196 (N_3196,N_2778,N_2961);
and U3197 (N_3197,N_2850,N_2937);
nor U3198 (N_3198,N_2804,N_2742);
or U3199 (N_3199,N_2433,N_2854);
xnor U3200 (N_3200,N_2397,N_2936);
nand U3201 (N_3201,N_2887,N_2851);
and U3202 (N_3202,N_2533,N_2451);
and U3203 (N_3203,N_2530,N_2806);
xnor U3204 (N_3204,N_2943,N_2733);
nor U3205 (N_3205,N_2940,N_2673);
or U3206 (N_3206,N_2250,N_2899);
nor U3207 (N_3207,N_2597,N_2970);
nand U3208 (N_3208,N_2400,N_2585);
xnor U3209 (N_3209,N_2263,N_2880);
xor U3210 (N_3210,N_2395,N_2561);
nor U3211 (N_3211,N_2994,N_2872);
xor U3212 (N_3212,N_2464,N_2262);
nor U3213 (N_3213,N_2862,N_2706);
and U3214 (N_3214,N_2276,N_2370);
nor U3215 (N_3215,N_2500,N_2251);
nor U3216 (N_3216,N_2612,N_2822);
or U3217 (N_3217,N_2525,N_2541);
and U3218 (N_3218,N_2410,N_2519);
nand U3219 (N_3219,N_2945,N_2308);
and U3220 (N_3220,N_2265,N_2770);
nor U3221 (N_3221,N_2685,N_2604);
xnor U3222 (N_3222,N_2847,N_2347);
and U3223 (N_3223,N_2702,N_2416);
or U3224 (N_3224,N_2950,N_2511);
xnor U3225 (N_3225,N_2496,N_2631);
xnor U3226 (N_3226,N_2848,N_2396);
or U3227 (N_3227,N_2392,N_2607);
xnor U3228 (N_3228,N_2621,N_2767);
or U3229 (N_3229,N_2952,N_2618);
or U3230 (N_3230,N_2603,N_2458);
and U3231 (N_3231,N_2388,N_2343);
xor U3232 (N_3232,N_2432,N_2413);
and U3233 (N_3233,N_2828,N_2639);
nor U3234 (N_3234,N_2995,N_2831);
or U3235 (N_3235,N_2403,N_2462);
nand U3236 (N_3236,N_2515,N_2765);
or U3237 (N_3237,N_2930,N_2321);
xnor U3238 (N_3238,N_2665,N_2897);
xnor U3239 (N_3239,N_2258,N_2948);
xnor U3240 (N_3240,N_2758,N_2698);
nor U3241 (N_3241,N_2629,N_2445);
nand U3242 (N_3242,N_2832,N_2905);
nor U3243 (N_3243,N_2332,N_2627);
and U3244 (N_3244,N_2287,N_2411);
xor U3245 (N_3245,N_2734,N_2297);
nor U3246 (N_3246,N_2548,N_2760);
xor U3247 (N_3247,N_2325,N_2918);
and U3248 (N_3248,N_2426,N_2619);
xnor U3249 (N_3249,N_2927,N_2965);
or U3250 (N_3250,N_2877,N_2870);
and U3251 (N_3251,N_2385,N_2960);
nor U3252 (N_3252,N_2715,N_2394);
xor U3253 (N_3253,N_2311,N_2598);
and U3254 (N_3254,N_2625,N_2352);
or U3255 (N_3255,N_2813,N_2586);
or U3256 (N_3256,N_2953,N_2711);
xor U3257 (N_3257,N_2465,N_2466);
and U3258 (N_3258,N_2826,N_2661);
nor U3259 (N_3259,N_2430,N_2990);
and U3260 (N_3260,N_2534,N_2421);
and U3261 (N_3261,N_2911,N_2299);
xnor U3262 (N_3262,N_2988,N_2280);
nor U3263 (N_3263,N_2550,N_2294);
xor U3264 (N_3264,N_2424,N_2376);
and U3265 (N_3265,N_2710,N_2439);
or U3266 (N_3266,N_2633,N_2891);
nor U3267 (N_3267,N_2992,N_2699);
nor U3268 (N_3268,N_2261,N_2834);
nor U3269 (N_3269,N_2393,N_2836);
xor U3270 (N_3270,N_2259,N_2367);
nand U3271 (N_3271,N_2805,N_2981);
nand U3272 (N_3272,N_2418,N_2926);
xnor U3273 (N_3273,N_2344,N_2731);
nor U3274 (N_3274,N_2284,N_2624);
xor U3275 (N_3275,N_2907,N_2348);
and U3276 (N_3276,N_2577,N_2713);
nand U3277 (N_3277,N_2781,N_2626);
nand U3278 (N_3278,N_2281,N_2684);
nand U3279 (N_3279,N_2374,N_2845);
nor U3280 (N_3280,N_2642,N_2982);
and U3281 (N_3281,N_2482,N_2456);
nor U3282 (N_3282,N_2743,N_2508);
and U3283 (N_3283,N_2517,N_2689);
xor U3284 (N_3284,N_2978,N_2371);
or U3285 (N_3285,N_2382,N_2449);
xnor U3286 (N_3286,N_2474,N_2819);
nor U3287 (N_3287,N_2313,N_2756);
nand U3288 (N_3288,N_2869,N_2991);
or U3289 (N_3289,N_2389,N_2824);
and U3290 (N_3290,N_2419,N_2497);
nor U3291 (N_3291,N_2708,N_2431);
nor U3292 (N_3292,N_2554,N_2319);
nand U3293 (N_3293,N_2579,N_2564);
and U3294 (N_3294,N_2589,N_2302);
and U3295 (N_3295,N_2384,N_2799);
nor U3296 (N_3296,N_2876,N_2391);
nor U3297 (N_3297,N_2473,N_2809);
nand U3298 (N_3298,N_2886,N_2502);
or U3299 (N_3299,N_2686,N_2472);
nor U3300 (N_3300,N_2815,N_2555);
nor U3301 (N_3301,N_2271,N_2757);
or U3302 (N_3302,N_2578,N_2956);
xor U3303 (N_3303,N_2855,N_2925);
xnor U3304 (N_3304,N_2440,N_2337);
nand U3305 (N_3305,N_2315,N_2980);
and U3306 (N_3306,N_2314,N_2798);
or U3307 (N_3307,N_2495,N_2415);
xor U3308 (N_3308,N_2504,N_2859);
or U3309 (N_3309,N_2682,N_2279);
or U3310 (N_3310,N_2428,N_2485);
and U3311 (N_3311,N_2531,N_2722);
nand U3312 (N_3312,N_2787,N_2915);
and U3313 (N_3313,N_2752,N_2662);
and U3314 (N_3314,N_2929,N_2871);
nand U3315 (N_3315,N_2609,N_2254);
and U3316 (N_3316,N_2823,N_2551);
xnor U3317 (N_3317,N_2398,N_2341);
or U3318 (N_3318,N_2769,N_2984);
nand U3319 (N_3319,N_2817,N_2914);
and U3320 (N_3320,N_2882,N_2777);
nor U3321 (N_3321,N_2520,N_2794);
and U3322 (N_3322,N_2825,N_2365);
and U3323 (N_3323,N_2968,N_2938);
or U3324 (N_3324,N_2282,N_2866);
nor U3325 (N_3325,N_2797,N_2829);
nand U3326 (N_3326,N_2487,N_2636);
or U3327 (N_3327,N_2696,N_2453);
or U3328 (N_3328,N_2298,N_2785);
and U3329 (N_3329,N_2681,N_2755);
nor U3330 (N_3330,N_2939,N_2793);
xor U3331 (N_3331,N_2429,N_2762);
nand U3332 (N_3332,N_2366,N_2875);
nor U3333 (N_3333,N_2523,N_2570);
nand U3334 (N_3334,N_2510,N_2486);
xnor U3335 (N_3335,N_2690,N_2427);
and U3336 (N_3336,N_2275,N_2966);
and U3337 (N_3337,N_2977,N_2727);
nor U3338 (N_3338,N_2878,N_2572);
xnor U3339 (N_3339,N_2738,N_2645);
nand U3340 (N_3340,N_2997,N_2724);
nand U3341 (N_3341,N_2267,N_2484);
or U3342 (N_3342,N_2810,N_2528);
nor U3343 (N_3343,N_2610,N_2644);
nor U3344 (N_3344,N_2441,N_2457);
or U3345 (N_3345,N_2414,N_2471);
or U3346 (N_3346,N_2723,N_2865);
or U3347 (N_3347,N_2306,N_2786);
nor U3348 (N_3348,N_2947,N_2979);
xor U3349 (N_3349,N_2446,N_2260);
or U3350 (N_3350,N_2542,N_2273);
nor U3351 (N_3351,N_2812,N_2571);
and U3352 (N_3352,N_2920,N_2655);
and U3353 (N_3353,N_2814,N_2335);
nor U3354 (N_3354,N_2349,N_2379);
or U3355 (N_3355,N_2985,N_2725);
and U3356 (N_3356,N_2749,N_2455);
nand U3357 (N_3357,N_2640,N_2983);
or U3358 (N_3358,N_2962,N_2841);
or U3359 (N_3359,N_2327,N_2773);
nand U3360 (N_3360,N_2595,N_2476);
and U3361 (N_3361,N_2693,N_2975);
nand U3362 (N_3362,N_2501,N_2718);
xor U3363 (N_3363,N_2469,N_2322);
nand U3364 (N_3364,N_2375,N_2969);
nand U3365 (N_3365,N_2553,N_2452);
and U3366 (N_3366,N_2320,N_2305);
and U3367 (N_3367,N_2581,N_2838);
nor U3368 (N_3368,N_2964,N_2660);
nand U3369 (N_3369,N_2291,N_2954);
or U3370 (N_3370,N_2425,N_2883);
xor U3371 (N_3371,N_2576,N_2401);
nor U3372 (N_3372,N_2295,N_2359);
nand U3373 (N_3373,N_2739,N_2653);
and U3374 (N_3374,N_2358,N_2821);
or U3375 (N_3375,N_2638,N_2654);
or U3376 (N_3376,N_2882,N_2337);
or U3377 (N_3377,N_2857,N_2567);
and U3378 (N_3378,N_2763,N_2303);
and U3379 (N_3379,N_2891,N_2945);
and U3380 (N_3380,N_2594,N_2782);
nand U3381 (N_3381,N_2949,N_2937);
xor U3382 (N_3382,N_2569,N_2433);
xnor U3383 (N_3383,N_2485,N_2776);
xor U3384 (N_3384,N_2702,N_2399);
nor U3385 (N_3385,N_2389,N_2956);
or U3386 (N_3386,N_2332,N_2727);
nand U3387 (N_3387,N_2650,N_2938);
or U3388 (N_3388,N_2982,N_2887);
xnor U3389 (N_3389,N_2598,N_2970);
nor U3390 (N_3390,N_2959,N_2261);
nand U3391 (N_3391,N_2338,N_2663);
nand U3392 (N_3392,N_2902,N_2887);
xnor U3393 (N_3393,N_2432,N_2927);
nor U3394 (N_3394,N_2826,N_2635);
xnor U3395 (N_3395,N_2798,N_2599);
nand U3396 (N_3396,N_2556,N_2588);
or U3397 (N_3397,N_2524,N_2457);
xor U3398 (N_3398,N_2460,N_2996);
nand U3399 (N_3399,N_2894,N_2261);
nor U3400 (N_3400,N_2979,N_2582);
nand U3401 (N_3401,N_2389,N_2788);
and U3402 (N_3402,N_2685,N_2520);
and U3403 (N_3403,N_2813,N_2920);
nand U3404 (N_3404,N_2640,N_2436);
xnor U3405 (N_3405,N_2879,N_2449);
xor U3406 (N_3406,N_2998,N_2600);
and U3407 (N_3407,N_2817,N_2563);
and U3408 (N_3408,N_2276,N_2670);
or U3409 (N_3409,N_2706,N_2573);
or U3410 (N_3410,N_2739,N_2635);
or U3411 (N_3411,N_2489,N_2560);
nand U3412 (N_3412,N_2770,N_2347);
or U3413 (N_3413,N_2901,N_2874);
nand U3414 (N_3414,N_2264,N_2433);
xor U3415 (N_3415,N_2685,N_2468);
nor U3416 (N_3416,N_2263,N_2904);
or U3417 (N_3417,N_2919,N_2389);
nand U3418 (N_3418,N_2720,N_2464);
and U3419 (N_3419,N_2923,N_2430);
nor U3420 (N_3420,N_2474,N_2575);
nor U3421 (N_3421,N_2465,N_2326);
nor U3422 (N_3422,N_2631,N_2773);
and U3423 (N_3423,N_2269,N_2985);
and U3424 (N_3424,N_2400,N_2390);
and U3425 (N_3425,N_2719,N_2411);
nand U3426 (N_3426,N_2966,N_2905);
and U3427 (N_3427,N_2439,N_2466);
xnor U3428 (N_3428,N_2994,N_2439);
or U3429 (N_3429,N_2830,N_2355);
nand U3430 (N_3430,N_2850,N_2677);
and U3431 (N_3431,N_2589,N_2340);
or U3432 (N_3432,N_2720,N_2667);
nor U3433 (N_3433,N_2476,N_2464);
nand U3434 (N_3434,N_2795,N_2550);
nor U3435 (N_3435,N_2833,N_2258);
xnor U3436 (N_3436,N_2716,N_2505);
nor U3437 (N_3437,N_2272,N_2723);
nand U3438 (N_3438,N_2788,N_2469);
and U3439 (N_3439,N_2695,N_2322);
xor U3440 (N_3440,N_2271,N_2767);
nor U3441 (N_3441,N_2792,N_2449);
nand U3442 (N_3442,N_2864,N_2886);
nor U3443 (N_3443,N_2422,N_2508);
nand U3444 (N_3444,N_2577,N_2782);
xnor U3445 (N_3445,N_2322,N_2881);
or U3446 (N_3446,N_2529,N_2322);
or U3447 (N_3447,N_2489,N_2415);
or U3448 (N_3448,N_2356,N_2723);
nor U3449 (N_3449,N_2560,N_2698);
xnor U3450 (N_3450,N_2287,N_2426);
or U3451 (N_3451,N_2253,N_2472);
nand U3452 (N_3452,N_2483,N_2826);
xor U3453 (N_3453,N_2525,N_2824);
and U3454 (N_3454,N_2568,N_2904);
or U3455 (N_3455,N_2830,N_2564);
nand U3456 (N_3456,N_2419,N_2960);
or U3457 (N_3457,N_2411,N_2277);
nand U3458 (N_3458,N_2965,N_2854);
nand U3459 (N_3459,N_2352,N_2727);
xor U3460 (N_3460,N_2853,N_2955);
xor U3461 (N_3461,N_2631,N_2998);
and U3462 (N_3462,N_2374,N_2284);
and U3463 (N_3463,N_2411,N_2959);
and U3464 (N_3464,N_2901,N_2319);
nand U3465 (N_3465,N_2550,N_2830);
nand U3466 (N_3466,N_2745,N_2267);
xnor U3467 (N_3467,N_2270,N_2512);
nand U3468 (N_3468,N_2616,N_2927);
xnor U3469 (N_3469,N_2837,N_2811);
and U3470 (N_3470,N_2876,N_2302);
nand U3471 (N_3471,N_2397,N_2998);
xor U3472 (N_3472,N_2699,N_2480);
nand U3473 (N_3473,N_2972,N_2980);
or U3474 (N_3474,N_2783,N_2795);
xor U3475 (N_3475,N_2569,N_2264);
and U3476 (N_3476,N_2538,N_2935);
xor U3477 (N_3477,N_2694,N_2612);
xnor U3478 (N_3478,N_2974,N_2579);
nor U3479 (N_3479,N_2962,N_2882);
nor U3480 (N_3480,N_2504,N_2441);
and U3481 (N_3481,N_2408,N_2579);
nor U3482 (N_3482,N_2599,N_2551);
nand U3483 (N_3483,N_2884,N_2336);
xor U3484 (N_3484,N_2507,N_2790);
and U3485 (N_3485,N_2314,N_2550);
or U3486 (N_3486,N_2919,N_2992);
or U3487 (N_3487,N_2509,N_2763);
xor U3488 (N_3488,N_2320,N_2917);
nand U3489 (N_3489,N_2860,N_2397);
or U3490 (N_3490,N_2878,N_2976);
xnor U3491 (N_3491,N_2921,N_2737);
xnor U3492 (N_3492,N_2539,N_2642);
nor U3493 (N_3493,N_2498,N_2263);
and U3494 (N_3494,N_2929,N_2641);
nand U3495 (N_3495,N_2482,N_2442);
nor U3496 (N_3496,N_2798,N_2791);
nor U3497 (N_3497,N_2753,N_2580);
xnor U3498 (N_3498,N_2802,N_2914);
or U3499 (N_3499,N_2887,N_2613);
xor U3500 (N_3500,N_2322,N_2604);
xnor U3501 (N_3501,N_2516,N_2416);
nand U3502 (N_3502,N_2387,N_2675);
or U3503 (N_3503,N_2742,N_2580);
xnor U3504 (N_3504,N_2711,N_2360);
xnor U3505 (N_3505,N_2330,N_2831);
nand U3506 (N_3506,N_2787,N_2319);
xor U3507 (N_3507,N_2483,N_2701);
nand U3508 (N_3508,N_2397,N_2425);
nor U3509 (N_3509,N_2348,N_2996);
or U3510 (N_3510,N_2367,N_2318);
nand U3511 (N_3511,N_2620,N_2894);
nor U3512 (N_3512,N_2374,N_2463);
or U3513 (N_3513,N_2810,N_2787);
nand U3514 (N_3514,N_2590,N_2945);
and U3515 (N_3515,N_2978,N_2587);
or U3516 (N_3516,N_2561,N_2339);
nor U3517 (N_3517,N_2355,N_2330);
xor U3518 (N_3518,N_2900,N_2668);
nor U3519 (N_3519,N_2724,N_2892);
or U3520 (N_3520,N_2804,N_2600);
and U3521 (N_3521,N_2279,N_2320);
nor U3522 (N_3522,N_2628,N_2633);
nor U3523 (N_3523,N_2610,N_2572);
nor U3524 (N_3524,N_2973,N_2771);
or U3525 (N_3525,N_2310,N_2430);
and U3526 (N_3526,N_2520,N_2514);
xnor U3527 (N_3527,N_2787,N_2738);
xor U3528 (N_3528,N_2291,N_2457);
or U3529 (N_3529,N_2308,N_2282);
nand U3530 (N_3530,N_2417,N_2591);
xor U3531 (N_3531,N_2577,N_2579);
nor U3532 (N_3532,N_2666,N_2952);
and U3533 (N_3533,N_2993,N_2974);
or U3534 (N_3534,N_2503,N_2425);
nor U3535 (N_3535,N_2703,N_2258);
and U3536 (N_3536,N_2604,N_2372);
xor U3537 (N_3537,N_2320,N_2251);
nand U3538 (N_3538,N_2532,N_2873);
nand U3539 (N_3539,N_2353,N_2842);
or U3540 (N_3540,N_2262,N_2924);
nor U3541 (N_3541,N_2475,N_2960);
and U3542 (N_3542,N_2503,N_2398);
nor U3543 (N_3543,N_2755,N_2743);
nor U3544 (N_3544,N_2986,N_2269);
or U3545 (N_3545,N_2266,N_2670);
xnor U3546 (N_3546,N_2427,N_2784);
nor U3547 (N_3547,N_2928,N_2334);
xnor U3548 (N_3548,N_2571,N_2787);
and U3549 (N_3549,N_2659,N_2483);
xnor U3550 (N_3550,N_2716,N_2868);
and U3551 (N_3551,N_2546,N_2773);
or U3552 (N_3552,N_2394,N_2365);
and U3553 (N_3553,N_2333,N_2991);
xor U3554 (N_3554,N_2766,N_2556);
nand U3555 (N_3555,N_2506,N_2660);
xnor U3556 (N_3556,N_2331,N_2725);
xnor U3557 (N_3557,N_2448,N_2811);
nand U3558 (N_3558,N_2591,N_2308);
xnor U3559 (N_3559,N_2544,N_2783);
or U3560 (N_3560,N_2310,N_2852);
or U3561 (N_3561,N_2594,N_2981);
nand U3562 (N_3562,N_2357,N_2288);
and U3563 (N_3563,N_2262,N_2339);
nor U3564 (N_3564,N_2303,N_2379);
and U3565 (N_3565,N_2293,N_2328);
nor U3566 (N_3566,N_2888,N_2272);
and U3567 (N_3567,N_2716,N_2684);
or U3568 (N_3568,N_2304,N_2368);
xnor U3569 (N_3569,N_2507,N_2946);
and U3570 (N_3570,N_2992,N_2573);
nand U3571 (N_3571,N_2954,N_2507);
xor U3572 (N_3572,N_2565,N_2717);
nor U3573 (N_3573,N_2335,N_2658);
xnor U3574 (N_3574,N_2910,N_2609);
xor U3575 (N_3575,N_2908,N_2374);
xnor U3576 (N_3576,N_2808,N_2448);
and U3577 (N_3577,N_2568,N_2623);
xnor U3578 (N_3578,N_2369,N_2814);
xnor U3579 (N_3579,N_2327,N_2507);
nor U3580 (N_3580,N_2839,N_2292);
xnor U3581 (N_3581,N_2803,N_2681);
nand U3582 (N_3582,N_2251,N_2687);
xnor U3583 (N_3583,N_2830,N_2874);
nand U3584 (N_3584,N_2889,N_2929);
or U3585 (N_3585,N_2423,N_2835);
nor U3586 (N_3586,N_2841,N_2958);
nor U3587 (N_3587,N_2545,N_2824);
and U3588 (N_3588,N_2747,N_2999);
nand U3589 (N_3589,N_2843,N_2443);
xnor U3590 (N_3590,N_2779,N_2757);
and U3591 (N_3591,N_2997,N_2785);
nand U3592 (N_3592,N_2638,N_2328);
nor U3593 (N_3593,N_2917,N_2797);
and U3594 (N_3594,N_2608,N_2877);
or U3595 (N_3595,N_2879,N_2940);
or U3596 (N_3596,N_2785,N_2772);
nor U3597 (N_3597,N_2607,N_2469);
xnor U3598 (N_3598,N_2396,N_2962);
xor U3599 (N_3599,N_2418,N_2448);
and U3600 (N_3600,N_2915,N_2709);
xor U3601 (N_3601,N_2672,N_2363);
and U3602 (N_3602,N_2414,N_2413);
and U3603 (N_3603,N_2371,N_2256);
or U3604 (N_3604,N_2813,N_2541);
xnor U3605 (N_3605,N_2773,N_2484);
nand U3606 (N_3606,N_2344,N_2845);
nand U3607 (N_3607,N_2942,N_2914);
nor U3608 (N_3608,N_2859,N_2835);
and U3609 (N_3609,N_2467,N_2560);
or U3610 (N_3610,N_2829,N_2876);
nand U3611 (N_3611,N_2326,N_2350);
or U3612 (N_3612,N_2492,N_2833);
xnor U3613 (N_3613,N_2402,N_2323);
nor U3614 (N_3614,N_2715,N_2377);
nand U3615 (N_3615,N_2311,N_2551);
nor U3616 (N_3616,N_2980,N_2932);
xnor U3617 (N_3617,N_2330,N_2400);
and U3618 (N_3618,N_2400,N_2775);
nand U3619 (N_3619,N_2399,N_2650);
xor U3620 (N_3620,N_2476,N_2902);
nor U3621 (N_3621,N_2736,N_2707);
xor U3622 (N_3622,N_2339,N_2445);
or U3623 (N_3623,N_2632,N_2404);
nor U3624 (N_3624,N_2780,N_2985);
nand U3625 (N_3625,N_2373,N_2855);
nand U3626 (N_3626,N_2560,N_2753);
nor U3627 (N_3627,N_2515,N_2550);
nor U3628 (N_3628,N_2438,N_2451);
and U3629 (N_3629,N_2790,N_2695);
and U3630 (N_3630,N_2286,N_2400);
or U3631 (N_3631,N_2585,N_2817);
and U3632 (N_3632,N_2985,N_2266);
or U3633 (N_3633,N_2571,N_2592);
xor U3634 (N_3634,N_2619,N_2739);
nand U3635 (N_3635,N_2361,N_2523);
nand U3636 (N_3636,N_2925,N_2285);
and U3637 (N_3637,N_2941,N_2917);
nor U3638 (N_3638,N_2818,N_2753);
nor U3639 (N_3639,N_2418,N_2699);
nor U3640 (N_3640,N_2303,N_2940);
nor U3641 (N_3641,N_2278,N_2788);
nor U3642 (N_3642,N_2504,N_2591);
xor U3643 (N_3643,N_2441,N_2425);
nor U3644 (N_3644,N_2810,N_2757);
nor U3645 (N_3645,N_2391,N_2561);
or U3646 (N_3646,N_2459,N_2470);
or U3647 (N_3647,N_2432,N_2871);
nand U3648 (N_3648,N_2638,N_2836);
xnor U3649 (N_3649,N_2530,N_2911);
nand U3650 (N_3650,N_2928,N_2752);
xnor U3651 (N_3651,N_2707,N_2764);
xor U3652 (N_3652,N_2555,N_2534);
or U3653 (N_3653,N_2748,N_2530);
nand U3654 (N_3654,N_2936,N_2528);
xor U3655 (N_3655,N_2380,N_2547);
and U3656 (N_3656,N_2484,N_2756);
nor U3657 (N_3657,N_2924,N_2302);
xor U3658 (N_3658,N_2779,N_2858);
or U3659 (N_3659,N_2610,N_2992);
xor U3660 (N_3660,N_2416,N_2558);
nand U3661 (N_3661,N_2985,N_2574);
nor U3662 (N_3662,N_2614,N_2360);
nand U3663 (N_3663,N_2736,N_2411);
or U3664 (N_3664,N_2291,N_2894);
or U3665 (N_3665,N_2641,N_2904);
and U3666 (N_3666,N_2837,N_2979);
nand U3667 (N_3667,N_2256,N_2815);
nand U3668 (N_3668,N_2863,N_2267);
nor U3669 (N_3669,N_2920,N_2562);
nor U3670 (N_3670,N_2900,N_2645);
xnor U3671 (N_3671,N_2259,N_2543);
or U3672 (N_3672,N_2475,N_2283);
nand U3673 (N_3673,N_2784,N_2420);
nand U3674 (N_3674,N_2881,N_2868);
and U3675 (N_3675,N_2905,N_2722);
or U3676 (N_3676,N_2938,N_2358);
or U3677 (N_3677,N_2881,N_2967);
and U3678 (N_3678,N_2536,N_2694);
nand U3679 (N_3679,N_2828,N_2525);
nand U3680 (N_3680,N_2551,N_2537);
or U3681 (N_3681,N_2355,N_2429);
and U3682 (N_3682,N_2503,N_2378);
or U3683 (N_3683,N_2271,N_2922);
or U3684 (N_3684,N_2882,N_2420);
nor U3685 (N_3685,N_2663,N_2747);
nor U3686 (N_3686,N_2289,N_2992);
and U3687 (N_3687,N_2690,N_2644);
nor U3688 (N_3688,N_2372,N_2492);
and U3689 (N_3689,N_2606,N_2934);
nor U3690 (N_3690,N_2409,N_2572);
nand U3691 (N_3691,N_2766,N_2696);
nor U3692 (N_3692,N_2641,N_2997);
or U3693 (N_3693,N_2293,N_2395);
nand U3694 (N_3694,N_2407,N_2321);
nor U3695 (N_3695,N_2307,N_2518);
and U3696 (N_3696,N_2375,N_2496);
nand U3697 (N_3697,N_2522,N_2996);
and U3698 (N_3698,N_2787,N_2762);
nand U3699 (N_3699,N_2877,N_2678);
xor U3700 (N_3700,N_2282,N_2912);
or U3701 (N_3701,N_2530,N_2351);
nand U3702 (N_3702,N_2743,N_2820);
nor U3703 (N_3703,N_2728,N_2344);
nand U3704 (N_3704,N_2471,N_2289);
or U3705 (N_3705,N_2524,N_2827);
nor U3706 (N_3706,N_2631,N_2571);
xor U3707 (N_3707,N_2563,N_2886);
nor U3708 (N_3708,N_2311,N_2829);
nand U3709 (N_3709,N_2613,N_2554);
or U3710 (N_3710,N_2719,N_2610);
or U3711 (N_3711,N_2442,N_2512);
and U3712 (N_3712,N_2607,N_2534);
or U3713 (N_3713,N_2554,N_2888);
or U3714 (N_3714,N_2952,N_2600);
and U3715 (N_3715,N_2825,N_2872);
nor U3716 (N_3716,N_2688,N_2909);
nor U3717 (N_3717,N_2790,N_2996);
nand U3718 (N_3718,N_2453,N_2254);
nand U3719 (N_3719,N_2858,N_2476);
nand U3720 (N_3720,N_2606,N_2260);
and U3721 (N_3721,N_2349,N_2687);
nor U3722 (N_3722,N_2592,N_2313);
and U3723 (N_3723,N_2977,N_2768);
nor U3724 (N_3724,N_2800,N_2714);
or U3725 (N_3725,N_2466,N_2648);
xor U3726 (N_3726,N_2858,N_2968);
or U3727 (N_3727,N_2401,N_2480);
xor U3728 (N_3728,N_2261,N_2761);
nand U3729 (N_3729,N_2631,N_2348);
nand U3730 (N_3730,N_2751,N_2998);
nand U3731 (N_3731,N_2373,N_2269);
nor U3732 (N_3732,N_2618,N_2686);
or U3733 (N_3733,N_2882,N_2490);
and U3734 (N_3734,N_2953,N_2442);
or U3735 (N_3735,N_2997,N_2795);
and U3736 (N_3736,N_2990,N_2455);
nor U3737 (N_3737,N_2426,N_2936);
or U3738 (N_3738,N_2296,N_2607);
nand U3739 (N_3739,N_2831,N_2567);
nor U3740 (N_3740,N_2673,N_2332);
nand U3741 (N_3741,N_2325,N_2453);
and U3742 (N_3742,N_2983,N_2707);
xor U3743 (N_3743,N_2537,N_2652);
nor U3744 (N_3744,N_2254,N_2505);
and U3745 (N_3745,N_2478,N_2268);
and U3746 (N_3746,N_2684,N_2994);
nor U3747 (N_3747,N_2925,N_2711);
nor U3748 (N_3748,N_2593,N_2834);
nor U3749 (N_3749,N_2714,N_2396);
nor U3750 (N_3750,N_3576,N_3545);
xor U3751 (N_3751,N_3726,N_3607);
nand U3752 (N_3752,N_3254,N_3094);
or U3753 (N_3753,N_3736,N_3089);
xor U3754 (N_3754,N_3129,N_3009);
xor U3755 (N_3755,N_3642,N_3533);
and U3756 (N_3756,N_3054,N_3543);
nand U3757 (N_3757,N_3041,N_3537);
xnor U3758 (N_3758,N_3738,N_3130);
xnor U3759 (N_3759,N_3617,N_3201);
or U3760 (N_3760,N_3683,N_3058);
xnor U3761 (N_3761,N_3223,N_3444);
nor U3762 (N_3762,N_3316,N_3463);
xnor U3763 (N_3763,N_3399,N_3148);
nand U3764 (N_3764,N_3234,N_3556);
nand U3765 (N_3765,N_3423,N_3300);
and U3766 (N_3766,N_3220,N_3559);
and U3767 (N_3767,N_3407,N_3066);
nand U3768 (N_3768,N_3677,N_3579);
and U3769 (N_3769,N_3627,N_3247);
and U3770 (N_3770,N_3048,N_3561);
or U3771 (N_3771,N_3386,N_3394);
and U3772 (N_3772,N_3601,N_3289);
or U3773 (N_3773,N_3733,N_3389);
nor U3774 (N_3774,N_3169,N_3431);
nand U3775 (N_3775,N_3266,N_3635);
or U3776 (N_3776,N_3060,N_3575);
or U3777 (N_3777,N_3645,N_3414);
xor U3778 (N_3778,N_3720,N_3078);
nand U3779 (N_3779,N_3728,N_3090);
xor U3780 (N_3780,N_3013,N_3430);
xor U3781 (N_3781,N_3314,N_3737);
nor U3782 (N_3782,N_3401,N_3465);
nand U3783 (N_3783,N_3320,N_3290);
xor U3784 (N_3784,N_3714,N_3517);
nor U3785 (N_3785,N_3330,N_3236);
xor U3786 (N_3786,N_3040,N_3535);
nand U3787 (N_3787,N_3364,N_3433);
nor U3788 (N_3788,N_3280,N_3570);
nor U3789 (N_3789,N_3075,N_3206);
or U3790 (N_3790,N_3719,N_3388);
nand U3791 (N_3791,N_3099,N_3208);
nand U3792 (N_3792,N_3548,N_3251);
nand U3793 (N_3793,N_3055,N_3161);
and U3794 (N_3794,N_3634,N_3437);
and U3795 (N_3795,N_3422,N_3195);
nor U3796 (N_3796,N_3371,N_3313);
nor U3797 (N_3797,N_3349,N_3295);
and U3798 (N_3798,N_3178,N_3176);
nor U3799 (N_3799,N_3032,N_3385);
xnor U3800 (N_3800,N_3049,N_3331);
xnor U3801 (N_3801,N_3270,N_3187);
and U3802 (N_3802,N_3566,N_3310);
xnor U3803 (N_3803,N_3749,N_3411);
xor U3804 (N_3804,N_3588,N_3450);
or U3805 (N_3805,N_3029,N_3079);
xnor U3806 (N_3806,N_3492,N_3328);
nor U3807 (N_3807,N_3097,N_3088);
xor U3808 (N_3808,N_3586,N_3235);
and U3809 (N_3809,N_3644,N_3151);
xnor U3810 (N_3810,N_3037,N_3282);
nand U3811 (N_3811,N_3549,N_3268);
and U3812 (N_3812,N_3360,N_3044);
and U3813 (N_3813,N_3214,N_3038);
nor U3814 (N_3814,N_3226,N_3231);
nand U3815 (N_3815,N_3536,N_3397);
nor U3816 (N_3816,N_3370,N_3014);
and U3817 (N_3817,N_3315,N_3229);
nand U3818 (N_3818,N_3356,N_3686);
xor U3819 (N_3819,N_3589,N_3082);
and U3820 (N_3820,N_3294,N_3241);
and U3821 (N_3821,N_3018,N_3454);
or U3822 (N_3822,N_3189,N_3653);
or U3823 (N_3823,N_3269,N_3134);
and U3824 (N_3824,N_3352,N_3580);
nor U3825 (N_3825,N_3516,N_3552);
xor U3826 (N_3826,N_3194,N_3396);
xor U3827 (N_3827,N_3286,N_3500);
or U3828 (N_3828,N_3156,N_3363);
xnor U3829 (N_3829,N_3664,N_3059);
xor U3830 (N_3830,N_3168,N_3404);
nand U3831 (N_3831,N_3452,N_3680);
nor U3832 (N_3832,N_3626,N_3693);
or U3833 (N_3833,N_3419,N_3367);
nor U3834 (N_3834,N_3380,N_3682);
or U3835 (N_3835,N_3460,N_3581);
or U3836 (N_3836,N_3424,N_3563);
or U3837 (N_3837,N_3152,N_3636);
or U3838 (N_3838,N_3687,N_3621);
and U3839 (N_3839,N_3122,N_3184);
nor U3840 (N_3840,N_3615,N_3470);
nor U3841 (N_3841,N_3354,N_3696);
nor U3842 (N_3842,N_3056,N_3299);
xor U3843 (N_3843,N_3068,N_3409);
xnor U3844 (N_3844,N_3429,N_3622);
nand U3845 (N_3845,N_3408,N_3468);
nor U3846 (N_3846,N_3547,N_3724);
nand U3847 (N_3847,N_3709,N_3238);
xnor U3848 (N_3848,N_3637,N_3233);
nor U3849 (N_3849,N_3115,N_3618);
or U3850 (N_3850,N_3106,N_3670);
nor U3851 (N_3851,N_3390,N_3623);
nand U3852 (N_3852,N_3193,N_3739);
and U3853 (N_3853,N_3480,N_3348);
nor U3854 (N_3854,N_3554,N_3139);
nor U3855 (N_3855,N_3436,N_3112);
nor U3856 (N_3856,N_3077,N_3024);
nor U3857 (N_3857,N_3522,N_3103);
nand U3858 (N_3858,N_3309,N_3050);
and U3859 (N_3859,N_3641,N_3610);
nor U3860 (N_3860,N_3676,N_3272);
xnor U3861 (N_3861,N_3159,N_3204);
and U3862 (N_3862,N_3126,N_3180);
nor U3863 (N_3863,N_3123,N_3202);
xor U3864 (N_3864,N_3303,N_3661);
nand U3865 (N_3865,N_3023,N_3649);
nor U3866 (N_3866,N_3695,N_3080);
or U3867 (N_3867,N_3592,N_3509);
or U3868 (N_3868,N_3342,N_3368);
nor U3869 (N_3869,N_3069,N_3132);
xor U3870 (N_3870,N_3485,N_3101);
and U3871 (N_3871,N_3667,N_3525);
xnor U3872 (N_3872,N_3604,N_3486);
or U3873 (N_3873,N_3074,N_3650);
xnor U3874 (N_3874,N_3491,N_3643);
or U3875 (N_3875,N_3387,N_3353);
and U3876 (N_3876,N_3108,N_3438);
xnor U3877 (N_3877,N_3402,N_3476);
nand U3878 (N_3878,N_3716,N_3250);
and U3879 (N_3879,N_3662,N_3495);
nor U3880 (N_3880,N_3551,N_3731);
and U3881 (N_3881,N_3020,N_3347);
nand U3882 (N_3882,N_3003,N_3712);
nand U3883 (N_3883,N_3186,N_3471);
xor U3884 (N_3884,N_3141,N_3256);
or U3885 (N_3885,N_3301,N_3513);
nor U3886 (N_3886,N_3200,N_3374);
and U3887 (N_3887,N_3598,N_3420);
nor U3888 (N_3888,N_3199,N_3067);
nor U3889 (N_3889,N_3605,N_3116);
and U3890 (N_3890,N_3619,N_3369);
nand U3891 (N_3891,N_3242,N_3722);
nor U3892 (N_3892,N_3669,N_3361);
or U3893 (N_3893,N_3191,N_3445);
nand U3894 (N_3894,N_3705,N_3277);
and U3895 (N_3895,N_3744,N_3603);
nand U3896 (N_3896,N_3703,N_3497);
or U3897 (N_3897,N_3150,N_3616);
or U3898 (N_3898,N_3560,N_3681);
xor U3899 (N_3899,N_3614,N_3612);
xor U3900 (N_3900,N_3594,N_3036);
nor U3901 (N_3901,N_3217,N_3655);
or U3902 (N_3902,N_3671,N_3568);
nor U3903 (N_3903,N_3087,N_3392);
or U3904 (N_3904,N_3698,N_3222);
or U3905 (N_3905,N_3104,N_3708);
xor U3906 (N_3906,N_3324,N_3039);
or U3907 (N_3907,N_3228,N_3591);
nor U3908 (N_3908,N_3011,N_3219);
or U3909 (N_3909,N_3205,N_3167);
or U3910 (N_3910,N_3015,N_3262);
xor U3911 (N_3911,N_3413,N_3117);
nand U3912 (N_3912,N_3322,N_3110);
and U3913 (N_3913,N_3625,N_3273);
nor U3914 (N_3914,N_3073,N_3569);
and U3915 (N_3915,N_3439,N_3538);
xnor U3916 (N_3916,N_3210,N_3532);
nor U3917 (N_3917,N_3428,N_3479);
nor U3918 (N_3918,N_3658,N_3263);
xor U3919 (N_3919,N_3212,N_3453);
and U3920 (N_3920,N_3511,N_3578);
nand U3921 (N_3921,N_3028,N_3045);
xnor U3922 (N_3922,N_3499,N_3692);
or U3923 (N_3923,N_3629,N_3595);
xor U3924 (N_3924,N_3230,N_3248);
nand U3925 (N_3925,N_3145,N_3417);
nand U3926 (N_3926,N_3652,N_3083);
xnor U3927 (N_3927,N_3425,N_3672);
xor U3928 (N_3928,N_3391,N_3285);
and U3929 (N_3929,N_3466,N_3304);
and U3930 (N_3930,N_3244,N_3524);
and U3931 (N_3931,N_3031,N_3657);
nor U3932 (N_3932,N_3260,N_3179);
and U3933 (N_3933,N_3157,N_3172);
or U3934 (N_3934,N_3362,N_3196);
and U3935 (N_3935,N_3225,N_3227);
or U3936 (N_3936,N_3648,N_3442);
and U3937 (N_3937,N_3472,N_3490);
xnor U3938 (N_3938,N_3174,N_3613);
nand U3939 (N_3939,N_3035,N_3084);
nor U3940 (N_3940,N_3427,N_3656);
nor U3941 (N_3941,N_3384,N_3530);
nor U3942 (N_3942,N_3489,N_3734);
nor U3943 (N_3943,N_3091,N_3173);
and U3944 (N_3944,N_3701,N_3119);
nor U3945 (N_3945,N_3046,N_3507);
and U3946 (N_3946,N_3221,N_3383);
and U3947 (N_3947,N_3382,N_3582);
and U3948 (N_3948,N_3639,N_3001);
or U3949 (N_3949,N_3170,N_3093);
and U3950 (N_3950,N_3631,N_3654);
nand U3951 (N_3951,N_3715,N_3329);
nor U3952 (N_3952,N_3539,N_3240);
and U3953 (N_3953,N_3555,N_3451);
and U3954 (N_3954,N_3181,N_3732);
nor U3955 (N_3955,N_3171,N_3307);
and U3956 (N_3956,N_3550,N_3688);
or U3957 (N_3957,N_3518,N_3574);
and U3958 (N_3958,N_3135,N_3502);
xnor U3959 (N_3959,N_3593,N_3081);
or U3960 (N_3960,N_3042,N_3526);
nor U3961 (N_3961,N_3432,N_3455);
nor U3962 (N_3962,N_3558,N_3577);
and U3963 (N_3963,N_3585,N_3350);
or U3964 (N_3964,N_3335,N_3124);
and U3965 (N_3965,N_3164,N_3140);
xor U3966 (N_3966,N_3209,N_3332);
or U3967 (N_3967,N_3506,N_3085);
nor U3968 (N_3968,N_3611,N_3211);
nor U3969 (N_3969,N_3323,N_3718);
nand U3970 (N_3970,N_3052,N_3183);
nor U3971 (N_3971,N_3488,N_3447);
xor U3972 (N_3972,N_3267,N_3410);
xnor U3973 (N_3973,N_3512,N_3632);
nand U3974 (N_3974,N_3665,N_3062);
and U3975 (N_3975,N_3478,N_3334);
nand U3976 (N_3976,N_3337,N_3487);
xor U3977 (N_3977,N_3684,N_3441);
xnor U3978 (N_3978,N_3344,N_3449);
xnor U3979 (N_3979,N_3540,N_3072);
nand U3980 (N_3980,N_3146,N_3587);
xnor U3981 (N_3981,N_3065,N_3531);
or U3982 (N_3982,N_3076,N_3608);
xnor U3983 (N_3983,N_3203,N_3259);
or U3984 (N_3984,N_3375,N_3275);
nand U3985 (N_3985,N_3448,N_3022);
or U3986 (N_3986,N_3306,N_3061);
nand U3987 (N_3987,N_3128,N_3546);
and U3988 (N_3988,N_3057,N_3120);
or U3989 (N_3989,N_3457,N_3702);
xnor U3990 (N_3990,N_3748,N_3249);
nand U3991 (N_3991,N_3679,N_3373);
xnor U3992 (N_3992,N_3366,N_3175);
nor U3993 (N_3993,N_3659,N_3529);
and U3994 (N_3994,N_3121,N_3185);
nor U3995 (N_3995,N_3005,N_3494);
or U3996 (N_3996,N_3070,N_3276);
or U3997 (N_3997,N_3102,N_3302);
nand U3998 (N_3998,N_3508,N_3343);
or U3999 (N_3999,N_3421,N_3160);
nor U4000 (N_4000,N_3572,N_3503);
xor U4001 (N_4001,N_3137,N_3026);
or U4002 (N_4002,N_3461,N_3237);
and U4003 (N_4003,N_3745,N_3271);
nor U4004 (N_4004,N_3138,N_3707);
and U4005 (N_4005,N_3341,N_3136);
or U4006 (N_4006,N_3400,N_3198);
or U4007 (N_4007,N_3673,N_3747);
nor U4008 (N_4008,N_3590,N_3190);
nand U4009 (N_4009,N_3215,N_3691);
nand U4010 (N_4010,N_3006,N_3469);
or U4011 (N_4011,N_3064,N_3446);
nor U4012 (N_4012,N_3142,N_3327);
xor U4013 (N_4013,N_3154,N_3418);
nand U4014 (N_4014,N_3111,N_3165);
xor U4015 (N_4015,N_3440,N_3412);
or U4016 (N_4016,N_3562,N_3007);
or U4017 (N_4017,N_3246,N_3188);
xnor U4018 (N_4018,N_3381,N_3265);
xor U4019 (N_4019,N_3321,N_3646);
nand U4020 (N_4020,N_3741,N_3027);
xnor U4021 (N_4021,N_3207,N_3434);
nor U4022 (N_4022,N_3378,N_3264);
xnor U4023 (N_4023,N_3481,N_3501);
nor U4024 (N_4024,N_3326,N_3542);
xor U4025 (N_4025,N_3279,N_3257);
nand U4026 (N_4026,N_3125,N_3034);
nand U4027 (N_4027,N_3395,N_3729);
nand U4028 (N_4028,N_3192,N_3131);
nand U4029 (N_4029,N_3483,N_3095);
nand U4030 (N_4030,N_3177,N_3651);
nor U4031 (N_4031,N_3700,N_3514);
and U4032 (N_4032,N_3443,N_3710);
xnor U4033 (N_4033,N_3435,N_3092);
and U4034 (N_4034,N_3458,N_3298);
or U4035 (N_4035,N_3505,N_3305);
or U4036 (N_4036,N_3398,N_3030);
nand U4037 (N_4037,N_3484,N_3357);
xor U4038 (N_4038,N_3515,N_3312);
nor U4039 (N_4039,N_3105,N_3377);
nand U4040 (N_4040,N_3415,N_3292);
nor U4041 (N_4041,N_3606,N_3406);
xor U4042 (N_4042,N_3287,N_3359);
and U4043 (N_4043,N_3063,N_3100);
xnor U4044 (N_4044,N_3699,N_3735);
and U4045 (N_4045,N_3118,N_3557);
xor U4046 (N_4046,N_3182,N_3743);
nand U4047 (N_4047,N_3033,N_3475);
nor U4048 (N_4048,N_3213,N_3721);
and U4049 (N_4049,N_3496,N_3467);
and U4050 (N_4050,N_3153,N_3010);
xnor U4051 (N_4051,N_3723,N_3746);
nor U4052 (N_4052,N_3000,N_3544);
or U4053 (N_4053,N_3311,N_3288);
and U4054 (N_4054,N_3628,N_3086);
nor U4055 (N_4055,N_3678,N_3053);
and U4056 (N_4056,N_3109,N_3197);
nor U4057 (N_4057,N_3143,N_3583);
xnor U4058 (N_4058,N_3527,N_3564);
xnor U4059 (N_4059,N_3293,N_3346);
nor U4060 (N_4060,N_3163,N_3071);
or U4061 (N_4061,N_3459,N_3640);
and U4062 (N_4062,N_3573,N_3633);
nor U4063 (N_4063,N_3602,N_3740);
nor U4064 (N_4064,N_3283,N_3528);
or U4065 (N_4065,N_3666,N_3426);
nor U4066 (N_4066,N_3498,N_3553);
xnor U4067 (N_4067,N_3638,N_3008);
and U4068 (N_4068,N_3243,N_3252);
nand U4069 (N_4069,N_3534,N_3253);
nor U4070 (N_4070,N_3493,N_3351);
xnor U4071 (N_4071,N_3376,N_3218);
xor U4072 (N_4072,N_3224,N_3694);
or U4073 (N_4073,N_3372,N_3098);
and U4074 (N_4074,N_3245,N_3147);
and U4075 (N_4075,N_3620,N_3308);
and U4076 (N_4076,N_3477,N_3297);
nor U4077 (N_4077,N_3336,N_3405);
xnor U4078 (N_4078,N_3600,N_3379);
nand U4079 (N_4079,N_3403,N_3675);
nor U4080 (N_4080,N_3663,N_3519);
nor U4081 (N_4081,N_3599,N_3239);
or U4082 (N_4082,N_3624,N_3144);
xnor U4083 (N_4083,N_3510,N_3155);
or U4084 (N_4084,N_3365,N_3630);
xor U4085 (N_4085,N_3133,N_3473);
nand U4086 (N_4086,N_3149,N_3284);
nor U4087 (N_4087,N_3004,N_3043);
xor U4088 (N_4088,N_3660,N_3565);
nor U4089 (N_4089,N_3017,N_3355);
and U4090 (N_4090,N_3674,N_3345);
nor U4091 (N_4091,N_3019,N_3520);
and U4092 (N_4092,N_3456,N_3216);
and U4093 (N_4093,N_3462,N_3107);
xnor U4094 (N_4094,N_3278,N_3571);
nor U4095 (N_4095,N_3158,N_3647);
or U4096 (N_4096,N_3296,N_3711);
and U4097 (N_4097,N_3333,N_3725);
xnor U4098 (N_4098,N_3523,N_3464);
xor U4099 (N_4099,N_3704,N_3012);
nand U4100 (N_4100,N_3166,N_3317);
and U4101 (N_4101,N_3697,N_3325);
nand U4102 (N_4102,N_3114,N_3258);
or U4103 (N_4103,N_3358,N_3339);
or U4104 (N_4104,N_3541,N_3730);
nor U4105 (N_4105,N_3690,N_3597);
and U4106 (N_4106,N_3742,N_3002);
nand U4107 (N_4107,N_3596,N_3319);
or U4108 (N_4108,N_3255,N_3416);
nand U4109 (N_4109,N_3609,N_3504);
and U4110 (N_4110,N_3706,N_3291);
or U4111 (N_4111,N_3021,N_3051);
or U4112 (N_4112,N_3025,N_3713);
or U4113 (N_4113,N_3096,N_3474);
xnor U4114 (N_4114,N_3567,N_3261);
nand U4115 (N_4115,N_3685,N_3689);
nand U4116 (N_4116,N_3668,N_3340);
or U4117 (N_4117,N_3127,N_3162);
and U4118 (N_4118,N_3274,N_3717);
xor U4119 (N_4119,N_3393,N_3482);
nand U4120 (N_4120,N_3281,N_3047);
xor U4121 (N_4121,N_3016,N_3727);
nand U4122 (N_4122,N_3318,N_3521);
nand U4123 (N_4123,N_3232,N_3584);
nor U4124 (N_4124,N_3113,N_3338);
nand U4125 (N_4125,N_3739,N_3684);
nor U4126 (N_4126,N_3380,N_3119);
nand U4127 (N_4127,N_3702,N_3059);
or U4128 (N_4128,N_3333,N_3313);
and U4129 (N_4129,N_3688,N_3332);
nand U4130 (N_4130,N_3309,N_3637);
and U4131 (N_4131,N_3259,N_3396);
nand U4132 (N_4132,N_3217,N_3197);
and U4133 (N_4133,N_3454,N_3360);
nand U4134 (N_4134,N_3002,N_3411);
nor U4135 (N_4135,N_3073,N_3543);
xnor U4136 (N_4136,N_3552,N_3052);
and U4137 (N_4137,N_3019,N_3443);
xnor U4138 (N_4138,N_3329,N_3623);
nor U4139 (N_4139,N_3591,N_3621);
nand U4140 (N_4140,N_3200,N_3339);
xor U4141 (N_4141,N_3222,N_3395);
nand U4142 (N_4142,N_3169,N_3187);
xor U4143 (N_4143,N_3081,N_3046);
or U4144 (N_4144,N_3407,N_3656);
or U4145 (N_4145,N_3652,N_3141);
nand U4146 (N_4146,N_3277,N_3458);
xnor U4147 (N_4147,N_3393,N_3700);
xor U4148 (N_4148,N_3380,N_3254);
nand U4149 (N_4149,N_3566,N_3409);
nor U4150 (N_4150,N_3618,N_3568);
nand U4151 (N_4151,N_3712,N_3531);
and U4152 (N_4152,N_3080,N_3050);
nand U4153 (N_4153,N_3530,N_3354);
and U4154 (N_4154,N_3639,N_3589);
nor U4155 (N_4155,N_3196,N_3524);
and U4156 (N_4156,N_3127,N_3356);
nand U4157 (N_4157,N_3034,N_3452);
or U4158 (N_4158,N_3329,N_3612);
or U4159 (N_4159,N_3298,N_3018);
nor U4160 (N_4160,N_3320,N_3253);
and U4161 (N_4161,N_3231,N_3417);
and U4162 (N_4162,N_3276,N_3746);
nand U4163 (N_4163,N_3032,N_3298);
xor U4164 (N_4164,N_3532,N_3444);
and U4165 (N_4165,N_3090,N_3419);
and U4166 (N_4166,N_3615,N_3610);
nand U4167 (N_4167,N_3448,N_3369);
or U4168 (N_4168,N_3046,N_3329);
xnor U4169 (N_4169,N_3427,N_3673);
or U4170 (N_4170,N_3174,N_3039);
nand U4171 (N_4171,N_3270,N_3677);
xnor U4172 (N_4172,N_3160,N_3148);
nand U4173 (N_4173,N_3168,N_3376);
nor U4174 (N_4174,N_3459,N_3068);
or U4175 (N_4175,N_3596,N_3628);
nor U4176 (N_4176,N_3591,N_3729);
nand U4177 (N_4177,N_3261,N_3644);
or U4178 (N_4178,N_3073,N_3672);
nand U4179 (N_4179,N_3527,N_3742);
nor U4180 (N_4180,N_3403,N_3027);
and U4181 (N_4181,N_3615,N_3641);
or U4182 (N_4182,N_3376,N_3002);
or U4183 (N_4183,N_3708,N_3031);
and U4184 (N_4184,N_3552,N_3234);
nor U4185 (N_4185,N_3041,N_3545);
or U4186 (N_4186,N_3000,N_3358);
nand U4187 (N_4187,N_3655,N_3152);
and U4188 (N_4188,N_3678,N_3572);
or U4189 (N_4189,N_3284,N_3313);
or U4190 (N_4190,N_3458,N_3240);
nand U4191 (N_4191,N_3575,N_3615);
nor U4192 (N_4192,N_3005,N_3327);
and U4193 (N_4193,N_3168,N_3132);
nor U4194 (N_4194,N_3298,N_3171);
nand U4195 (N_4195,N_3541,N_3164);
and U4196 (N_4196,N_3230,N_3738);
or U4197 (N_4197,N_3633,N_3044);
and U4198 (N_4198,N_3690,N_3723);
and U4199 (N_4199,N_3604,N_3466);
or U4200 (N_4200,N_3160,N_3672);
nor U4201 (N_4201,N_3037,N_3642);
and U4202 (N_4202,N_3746,N_3585);
nand U4203 (N_4203,N_3293,N_3020);
or U4204 (N_4204,N_3667,N_3264);
nor U4205 (N_4205,N_3682,N_3080);
nand U4206 (N_4206,N_3602,N_3106);
or U4207 (N_4207,N_3353,N_3078);
nand U4208 (N_4208,N_3571,N_3360);
xnor U4209 (N_4209,N_3302,N_3019);
nor U4210 (N_4210,N_3320,N_3373);
nor U4211 (N_4211,N_3657,N_3295);
nor U4212 (N_4212,N_3403,N_3445);
and U4213 (N_4213,N_3699,N_3223);
nor U4214 (N_4214,N_3447,N_3546);
xnor U4215 (N_4215,N_3746,N_3548);
and U4216 (N_4216,N_3624,N_3074);
nor U4217 (N_4217,N_3245,N_3254);
or U4218 (N_4218,N_3545,N_3478);
xor U4219 (N_4219,N_3131,N_3468);
xnor U4220 (N_4220,N_3738,N_3343);
xor U4221 (N_4221,N_3021,N_3298);
and U4222 (N_4222,N_3379,N_3448);
nand U4223 (N_4223,N_3497,N_3552);
and U4224 (N_4224,N_3596,N_3563);
xor U4225 (N_4225,N_3202,N_3480);
xnor U4226 (N_4226,N_3549,N_3128);
and U4227 (N_4227,N_3038,N_3246);
nand U4228 (N_4228,N_3224,N_3115);
and U4229 (N_4229,N_3423,N_3028);
nand U4230 (N_4230,N_3367,N_3304);
xnor U4231 (N_4231,N_3124,N_3408);
or U4232 (N_4232,N_3061,N_3005);
xnor U4233 (N_4233,N_3080,N_3680);
xor U4234 (N_4234,N_3004,N_3293);
nand U4235 (N_4235,N_3339,N_3685);
nor U4236 (N_4236,N_3404,N_3647);
xor U4237 (N_4237,N_3042,N_3668);
nand U4238 (N_4238,N_3095,N_3283);
xnor U4239 (N_4239,N_3613,N_3493);
nand U4240 (N_4240,N_3371,N_3517);
and U4241 (N_4241,N_3513,N_3376);
nand U4242 (N_4242,N_3313,N_3137);
and U4243 (N_4243,N_3183,N_3286);
xor U4244 (N_4244,N_3417,N_3030);
nor U4245 (N_4245,N_3257,N_3556);
nor U4246 (N_4246,N_3690,N_3573);
or U4247 (N_4247,N_3271,N_3034);
and U4248 (N_4248,N_3342,N_3068);
xnor U4249 (N_4249,N_3144,N_3111);
nand U4250 (N_4250,N_3608,N_3691);
and U4251 (N_4251,N_3171,N_3591);
nor U4252 (N_4252,N_3340,N_3038);
and U4253 (N_4253,N_3384,N_3414);
nor U4254 (N_4254,N_3585,N_3712);
or U4255 (N_4255,N_3539,N_3364);
xor U4256 (N_4256,N_3676,N_3581);
or U4257 (N_4257,N_3349,N_3231);
nand U4258 (N_4258,N_3511,N_3690);
xnor U4259 (N_4259,N_3393,N_3525);
xor U4260 (N_4260,N_3064,N_3516);
or U4261 (N_4261,N_3684,N_3342);
xor U4262 (N_4262,N_3142,N_3118);
nor U4263 (N_4263,N_3513,N_3609);
and U4264 (N_4264,N_3581,N_3635);
nand U4265 (N_4265,N_3540,N_3188);
nand U4266 (N_4266,N_3720,N_3060);
nor U4267 (N_4267,N_3443,N_3284);
and U4268 (N_4268,N_3002,N_3113);
nand U4269 (N_4269,N_3293,N_3091);
nor U4270 (N_4270,N_3363,N_3115);
and U4271 (N_4271,N_3188,N_3148);
or U4272 (N_4272,N_3009,N_3418);
and U4273 (N_4273,N_3352,N_3586);
nor U4274 (N_4274,N_3329,N_3146);
xnor U4275 (N_4275,N_3133,N_3511);
nor U4276 (N_4276,N_3745,N_3191);
xor U4277 (N_4277,N_3242,N_3554);
xnor U4278 (N_4278,N_3114,N_3671);
xor U4279 (N_4279,N_3377,N_3142);
xor U4280 (N_4280,N_3201,N_3687);
xor U4281 (N_4281,N_3749,N_3730);
and U4282 (N_4282,N_3144,N_3203);
and U4283 (N_4283,N_3070,N_3253);
nand U4284 (N_4284,N_3185,N_3112);
nand U4285 (N_4285,N_3361,N_3649);
or U4286 (N_4286,N_3211,N_3356);
xnor U4287 (N_4287,N_3576,N_3713);
or U4288 (N_4288,N_3229,N_3658);
or U4289 (N_4289,N_3321,N_3519);
nand U4290 (N_4290,N_3748,N_3636);
nand U4291 (N_4291,N_3246,N_3682);
or U4292 (N_4292,N_3451,N_3558);
nand U4293 (N_4293,N_3653,N_3561);
and U4294 (N_4294,N_3169,N_3111);
nand U4295 (N_4295,N_3421,N_3739);
and U4296 (N_4296,N_3471,N_3392);
or U4297 (N_4297,N_3140,N_3421);
nand U4298 (N_4298,N_3734,N_3063);
xor U4299 (N_4299,N_3052,N_3335);
or U4300 (N_4300,N_3316,N_3128);
or U4301 (N_4301,N_3268,N_3196);
xor U4302 (N_4302,N_3209,N_3491);
nand U4303 (N_4303,N_3164,N_3721);
nor U4304 (N_4304,N_3669,N_3271);
xor U4305 (N_4305,N_3603,N_3459);
nand U4306 (N_4306,N_3354,N_3706);
nor U4307 (N_4307,N_3682,N_3305);
or U4308 (N_4308,N_3179,N_3242);
or U4309 (N_4309,N_3389,N_3554);
nor U4310 (N_4310,N_3247,N_3290);
or U4311 (N_4311,N_3584,N_3701);
nor U4312 (N_4312,N_3080,N_3406);
nor U4313 (N_4313,N_3092,N_3482);
nand U4314 (N_4314,N_3072,N_3415);
or U4315 (N_4315,N_3440,N_3617);
and U4316 (N_4316,N_3616,N_3069);
xnor U4317 (N_4317,N_3423,N_3710);
or U4318 (N_4318,N_3277,N_3518);
and U4319 (N_4319,N_3436,N_3055);
nand U4320 (N_4320,N_3138,N_3109);
nor U4321 (N_4321,N_3250,N_3188);
nand U4322 (N_4322,N_3554,N_3598);
or U4323 (N_4323,N_3585,N_3311);
nor U4324 (N_4324,N_3089,N_3311);
nor U4325 (N_4325,N_3019,N_3536);
xor U4326 (N_4326,N_3569,N_3529);
and U4327 (N_4327,N_3325,N_3061);
xnor U4328 (N_4328,N_3046,N_3442);
nand U4329 (N_4329,N_3474,N_3203);
or U4330 (N_4330,N_3745,N_3269);
or U4331 (N_4331,N_3574,N_3187);
nand U4332 (N_4332,N_3730,N_3103);
or U4333 (N_4333,N_3539,N_3037);
or U4334 (N_4334,N_3224,N_3029);
or U4335 (N_4335,N_3585,N_3018);
nand U4336 (N_4336,N_3563,N_3005);
nand U4337 (N_4337,N_3733,N_3142);
xor U4338 (N_4338,N_3626,N_3204);
nor U4339 (N_4339,N_3437,N_3085);
and U4340 (N_4340,N_3467,N_3748);
xor U4341 (N_4341,N_3188,N_3625);
nor U4342 (N_4342,N_3197,N_3513);
and U4343 (N_4343,N_3588,N_3464);
and U4344 (N_4344,N_3732,N_3145);
nor U4345 (N_4345,N_3357,N_3371);
or U4346 (N_4346,N_3722,N_3400);
nand U4347 (N_4347,N_3657,N_3522);
nor U4348 (N_4348,N_3197,N_3083);
nand U4349 (N_4349,N_3044,N_3344);
nor U4350 (N_4350,N_3106,N_3175);
and U4351 (N_4351,N_3180,N_3014);
nand U4352 (N_4352,N_3189,N_3342);
nand U4353 (N_4353,N_3120,N_3522);
nor U4354 (N_4354,N_3730,N_3487);
nor U4355 (N_4355,N_3329,N_3604);
or U4356 (N_4356,N_3711,N_3106);
xor U4357 (N_4357,N_3231,N_3108);
xnor U4358 (N_4358,N_3015,N_3252);
nor U4359 (N_4359,N_3475,N_3488);
nand U4360 (N_4360,N_3315,N_3234);
nor U4361 (N_4361,N_3239,N_3000);
xor U4362 (N_4362,N_3207,N_3545);
and U4363 (N_4363,N_3695,N_3217);
and U4364 (N_4364,N_3066,N_3337);
xor U4365 (N_4365,N_3109,N_3686);
nor U4366 (N_4366,N_3510,N_3735);
or U4367 (N_4367,N_3130,N_3419);
and U4368 (N_4368,N_3433,N_3166);
xnor U4369 (N_4369,N_3744,N_3342);
and U4370 (N_4370,N_3478,N_3456);
or U4371 (N_4371,N_3298,N_3418);
or U4372 (N_4372,N_3627,N_3429);
or U4373 (N_4373,N_3371,N_3646);
xor U4374 (N_4374,N_3178,N_3276);
and U4375 (N_4375,N_3570,N_3010);
and U4376 (N_4376,N_3592,N_3018);
and U4377 (N_4377,N_3115,N_3372);
xnor U4378 (N_4378,N_3070,N_3001);
nor U4379 (N_4379,N_3059,N_3636);
nor U4380 (N_4380,N_3553,N_3304);
nand U4381 (N_4381,N_3590,N_3484);
or U4382 (N_4382,N_3189,N_3512);
and U4383 (N_4383,N_3462,N_3274);
nand U4384 (N_4384,N_3628,N_3134);
or U4385 (N_4385,N_3224,N_3268);
or U4386 (N_4386,N_3546,N_3411);
and U4387 (N_4387,N_3456,N_3301);
xnor U4388 (N_4388,N_3053,N_3024);
nor U4389 (N_4389,N_3473,N_3653);
nor U4390 (N_4390,N_3623,N_3420);
and U4391 (N_4391,N_3591,N_3571);
nor U4392 (N_4392,N_3541,N_3286);
and U4393 (N_4393,N_3176,N_3098);
or U4394 (N_4394,N_3124,N_3539);
xor U4395 (N_4395,N_3118,N_3720);
nand U4396 (N_4396,N_3272,N_3094);
or U4397 (N_4397,N_3128,N_3286);
xor U4398 (N_4398,N_3355,N_3461);
and U4399 (N_4399,N_3474,N_3562);
xor U4400 (N_4400,N_3318,N_3526);
xor U4401 (N_4401,N_3198,N_3661);
and U4402 (N_4402,N_3722,N_3505);
nor U4403 (N_4403,N_3709,N_3276);
or U4404 (N_4404,N_3292,N_3372);
nand U4405 (N_4405,N_3018,N_3500);
or U4406 (N_4406,N_3279,N_3713);
nor U4407 (N_4407,N_3326,N_3538);
or U4408 (N_4408,N_3661,N_3442);
and U4409 (N_4409,N_3242,N_3013);
nand U4410 (N_4410,N_3009,N_3017);
and U4411 (N_4411,N_3544,N_3229);
xnor U4412 (N_4412,N_3290,N_3381);
or U4413 (N_4413,N_3674,N_3587);
nor U4414 (N_4414,N_3682,N_3261);
xnor U4415 (N_4415,N_3702,N_3695);
and U4416 (N_4416,N_3219,N_3728);
and U4417 (N_4417,N_3563,N_3477);
xor U4418 (N_4418,N_3681,N_3270);
nand U4419 (N_4419,N_3431,N_3123);
or U4420 (N_4420,N_3444,N_3432);
xnor U4421 (N_4421,N_3069,N_3442);
nor U4422 (N_4422,N_3365,N_3150);
or U4423 (N_4423,N_3467,N_3153);
nand U4424 (N_4424,N_3563,N_3327);
nor U4425 (N_4425,N_3733,N_3448);
nand U4426 (N_4426,N_3470,N_3190);
nand U4427 (N_4427,N_3177,N_3681);
and U4428 (N_4428,N_3477,N_3421);
xnor U4429 (N_4429,N_3708,N_3605);
and U4430 (N_4430,N_3450,N_3683);
or U4431 (N_4431,N_3046,N_3483);
xnor U4432 (N_4432,N_3448,N_3337);
or U4433 (N_4433,N_3594,N_3338);
nor U4434 (N_4434,N_3212,N_3074);
nor U4435 (N_4435,N_3505,N_3693);
nor U4436 (N_4436,N_3577,N_3163);
and U4437 (N_4437,N_3619,N_3140);
and U4438 (N_4438,N_3332,N_3122);
and U4439 (N_4439,N_3632,N_3198);
nand U4440 (N_4440,N_3485,N_3638);
nor U4441 (N_4441,N_3446,N_3163);
xnor U4442 (N_4442,N_3463,N_3624);
nand U4443 (N_4443,N_3726,N_3240);
nand U4444 (N_4444,N_3425,N_3126);
or U4445 (N_4445,N_3064,N_3367);
and U4446 (N_4446,N_3225,N_3725);
or U4447 (N_4447,N_3563,N_3676);
or U4448 (N_4448,N_3663,N_3385);
nand U4449 (N_4449,N_3398,N_3630);
nand U4450 (N_4450,N_3574,N_3641);
xnor U4451 (N_4451,N_3597,N_3688);
nor U4452 (N_4452,N_3723,N_3467);
and U4453 (N_4453,N_3294,N_3617);
or U4454 (N_4454,N_3305,N_3139);
and U4455 (N_4455,N_3731,N_3496);
nand U4456 (N_4456,N_3103,N_3337);
nor U4457 (N_4457,N_3432,N_3495);
xor U4458 (N_4458,N_3190,N_3568);
nor U4459 (N_4459,N_3046,N_3161);
and U4460 (N_4460,N_3515,N_3465);
xor U4461 (N_4461,N_3487,N_3671);
nor U4462 (N_4462,N_3489,N_3129);
xor U4463 (N_4463,N_3142,N_3438);
nor U4464 (N_4464,N_3067,N_3617);
or U4465 (N_4465,N_3101,N_3354);
nand U4466 (N_4466,N_3184,N_3094);
xor U4467 (N_4467,N_3515,N_3473);
or U4468 (N_4468,N_3159,N_3036);
xor U4469 (N_4469,N_3457,N_3132);
nand U4470 (N_4470,N_3053,N_3009);
or U4471 (N_4471,N_3543,N_3112);
and U4472 (N_4472,N_3117,N_3313);
xnor U4473 (N_4473,N_3365,N_3377);
or U4474 (N_4474,N_3690,N_3152);
and U4475 (N_4475,N_3166,N_3559);
nand U4476 (N_4476,N_3334,N_3588);
or U4477 (N_4477,N_3720,N_3444);
xnor U4478 (N_4478,N_3280,N_3310);
and U4479 (N_4479,N_3315,N_3496);
nor U4480 (N_4480,N_3298,N_3120);
nand U4481 (N_4481,N_3112,N_3463);
nor U4482 (N_4482,N_3499,N_3077);
or U4483 (N_4483,N_3064,N_3355);
nor U4484 (N_4484,N_3635,N_3128);
xnor U4485 (N_4485,N_3218,N_3713);
or U4486 (N_4486,N_3701,N_3071);
xor U4487 (N_4487,N_3244,N_3044);
nor U4488 (N_4488,N_3120,N_3724);
nor U4489 (N_4489,N_3263,N_3266);
nor U4490 (N_4490,N_3268,N_3074);
nand U4491 (N_4491,N_3321,N_3729);
or U4492 (N_4492,N_3178,N_3401);
nor U4493 (N_4493,N_3138,N_3015);
nor U4494 (N_4494,N_3457,N_3015);
xnor U4495 (N_4495,N_3394,N_3046);
nor U4496 (N_4496,N_3307,N_3228);
xnor U4497 (N_4497,N_3448,N_3122);
or U4498 (N_4498,N_3258,N_3476);
nand U4499 (N_4499,N_3273,N_3201);
and U4500 (N_4500,N_4100,N_3865);
nand U4501 (N_4501,N_4035,N_4152);
nand U4502 (N_4502,N_4202,N_4346);
nor U4503 (N_4503,N_4066,N_4015);
or U4504 (N_4504,N_4394,N_4382);
and U4505 (N_4505,N_3833,N_4248);
and U4506 (N_4506,N_4338,N_4377);
or U4507 (N_4507,N_4411,N_4033);
and U4508 (N_4508,N_4439,N_4206);
nor U4509 (N_4509,N_3774,N_3921);
nand U4510 (N_4510,N_4457,N_4291);
and U4511 (N_4511,N_3803,N_4469);
xor U4512 (N_4512,N_4437,N_3913);
and U4513 (N_4513,N_4296,N_4478);
and U4514 (N_4514,N_4375,N_3871);
nand U4515 (N_4515,N_3794,N_4150);
xor U4516 (N_4516,N_3769,N_3973);
xnor U4517 (N_4517,N_3952,N_3999);
xor U4518 (N_4518,N_4396,N_3885);
xnor U4519 (N_4519,N_3998,N_4170);
nand U4520 (N_4520,N_3970,N_3848);
nand U4521 (N_4521,N_4371,N_4062);
xor U4522 (N_4522,N_4395,N_4246);
nand U4523 (N_4523,N_4118,N_4089);
or U4524 (N_4524,N_4332,N_4417);
nand U4525 (N_4525,N_4413,N_4078);
xnor U4526 (N_4526,N_4330,N_4186);
and U4527 (N_4527,N_3785,N_4096);
xor U4528 (N_4528,N_4091,N_4435);
nand U4529 (N_4529,N_4389,N_4086);
or U4530 (N_4530,N_4381,N_4353);
nor U4531 (N_4531,N_4260,N_4324);
and U4532 (N_4532,N_3934,N_4017);
and U4533 (N_4533,N_3975,N_3855);
and U4534 (N_4534,N_3856,N_4159);
or U4535 (N_4535,N_3840,N_4074);
xnor U4536 (N_4536,N_3897,N_4221);
nand U4537 (N_4537,N_4155,N_4300);
nor U4538 (N_4538,N_3882,N_4178);
xor U4539 (N_4539,N_4168,N_4490);
or U4540 (N_4540,N_4347,N_4426);
or U4541 (N_4541,N_3990,N_4295);
or U4542 (N_4542,N_3910,N_3839);
and U4543 (N_4543,N_4354,N_4459);
xnor U4544 (N_4544,N_4303,N_4321);
xnor U4545 (N_4545,N_4356,N_4214);
nand U4546 (N_4546,N_4323,N_4290);
nand U4547 (N_4547,N_4129,N_4320);
or U4548 (N_4548,N_4113,N_4101);
or U4549 (N_4549,N_4174,N_4053);
or U4550 (N_4550,N_4005,N_4122);
nor U4551 (N_4551,N_4414,N_3821);
and U4552 (N_4552,N_4080,N_4494);
nor U4553 (N_4553,N_3945,N_4355);
or U4554 (N_4554,N_4154,N_4238);
nor U4555 (N_4555,N_4183,N_3901);
and U4556 (N_4556,N_3877,N_3963);
nor U4557 (N_4557,N_4404,N_4376);
nor U4558 (N_4558,N_4307,N_4442);
or U4559 (N_4559,N_3888,N_3964);
and U4560 (N_4560,N_4102,N_3811);
xor U4561 (N_4561,N_3827,N_4189);
nor U4562 (N_4562,N_3971,N_4384);
nand U4563 (N_4563,N_4399,N_3889);
or U4564 (N_4564,N_4172,N_3987);
xnor U4565 (N_4565,N_3854,N_4367);
or U4566 (N_4566,N_4232,N_3908);
and U4567 (N_4567,N_4109,N_4265);
xor U4568 (N_4568,N_4099,N_4194);
nand U4569 (N_4569,N_4120,N_4054);
or U4570 (N_4570,N_4224,N_3923);
nor U4571 (N_4571,N_4107,N_3789);
nand U4572 (N_4572,N_3767,N_4406);
or U4573 (N_4573,N_3974,N_3801);
or U4574 (N_4574,N_4019,N_3866);
or U4575 (N_4575,N_4496,N_3804);
or U4576 (N_4576,N_4177,N_4464);
nor U4577 (N_4577,N_3935,N_4081);
or U4578 (N_4578,N_4234,N_4403);
nor U4579 (N_4579,N_4423,N_4402);
and U4580 (N_4580,N_4067,N_4361);
nand U4581 (N_4581,N_4002,N_4249);
or U4582 (N_4582,N_3860,N_3956);
or U4583 (N_4583,N_4216,N_4123);
xnor U4584 (N_4584,N_3850,N_4344);
and U4585 (N_4585,N_4133,N_4227);
or U4586 (N_4586,N_4491,N_3788);
xnor U4587 (N_4587,N_3916,N_4463);
nor U4588 (N_4588,N_4008,N_4124);
and U4589 (N_4589,N_4110,N_4387);
and U4590 (N_4590,N_4497,N_4313);
nor U4591 (N_4591,N_4079,N_4433);
nor U4592 (N_4592,N_3812,N_4283);
and U4593 (N_4593,N_4446,N_4372);
xor U4594 (N_4594,N_4378,N_4336);
xnor U4595 (N_4595,N_4201,N_4495);
nor U4596 (N_4596,N_4476,N_4370);
or U4597 (N_4597,N_4203,N_4340);
nand U4598 (N_4598,N_4309,N_3802);
nor U4599 (N_4599,N_4187,N_3797);
xnor U4600 (N_4600,N_3845,N_4251);
nand U4601 (N_4601,N_4266,N_3842);
nor U4602 (N_4602,N_3890,N_4195);
nand U4603 (N_4603,N_4181,N_3881);
nor U4604 (N_4604,N_3816,N_3776);
or U4605 (N_4605,N_4220,N_3787);
xnor U4606 (N_4606,N_3920,N_4032);
xor U4607 (N_4607,N_4140,N_3783);
and U4608 (N_4608,N_3817,N_4358);
nor U4609 (N_4609,N_4487,N_3924);
and U4610 (N_4610,N_4114,N_4279);
and U4611 (N_4611,N_3981,N_4072);
xor U4612 (N_4612,N_3810,N_3884);
xor U4613 (N_4613,N_3809,N_3763);
and U4614 (N_4614,N_4157,N_4176);
and U4615 (N_4615,N_3828,N_4304);
nor U4616 (N_4616,N_4134,N_4432);
nor U4617 (N_4617,N_4191,N_4341);
xnor U4618 (N_4618,N_4209,N_4185);
and U4619 (N_4619,N_4352,N_4342);
or U4620 (N_4620,N_4103,N_4012);
or U4621 (N_4621,N_3967,N_3902);
or U4622 (N_4622,N_4180,N_4379);
nor U4623 (N_4623,N_4418,N_3903);
and U4624 (N_4624,N_4470,N_3954);
or U4625 (N_4625,N_4455,N_4410);
or U4626 (N_4626,N_4294,N_4121);
nand U4627 (N_4627,N_4284,N_3800);
xnor U4628 (N_4628,N_4310,N_3868);
xor U4629 (N_4629,N_4373,N_4095);
nand U4630 (N_4630,N_3972,N_3886);
or U4631 (N_4631,N_4253,N_3823);
nor U4632 (N_4632,N_3754,N_4037);
nor U4633 (N_4633,N_3909,N_3843);
nand U4634 (N_4634,N_4151,N_3872);
nand U4635 (N_4635,N_4474,N_4024);
xor U4636 (N_4636,N_3977,N_3892);
nor U4637 (N_4637,N_3859,N_4050);
nand U4638 (N_4638,N_3777,N_4198);
nor U4639 (N_4639,N_4480,N_4473);
and U4640 (N_4640,N_3922,N_3757);
xnor U4641 (N_4641,N_4128,N_3837);
and U4642 (N_4642,N_4380,N_4302);
nor U4643 (N_4643,N_4041,N_3782);
nand U4644 (N_4644,N_3953,N_4065);
xor U4645 (N_4645,N_4275,N_3781);
or U4646 (N_4646,N_3768,N_4021);
or U4647 (N_4647,N_4475,N_4293);
xor U4648 (N_4648,N_4398,N_4166);
xnor U4649 (N_4649,N_4282,N_4038);
nand U4650 (N_4650,N_4343,N_4142);
xnor U4651 (N_4651,N_4093,N_3926);
nand U4652 (N_4652,N_3969,N_4222);
nor U4653 (N_4653,N_3948,N_3805);
or U4654 (N_4654,N_4499,N_4044);
and U4655 (N_4655,N_3899,N_3978);
nor U4656 (N_4656,N_3820,N_3991);
and U4657 (N_4657,N_3929,N_3876);
xor U4658 (N_4658,N_4141,N_3771);
nor U4659 (N_4659,N_4368,N_3799);
or U4660 (N_4660,N_4472,N_3928);
xnor U4661 (N_4661,N_3786,N_4374);
xnor U4662 (N_4662,N_3944,N_4448);
or U4663 (N_4663,N_4068,N_3939);
nor U4664 (N_4664,N_4301,N_4257);
nand U4665 (N_4665,N_3949,N_4467);
or U4666 (N_4666,N_4034,N_4058);
or U4667 (N_4667,N_4173,N_4261);
and U4668 (N_4668,N_4149,N_4167);
and U4669 (N_4669,N_4441,N_4126);
nand U4670 (N_4670,N_3792,N_4022);
xor U4671 (N_4671,N_4011,N_3942);
nand U4672 (N_4672,N_4366,N_4390);
nand U4673 (N_4673,N_4046,N_4468);
or U4674 (N_4674,N_4436,N_4327);
and U4675 (N_4675,N_4077,N_4461);
or U4676 (N_4676,N_4083,N_4042);
nor U4677 (N_4677,N_3806,N_4229);
or U4678 (N_4678,N_3849,N_3857);
nor U4679 (N_4679,N_4345,N_4292);
and U4680 (N_4680,N_4444,N_4429);
nand U4681 (N_4681,N_4447,N_3793);
and U4682 (N_4682,N_4485,N_3822);
nand U4683 (N_4683,N_3951,N_3994);
nor U4684 (N_4684,N_3755,N_3915);
nand U4685 (N_4685,N_4088,N_3958);
xor U4686 (N_4686,N_4269,N_4409);
nor U4687 (N_4687,N_3966,N_3895);
and U4688 (N_4688,N_4277,N_4287);
nand U4689 (N_4689,N_4393,N_4138);
and U4690 (N_4690,N_4148,N_4351);
nand U4691 (N_4691,N_4207,N_4252);
or U4692 (N_4692,N_4049,N_3959);
and U4693 (N_4693,N_4117,N_3982);
or U4694 (N_4694,N_3904,N_4223);
nand U4695 (N_4695,N_4348,N_4235);
or U4696 (N_4696,N_4482,N_4061);
xor U4697 (N_4697,N_3984,N_4000);
or U4698 (N_4698,N_4001,N_4360);
xnor U4699 (N_4699,N_4274,N_3780);
or U4700 (N_4700,N_3818,N_3896);
nand U4701 (N_4701,N_4225,N_4272);
nor U4702 (N_4702,N_3983,N_3878);
xor U4703 (N_4703,N_4190,N_3838);
or U4704 (N_4704,N_4306,N_3830);
nand U4705 (N_4705,N_4145,N_4127);
nor U4706 (N_4706,N_3778,N_4048);
and U4707 (N_4707,N_4416,N_4014);
and U4708 (N_4708,N_3869,N_3879);
xor U4709 (N_4709,N_4483,N_3927);
nor U4710 (N_4710,N_3918,N_4314);
xnor U4711 (N_4711,N_4239,N_3796);
or U4712 (N_4712,N_4132,N_3940);
or U4713 (N_4713,N_3961,N_4493);
nand U4714 (N_4714,N_4450,N_4026);
and U4715 (N_4715,N_4419,N_4299);
nor U4716 (N_4716,N_3996,N_3824);
xor U4717 (N_4717,N_3965,N_4215);
and U4718 (N_4718,N_3985,N_4449);
nand U4719 (N_4719,N_4063,N_3751);
nor U4720 (N_4720,N_4060,N_4454);
nor U4721 (N_4721,N_3989,N_3853);
and U4722 (N_4722,N_3773,N_3852);
nor U4723 (N_4723,N_4161,N_3914);
nand U4724 (N_4724,N_4388,N_4137);
nor U4725 (N_4725,N_3766,N_3832);
nor U4726 (N_4726,N_4339,N_4421);
nor U4727 (N_4727,N_4059,N_3846);
and U4728 (N_4728,N_4064,N_4247);
nand U4729 (N_4729,N_4465,N_4076);
or U4730 (N_4730,N_3941,N_4164);
nor U4731 (N_4731,N_3867,N_3863);
nor U4732 (N_4732,N_4385,N_4407);
nand U4733 (N_4733,N_3932,N_4263);
nor U4734 (N_4734,N_4090,N_3988);
xnor U4735 (N_4735,N_4092,N_4255);
nor U4736 (N_4736,N_4028,N_3947);
nor U4737 (N_4737,N_4318,N_4010);
nor U4738 (N_4738,N_4007,N_4193);
nor U4739 (N_4739,N_4219,N_3912);
nand U4740 (N_4740,N_4097,N_4075);
nand U4741 (N_4741,N_3992,N_4040);
and U4742 (N_4742,N_3825,N_4271);
xor U4743 (N_4743,N_4245,N_4428);
nor U4744 (N_4744,N_4315,N_4213);
or U4745 (N_4745,N_4452,N_4392);
and U4746 (N_4746,N_4211,N_4242);
nand U4747 (N_4747,N_4451,N_4111);
nand U4748 (N_4748,N_4184,N_3874);
and U4749 (N_4749,N_3829,N_4051);
nor U4750 (N_4750,N_4333,N_3772);
and U4751 (N_4751,N_3936,N_4073);
or U4752 (N_4752,N_3887,N_4427);
or U4753 (N_4753,N_4188,N_4036);
and U4754 (N_4754,N_3957,N_3814);
nand U4755 (N_4755,N_3993,N_3834);
and U4756 (N_4756,N_4175,N_3925);
nand U4757 (N_4757,N_3795,N_4130);
xnor U4758 (N_4758,N_4391,N_4350);
and U4759 (N_4759,N_3898,N_3960);
nor U4760 (N_4760,N_3907,N_4278);
nand U4761 (N_4761,N_4230,N_3819);
xor U4762 (N_4762,N_4316,N_4143);
nor U4763 (N_4763,N_4329,N_3919);
or U4764 (N_4764,N_4105,N_4259);
nor U4765 (N_4765,N_4025,N_3791);
or U4766 (N_4766,N_4045,N_3826);
nor U4767 (N_4767,N_4481,N_3986);
nor U4768 (N_4768,N_3761,N_4359);
nor U4769 (N_4769,N_4453,N_4244);
and U4770 (N_4770,N_4362,N_4094);
and U4771 (N_4771,N_3862,N_4285);
and U4772 (N_4772,N_4386,N_3851);
xnor U4773 (N_4773,N_4165,N_4276);
and U4774 (N_4774,N_4228,N_4240);
and U4775 (N_4775,N_4205,N_4196);
xnor U4776 (N_4776,N_4013,N_4163);
and U4777 (N_4777,N_4136,N_4311);
or U4778 (N_4778,N_3893,N_4357);
and U4779 (N_4779,N_4256,N_4322);
or U4780 (N_4780,N_4312,N_3784);
nand U4781 (N_4781,N_4069,N_4270);
xor U4782 (N_4782,N_4331,N_4115);
nand U4783 (N_4783,N_3880,N_4200);
nand U4784 (N_4784,N_4484,N_4489);
nor U4785 (N_4785,N_4273,N_4006);
or U4786 (N_4786,N_4208,N_3765);
nor U4787 (N_4787,N_4082,N_3758);
nor U4788 (N_4788,N_4231,N_3938);
nand U4789 (N_4789,N_4139,N_4363);
nor U4790 (N_4790,N_4262,N_4456);
xor U4791 (N_4791,N_4243,N_4488);
or U4792 (N_4792,N_4365,N_3753);
xnor U4793 (N_4793,N_4158,N_4317);
nand U4794 (N_4794,N_4405,N_4305);
and U4795 (N_4795,N_4422,N_4197);
or U4796 (N_4796,N_4460,N_4003);
and U4797 (N_4797,N_3813,N_4281);
nor U4798 (N_4798,N_3955,N_3917);
or U4799 (N_4799,N_4171,N_3980);
xor U4800 (N_4800,N_4412,N_4018);
xnor U4801 (N_4801,N_4280,N_3775);
xnor U4802 (N_4802,N_3808,N_3807);
xnor U4803 (N_4803,N_3798,N_4369);
and U4804 (N_4804,N_4334,N_3979);
nor U4805 (N_4805,N_4264,N_4179);
xnor U4806 (N_4806,N_4135,N_3883);
and U4807 (N_4807,N_4267,N_3762);
nor U4808 (N_4808,N_4192,N_3759);
xnor U4809 (N_4809,N_4288,N_4182);
nand U4810 (N_4810,N_4098,N_4349);
nand U4811 (N_4811,N_4431,N_4400);
xor U4812 (N_4812,N_4218,N_3937);
and U4813 (N_4813,N_4210,N_3844);
xnor U4814 (N_4814,N_4029,N_4112);
xor U4815 (N_4815,N_4438,N_3875);
and U4816 (N_4816,N_3946,N_4057);
and U4817 (N_4817,N_4087,N_4108);
xnor U4818 (N_4818,N_3756,N_3861);
or U4819 (N_4819,N_3906,N_4116);
xnor U4820 (N_4820,N_3760,N_3815);
xnor U4821 (N_4821,N_3750,N_4401);
nand U4822 (N_4822,N_4415,N_4047);
xor U4823 (N_4823,N_4425,N_3931);
xnor U4824 (N_4824,N_4477,N_4268);
and U4825 (N_4825,N_3858,N_4420);
or U4826 (N_4826,N_4237,N_4297);
or U4827 (N_4827,N_3841,N_3911);
xor U4828 (N_4828,N_4030,N_4325);
or U4829 (N_4829,N_4479,N_4217);
xor U4830 (N_4830,N_3770,N_4408);
nand U4831 (N_4831,N_3836,N_4199);
nand U4832 (N_4832,N_4212,N_4462);
nor U4833 (N_4833,N_4434,N_4052);
and U4834 (N_4834,N_4430,N_4043);
nand U4835 (N_4835,N_4085,N_3891);
nor U4836 (N_4836,N_4498,N_4055);
nor U4837 (N_4837,N_4492,N_4308);
xnor U4838 (N_4838,N_3930,N_4236);
nor U4839 (N_4839,N_4337,N_4233);
nand U4840 (N_4840,N_4286,N_3997);
nand U4841 (N_4841,N_4250,N_3847);
or U4842 (N_4842,N_4466,N_3950);
nand U4843 (N_4843,N_4471,N_4004);
nor U4844 (N_4844,N_3779,N_3864);
and U4845 (N_4845,N_4119,N_3831);
and U4846 (N_4846,N_4146,N_4131);
xnor U4847 (N_4847,N_4027,N_3764);
nand U4848 (N_4848,N_4147,N_4023);
and U4849 (N_4849,N_4169,N_3870);
nor U4850 (N_4850,N_4397,N_4056);
nor U4851 (N_4851,N_3894,N_4445);
and U4852 (N_4852,N_3873,N_3790);
and U4853 (N_4853,N_4016,N_3968);
nand U4854 (N_4854,N_4226,N_3900);
xnor U4855 (N_4855,N_3943,N_4424);
xnor U4856 (N_4856,N_4104,N_4084);
or U4857 (N_4857,N_4326,N_4298);
and U4858 (N_4858,N_4335,N_4458);
xor U4859 (N_4859,N_4039,N_4486);
and U4860 (N_4860,N_4319,N_4144);
nand U4861 (N_4861,N_4328,N_4071);
nor U4862 (N_4862,N_4254,N_4160);
xnor U4863 (N_4863,N_4153,N_4440);
nand U4864 (N_4864,N_4031,N_4364);
xnor U4865 (N_4865,N_4258,N_4070);
nor U4866 (N_4866,N_3976,N_4009);
and U4867 (N_4867,N_3752,N_3962);
nand U4868 (N_4868,N_4289,N_4125);
xnor U4869 (N_4869,N_4204,N_3933);
or U4870 (N_4870,N_4443,N_4156);
nand U4871 (N_4871,N_4020,N_4106);
or U4872 (N_4872,N_3995,N_4241);
and U4873 (N_4873,N_4383,N_3905);
xor U4874 (N_4874,N_3835,N_4162);
and U4875 (N_4875,N_4078,N_4287);
nor U4876 (N_4876,N_3769,N_3927);
and U4877 (N_4877,N_4230,N_4165);
or U4878 (N_4878,N_3937,N_4418);
nand U4879 (N_4879,N_4071,N_4237);
or U4880 (N_4880,N_4215,N_3784);
nor U4881 (N_4881,N_4161,N_3753);
nand U4882 (N_4882,N_4177,N_3977);
or U4883 (N_4883,N_4066,N_3928);
or U4884 (N_4884,N_3878,N_4093);
xor U4885 (N_4885,N_4469,N_4050);
or U4886 (N_4886,N_4127,N_3780);
nor U4887 (N_4887,N_4150,N_4124);
or U4888 (N_4888,N_4136,N_4330);
or U4889 (N_4889,N_4060,N_4370);
and U4890 (N_4890,N_4344,N_3947);
nor U4891 (N_4891,N_3828,N_3993);
or U4892 (N_4892,N_4237,N_3876);
or U4893 (N_4893,N_3906,N_4160);
and U4894 (N_4894,N_4487,N_4107);
nand U4895 (N_4895,N_3960,N_3951);
nand U4896 (N_4896,N_4237,N_4466);
and U4897 (N_4897,N_3929,N_3775);
or U4898 (N_4898,N_3884,N_4474);
nor U4899 (N_4899,N_3867,N_4252);
and U4900 (N_4900,N_4314,N_3763);
xnor U4901 (N_4901,N_4472,N_4211);
nand U4902 (N_4902,N_4251,N_4256);
or U4903 (N_4903,N_4138,N_3770);
xnor U4904 (N_4904,N_4475,N_4252);
nor U4905 (N_4905,N_4004,N_3806);
nor U4906 (N_4906,N_4211,N_4117);
or U4907 (N_4907,N_4171,N_3849);
and U4908 (N_4908,N_4142,N_4226);
nor U4909 (N_4909,N_4158,N_4474);
or U4910 (N_4910,N_3884,N_4486);
or U4911 (N_4911,N_4026,N_4286);
and U4912 (N_4912,N_4317,N_4030);
xor U4913 (N_4913,N_3763,N_4397);
nand U4914 (N_4914,N_4368,N_4200);
nor U4915 (N_4915,N_3986,N_4100);
nor U4916 (N_4916,N_4087,N_3758);
and U4917 (N_4917,N_4295,N_4411);
nor U4918 (N_4918,N_4107,N_4338);
and U4919 (N_4919,N_4030,N_4456);
nor U4920 (N_4920,N_4067,N_3924);
nor U4921 (N_4921,N_4042,N_4125);
nand U4922 (N_4922,N_3786,N_4075);
nand U4923 (N_4923,N_4088,N_3864);
xor U4924 (N_4924,N_4092,N_4366);
and U4925 (N_4925,N_3957,N_4311);
xor U4926 (N_4926,N_3779,N_4177);
nor U4927 (N_4927,N_4118,N_3823);
xnor U4928 (N_4928,N_3753,N_4415);
xor U4929 (N_4929,N_4429,N_4383);
and U4930 (N_4930,N_4452,N_4362);
or U4931 (N_4931,N_4377,N_4462);
and U4932 (N_4932,N_4177,N_3927);
xnor U4933 (N_4933,N_4246,N_4260);
nor U4934 (N_4934,N_3984,N_4094);
or U4935 (N_4935,N_3770,N_4302);
and U4936 (N_4936,N_4338,N_3915);
nor U4937 (N_4937,N_4189,N_4275);
nand U4938 (N_4938,N_3799,N_3921);
xnor U4939 (N_4939,N_4017,N_3800);
nor U4940 (N_4940,N_3950,N_4155);
and U4941 (N_4941,N_3750,N_4356);
nor U4942 (N_4942,N_3914,N_3930);
xnor U4943 (N_4943,N_3891,N_4268);
or U4944 (N_4944,N_4079,N_4458);
or U4945 (N_4945,N_4416,N_3888);
or U4946 (N_4946,N_4297,N_4296);
or U4947 (N_4947,N_3761,N_4229);
or U4948 (N_4948,N_4227,N_3881);
and U4949 (N_4949,N_4482,N_4324);
and U4950 (N_4950,N_4063,N_4413);
and U4951 (N_4951,N_3862,N_3854);
or U4952 (N_4952,N_4079,N_4160);
xor U4953 (N_4953,N_3780,N_4363);
xnor U4954 (N_4954,N_3764,N_4192);
or U4955 (N_4955,N_4367,N_3841);
xor U4956 (N_4956,N_4393,N_4383);
or U4957 (N_4957,N_3992,N_3888);
nor U4958 (N_4958,N_3844,N_3791);
or U4959 (N_4959,N_4327,N_4032);
and U4960 (N_4960,N_3941,N_3764);
nor U4961 (N_4961,N_3766,N_4497);
or U4962 (N_4962,N_4188,N_4148);
xnor U4963 (N_4963,N_3778,N_4451);
nor U4964 (N_4964,N_4322,N_3867);
and U4965 (N_4965,N_3963,N_4107);
xor U4966 (N_4966,N_4349,N_3865);
or U4967 (N_4967,N_4347,N_4131);
xnor U4968 (N_4968,N_4167,N_4341);
and U4969 (N_4969,N_3926,N_3822);
nor U4970 (N_4970,N_3872,N_3759);
nor U4971 (N_4971,N_4039,N_3924);
and U4972 (N_4972,N_4172,N_4392);
xor U4973 (N_4973,N_4396,N_4221);
and U4974 (N_4974,N_4123,N_4159);
or U4975 (N_4975,N_4442,N_4489);
nand U4976 (N_4976,N_4148,N_4158);
xnor U4977 (N_4977,N_4059,N_4000);
nand U4978 (N_4978,N_3867,N_4345);
and U4979 (N_4979,N_3957,N_4101);
and U4980 (N_4980,N_3946,N_4389);
nor U4981 (N_4981,N_3770,N_3847);
nand U4982 (N_4982,N_4207,N_4483);
xnor U4983 (N_4983,N_4189,N_3877);
or U4984 (N_4984,N_4404,N_4457);
or U4985 (N_4985,N_4083,N_4491);
nor U4986 (N_4986,N_4158,N_4335);
and U4987 (N_4987,N_4494,N_4251);
nand U4988 (N_4988,N_4180,N_3881);
and U4989 (N_4989,N_3905,N_4186);
or U4990 (N_4990,N_4413,N_3809);
nor U4991 (N_4991,N_4274,N_4052);
or U4992 (N_4992,N_4225,N_4140);
xnor U4993 (N_4993,N_4097,N_4021);
xnor U4994 (N_4994,N_4014,N_4288);
or U4995 (N_4995,N_3822,N_4293);
nor U4996 (N_4996,N_3770,N_3915);
xor U4997 (N_4997,N_4218,N_3999);
nor U4998 (N_4998,N_3890,N_4335);
and U4999 (N_4999,N_4205,N_4013);
nand U5000 (N_5000,N_3990,N_4409);
and U5001 (N_5001,N_4472,N_4413);
nor U5002 (N_5002,N_3982,N_4482);
nor U5003 (N_5003,N_4231,N_4102);
nor U5004 (N_5004,N_3803,N_4098);
or U5005 (N_5005,N_4035,N_3786);
and U5006 (N_5006,N_4007,N_4126);
and U5007 (N_5007,N_3751,N_4134);
or U5008 (N_5008,N_3783,N_4278);
xor U5009 (N_5009,N_4232,N_4337);
xnor U5010 (N_5010,N_4415,N_4241);
nor U5011 (N_5011,N_4401,N_4185);
and U5012 (N_5012,N_4173,N_4013);
xnor U5013 (N_5013,N_3842,N_4040);
xnor U5014 (N_5014,N_4229,N_4017);
and U5015 (N_5015,N_3837,N_4440);
nor U5016 (N_5016,N_4100,N_3872);
or U5017 (N_5017,N_4413,N_4409);
and U5018 (N_5018,N_4243,N_4366);
xnor U5019 (N_5019,N_4007,N_3794);
nand U5020 (N_5020,N_3804,N_4260);
nor U5021 (N_5021,N_3765,N_4226);
and U5022 (N_5022,N_4174,N_4325);
nand U5023 (N_5023,N_4046,N_4454);
and U5024 (N_5024,N_4457,N_3931);
xnor U5025 (N_5025,N_3823,N_4073);
nand U5026 (N_5026,N_4466,N_4322);
or U5027 (N_5027,N_4409,N_3948);
or U5028 (N_5028,N_3960,N_4317);
nor U5029 (N_5029,N_3794,N_4448);
or U5030 (N_5030,N_3909,N_4067);
nand U5031 (N_5031,N_3895,N_4099);
or U5032 (N_5032,N_4433,N_4105);
xnor U5033 (N_5033,N_3884,N_4216);
xor U5034 (N_5034,N_4044,N_3779);
nand U5035 (N_5035,N_3858,N_4204);
and U5036 (N_5036,N_3913,N_4174);
xor U5037 (N_5037,N_4374,N_3926);
and U5038 (N_5038,N_4442,N_4472);
or U5039 (N_5039,N_3800,N_4041);
xnor U5040 (N_5040,N_4304,N_3872);
and U5041 (N_5041,N_4042,N_3997);
and U5042 (N_5042,N_4441,N_4311);
and U5043 (N_5043,N_4168,N_4039);
or U5044 (N_5044,N_4151,N_3813);
xor U5045 (N_5045,N_3757,N_4089);
nor U5046 (N_5046,N_4490,N_3892);
nand U5047 (N_5047,N_4282,N_3791);
or U5048 (N_5048,N_4087,N_3790);
and U5049 (N_5049,N_3848,N_3950);
and U5050 (N_5050,N_3774,N_4076);
and U5051 (N_5051,N_4319,N_4068);
xnor U5052 (N_5052,N_4458,N_3750);
or U5053 (N_5053,N_4284,N_3936);
and U5054 (N_5054,N_4169,N_4366);
and U5055 (N_5055,N_4025,N_3847);
and U5056 (N_5056,N_4437,N_4230);
xor U5057 (N_5057,N_3958,N_3887);
nor U5058 (N_5058,N_4236,N_3806);
and U5059 (N_5059,N_3928,N_4179);
or U5060 (N_5060,N_3750,N_4267);
or U5061 (N_5061,N_4114,N_4455);
and U5062 (N_5062,N_4444,N_4024);
nand U5063 (N_5063,N_3950,N_4126);
or U5064 (N_5064,N_4103,N_3751);
xnor U5065 (N_5065,N_3871,N_4302);
nand U5066 (N_5066,N_4041,N_4158);
and U5067 (N_5067,N_3958,N_4261);
and U5068 (N_5068,N_4202,N_3842);
xor U5069 (N_5069,N_3863,N_4059);
nor U5070 (N_5070,N_3879,N_3867);
xor U5071 (N_5071,N_3773,N_4267);
xnor U5072 (N_5072,N_3918,N_3776);
xnor U5073 (N_5073,N_3938,N_4056);
or U5074 (N_5074,N_4073,N_4225);
or U5075 (N_5075,N_3961,N_4457);
or U5076 (N_5076,N_4122,N_4421);
or U5077 (N_5077,N_4465,N_3939);
or U5078 (N_5078,N_4176,N_4170);
nor U5079 (N_5079,N_4179,N_4352);
and U5080 (N_5080,N_4057,N_4468);
or U5081 (N_5081,N_3960,N_3933);
xnor U5082 (N_5082,N_4223,N_4471);
nand U5083 (N_5083,N_4374,N_4278);
or U5084 (N_5084,N_4359,N_4056);
and U5085 (N_5085,N_4370,N_4435);
nand U5086 (N_5086,N_3893,N_4384);
xnor U5087 (N_5087,N_4374,N_4000);
nand U5088 (N_5088,N_4442,N_4339);
or U5089 (N_5089,N_4104,N_4018);
nor U5090 (N_5090,N_4053,N_4292);
or U5091 (N_5091,N_4402,N_3935);
xnor U5092 (N_5092,N_4208,N_4043);
nand U5093 (N_5093,N_4175,N_4398);
nor U5094 (N_5094,N_4072,N_3841);
nand U5095 (N_5095,N_3818,N_4301);
xor U5096 (N_5096,N_4034,N_4409);
or U5097 (N_5097,N_3794,N_3826);
nor U5098 (N_5098,N_4033,N_3781);
nor U5099 (N_5099,N_4231,N_3811);
nor U5100 (N_5100,N_3837,N_4443);
xnor U5101 (N_5101,N_4149,N_3974);
and U5102 (N_5102,N_4391,N_3854);
or U5103 (N_5103,N_4133,N_4180);
or U5104 (N_5104,N_4204,N_4468);
nor U5105 (N_5105,N_4084,N_3859);
nand U5106 (N_5106,N_4398,N_3848);
nor U5107 (N_5107,N_4117,N_4493);
and U5108 (N_5108,N_4211,N_4495);
and U5109 (N_5109,N_3907,N_4022);
nand U5110 (N_5110,N_3911,N_4381);
or U5111 (N_5111,N_4335,N_3923);
and U5112 (N_5112,N_3829,N_4019);
nand U5113 (N_5113,N_4218,N_4280);
and U5114 (N_5114,N_3974,N_4254);
nand U5115 (N_5115,N_3848,N_3751);
nor U5116 (N_5116,N_3816,N_3759);
or U5117 (N_5117,N_4041,N_4404);
xnor U5118 (N_5118,N_4222,N_4471);
xor U5119 (N_5119,N_4076,N_4005);
and U5120 (N_5120,N_4146,N_3970);
nor U5121 (N_5121,N_4266,N_3838);
xor U5122 (N_5122,N_4140,N_4272);
nor U5123 (N_5123,N_4449,N_3902);
and U5124 (N_5124,N_3836,N_4230);
nor U5125 (N_5125,N_4329,N_4265);
or U5126 (N_5126,N_4203,N_4029);
xor U5127 (N_5127,N_3896,N_3970);
or U5128 (N_5128,N_3823,N_4481);
and U5129 (N_5129,N_3973,N_4151);
nand U5130 (N_5130,N_4385,N_4090);
or U5131 (N_5131,N_3891,N_4488);
or U5132 (N_5132,N_4040,N_3895);
nor U5133 (N_5133,N_4484,N_3838);
xnor U5134 (N_5134,N_3924,N_3970);
nor U5135 (N_5135,N_3918,N_4405);
xnor U5136 (N_5136,N_4165,N_4348);
or U5137 (N_5137,N_4368,N_4329);
xnor U5138 (N_5138,N_3920,N_4157);
and U5139 (N_5139,N_3963,N_4164);
and U5140 (N_5140,N_4339,N_3791);
or U5141 (N_5141,N_3813,N_3956);
nor U5142 (N_5142,N_3921,N_4120);
or U5143 (N_5143,N_4486,N_4041);
xnor U5144 (N_5144,N_3844,N_3777);
xor U5145 (N_5145,N_4214,N_4439);
nor U5146 (N_5146,N_3796,N_3861);
and U5147 (N_5147,N_4063,N_4254);
nand U5148 (N_5148,N_3806,N_4084);
nand U5149 (N_5149,N_4043,N_3964);
and U5150 (N_5150,N_4188,N_3854);
xnor U5151 (N_5151,N_4052,N_4019);
or U5152 (N_5152,N_4020,N_4130);
nor U5153 (N_5153,N_3898,N_3844);
and U5154 (N_5154,N_3937,N_4212);
and U5155 (N_5155,N_4229,N_3890);
xor U5156 (N_5156,N_4141,N_4405);
and U5157 (N_5157,N_4106,N_4414);
and U5158 (N_5158,N_4353,N_4023);
and U5159 (N_5159,N_3760,N_3954);
and U5160 (N_5160,N_3855,N_4071);
or U5161 (N_5161,N_4121,N_4334);
nor U5162 (N_5162,N_3937,N_3851);
xnor U5163 (N_5163,N_4468,N_4436);
nand U5164 (N_5164,N_4230,N_3999);
xor U5165 (N_5165,N_4052,N_3817);
nor U5166 (N_5166,N_4337,N_4115);
xor U5167 (N_5167,N_3810,N_4233);
or U5168 (N_5168,N_4282,N_3886);
xnor U5169 (N_5169,N_3842,N_4070);
and U5170 (N_5170,N_4035,N_4250);
or U5171 (N_5171,N_3784,N_4127);
and U5172 (N_5172,N_3988,N_4069);
and U5173 (N_5173,N_4145,N_4458);
and U5174 (N_5174,N_4146,N_4173);
and U5175 (N_5175,N_4210,N_4232);
and U5176 (N_5176,N_4467,N_3801);
or U5177 (N_5177,N_3943,N_3822);
xnor U5178 (N_5178,N_4301,N_4343);
nand U5179 (N_5179,N_3801,N_4119);
nor U5180 (N_5180,N_4013,N_4456);
nor U5181 (N_5181,N_3991,N_4196);
nand U5182 (N_5182,N_4138,N_4218);
xor U5183 (N_5183,N_3970,N_4026);
and U5184 (N_5184,N_4461,N_4431);
xor U5185 (N_5185,N_4063,N_4032);
nand U5186 (N_5186,N_3804,N_4190);
nand U5187 (N_5187,N_4141,N_4377);
and U5188 (N_5188,N_4169,N_3900);
or U5189 (N_5189,N_3890,N_4328);
or U5190 (N_5190,N_3917,N_4166);
and U5191 (N_5191,N_4469,N_4295);
xnor U5192 (N_5192,N_3971,N_4424);
xor U5193 (N_5193,N_4128,N_4371);
nor U5194 (N_5194,N_4090,N_4394);
or U5195 (N_5195,N_3984,N_4035);
or U5196 (N_5196,N_3957,N_4314);
or U5197 (N_5197,N_4176,N_4383);
xnor U5198 (N_5198,N_3751,N_4387);
or U5199 (N_5199,N_4437,N_3878);
xor U5200 (N_5200,N_3876,N_4461);
xnor U5201 (N_5201,N_4177,N_3961);
and U5202 (N_5202,N_3939,N_4142);
nor U5203 (N_5203,N_3832,N_3849);
or U5204 (N_5204,N_4069,N_4090);
nand U5205 (N_5205,N_3809,N_4339);
nor U5206 (N_5206,N_4193,N_4289);
nand U5207 (N_5207,N_3907,N_4405);
xor U5208 (N_5208,N_4290,N_4375);
nand U5209 (N_5209,N_4178,N_4031);
nand U5210 (N_5210,N_4112,N_4129);
and U5211 (N_5211,N_4166,N_4316);
and U5212 (N_5212,N_4111,N_4425);
and U5213 (N_5213,N_4492,N_3926);
or U5214 (N_5214,N_3941,N_4076);
nand U5215 (N_5215,N_4482,N_3894);
nand U5216 (N_5216,N_4355,N_3931);
or U5217 (N_5217,N_4271,N_4479);
nand U5218 (N_5218,N_4246,N_4020);
nor U5219 (N_5219,N_4090,N_4343);
and U5220 (N_5220,N_4408,N_4156);
nor U5221 (N_5221,N_3891,N_4230);
and U5222 (N_5222,N_4025,N_4482);
nor U5223 (N_5223,N_4442,N_3865);
nand U5224 (N_5224,N_4360,N_3946);
xnor U5225 (N_5225,N_4341,N_3884);
or U5226 (N_5226,N_4382,N_4381);
or U5227 (N_5227,N_4287,N_3766);
nor U5228 (N_5228,N_4083,N_4208);
and U5229 (N_5229,N_3879,N_3825);
xor U5230 (N_5230,N_4399,N_4058);
or U5231 (N_5231,N_4066,N_4291);
and U5232 (N_5232,N_4484,N_4275);
or U5233 (N_5233,N_4275,N_3838);
nor U5234 (N_5234,N_4001,N_4129);
nand U5235 (N_5235,N_3927,N_4407);
and U5236 (N_5236,N_4220,N_3941);
nor U5237 (N_5237,N_4184,N_3827);
nor U5238 (N_5238,N_3803,N_4317);
or U5239 (N_5239,N_3762,N_3816);
xor U5240 (N_5240,N_4428,N_4407);
and U5241 (N_5241,N_4277,N_3906);
or U5242 (N_5242,N_3976,N_3845);
nand U5243 (N_5243,N_4498,N_3991);
or U5244 (N_5244,N_3760,N_4362);
nor U5245 (N_5245,N_4242,N_4038);
or U5246 (N_5246,N_4235,N_4288);
nand U5247 (N_5247,N_4368,N_4165);
xnor U5248 (N_5248,N_4156,N_4453);
xor U5249 (N_5249,N_4019,N_4009);
and U5250 (N_5250,N_4953,N_4855);
and U5251 (N_5251,N_4709,N_4558);
or U5252 (N_5252,N_4889,N_4924);
nor U5253 (N_5253,N_4574,N_5091);
nor U5254 (N_5254,N_4506,N_4861);
and U5255 (N_5255,N_4962,N_4965);
nor U5256 (N_5256,N_5019,N_4579);
xor U5257 (N_5257,N_5155,N_5237);
nand U5258 (N_5258,N_4763,N_4777);
nor U5259 (N_5259,N_4616,N_4720);
xor U5260 (N_5260,N_4689,N_4987);
nand U5261 (N_5261,N_5000,N_4839);
nor U5262 (N_5262,N_4974,N_4882);
nand U5263 (N_5263,N_4698,N_5226);
xnor U5264 (N_5264,N_5097,N_4624);
or U5265 (N_5265,N_4840,N_5101);
nor U5266 (N_5266,N_4678,N_4617);
and U5267 (N_5267,N_5141,N_4576);
nor U5268 (N_5268,N_5061,N_4542);
nor U5269 (N_5269,N_5013,N_4550);
nand U5270 (N_5270,N_5190,N_5107);
or U5271 (N_5271,N_4809,N_5017);
nor U5272 (N_5272,N_4926,N_4897);
and U5273 (N_5273,N_4896,N_4937);
and U5274 (N_5274,N_4853,N_4806);
nor U5275 (N_5275,N_4780,N_5193);
nor U5276 (N_5276,N_4788,N_5129);
nor U5277 (N_5277,N_4728,N_4641);
xor U5278 (N_5278,N_5041,N_4673);
and U5279 (N_5279,N_5059,N_5029);
and U5280 (N_5280,N_4836,N_5021);
nand U5281 (N_5281,N_4925,N_4905);
or U5282 (N_5282,N_4607,N_4969);
nor U5283 (N_5283,N_4818,N_4943);
nand U5284 (N_5284,N_4612,N_4930);
xor U5285 (N_5285,N_5120,N_5229);
nand U5286 (N_5286,N_5007,N_5036);
and U5287 (N_5287,N_5157,N_4770);
or U5288 (N_5288,N_4663,N_4767);
nor U5289 (N_5289,N_4580,N_5216);
or U5290 (N_5290,N_4939,N_4980);
nor U5291 (N_5291,N_4595,N_4927);
or U5292 (N_5292,N_5067,N_5015);
and U5293 (N_5293,N_4594,N_5108);
or U5294 (N_5294,N_5242,N_5234);
or U5295 (N_5295,N_4560,N_5196);
or U5296 (N_5296,N_4998,N_4913);
nor U5297 (N_5297,N_4816,N_5240);
nor U5298 (N_5298,N_5016,N_4691);
nor U5299 (N_5299,N_4752,N_4803);
xnor U5300 (N_5300,N_5047,N_4845);
nand U5301 (N_5301,N_5056,N_4511);
nand U5302 (N_5302,N_5011,N_4584);
nor U5303 (N_5303,N_4958,N_4894);
or U5304 (N_5304,N_4512,N_4971);
nand U5305 (N_5305,N_5084,N_4810);
xor U5306 (N_5306,N_5184,N_4537);
and U5307 (N_5307,N_5124,N_4849);
and U5308 (N_5308,N_5208,N_5106);
or U5309 (N_5309,N_4835,N_4957);
xnor U5310 (N_5310,N_4976,N_4597);
nand U5311 (N_5311,N_5116,N_5055);
xor U5312 (N_5312,N_5249,N_5039);
nor U5313 (N_5313,N_5200,N_4885);
xor U5314 (N_5314,N_4898,N_5026);
nor U5315 (N_5315,N_4887,N_4961);
xnor U5316 (N_5316,N_5148,N_4539);
or U5317 (N_5317,N_4640,N_4915);
or U5318 (N_5318,N_4750,N_4815);
nor U5319 (N_5319,N_4546,N_5113);
and U5320 (N_5320,N_5149,N_4644);
xnor U5321 (N_5321,N_4572,N_4951);
xor U5322 (N_5322,N_5225,N_5128);
nand U5323 (N_5323,N_4982,N_4592);
or U5324 (N_5324,N_4578,N_4726);
and U5325 (N_5325,N_4547,N_4510);
nand U5326 (N_5326,N_5075,N_5009);
and U5327 (N_5327,N_4602,N_4825);
and U5328 (N_5328,N_4970,N_4633);
or U5329 (N_5329,N_4844,N_4850);
xor U5330 (N_5330,N_5144,N_4710);
or U5331 (N_5331,N_4636,N_4846);
nand U5332 (N_5332,N_5146,N_4817);
xnor U5333 (N_5333,N_4757,N_4876);
xnor U5334 (N_5334,N_4877,N_5025);
or U5335 (N_5335,N_5086,N_4901);
and U5336 (N_5336,N_5223,N_4851);
nand U5337 (N_5337,N_4609,N_4591);
xor U5338 (N_5338,N_4541,N_4860);
xnor U5339 (N_5339,N_4766,N_5058);
xor U5340 (N_5340,N_4833,N_4517);
nor U5341 (N_5341,N_5005,N_4749);
xnor U5342 (N_5342,N_5048,N_5188);
xnor U5343 (N_5343,N_5186,N_4929);
xnor U5344 (N_5344,N_4518,N_4563);
and U5345 (N_5345,N_5241,N_4588);
xnor U5346 (N_5346,N_4956,N_5228);
or U5347 (N_5347,N_4813,N_4514);
xnor U5348 (N_5348,N_4694,N_4559);
or U5349 (N_5349,N_5032,N_4564);
nand U5350 (N_5350,N_5217,N_4964);
xnor U5351 (N_5351,N_5177,N_4590);
and U5352 (N_5352,N_4676,N_4714);
xnor U5353 (N_5353,N_4758,N_5053);
or U5354 (N_5354,N_4683,N_4543);
nand U5355 (N_5355,N_5050,N_4865);
and U5356 (N_5356,N_4508,N_4827);
xor U5357 (N_5357,N_5100,N_5233);
nand U5358 (N_5358,N_4988,N_5038);
nor U5359 (N_5359,N_4808,N_5137);
or U5360 (N_5360,N_4565,N_4880);
nand U5361 (N_5361,N_4776,N_5165);
nor U5362 (N_5362,N_5199,N_5248);
nor U5363 (N_5363,N_5238,N_5060);
and U5364 (N_5364,N_4661,N_5081);
xnor U5365 (N_5365,N_4871,N_4621);
xor U5366 (N_5366,N_4613,N_4812);
nor U5367 (N_5367,N_4682,N_5030);
or U5368 (N_5368,N_4799,N_4742);
nand U5369 (N_5369,N_5201,N_4669);
nand U5370 (N_5370,N_4679,N_5145);
nand U5371 (N_5371,N_4891,N_4955);
nand U5372 (N_5372,N_4606,N_5161);
nor U5373 (N_5373,N_4945,N_4680);
nand U5374 (N_5374,N_4746,N_4549);
nor U5375 (N_5375,N_4522,N_4843);
nand U5376 (N_5376,N_5246,N_4646);
or U5377 (N_5377,N_4852,N_4700);
xnor U5378 (N_5378,N_4823,N_5134);
nor U5379 (N_5379,N_5002,N_4548);
nand U5380 (N_5380,N_4762,N_4906);
xnor U5381 (N_5381,N_4918,N_5087);
xor U5382 (N_5382,N_4703,N_4977);
or U5383 (N_5383,N_4736,N_4931);
or U5384 (N_5384,N_5118,N_5189);
or U5385 (N_5385,N_4890,N_4536);
and U5386 (N_5386,N_4625,N_5232);
nand U5387 (N_5387,N_4618,N_4715);
or U5388 (N_5388,N_5221,N_4768);
xor U5389 (N_5389,N_4996,N_4598);
or U5390 (N_5390,N_5173,N_4793);
and U5391 (N_5391,N_4527,N_5207);
nor U5392 (N_5392,N_4556,N_4596);
nor U5393 (N_5393,N_4902,N_4893);
nand U5394 (N_5394,N_5230,N_4960);
and U5395 (N_5395,N_5150,N_5172);
nor U5396 (N_5396,N_5180,N_5136);
nor U5397 (N_5397,N_5210,N_4687);
or U5398 (N_5398,N_4681,N_5044);
nand U5399 (N_5399,N_5235,N_4668);
nand U5400 (N_5400,N_5244,N_5219);
xor U5401 (N_5401,N_4630,N_4791);
or U5402 (N_5402,N_4677,N_5057);
or U5403 (N_5403,N_5010,N_4652);
nand U5404 (N_5404,N_4811,N_5103);
nor U5405 (N_5405,N_4684,N_5072);
and U5406 (N_5406,N_5176,N_5153);
nor U5407 (N_5407,N_4944,N_4520);
or U5408 (N_5408,N_5159,N_4557);
or U5409 (N_5409,N_5117,N_4582);
or U5410 (N_5410,N_5212,N_5227);
xnor U5411 (N_5411,N_4761,N_5215);
nor U5412 (N_5412,N_5003,N_4695);
or U5413 (N_5413,N_4690,N_4631);
nand U5414 (N_5414,N_5195,N_5096);
nand U5415 (N_5415,N_5224,N_4748);
or U5416 (N_5416,N_4783,N_4935);
xnor U5417 (N_5417,N_5236,N_4718);
nand U5418 (N_5418,N_4934,N_4722);
or U5419 (N_5419,N_4528,N_4516);
nor U5420 (N_5420,N_5183,N_4747);
or U5421 (N_5421,N_4830,N_4721);
nand U5422 (N_5422,N_5079,N_5122);
nand U5423 (N_5423,N_4858,N_4587);
or U5424 (N_5424,N_4525,N_4910);
or U5425 (N_5425,N_4983,N_5066);
and U5426 (N_5426,N_4706,N_5247);
and U5427 (N_5427,N_4637,N_5074);
nand U5428 (N_5428,N_4868,N_4660);
and U5429 (N_5429,N_5191,N_5119);
and U5430 (N_5430,N_4778,N_5004);
and U5431 (N_5431,N_4735,N_5023);
nand U5432 (N_5432,N_4814,N_4538);
nand U5433 (N_5433,N_5008,N_4928);
or U5434 (N_5434,N_5109,N_4568);
nor U5435 (N_5435,N_5206,N_4821);
nor U5436 (N_5436,N_5064,N_4664);
xnor U5437 (N_5437,N_5063,N_4730);
xor U5438 (N_5438,N_4738,N_4649);
nand U5439 (N_5439,N_4501,N_5139);
xor U5440 (N_5440,N_5218,N_4942);
nor U5441 (N_5441,N_5104,N_4966);
or U5442 (N_5442,N_4686,N_4984);
nor U5443 (N_5443,N_4632,N_4604);
xor U5444 (N_5444,N_4719,N_5222);
or U5445 (N_5445,N_5166,N_4696);
nand U5446 (N_5446,N_4507,N_4530);
or U5447 (N_5447,N_4932,N_4751);
xnor U5448 (N_5448,N_4754,N_5178);
nor U5449 (N_5449,N_4713,N_4771);
nor U5450 (N_5450,N_4899,N_4645);
nor U5451 (N_5451,N_4653,N_4985);
nand U5452 (N_5452,N_4992,N_5174);
and U5453 (N_5453,N_4724,N_4544);
xor U5454 (N_5454,N_4941,N_4567);
nor U5455 (N_5455,N_4732,N_4659);
nand U5456 (N_5456,N_4794,N_5088);
and U5457 (N_5457,N_4699,N_4531);
xnor U5458 (N_5458,N_5220,N_4864);
xor U5459 (N_5459,N_4500,N_4975);
nor U5460 (N_5460,N_4725,N_4755);
and U5461 (N_5461,N_5147,N_4600);
and U5462 (N_5462,N_4523,N_4873);
or U5463 (N_5463,N_4716,N_4671);
nor U5464 (N_5464,N_4781,N_5167);
nor U5465 (N_5465,N_4705,N_4667);
and U5466 (N_5466,N_4634,N_4765);
and U5467 (N_5467,N_4727,N_5018);
nor U5468 (N_5468,N_4981,N_4862);
nand U5469 (N_5469,N_4672,N_4739);
nand U5470 (N_5470,N_4842,N_5115);
nor U5471 (N_5471,N_4949,N_4533);
nor U5472 (N_5472,N_4648,N_5132);
and U5473 (N_5473,N_5027,N_4570);
and U5474 (N_5474,N_5049,N_4702);
nand U5475 (N_5475,N_5090,N_4911);
or U5476 (N_5476,N_4874,N_5205);
or U5477 (N_5477,N_4697,N_4787);
nand U5478 (N_5478,N_4968,N_5089);
xnor U5479 (N_5479,N_4566,N_5182);
or U5480 (N_5480,N_4756,N_4764);
xor U5481 (N_5481,N_4581,N_4622);
nand U5482 (N_5482,N_5211,N_4888);
or U5483 (N_5483,N_4909,N_5214);
nand U5484 (N_5484,N_5133,N_4804);
nand U5485 (N_5485,N_5065,N_4993);
xnor U5486 (N_5486,N_4784,N_5245);
and U5487 (N_5487,N_5187,N_4513);
nand U5488 (N_5488,N_4740,N_5168);
nand U5489 (N_5489,N_5231,N_4805);
nand U5490 (N_5490,N_4774,N_4922);
xor U5491 (N_5491,N_5105,N_4800);
nor U5492 (N_5492,N_4963,N_5158);
and U5493 (N_5493,N_5121,N_4997);
nor U5494 (N_5494,N_4526,N_5152);
nand U5495 (N_5495,N_5082,N_4940);
nor U5496 (N_5496,N_4524,N_4674);
nand U5497 (N_5497,N_5125,N_4995);
nor U5498 (N_5498,N_4731,N_4773);
or U5499 (N_5499,N_4647,N_4532);
nor U5500 (N_5500,N_5024,N_4665);
or U5501 (N_5501,N_4886,N_4881);
and U5502 (N_5502,N_4838,N_4837);
nor U5503 (N_5503,N_5111,N_5154);
or U5504 (N_5504,N_5164,N_4701);
nand U5505 (N_5505,N_4847,N_5102);
xnor U5506 (N_5506,N_4519,N_4503);
or U5507 (N_5507,N_4900,N_5012);
or U5508 (N_5508,N_4610,N_4743);
and U5509 (N_5509,N_4662,N_5006);
and U5510 (N_5510,N_4575,N_4947);
or U5511 (N_5511,N_4895,N_5123);
and U5512 (N_5512,N_4552,N_5098);
or U5513 (N_5513,N_4952,N_4651);
nand U5514 (N_5514,N_5020,N_5179);
or U5515 (N_5515,N_5204,N_5209);
nor U5516 (N_5516,N_5143,N_4919);
or U5517 (N_5517,N_4638,N_4903);
or U5518 (N_5518,N_4994,N_4920);
nand U5519 (N_5519,N_4571,N_5068);
nand U5520 (N_5520,N_4535,N_4848);
nand U5521 (N_5521,N_5151,N_4789);
nor U5522 (N_5522,N_4655,N_4569);
nand U5523 (N_5523,N_5110,N_4628);
xnor U5524 (N_5524,N_5046,N_4619);
nand U5525 (N_5525,N_4946,N_4834);
xnor U5526 (N_5526,N_5052,N_5138);
and U5527 (N_5527,N_4938,N_4807);
xnor U5528 (N_5528,N_4870,N_5175);
nand U5529 (N_5529,N_5043,N_4561);
nor U5530 (N_5530,N_4635,N_4769);
xor U5531 (N_5531,N_4658,N_4795);
or U5532 (N_5532,N_4967,N_4933);
xor U5533 (N_5533,N_5156,N_4954);
xnor U5534 (N_5534,N_4826,N_4989);
and U5535 (N_5535,N_4917,N_5071);
nand U5536 (N_5536,N_4921,N_4883);
nand U5537 (N_5537,N_4841,N_4796);
and U5538 (N_5538,N_4586,N_4759);
nor U5539 (N_5539,N_4693,N_5181);
and U5540 (N_5540,N_4798,N_4875);
nand U5541 (N_5541,N_4540,N_4712);
or U5542 (N_5542,N_4892,N_4999);
xnor U5543 (N_5543,N_4914,N_4611);
nand U5544 (N_5544,N_4792,N_4573);
nand U5545 (N_5545,N_5203,N_5239);
nor U5546 (N_5546,N_4990,N_5140);
or U5547 (N_5547,N_4577,N_5045);
and U5548 (N_5548,N_5092,N_5099);
and U5549 (N_5549,N_4863,N_4521);
and U5550 (N_5550,N_4551,N_5194);
nand U5551 (N_5551,N_5054,N_5095);
nand U5552 (N_5552,N_5077,N_5069);
nor U5553 (N_5553,N_5127,N_5131);
xor U5554 (N_5554,N_4912,N_5126);
nor U5555 (N_5555,N_5202,N_4904);
xnor U5556 (N_5556,N_4553,N_5142);
or U5557 (N_5557,N_5051,N_5185);
nor U5558 (N_5558,N_5080,N_4786);
or U5559 (N_5559,N_4878,N_4737);
xnor U5560 (N_5560,N_5169,N_4802);
or U5561 (N_5561,N_4979,N_5213);
xnor U5562 (N_5562,N_4908,N_5170);
nor U5563 (N_5563,N_4936,N_4654);
or U5564 (N_5564,N_5198,N_4643);
or U5565 (N_5565,N_4627,N_4688);
xnor U5566 (N_5566,N_4509,N_5083);
xnor U5567 (N_5567,N_4707,N_5130);
nor U5568 (N_5568,N_4603,N_5033);
or U5569 (N_5569,N_4907,N_5112);
or U5570 (N_5570,N_4708,N_4620);
nand U5571 (N_5571,N_4589,N_4505);
nor U5572 (N_5572,N_4593,N_4675);
or U5573 (N_5573,N_5085,N_4605);
nand U5574 (N_5574,N_5062,N_5022);
xor U5575 (N_5575,N_4642,N_5040);
and U5576 (N_5576,N_4650,N_4639);
nor U5577 (N_5577,N_4884,N_4583);
nand U5578 (N_5578,N_4504,N_4623);
xnor U5579 (N_5579,N_4854,N_4879);
or U5580 (N_5580,N_4948,N_5001);
xnor U5581 (N_5581,N_4692,N_4866);
xor U5582 (N_5582,N_4723,N_4829);
nor U5583 (N_5583,N_5160,N_5028);
nor U5584 (N_5584,N_4986,N_4615);
and U5585 (N_5585,N_5070,N_5014);
and U5586 (N_5586,N_4554,N_4729);
or U5587 (N_5587,N_4785,N_4831);
nand U5588 (N_5588,N_4832,N_4562);
or U5589 (N_5589,N_4626,N_5078);
and U5590 (N_5590,N_4820,N_4991);
and U5591 (N_5591,N_4608,N_5042);
nand U5592 (N_5592,N_4741,N_4869);
nand U5593 (N_5593,N_5162,N_4502);
nor U5594 (N_5594,N_4599,N_4711);
nor U5595 (N_5595,N_4545,N_5197);
xor U5596 (N_5596,N_4857,N_5031);
xor U5597 (N_5597,N_4782,N_4828);
or U5598 (N_5598,N_4601,N_4822);
xor U5599 (N_5599,N_4779,N_4585);
or U5600 (N_5600,N_4717,N_4923);
xnor U5601 (N_5601,N_5171,N_4760);
xnor U5602 (N_5602,N_4733,N_4872);
nor U5603 (N_5603,N_5073,N_5037);
xnor U5604 (N_5604,N_4950,N_4753);
or U5605 (N_5605,N_5135,N_4801);
nor U5606 (N_5606,N_4685,N_4555);
nand U5607 (N_5607,N_4775,N_4856);
or U5608 (N_5608,N_5094,N_4772);
and U5609 (N_5609,N_5034,N_4534);
and U5610 (N_5610,N_4867,N_4734);
xor U5611 (N_5611,N_5163,N_4656);
nor U5612 (N_5612,N_4529,N_5035);
xor U5613 (N_5613,N_4973,N_4859);
nor U5614 (N_5614,N_4629,N_5114);
or U5615 (N_5615,N_5192,N_5093);
xnor U5616 (N_5616,N_4916,N_5243);
xor U5617 (N_5617,N_4515,N_4657);
or U5618 (N_5618,N_4670,N_4790);
or U5619 (N_5619,N_4666,N_4744);
xnor U5620 (N_5620,N_4959,N_4819);
xnor U5621 (N_5621,N_4797,N_4972);
nand U5622 (N_5622,N_4824,N_4745);
nor U5623 (N_5623,N_4978,N_5076);
nand U5624 (N_5624,N_4614,N_4704);
and U5625 (N_5625,N_5139,N_4777);
or U5626 (N_5626,N_5026,N_4958);
or U5627 (N_5627,N_4778,N_4520);
nor U5628 (N_5628,N_4708,N_4727);
nor U5629 (N_5629,N_4535,N_5019);
nand U5630 (N_5630,N_4501,N_4623);
xor U5631 (N_5631,N_4741,N_4862);
and U5632 (N_5632,N_5144,N_5211);
nand U5633 (N_5633,N_4811,N_4779);
and U5634 (N_5634,N_4990,N_4888);
xnor U5635 (N_5635,N_4628,N_5025);
or U5636 (N_5636,N_5049,N_5100);
or U5637 (N_5637,N_5095,N_4564);
xor U5638 (N_5638,N_4649,N_5209);
or U5639 (N_5639,N_4958,N_4774);
nor U5640 (N_5640,N_4661,N_4924);
xor U5641 (N_5641,N_4707,N_4516);
and U5642 (N_5642,N_5069,N_4849);
xnor U5643 (N_5643,N_4688,N_5029);
or U5644 (N_5644,N_4976,N_4811);
and U5645 (N_5645,N_4776,N_4920);
nand U5646 (N_5646,N_5048,N_5111);
or U5647 (N_5647,N_4787,N_4809);
nand U5648 (N_5648,N_4875,N_4882);
nand U5649 (N_5649,N_4870,N_5100);
and U5650 (N_5650,N_5030,N_4611);
and U5651 (N_5651,N_4610,N_4936);
nand U5652 (N_5652,N_5154,N_4916);
and U5653 (N_5653,N_4914,N_5232);
nor U5654 (N_5654,N_4524,N_5093);
nor U5655 (N_5655,N_4814,N_4828);
nand U5656 (N_5656,N_5136,N_5088);
and U5657 (N_5657,N_5140,N_5165);
and U5658 (N_5658,N_4544,N_4535);
xnor U5659 (N_5659,N_4953,N_4635);
xor U5660 (N_5660,N_4656,N_5036);
and U5661 (N_5661,N_5018,N_4990);
nand U5662 (N_5662,N_4847,N_4924);
nand U5663 (N_5663,N_5127,N_4529);
xnor U5664 (N_5664,N_4907,N_4518);
xor U5665 (N_5665,N_4650,N_4535);
xor U5666 (N_5666,N_5047,N_5099);
nor U5667 (N_5667,N_5206,N_5202);
nand U5668 (N_5668,N_4868,N_4995);
or U5669 (N_5669,N_5055,N_5064);
nand U5670 (N_5670,N_4626,N_4974);
xnor U5671 (N_5671,N_4992,N_4881);
or U5672 (N_5672,N_4887,N_4859);
xor U5673 (N_5673,N_4547,N_4748);
or U5674 (N_5674,N_5091,N_4738);
nor U5675 (N_5675,N_4566,N_5042);
nand U5676 (N_5676,N_4814,N_4774);
and U5677 (N_5677,N_4969,N_4576);
and U5678 (N_5678,N_5096,N_4603);
and U5679 (N_5679,N_5046,N_4947);
xor U5680 (N_5680,N_5176,N_4760);
nand U5681 (N_5681,N_4652,N_4743);
or U5682 (N_5682,N_4981,N_4551);
xnor U5683 (N_5683,N_5078,N_5173);
nand U5684 (N_5684,N_5106,N_4606);
nor U5685 (N_5685,N_5148,N_5006);
or U5686 (N_5686,N_5185,N_5151);
and U5687 (N_5687,N_4802,N_4757);
or U5688 (N_5688,N_4694,N_5204);
nand U5689 (N_5689,N_4642,N_4609);
and U5690 (N_5690,N_4985,N_5073);
or U5691 (N_5691,N_4502,N_4731);
nand U5692 (N_5692,N_4926,N_4947);
and U5693 (N_5693,N_4553,N_4711);
or U5694 (N_5694,N_5067,N_4676);
or U5695 (N_5695,N_4688,N_4523);
or U5696 (N_5696,N_4897,N_5168);
nor U5697 (N_5697,N_5026,N_4906);
xnor U5698 (N_5698,N_4809,N_4879);
nand U5699 (N_5699,N_5079,N_5068);
nor U5700 (N_5700,N_4865,N_4664);
and U5701 (N_5701,N_4605,N_5245);
xor U5702 (N_5702,N_5096,N_4866);
nand U5703 (N_5703,N_4510,N_5231);
nor U5704 (N_5704,N_5170,N_4867);
nand U5705 (N_5705,N_5019,N_4804);
xor U5706 (N_5706,N_4560,N_4772);
xnor U5707 (N_5707,N_4900,N_5033);
or U5708 (N_5708,N_4723,N_5122);
nor U5709 (N_5709,N_4675,N_5115);
nand U5710 (N_5710,N_4557,N_4932);
nor U5711 (N_5711,N_4678,N_4515);
xor U5712 (N_5712,N_4791,N_4705);
and U5713 (N_5713,N_5210,N_4733);
xor U5714 (N_5714,N_4941,N_4740);
nand U5715 (N_5715,N_4981,N_4725);
xor U5716 (N_5716,N_4622,N_4502);
and U5717 (N_5717,N_4880,N_5061);
nand U5718 (N_5718,N_5165,N_4936);
nor U5719 (N_5719,N_5125,N_5015);
or U5720 (N_5720,N_5089,N_4753);
nor U5721 (N_5721,N_4700,N_4797);
xor U5722 (N_5722,N_5207,N_4638);
or U5723 (N_5723,N_4670,N_4514);
or U5724 (N_5724,N_4589,N_5244);
or U5725 (N_5725,N_4611,N_5097);
nor U5726 (N_5726,N_5064,N_4943);
or U5727 (N_5727,N_4539,N_4945);
nand U5728 (N_5728,N_4652,N_4924);
nor U5729 (N_5729,N_5037,N_5087);
nand U5730 (N_5730,N_5125,N_5106);
nor U5731 (N_5731,N_4680,N_5200);
nor U5732 (N_5732,N_4716,N_4597);
xnor U5733 (N_5733,N_4530,N_4854);
or U5734 (N_5734,N_4914,N_4983);
nor U5735 (N_5735,N_4752,N_5112);
nor U5736 (N_5736,N_4621,N_4792);
nand U5737 (N_5737,N_5228,N_4595);
or U5738 (N_5738,N_4723,N_4561);
nor U5739 (N_5739,N_5024,N_4808);
nor U5740 (N_5740,N_5051,N_5056);
xor U5741 (N_5741,N_5098,N_5151);
xor U5742 (N_5742,N_4766,N_5232);
xor U5743 (N_5743,N_5067,N_5058);
or U5744 (N_5744,N_4981,N_4716);
or U5745 (N_5745,N_4982,N_4653);
nand U5746 (N_5746,N_4959,N_4801);
nor U5747 (N_5747,N_4691,N_4755);
and U5748 (N_5748,N_5057,N_4784);
and U5749 (N_5749,N_4977,N_5230);
and U5750 (N_5750,N_4777,N_4683);
and U5751 (N_5751,N_4710,N_4516);
xnor U5752 (N_5752,N_4708,N_5160);
xnor U5753 (N_5753,N_4552,N_5186);
nand U5754 (N_5754,N_4836,N_4877);
nor U5755 (N_5755,N_4698,N_5173);
nor U5756 (N_5756,N_5133,N_5152);
nand U5757 (N_5757,N_4548,N_4537);
xnor U5758 (N_5758,N_4859,N_4927);
xnor U5759 (N_5759,N_5050,N_4572);
and U5760 (N_5760,N_4840,N_5023);
nand U5761 (N_5761,N_4846,N_4896);
and U5762 (N_5762,N_4866,N_4799);
nor U5763 (N_5763,N_4630,N_4592);
or U5764 (N_5764,N_4876,N_4683);
nand U5765 (N_5765,N_5057,N_4905);
and U5766 (N_5766,N_5067,N_4516);
nand U5767 (N_5767,N_4703,N_4700);
and U5768 (N_5768,N_4685,N_4832);
and U5769 (N_5769,N_4655,N_5105);
xnor U5770 (N_5770,N_4758,N_4968);
xnor U5771 (N_5771,N_4599,N_4515);
and U5772 (N_5772,N_4768,N_5013);
nand U5773 (N_5773,N_5229,N_4963);
nor U5774 (N_5774,N_5069,N_5012);
or U5775 (N_5775,N_5244,N_4524);
or U5776 (N_5776,N_5101,N_5022);
nor U5777 (N_5777,N_4559,N_5096);
or U5778 (N_5778,N_5230,N_5126);
or U5779 (N_5779,N_5110,N_5143);
nand U5780 (N_5780,N_4864,N_5063);
xnor U5781 (N_5781,N_4863,N_5189);
xor U5782 (N_5782,N_4748,N_5134);
or U5783 (N_5783,N_4795,N_4918);
nand U5784 (N_5784,N_5129,N_5046);
and U5785 (N_5785,N_5056,N_4789);
nor U5786 (N_5786,N_5038,N_4501);
and U5787 (N_5787,N_5129,N_5089);
xor U5788 (N_5788,N_4826,N_4986);
and U5789 (N_5789,N_5012,N_4835);
xnor U5790 (N_5790,N_4846,N_5081);
nand U5791 (N_5791,N_5127,N_4550);
nor U5792 (N_5792,N_5237,N_5204);
and U5793 (N_5793,N_4870,N_5038);
and U5794 (N_5794,N_4572,N_4851);
nor U5795 (N_5795,N_4915,N_5008);
or U5796 (N_5796,N_5220,N_5121);
xor U5797 (N_5797,N_5018,N_4816);
xor U5798 (N_5798,N_4863,N_5135);
or U5799 (N_5799,N_4769,N_4910);
nor U5800 (N_5800,N_5135,N_5150);
nand U5801 (N_5801,N_5063,N_4646);
nand U5802 (N_5802,N_4987,N_4988);
nor U5803 (N_5803,N_4684,N_5161);
nor U5804 (N_5804,N_4646,N_4653);
xor U5805 (N_5805,N_4620,N_4627);
nand U5806 (N_5806,N_5224,N_4977);
nand U5807 (N_5807,N_4544,N_4633);
and U5808 (N_5808,N_4997,N_5067);
or U5809 (N_5809,N_4699,N_4601);
nand U5810 (N_5810,N_4952,N_5213);
nor U5811 (N_5811,N_4952,N_4784);
xnor U5812 (N_5812,N_4828,N_4619);
and U5813 (N_5813,N_5159,N_4572);
nor U5814 (N_5814,N_4739,N_4770);
xnor U5815 (N_5815,N_4986,N_4551);
and U5816 (N_5816,N_5075,N_5165);
and U5817 (N_5817,N_4506,N_5172);
nand U5818 (N_5818,N_4864,N_5116);
nand U5819 (N_5819,N_4529,N_4989);
nand U5820 (N_5820,N_4736,N_4944);
nand U5821 (N_5821,N_4658,N_5114);
xnor U5822 (N_5822,N_4554,N_4846);
nand U5823 (N_5823,N_5026,N_4828);
nor U5824 (N_5824,N_4957,N_4996);
nand U5825 (N_5825,N_5183,N_4634);
xnor U5826 (N_5826,N_4877,N_4618);
or U5827 (N_5827,N_4821,N_5226);
nor U5828 (N_5828,N_4682,N_5112);
xnor U5829 (N_5829,N_5244,N_4604);
and U5830 (N_5830,N_5213,N_4847);
xnor U5831 (N_5831,N_4595,N_4689);
nor U5832 (N_5832,N_5035,N_4757);
or U5833 (N_5833,N_4741,N_5007);
nor U5834 (N_5834,N_5128,N_5050);
or U5835 (N_5835,N_4651,N_5137);
nor U5836 (N_5836,N_5216,N_4509);
or U5837 (N_5837,N_4620,N_4803);
and U5838 (N_5838,N_4529,N_5173);
and U5839 (N_5839,N_4524,N_4623);
and U5840 (N_5840,N_5183,N_4567);
nor U5841 (N_5841,N_4898,N_5004);
nor U5842 (N_5842,N_4554,N_5231);
or U5843 (N_5843,N_5188,N_4587);
or U5844 (N_5844,N_5042,N_4586);
nor U5845 (N_5845,N_5177,N_4542);
or U5846 (N_5846,N_5229,N_4830);
xor U5847 (N_5847,N_4545,N_5099);
nand U5848 (N_5848,N_4828,N_5094);
or U5849 (N_5849,N_4559,N_4588);
nand U5850 (N_5850,N_5121,N_4862);
nor U5851 (N_5851,N_4801,N_5207);
nor U5852 (N_5852,N_5056,N_4775);
xnor U5853 (N_5853,N_4993,N_4775);
nor U5854 (N_5854,N_5071,N_4591);
and U5855 (N_5855,N_4943,N_4600);
or U5856 (N_5856,N_5196,N_4588);
nor U5857 (N_5857,N_4909,N_4816);
xor U5858 (N_5858,N_5086,N_4746);
and U5859 (N_5859,N_4911,N_5106);
nor U5860 (N_5860,N_4716,N_4781);
nand U5861 (N_5861,N_4948,N_5047);
or U5862 (N_5862,N_5159,N_5113);
xor U5863 (N_5863,N_4963,N_5029);
nand U5864 (N_5864,N_4994,N_5035);
nor U5865 (N_5865,N_4783,N_4656);
xor U5866 (N_5866,N_4836,N_5166);
xor U5867 (N_5867,N_4687,N_5148);
nor U5868 (N_5868,N_4908,N_5217);
nand U5869 (N_5869,N_4826,N_5016);
xor U5870 (N_5870,N_5125,N_4819);
nor U5871 (N_5871,N_4949,N_4539);
nand U5872 (N_5872,N_5018,N_5235);
or U5873 (N_5873,N_4750,N_5093);
xor U5874 (N_5874,N_5073,N_4644);
nor U5875 (N_5875,N_5240,N_4770);
xor U5876 (N_5876,N_4761,N_5007);
or U5877 (N_5877,N_4958,N_5166);
nor U5878 (N_5878,N_5018,N_4888);
nand U5879 (N_5879,N_5002,N_4691);
nor U5880 (N_5880,N_4599,N_5078);
nand U5881 (N_5881,N_5105,N_4544);
and U5882 (N_5882,N_5020,N_4508);
or U5883 (N_5883,N_4989,N_5086);
nor U5884 (N_5884,N_4632,N_4584);
xor U5885 (N_5885,N_5067,N_5091);
nand U5886 (N_5886,N_5231,N_5002);
or U5887 (N_5887,N_5056,N_5079);
nor U5888 (N_5888,N_4964,N_4522);
nand U5889 (N_5889,N_5037,N_4975);
nor U5890 (N_5890,N_4943,N_5248);
or U5891 (N_5891,N_4585,N_4983);
or U5892 (N_5892,N_4977,N_4867);
and U5893 (N_5893,N_4533,N_4683);
xor U5894 (N_5894,N_5073,N_5207);
or U5895 (N_5895,N_5237,N_4558);
and U5896 (N_5896,N_5141,N_4562);
or U5897 (N_5897,N_4566,N_4557);
nor U5898 (N_5898,N_4763,N_4934);
xor U5899 (N_5899,N_4835,N_5199);
nor U5900 (N_5900,N_4911,N_4950);
nor U5901 (N_5901,N_4900,N_4800);
and U5902 (N_5902,N_4595,N_4791);
nor U5903 (N_5903,N_4604,N_4649);
xnor U5904 (N_5904,N_5022,N_4728);
or U5905 (N_5905,N_4983,N_4734);
and U5906 (N_5906,N_4795,N_4526);
nand U5907 (N_5907,N_5065,N_4712);
and U5908 (N_5908,N_5011,N_4980);
xnor U5909 (N_5909,N_4625,N_4940);
xnor U5910 (N_5910,N_4794,N_5067);
and U5911 (N_5911,N_4994,N_4630);
nand U5912 (N_5912,N_4576,N_5148);
and U5913 (N_5913,N_4771,N_4532);
and U5914 (N_5914,N_5224,N_4961);
or U5915 (N_5915,N_4934,N_4928);
nor U5916 (N_5916,N_4853,N_4866);
xor U5917 (N_5917,N_4946,N_4627);
or U5918 (N_5918,N_5164,N_5245);
xnor U5919 (N_5919,N_4785,N_4846);
or U5920 (N_5920,N_5242,N_4712);
nor U5921 (N_5921,N_4614,N_5213);
or U5922 (N_5922,N_4608,N_4711);
xnor U5923 (N_5923,N_5064,N_5030);
xor U5924 (N_5924,N_4792,N_4860);
nand U5925 (N_5925,N_4781,N_5035);
or U5926 (N_5926,N_4665,N_4651);
nor U5927 (N_5927,N_4919,N_4590);
or U5928 (N_5928,N_4916,N_4820);
nor U5929 (N_5929,N_4808,N_4618);
and U5930 (N_5930,N_4802,N_4983);
and U5931 (N_5931,N_4581,N_4910);
nor U5932 (N_5932,N_4572,N_4664);
nand U5933 (N_5933,N_5226,N_5203);
and U5934 (N_5934,N_4539,N_4554);
xor U5935 (N_5935,N_5062,N_4935);
or U5936 (N_5936,N_4749,N_4772);
nand U5937 (N_5937,N_4905,N_4924);
and U5938 (N_5938,N_4830,N_5044);
xor U5939 (N_5939,N_4524,N_5224);
nand U5940 (N_5940,N_5182,N_4762);
xor U5941 (N_5941,N_4528,N_4602);
and U5942 (N_5942,N_4552,N_4779);
or U5943 (N_5943,N_4931,N_4842);
nand U5944 (N_5944,N_4884,N_4899);
nor U5945 (N_5945,N_4526,N_4744);
nand U5946 (N_5946,N_4894,N_4974);
or U5947 (N_5947,N_4569,N_4767);
or U5948 (N_5948,N_4929,N_4626);
and U5949 (N_5949,N_4898,N_5117);
nand U5950 (N_5950,N_4688,N_4569);
or U5951 (N_5951,N_4690,N_5029);
and U5952 (N_5952,N_5211,N_4926);
and U5953 (N_5953,N_4557,N_4875);
and U5954 (N_5954,N_4757,N_4874);
and U5955 (N_5955,N_5232,N_5121);
and U5956 (N_5956,N_4632,N_4571);
xnor U5957 (N_5957,N_4503,N_5070);
xnor U5958 (N_5958,N_5115,N_4674);
or U5959 (N_5959,N_4817,N_5233);
and U5960 (N_5960,N_4869,N_5194);
or U5961 (N_5961,N_5241,N_4816);
xnor U5962 (N_5962,N_4512,N_4501);
and U5963 (N_5963,N_5051,N_4664);
nand U5964 (N_5964,N_4758,N_4688);
and U5965 (N_5965,N_4845,N_5069);
and U5966 (N_5966,N_5110,N_4911);
nand U5967 (N_5967,N_4686,N_5046);
or U5968 (N_5968,N_4803,N_5029);
nand U5969 (N_5969,N_4839,N_4888);
or U5970 (N_5970,N_4763,N_4908);
or U5971 (N_5971,N_5163,N_4571);
nor U5972 (N_5972,N_5219,N_4978);
nand U5973 (N_5973,N_5139,N_5096);
xnor U5974 (N_5974,N_5162,N_5085);
and U5975 (N_5975,N_5063,N_4829);
or U5976 (N_5976,N_5046,N_4665);
and U5977 (N_5977,N_4848,N_4855);
nand U5978 (N_5978,N_4639,N_4848);
nand U5979 (N_5979,N_4578,N_4841);
nor U5980 (N_5980,N_5041,N_4682);
nor U5981 (N_5981,N_4778,N_4851);
or U5982 (N_5982,N_5025,N_4876);
nand U5983 (N_5983,N_5237,N_4806);
nor U5984 (N_5984,N_4672,N_4957);
nor U5985 (N_5985,N_5125,N_4552);
nand U5986 (N_5986,N_5233,N_4718);
or U5987 (N_5987,N_5188,N_5005);
nor U5988 (N_5988,N_4842,N_5114);
nor U5989 (N_5989,N_4932,N_4995);
nor U5990 (N_5990,N_5207,N_4685);
or U5991 (N_5991,N_5191,N_4592);
xnor U5992 (N_5992,N_5072,N_5242);
and U5993 (N_5993,N_4657,N_5157);
xor U5994 (N_5994,N_4943,N_4567);
xor U5995 (N_5995,N_4605,N_5101);
xnor U5996 (N_5996,N_4782,N_5037);
nand U5997 (N_5997,N_4502,N_4799);
xor U5998 (N_5998,N_4923,N_4656);
xor U5999 (N_5999,N_4757,N_5239);
or U6000 (N_6000,N_5475,N_5807);
xnor U6001 (N_6001,N_5579,N_5465);
and U6002 (N_6002,N_5435,N_5455);
and U6003 (N_6003,N_5392,N_5381);
or U6004 (N_6004,N_5756,N_5285);
nor U6005 (N_6005,N_5681,N_5943);
and U6006 (N_6006,N_5782,N_5798);
xor U6007 (N_6007,N_5634,N_5696);
nand U6008 (N_6008,N_5764,N_5910);
nor U6009 (N_6009,N_5480,N_5519);
and U6010 (N_6010,N_5427,N_5655);
and U6011 (N_6011,N_5532,N_5868);
nand U6012 (N_6012,N_5975,N_5441);
nor U6013 (N_6013,N_5436,N_5469);
and U6014 (N_6014,N_5330,N_5449);
nand U6015 (N_6015,N_5903,N_5640);
and U6016 (N_6016,N_5871,N_5405);
or U6017 (N_6017,N_5996,N_5929);
or U6018 (N_6018,N_5886,N_5918);
or U6019 (N_6019,N_5927,N_5725);
and U6020 (N_6020,N_5628,N_5810);
nor U6021 (N_6021,N_5793,N_5960);
or U6022 (N_6022,N_5522,N_5763);
nor U6023 (N_6023,N_5361,N_5269);
or U6024 (N_6024,N_5790,N_5332);
xnor U6025 (N_6025,N_5999,N_5397);
or U6026 (N_6026,N_5489,N_5765);
nor U6027 (N_6027,N_5732,N_5341);
xnor U6028 (N_6028,N_5561,N_5671);
and U6029 (N_6029,N_5598,N_5669);
or U6030 (N_6030,N_5797,N_5914);
nor U6031 (N_6031,N_5878,N_5733);
nand U6032 (N_6032,N_5576,N_5981);
xor U6033 (N_6033,N_5883,N_5746);
and U6034 (N_6034,N_5492,N_5823);
xor U6035 (N_6035,N_5656,N_5843);
and U6036 (N_6036,N_5761,N_5958);
nor U6037 (N_6037,N_5691,N_5390);
and U6038 (N_6038,N_5560,N_5808);
xor U6039 (N_6039,N_5700,N_5491);
or U6040 (N_6040,N_5302,N_5463);
or U6041 (N_6041,N_5288,N_5251);
xnor U6042 (N_6042,N_5428,N_5483);
and U6043 (N_6043,N_5722,N_5769);
nor U6044 (N_6044,N_5657,N_5425);
or U6045 (N_6045,N_5697,N_5688);
xnor U6046 (N_6046,N_5750,N_5266);
or U6047 (N_6047,N_5282,N_5580);
xnor U6048 (N_6048,N_5633,N_5500);
or U6049 (N_6049,N_5607,N_5401);
or U6050 (N_6050,N_5612,N_5378);
or U6051 (N_6051,N_5791,N_5521);
nor U6052 (N_6052,N_5415,N_5569);
and U6053 (N_6053,N_5389,N_5991);
nor U6054 (N_6054,N_5307,N_5711);
nand U6055 (N_6055,N_5759,N_5313);
and U6056 (N_6056,N_5841,N_5968);
nor U6057 (N_6057,N_5357,N_5388);
or U6058 (N_6058,N_5842,N_5873);
nor U6059 (N_6059,N_5311,N_5399);
xor U6060 (N_6060,N_5281,N_5358);
or U6061 (N_6061,N_5433,N_5424);
nand U6062 (N_6062,N_5507,N_5998);
and U6063 (N_6063,N_5801,N_5366);
nand U6064 (N_6064,N_5271,N_5546);
and U6065 (N_6065,N_5887,N_5961);
nor U6066 (N_6066,N_5595,N_5565);
xor U6067 (N_6067,N_5400,N_5987);
nand U6068 (N_6068,N_5942,N_5421);
and U6069 (N_6069,N_5408,N_5636);
or U6070 (N_6070,N_5740,N_5642);
nor U6071 (N_6071,N_5894,N_5846);
nand U6072 (N_6072,N_5516,N_5496);
nor U6073 (N_6073,N_5944,N_5438);
or U6074 (N_6074,N_5668,N_5789);
nor U6075 (N_6075,N_5992,N_5261);
nand U6076 (N_6076,N_5641,N_5803);
nand U6077 (N_6077,N_5515,N_5356);
or U6078 (N_6078,N_5979,N_5658);
xnor U6079 (N_6079,N_5348,N_5275);
and U6080 (N_6080,N_5833,N_5771);
or U6081 (N_6081,N_5673,N_5512);
nand U6082 (N_6082,N_5965,N_5335);
and U6083 (N_6083,N_5494,N_5360);
nand U6084 (N_6084,N_5646,N_5329);
xnor U6085 (N_6085,N_5613,N_5799);
nand U6086 (N_6086,N_5319,N_5384);
nor U6087 (N_6087,N_5826,N_5490);
nor U6088 (N_6088,N_5347,N_5953);
or U6089 (N_6089,N_5338,N_5616);
xnor U6090 (N_6090,N_5983,N_5638);
xor U6091 (N_6091,N_5581,N_5986);
xnor U6092 (N_6092,N_5343,N_5349);
xnor U6093 (N_6093,N_5306,N_5915);
nor U6094 (N_6094,N_5540,N_5362);
or U6095 (N_6095,N_5481,N_5555);
or U6096 (N_6096,N_5359,N_5539);
xor U6097 (N_6097,N_5821,N_5690);
nor U6098 (N_6098,N_5345,N_5312);
and U6099 (N_6099,N_5585,N_5908);
or U6100 (N_6100,N_5327,N_5370);
nor U6101 (N_6101,N_5395,N_5672);
xor U6102 (N_6102,N_5434,N_5809);
xor U6103 (N_6103,N_5670,N_5620);
nor U6104 (N_6104,N_5663,N_5501);
nor U6105 (N_6105,N_5704,N_5698);
and U6106 (N_6106,N_5604,N_5377);
xnor U6107 (N_6107,N_5351,N_5582);
xor U6108 (N_6108,N_5486,N_5605);
nand U6109 (N_6109,N_5568,N_5856);
nand U6110 (N_6110,N_5817,N_5255);
xor U6111 (N_6111,N_5818,N_5406);
xor U6112 (N_6112,N_5872,N_5694);
nor U6113 (N_6113,N_5280,N_5851);
nor U6114 (N_6114,N_5615,N_5660);
nor U6115 (N_6115,N_5296,N_5333);
nand U6116 (N_6116,N_5895,N_5713);
nand U6117 (N_6117,N_5250,N_5297);
xnor U6118 (N_6118,N_5837,N_5523);
or U6119 (N_6119,N_5447,N_5606);
xnor U6120 (N_6120,N_5890,N_5664);
or U6121 (N_6121,N_5778,N_5754);
xor U6122 (N_6122,N_5795,N_5334);
and U6123 (N_6123,N_5562,N_5462);
and U6124 (N_6124,N_5674,N_5477);
nand U6125 (N_6125,N_5665,N_5703);
nand U6126 (N_6126,N_5667,N_5577);
xnor U6127 (N_6127,N_5881,N_5687);
or U6128 (N_6128,N_5549,N_5547);
or U6129 (N_6129,N_5682,N_5721);
nor U6130 (N_6130,N_5830,N_5734);
and U6131 (N_6131,N_5744,N_5346);
nand U6132 (N_6132,N_5423,N_5932);
or U6133 (N_6133,N_5368,N_5310);
or U6134 (N_6134,N_5629,N_5344);
nor U6135 (N_6135,N_5928,N_5277);
nor U6136 (N_6136,N_5286,N_5858);
nor U6137 (N_6137,N_5289,N_5626);
or U6138 (N_6138,N_5644,N_5853);
or U6139 (N_6139,N_5325,N_5901);
nand U6140 (N_6140,N_5816,N_5743);
and U6141 (N_6141,N_5774,N_5314);
nand U6142 (N_6142,N_5749,N_5564);
or U6143 (N_6143,N_5315,N_5498);
xnor U6144 (N_6144,N_5430,N_5556);
or U6145 (N_6145,N_5410,N_5453);
and U6146 (N_6146,N_5573,N_5630);
nand U6147 (N_6147,N_5685,N_5534);
xnor U6148 (N_6148,N_5404,N_5859);
or U6149 (N_6149,N_5650,N_5773);
xor U6150 (N_6150,N_5326,N_5478);
and U6151 (N_6151,N_5884,N_5647);
xor U6152 (N_6152,N_5840,N_5331);
nor U6153 (N_6153,N_5493,N_5819);
xnor U6154 (N_6154,N_5416,N_5445);
nand U6155 (N_6155,N_5948,N_5941);
and U6156 (N_6156,N_5279,N_5679);
and U6157 (N_6157,N_5571,N_5552);
xor U6158 (N_6158,N_5768,N_5309);
xnor U6159 (N_6159,N_5848,N_5730);
and U6160 (N_6160,N_5900,N_5380);
or U6161 (N_6161,N_5814,N_5784);
nand U6162 (N_6162,N_5464,N_5301);
or U6163 (N_6163,N_5850,N_5383);
or U6164 (N_6164,N_5260,N_5363);
or U6165 (N_6165,N_5709,N_5382);
or U6166 (N_6166,N_5712,N_5468);
xnor U6167 (N_6167,N_5374,N_5542);
nand U6168 (N_6168,N_5731,N_5418);
xnor U6169 (N_6169,N_5533,N_5939);
nand U6170 (N_6170,N_5747,N_5340);
xor U6171 (N_6171,N_5551,N_5499);
and U6172 (N_6172,N_5940,N_5945);
xnor U6173 (N_6173,N_5320,N_5432);
nor U6174 (N_6174,N_5323,N_5758);
nand U6175 (N_6175,N_5662,N_5446);
nand U6176 (N_6176,N_5584,N_5708);
or U6177 (N_6177,N_5862,N_5502);
nand U6178 (N_6178,N_5632,N_5693);
and U6179 (N_6179,N_5590,N_5587);
xor U6180 (N_6180,N_5966,N_5511);
xnor U6181 (N_6181,N_5276,N_5457);
xor U6182 (N_6182,N_5291,N_5924);
xor U6183 (N_6183,N_5969,N_5263);
nor U6184 (N_6184,N_5505,N_5898);
nand U6185 (N_6185,N_5268,N_5411);
nor U6186 (N_6186,N_5920,N_5596);
and U6187 (N_6187,N_5867,N_5514);
xnor U6188 (N_6188,N_5906,N_5666);
and U6189 (N_6189,N_5300,N_5829);
nand U6190 (N_6190,N_5525,N_5484);
or U6191 (N_6191,N_5745,N_5369);
nor U6192 (N_6192,N_5802,N_5951);
nand U6193 (N_6193,N_5476,N_5394);
and U6194 (N_6194,N_5264,N_5470);
or U6195 (N_6195,N_5461,N_5426);
nor U6196 (N_6196,N_5787,N_5659);
and U6197 (N_6197,N_5957,N_5473);
nand U6198 (N_6198,N_5994,N_5550);
and U6199 (N_6199,N_5278,N_5931);
or U6200 (N_6200,N_5938,N_5917);
nand U6201 (N_6201,N_5838,N_5599);
or U6202 (N_6202,N_5376,N_5460);
or U6203 (N_6203,N_5839,N_5379);
or U6204 (N_6204,N_5706,N_5448);
and U6205 (N_6205,N_5592,N_5882);
nand U6206 (N_6206,N_5413,N_5825);
nor U6207 (N_6207,N_5788,N_5738);
nand U6208 (N_6208,N_5431,N_5964);
nor U6209 (N_6209,N_5267,N_5503);
or U6210 (N_6210,N_5274,N_5907);
xnor U6211 (N_6211,N_5583,N_5528);
nor U6212 (N_6212,N_5518,N_5935);
and U6213 (N_6213,N_5885,N_5365);
and U6214 (N_6214,N_5544,N_5252);
and U6215 (N_6215,N_5257,N_5482);
xnor U6216 (N_6216,N_5852,N_5328);
nor U6217 (N_6217,N_5923,N_5618);
or U6218 (N_6218,N_5701,N_5686);
and U6219 (N_6219,N_5272,N_5752);
nand U6220 (N_6220,N_5762,N_5471);
or U6221 (N_6221,N_5391,N_5517);
and U6222 (N_6222,N_5535,N_5813);
and U6223 (N_6223,N_5537,N_5678);
nor U6224 (N_6224,N_5982,N_5354);
nor U6225 (N_6225,N_5637,N_5287);
nand U6226 (N_6226,N_5324,N_5591);
nor U6227 (N_6227,N_5876,N_5429);
and U6228 (N_6228,N_5947,N_5985);
nand U6229 (N_6229,N_5407,N_5954);
nor U6230 (N_6230,N_5553,N_5995);
nand U6231 (N_6231,N_5724,N_5339);
and U6232 (N_6232,N_5558,N_5989);
nor U6233 (N_6233,N_5254,N_5689);
and U6234 (N_6234,N_5566,N_5949);
or U6235 (N_6235,N_5748,N_5624);
nor U6236 (N_6236,N_5993,N_5364);
nor U6237 (N_6237,N_5531,N_5290);
xnor U6238 (N_6238,N_5880,N_5892);
nand U6239 (N_6239,N_5770,N_5609);
nand U6240 (N_6240,N_5972,N_5834);
nand U6241 (N_6241,N_5353,N_5575);
nand U6242 (N_6242,N_5912,N_5265);
nand U6243 (N_6243,N_5815,N_5653);
and U6244 (N_6244,N_5718,N_5506);
xnor U6245 (N_6245,N_5946,N_5610);
xnor U6246 (N_6246,N_5766,N_5717);
and U6247 (N_6247,N_5726,N_5779);
and U6248 (N_6248,N_5710,N_5916);
and U6249 (N_6249,N_5299,N_5574);
and U6250 (N_6250,N_5488,N_5772);
xor U6251 (N_6251,N_5497,N_5661);
and U6252 (N_6252,N_5875,N_5648);
or U6253 (N_6253,N_5716,N_5757);
xor U6254 (N_6254,N_5896,N_5594);
or U6255 (N_6255,N_5893,N_5736);
xnor U6256 (N_6256,N_5836,N_5824);
or U6257 (N_6257,N_5835,N_5973);
and U6258 (N_6258,N_5372,N_5877);
nand U6259 (N_6259,N_5753,N_5352);
and U6260 (N_6260,N_5403,N_5990);
and U6261 (N_6261,N_5619,N_5723);
and U6262 (N_6262,N_5922,N_5776);
nor U6263 (N_6263,N_5485,N_5371);
xor U6264 (N_6264,N_5977,N_5980);
xor U6265 (N_6265,N_5589,N_5467);
or U6266 (N_6266,N_5651,N_5337);
nor U6267 (N_6267,N_5997,N_5861);
nor U6268 (N_6268,N_5538,N_5355);
nand U6269 (N_6269,N_5393,N_5913);
nand U6270 (N_6270,N_5775,N_5563);
xor U6271 (N_6271,N_5611,N_5976);
xor U6272 (N_6272,N_5812,N_5603);
or U6273 (N_6273,N_5419,N_5737);
xor U6274 (N_6274,N_5739,N_5777);
xnor U6275 (N_6275,N_5847,N_5262);
xor U6276 (N_6276,N_5675,N_5963);
and U6277 (N_6277,N_5909,N_5600);
or U6278 (N_6278,N_5458,N_5904);
or U6279 (N_6279,N_5865,N_5298);
xnor U6280 (N_6280,N_5959,N_5783);
nor U6281 (N_6281,N_5845,N_5714);
and U6282 (N_6282,N_5936,N_5617);
nand U6283 (N_6283,N_5934,N_5741);
nand U6284 (N_6284,N_5373,N_5548);
xor U6285 (N_6285,N_5530,N_5614);
xor U6286 (N_6286,N_5677,N_5316);
xnor U6287 (N_6287,N_5479,N_5627);
and U6288 (N_6288,N_5857,N_5412);
and U6289 (N_6289,N_5495,N_5336);
and U6290 (N_6290,N_5889,N_5524);
or U6291 (N_6291,N_5970,N_5863);
or U6292 (N_6292,N_5956,N_5402);
or U6293 (N_6293,N_5827,N_5926);
and U6294 (N_6294,N_5707,N_5367);
nor U6295 (N_6295,N_5444,N_5805);
nand U6296 (N_6296,N_5385,N_5317);
or U6297 (N_6297,N_5396,N_5719);
nand U6298 (N_6298,N_5294,N_5806);
nand U6299 (N_6299,N_5652,N_5273);
nor U6300 (N_6300,N_5578,N_5705);
or U6301 (N_6301,N_5414,N_5398);
and U6302 (N_6302,N_5601,N_5526);
and U6303 (N_6303,N_5735,N_5304);
or U6304 (N_6304,N_5962,N_5536);
nand U6305 (N_6305,N_5293,N_5459);
xor U6306 (N_6306,N_5342,N_5676);
xnor U6307 (N_6307,N_5925,N_5621);
xnor U6308 (N_6308,N_5452,N_5699);
and U6309 (N_6309,N_5792,N_5796);
or U6310 (N_6310,N_5950,N_5466);
nand U6311 (N_6311,N_5794,N_5937);
xnor U6312 (N_6312,N_5639,N_5854);
or U6313 (N_6313,N_5680,N_5866);
xor U6314 (N_6314,N_5767,N_5683);
and U6315 (N_6315,N_5545,N_5849);
xnor U6316 (N_6316,N_5695,N_5978);
or U6317 (N_6317,N_5828,N_5322);
or U6318 (N_6318,N_5897,N_5955);
nor U6319 (N_6319,N_5780,N_5510);
xnor U6320 (N_6320,N_5559,N_5645);
or U6321 (N_6321,N_5284,N_5729);
xnor U6322 (N_6322,N_5258,N_5684);
xnor U6323 (N_6323,N_5420,N_5860);
nand U6324 (N_6324,N_5557,N_5387);
nand U6325 (N_6325,N_5456,N_5487);
or U6326 (N_6326,N_5513,N_5832);
nor U6327 (N_6327,N_5508,N_5654);
nor U6328 (N_6328,N_5259,N_5622);
nor U6329 (N_6329,N_5831,N_5952);
nand U6330 (N_6330,N_5899,N_5715);
and U6331 (N_6331,N_5870,N_5844);
nand U6332 (N_6332,N_5804,N_5727);
and U6333 (N_6333,N_5375,N_5879);
or U6334 (N_6334,N_5295,N_5454);
nor U6335 (N_6335,N_5567,N_5439);
and U6336 (N_6336,N_5292,N_5509);
or U6337 (N_6337,N_5588,N_5635);
nand U6338 (N_6338,N_5305,N_5504);
xnor U6339 (N_6339,N_5570,N_5720);
nand U6340 (N_6340,N_5527,N_5541);
and U6341 (N_6341,N_5303,N_5974);
and U6342 (N_6342,N_5386,N_5921);
and U6343 (N_6343,N_5800,N_5820);
and U6344 (N_6344,N_5520,N_5417);
xor U6345 (N_6345,N_5321,N_5649);
or U6346 (N_6346,N_5785,N_5643);
or U6347 (N_6347,N_5554,N_5760);
or U6348 (N_6348,N_5911,N_5450);
and U6349 (N_6349,N_5308,N_5751);
nor U6350 (N_6350,N_5409,N_5443);
and U6351 (N_6351,N_5888,N_5692);
or U6352 (N_6352,N_5318,N_5855);
nor U6353 (N_6353,N_5529,N_5602);
and U6354 (N_6354,N_5728,N_5781);
or U6355 (N_6355,N_5472,N_5350);
and U6356 (N_6356,N_5256,N_5442);
or U6357 (N_6357,N_5967,N_5869);
nand U6358 (N_6358,N_5742,N_5593);
xnor U6359 (N_6359,N_5422,N_5930);
nor U6360 (N_6360,N_5437,N_5440);
nor U6361 (N_6361,N_5874,N_5984);
nand U6362 (N_6362,N_5811,N_5786);
or U6363 (N_6363,N_5919,N_5572);
nor U6364 (N_6364,N_5597,N_5822);
nor U6365 (N_6365,N_5253,N_5891);
and U6366 (N_6366,N_5933,N_5905);
nand U6367 (N_6367,N_5702,N_5543);
and U6368 (N_6368,N_5755,N_5631);
nor U6369 (N_6369,N_5902,N_5988);
and U6370 (N_6370,N_5270,N_5625);
nor U6371 (N_6371,N_5864,N_5474);
and U6372 (N_6372,N_5608,N_5283);
nor U6373 (N_6373,N_5623,N_5586);
and U6374 (N_6374,N_5971,N_5451);
nor U6375 (N_6375,N_5821,N_5452);
xnor U6376 (N_6376,N_5875,N_5472);
nand U6377 (N_6377,N_5436,N_5757);
nand U6378 (N_6378,N_5747,N_5574);
and U6379 (N_6379,N_5703,N_5758);
or U6380 (N_6380,N_5825,N_5670);
or U6381 (N_6381,N_5507,N_5790);
and U6382 (N_6382,N_5483,N_5469);
xnor U6383 (N_6383,N_5634,N_5967);
and U6384 (N_6384,N_5285,N_5984);
and U6385 (N_6385,N_5430,N_5900);
and U6386 (N_6386,N_5925,N_5253);
xnor U6387 (N_6387,N_5466,N_5684);
nor U6388 (N_6388,N_5675,N_5302);
nor U6389 (N_6389,N_5355,N_5882);
and U6390 (N_6390,N_5470,N_5282);
or U6391 (N_6391,N_5308,N_5510);
and U6392 (N_6392,N_5769,N_5348);
xnor U6393 (N_6393,N_5552,N_5734);
nand U6394 (N_6394,N_5563,N_5508);
xor U6395 (N_6395,N_5386,N_5422);
or U6396 (N_6396,N_5962,N_5848);
nor U6397 (N_6397,N_5606,N_5974);
and U6398 (N_6398,N_5393,N_5576);
and U6399 (N_6399,N_5565,N_5974);
and U6400 (N_6400,N_5448,N_5675);
nand U6401 (N_6401,N_5974,N_5889);
nand U6402 (N_6402,N_5882,N_5771);
and U6403 (N_6403,N_5756,N_5738);
or U6404 (N_6404,N_5325,N_5957);
and U6405 (N_6405,N_5957,N_5460);
nor U6406 (N_6406,N_5263,N_5634);
and U6407 (N_6407,N_5424,N_5549);
nor U6408 (N_6408,N_5367,N_5328);
nor U6409 (N_6409,N_5660,N_5364);
xnor U6410 (N_6410,N_5930,N_5987);
nand U6411 (N_6411,N_5939,N_5322);
and U6412 (N_6412,N_5954,N_5660);
nor U6413 (N_6413,N_5568,N_5908);
xor U6414 (N_6414,N_5900,N_5713);
or U6415 (N_6415,N_5333,N_5407);
or U6416 (N_6416,N_5615,N_5901);
and U6417 (N_6417,N_5693,N_5720);
xor U6418 (N_6418,N_5388,N_5635);
or U6419 (N_6419,N_5768,N_5402);
and U6420 (N_6420,N_5956,N_5531);
or U6421 (N_6421,N_5835,N_5706);
nor U6422 (N_6422,N_5822,N_5579);
or U6423 (N_6423,N_5515,N_5400);
xnor U6424 (N_6424,N_5560,N_5859);
or U6425 (N_6425,N_5659,N_5384);
nor U6426 (N_6426,N_5870,N_5742);
xor U6427 (N_6427,N_5451,N_5763);
nand U6428 (N_6428,N_5379,N_5499);
nand U6429 (N_6429,N_5483,N_5819);
nor U6430 (N_6430,N_5521,N_5454);
nor U6431 (N_6431,N_5945,N_5275);
or U6432 (N_6432,N_5997,N_5451);
and U6433 (N_6433,N_5839,N_5754);
nand U6434 (N_6434,N_5578,N_5746);
and U6435 (N_6435,N_5863,N_5445);
and U6436 (N_6436,N_5457,N_5624);
nor U6437 (N_6437,N_5683,N_5917);
nor U6438 (N_6438,N_5468,N_5335);
nor U6439 (N_6439,N_5449,N_5318);
and U6440 (N_6440,N_5555,N_5347);
nor U6441 (N_6441,N_5457,N_5600);
and U6442 (N_6442,N_5402,N_5867);
nor U6443 (N_6443,N_5541,N_5629);
nor U6444 (N_6444,N_5928,N_5967);
nand U6445 (N_6445,N_5872,N_5823);
nor U6446 (N_6446,N_5421,N_5541);
nor U6447 (N_6447,N_5689,N_5569);
nand U6448 (N_6448,N_5748,N_5812);
nand U6449 (N_6449,N_5655,N_5630);
xor U6450 (N_6450,N_5728,N_5567);
or U6451 (N_6451,N_5298,N_5740);
and U6452 (N_6452,N_5359,N_5730);
nor U6453 (N_6453,N_5595,N_5274);
nand U6454 (N_6454,N_5832,N_5323);
nor U6455 (N_6455,N_5849,N_5855);
xnor U6456 (N_6456,N_5332,N_5500);
and U6457 (N_6457,N_5434,N_5298);
or U6458 (N_6458,N_5820,N_5554);
and U6459 (N_6459,N_5642,N_5324);
and U6460 (N_6460,N_5594,N_5925);
xor U6461 (N_6461,N_5843,N_5982);
nand U6462 (N_6462,N_5766,N_5284);
xor U6463 (N_6463,N_5360,N_5461);
nand U6464 (N_6464,N_5690,N_5947);
and U6465 (N_6465,N_5647,N_5365);
xor U6466 (N_6466,N_5438,N_5514);
nor U6467 (N_6467,N_5883,N_5434);
xnor U6468 (N_6468,N_5663,N_5581);
and U6469 (N_6469,N_5608,N_5327);
nor U6470 (N_6470,N_5534,N_5294);
nand U6471 (N_6471,N_5884,N_5300);
xnor U6472 (N_6472,N_5809,N_5851);
or U6473 (N_6473,N_5423,N_5567);
xnor U6474 (N_6474,N_5552,N_5510);
or U6475 (N_6475,N_5717,N_5537);
and U6476 (N_6476,N_5673,N_5394);
xnor U6477 (N_6477,N_5284,N_5753);
nand U6478 (N_6478,N_5874,N_5367);
nand U6479 (N_6479,N_5377,N_5650);
xor U6480 (N_6480,N_5462,N_5571);
xnor U6481 (N_6481,N_5755,N_5531);
or U6482 (N_6482,N_5742,N_5441);
and U6483 (N_6483,N_5807,N_5654);
xor U6484 (N_6484,N_5755,N_5487);
xor U6485 (N_6485,N_5646,N_5648);
and U6486 (N_6486,N_5438,N_5783);
nor U6487 (N_6487,N_5881,N_5417);
and U6488 (N_6488,N_5389,N_5484);
nand U6489 (N_6489,N_5320,N_5311);
nor U6490 (N_6490,N_5501,N_5459);
xnor U6491 (N_6491,N_5954,N_5460);
nand U6492 (N_6492,N_5259,N_5976);
xnor U6493 (N_6493,N_5616,N_5263);
xor U6494 (N_6494,N_5501,N_5433);
nor U6495 (N_6495,N_5799,N_5827);
nand U6496 (N_6496,N_5517,N_5635);
nand U6497 (N_6497,N_5430,N_5418);
and U6498 (N_6498,N_5731,N_5642);
nand U6499 (N_6499,N_5359,N_5312);
and U6500 (N_6500,N_5360,N_5939);
nand U6501 (N_6501,N_5273,N_5525);
and U6502 (N_6502,N_5853,N_5368);
xor U6503 (N_6503,N_5809,N_5994);
or U6504 (N_6504,N_5815,N_5252);
and U6505 (N_6505,N_5666,N_5843);
nand U6506 (N_6506,N_5423,N_5788);
nand U6507 (N_6507,N_5584,N_5497);
nand U6508 (N_6508,N_5968,N_5328);
nor U6509 (N_6509,N_5701,N_5535);
nor U6510 (N_6510,N_5853,N_5915);
nor U6511 (N_6511,N_5312,N_5859);
or U6512 (N_6512,N_5496,N_5675);
and U6513 (N_6513,N_5826,N_5824);
nand U6514 (N_6514,N_5994,N_5882);
nor U6515 (N_6515,N_5519,N_5259);
nand U6516 (N_6516,N_5512,N_5473);
or U6517 (N_6517,N_5657,N_5770);
and U6518 (N_6518,N_5319,N_5900);
and U6519 (N_6519,N_5590,N_5731);
or U6520 (N_6520,N_5714,N_5563);
and U6521 (N_6521,N_5789,N_5300);
nor U6522 (N_6522,N_5644,N_5404);
nand U6523 (N_6523,N_5959,N_5561);
or U6524 (N_6524,N_5280,N_5716);
xnor U6525 (N_6525,N_5260,N_5990);
xnor U6526 (N_6526,N_5978,N_5667);
xnor U6527 (N_6527,N_5403,N_5498);
or U6528 (N_6528,N_5569,N_5657);
nor U6529 (N_6529,N_5933,N_5732);
and U6530 (N_6530,N_5700,N_5816);
nand U6531 (N_6531,N_5890,N_5586);
nor U6532 (N_6532,N_5467,N_5778);
nand U6533 (N_6533,N_5467,N_5265);
nand U6534 (N_6534,N_5871,N_5461);
nor U6535 (N_6535,N_5471,N_5368);
or U6536 (N_6536,N_5972,N_5879);
nand U6537 (N_6537,N_5456,N_5969);
nand U6538 (N_6538,N_5874,N_5919);
or U6539 (N_6539,N_5474,N_5622);
and U6540 (N_6540,N_5270,N_5464);
xor U6541 (N_6541,N_5945,N_5344);
or U6542 (N_6542,N_5891,N_5888);
or U6543 (N_6543,N_5300,N_5538);
xor U6544 (N_6544,N_5675,N_5622);
xnor U6545 (N_6545,N_5980,N_5313);
and U6546 (N_6546,N_5791,N_5362);
or U6547 (N_6547,N_5405,N_5438);
and U6548 (N_6548,N_5792,N_5491);
nor U6549 (N_6549,N_5351,N_5815);
nor U6550 (N_6550,N_5651,N_5279);
nand U6551 (N_6551,N_5790,N_5952);
xor U6552 (N_6552,N_5976,N_5253);
nand U6553 (N_6553,N_5383,N_5750);
or U6554 (N_6554,N_5436,N_5742);
or U6555 (N_6555,N_5291,N_5985);
nor U6556 (N_6556,N_5723,N_5668);
and U6557 (N_6557,N_5982,N_5924);
and U6558 (N_6558,N_5904,N_5442);
and U6559 (N_6559,N_5712,N_5261);
nor U6560 (N_6560,N_5958,N_5886);
and U6561 (N_6561,N_5994,N_5716);
or U6562 (N_6562,N_5565,N_5458);
nor U6563 (N_6563,N_5374,N_5289);
nand U6564 (N_6564,N_5505,N_5552);
or U6565 (N_6565,N_5318,N_5893);
and U6566 (N_6566,N_5395,N_5806);
xnor U6567 (N_6567,N_5862,N_5317);
and U6568 (N_6568,N_5600,N_5679);
nand U6569 (N_6569,N_5518,N_5640);
or U6570 (N_6570,N_5532,N_5323);
and U6571 (N_6571,N_5447,N_5803);
nor U6572 (N_6572,N_5523,N_5487);
nor U6573 (N_6573,N_5464,N_5300);
or U6574 (N_6574,N_5559,N_5913);
nand U6575 (N_6575,N_5698,N_5554);
nand U6576 (N_6576,N_5948,N_5576);
nand U6577 (N_6577,N_5574,N_5816);
and U6578 (N_6578,N_5433,N_5927);
xnor U6579 (N_6579,N_5954,N_5566);
and U6580 (N_6580,N_5443,N_5696);
or U6581 (N_6581,N_5354,N_5823);
and U6582 (N_6582,N_5254,N_5870);
xor U6583 (N_6583,N_5361,N_5805);
nor U6584 (N_6584,N_5251,N_5642);
nor U6585 (N_6585,N_5498,N_5288);
xor U6586 (N_6586,N_5844,N_5455);
nand U6587 (N_6587,N_5576,N_5805);
or U6588 (N_6588,N_5540,N_5938);
nor U6589 (N_6589,N_5531,N_5298);
nand U6590 (N_6590,N_5818,N_5862);
or U6591 (N_6591,N_5879,N_5585);
xnor U6592 (N_6592,N_5917,N_5884);
xnor U6593 (N_6593,N_5501,N_5526);
xnor U6594 (N_6594,N_5493,N_5710);
or U6595 (N_6595,N_5438,N_5897);
xnor U6596 (N_6596,N_5490,N_5537);
xnor U6597 (N_6597,N_5981,N_5499);
nand U6598 (N_6598,N_5394,N_5342);
nand U6599 (N_6599,N_5780,N_5303);
nor U6600 (N_6600,N_5676,N_5691);
xnor U6601 (N_6601,N_5798,N_5974);
nor U6602 (N_6602,N_5595,N_5419);
nand U6603 (N_6603,N_5424,N_5376);
or U6604 (N_6604,N_5638,N_5505);
nand U6605 (N_6605,N_5977,N_5523);
nand U6606 (N_6606,N_5825,N_5645);
or U6607 (N_6607,N_5589,N_5972);
or U6608 (N_6608,N_5532,N_5812);
or U6609 (N_6609,N_5344,N_5427);
or U6610 (N_6610,N_5577,N_5389);
xnor U6611 (N_6611,N_5828,N_5569);
or U6612 (N_6612,N_5691,N_5474);
xor U6613 (N_6613,N_5493,N_5643);
nand U6614 (N_6614,N_5290,N_5641);
and U6615 (N_6615,N_5337,N_5356);
nand U6616 (N_6616,N_5550,N_5488);
nand U6617 (N_6617,N_5846,N_5432);
xor U6618 (N_6618,N_5510,N_5389);
and U6619 (N_6619,N_5939,N_5586);
xnor U6620 (N_6620,N_5523,N_5779);
nand U6621 (N_6621,N_5589,N_5821);
or U6622 (N_6622,N_5883,N_5576);
or U6623 (N_6623,N_5790,N_5723);
or U6624 (N_6624,N_5713,N_5854);
nor U6625 (N_6625,N_5756,N_5375);
nor U6626 (N_6626,N_5825,N_5440);
and U6627 (N_6627,N_5857,N_5928);
nor U6628 (N_6628,N_5795,N_5818);
and U6629 (N_6629,N_5502,N_5749);
and U6630 (N_6630,N_5796,N_5324);
nor U6631 (N_6631,N_5989,N_5988);
and U6632 (N_6632,N_5926,N_5572);
or U6633 (N_6633,N_5631,N_5368);
nor U6634 (N_6634,N_5940,N_5631);
nand U6635 (N_6635,N_5880,N_5359);
and U6636 (N_6636,N_5888,N_5696);
xor U6637 (N_6637,N_5955,N_5929);
or U6638 (N_6638,N_5799,N_5676);
and U6639 (N_6639,N_5270,N_5532);
xor U6640 (N_6640,N_5345,N_5987);
xnor U6641 (N_6641,N_5542,N_5298);
nand U6642 (N_6642,N_5983,N_5548);
and U6643 (N_6643,N_5613,N_5320);
or U6644 (N_6644,N_5392,N_5267);
nor U6645 (N_6645,N_5538,N_5643);
nand U6646 (N_6646,N_5694,N_5908);
xnor U6647 (N_6647,N_5301,N_5730);
xnor U6648 (N_6648,N_5602,N_5324);
and U6649 (N_6649,N_5440,N_5750);
nor U6650 (N_6650,N_5432,N_5609);
nor U6651 (N_6651,N_5371,N_5514);
or U6652 (N_6652,N_5271,N_5543);
nor U6653 (N_6653,N_5360,N_5595);
xor U6654 (N_6654,N_5853,N_5979);
and U6655 (N_6655,N_5954,N_5900);
nand U6656 (N_6656,N_5441,N_5891);
and U6657 (N_6657,N_5659,N_5488);
nand U6658 (N_6658,N_5489,N_5768);
nor U6659 (N_6659,N_5848,N_5900);
nand U6660 (N_6660,N_5330,N_5581);
nor U6661 (N_6661,N_5855,N_5749);
nand U6662 (N_6662,N_5506,N_5281);
or U6663 (N_6663,N_5673,N_5596);
or U6664 (N_6664,N_5577,N_5964);
xnor U6665 (N_6665,N_5561,N_5781);
nor U6666 (N_6666,N_5319,N_5377);
or U6667 (N_6667,N_5927,N_5850);
xor U6668 (N_6668,N_5305,N_5464);
and U6669 (N_6669,N_5775,N_5357);
or U6670 (N_6670,N_5881,N_5321);
nand U6671 (N_6671,N_5765,N_5430);
nor U6672 (N_6672,N_5876,N_5378);
nand U6673 (N_6673,N_5342,N_5962);
xor U6674 (N_6674,N_5474,N_5280);
nor U6675 (N_6675,N_5609,N_5964);
nand U6676 (N_6676,N_5446,N_5739);
xor U6677 (N_6677,N_5758,N_5402);
and U6678 (N_6678,N_5376,N_5998);
nand U6679 (N_6679,N_5582,N_5468);
or U6680 (N_6680,N_5621,N_5425);
nor U6681 (N_6681,N_5524,N_5626);
and U6682 (N_6682,N_5404,N_5713);
xor U6683 (N_6683,N_5495,N_5437);
nor U6684 (N_6684,N_5297,N_5849);
xnor U6685 (N_6685,N_5492,N_5881);
nand U6686 (N_6686,N_5455,N_5945);
nand U6687 (N_6687,N_5289,N_5305);
nand U6688 (N_6688,N_5679,N_5628);
xnor U6689 (N_6689,N_5297,N_5453);
or U6690 (N_6690,N_5769,N_5566);
or U6691 (N_6691,N_5347,N_5906);
nand U6692 (N_6692,N_5349,N_5586);
xnor U6693 (N_6693,N_5751,N_5693);
or U6694 (N_6694,N_5961,N_5829);
xor U6695 (N_6695,N_5992,N_5553);
nand U6696 (N_6696,N_5563,N_5605);
xor U6697 (N_6697,N_5557,N_5708);
nand U6698 (N_6698,N_5945,N_5597);
nor U6699 (N_6699,N_5337,N_5909);
nor U6700 (N_6700,N_5873,N_5652);
nor U6701 (N_6701,N_5834,N_5487);
or U6702 (N_6702,N_5683,N_5674);
nor U6703 (N_6703,N_5501,N_5471);
nand U6704 (N_6704,N_5612,N_5903);
or U6705 (N_6705,N_5909,N_5911);
nand U6706 (N_6706,N_5778,N_5992);
nand U6707 (N_6707,N_5617,N_5697);
nand U6708 (N_6708,N_5659,N_5418);
xor U6709 (N_6709,N_5375,N_5302);
nor U6710 (N_6710,N_5914,N_5281);
nand U6711 (N_6711,N_5488,N_5802);
xnor U6712 (N_6712,N_5845,N_5266);
or U6713 (N_6713,N_5930,N_5956);
nand U6714 (N_6714,N_5991,N_5573);
xor U6715 (N_6715,N_5704,N_5864);
xnor U6716 (N_6716,N_5289,N_5927);
and U6717 (N_6717,N_5926,N_5630);
nand U6718 (N_6718,N_5604,N_5987);
or U6719 (N_6719,N_5691,N_5331);
or U6720 (N_6720,N_5268,N_5571);
nor U6721 (N_6721,N_5897,N_5551);
nor U6722 (N_6722,N_5428,N_5288);
or U6723 (N_6723,N_5527,N_5262);
nand U6724 (N_6724,N_5451,N_5538);
or U6725 (N_6725,N_5556,N_5279);
and U6726 (N_6726,N_5334,N_5268);
nand U6727 (N_6727,N_5963,N_5288);
and U6728 (N_6728,N_5647,N_5824);
or U6729 (N_6729,N_5992,N_5812);
and U6730 (N_6730,N_5484,N_5842);
or U6731 (N_6731,N_5674,N_5592);
xnor U6732 (N_6732,N_5701,N_5373);
nor U6733 (N_6733,N_5515,N_5800);
nor U6734 (N_6734,N_5250,N_5859);
nor U6735 (N_6735,N_5624,N_5502);
or U6736 (N_6736,N_5346,N_5442);
and U6737 (N_6737,N_5764,N_5408);
nor U6738 (N_6738,N_5261,N_5316);
xnor U6739 (N_6739,N_5276,N_5339);
xnor U6740 (N_6740,N_5965,N_5865);
xnor U6741 (N_6741,N_5467,N_5969);
nand U6742 (N_6742,N_5295,N_5997);
and U6743 (N_6743,N_5482,N_5970);
or U6744 (N_6744,N_5800,N_5845);
nor U6745 (N_6745,N_5584,N_5665);
or U6746 (N_6746,N_5901,N_5460);
nor U6747 (N_6747,N_5298,N_5867);
and U6748 (N_6748,N_5461,N_5678);
nand U6749 (N_6749,N_5732,N_5448);
nand U6750 (N_6750,N_6506,N_6582);
or U6751 (N_6751,N_6522,N_6235);
and U6752 (N_6752,N_6127,N_6330);
or U6753 (N_6753,N_6473,N_6301);
xnor U6754 (N_6754,N_6497,N_6526);
xor U6755 (N_6755,N_6270,N_6173);
nor U6756 (N_6756,N_6281,N_6385);
nor U6757 (N_6757,N_6575,N_6293);
xnor U6758 (N_6758,N_6300,N_6544);
nor U6759 (N_6759,N_6104,N_6248);
and U6760 (N_6760,N_6749,N_6653);
xor U6761 (N_6761,N_6186,N_6490);
and U6762 (N_6762,N_6311,N_6714);
and U6763 (N_6763,N_6643,N_6294);
nand U6764 (N_6764,N_6721,N_6552);
xor U6765 (N_6765,N_6456,N_6292);
nor U6766 (N_6766,N_6282,N_6010);
or U6767 (N_6767,N_6548,N_6433);
nand U6768 (N_6768,N_6727,N_6478);
xor U6769 (N_6769,N_6740,N_6629);
nand U6770 (N_6770,N_6233,N_6267);
xor U6771 (N_6771,N_6291,N_6567);
nand U6772 (N_6772,N_6082,N_6635);
and U6773 (N_6773,N_6482,N_6332);
xnor U6774 (N_6774,N_6670,N_6435);
nor U6775 (N_6775,N_6425,N_6346);
and U6776 (N_6776,N_6023,N_6373);
nand U6777 (N_6777,N_6144,N_6626);
nand U6778 (N_6778,N_6171,N_6241);
nand U6779 (N_6779,N_6296,N_6344);
xnor U6780 (N_6780,N_6187,N_6095);
nor U6781 (N_6781,N_6487,N_6299);
nor U6782 (N_6782,N_6628,N_6302);
nand U6783 (N_6783,N_6663,N_6045);
nand U6784 (N_6784,N_6091,N_6690);
and U6785 (N_6785,N_6021,N_6466);
and U6786 (N_6786,N_6258,N_6035);
xnor U6787 (N_6787,N_6207,N_6540);
nand U6788 (N_6788,N_6313,N_6122);
nand U6789 (N_6789,N_6170,N_6381);
nor U6790 (N_6790,N_6288,N_6659);
or U6791 (N_6791,N_6674,N_6504);
xor U6792 (N_6792,N_6115,N_6521);
and U6793 (N_6793,N_6362,N_6137);
or U6794 (N_6794,N_6649,N_6340);
or U6795 (N_6795,N_6725,N_6076);
nand U6796 (N_6796,N_6471,N_6185);
xnor U6797 (N_6797,N_6680,N_6246);
or U6798 (N_6798,N_6616,N_6275);
or U6799 (N_6799,N_6220,N_6215);
or U6800 (N_6800,N_6537,N_6426);
or U6801 (N_6801,N_6046,N_6372);
or U6802 (N_6802,N_6618,N_6297);
xnor U6803 (N_6803,N_6676,N_6534);
and U6804 (N_6804,N_6550,N_6577);
nand U6805 (N_6805,N_6324,N_6156);
or U6806 (N_6806,N_6198,N_6119);
nand U6807 (N_6807,N_6648,N_6142);
nand U6808 (N_6808,N_6056,N_6129);
nor U6809 (N_6809,N_6160,N_6025);
nand U6810 (N_6810,N_6625,N_6243);
nor U6811 (N_6811,N_6708,N_6084);
and U6812 (N_6812,N_6563,N_6146);
and U6813 (N_6813,N_6568,N_6510);
xnor U6814 (N_6814,N_6486,N_6274);
and U6815 (N_6815,N_6419,N_6431);
nand U6816 (N_6816,N_6543,N_6624);
nor U6817 (N_6817,N_6672,N_6650);
and U6818 (N_6818,N_6581,N_6099);
or U6819 (N_6819,N_6238,N_6304);
nor U6820 (N_6820,N_6579,N_6469);
nor U6821 (N_6821,N_6070,N_6283);
or U6822 (N_6822,N_6237,N_6354);
nor U6823 (N_6823,N_6605,N_6453);
and U6824 (N_6824,N_6610,N_6403);
or U6825 (N_6825,N_6081,N_6131);
xor U6826 (N_6826,N_6613,N_6062);
and U6827 (N_6827,N_6107,N_6517);
and U6828 (N_6828,N_6390,N_6150);
or U6829 (N_6829,N_6580,N_6097);
nand U6830 (N_6830,N_6361,N_6379);
nor U6831 (N_6831,N_6323,N_6639);
xnor U6832 (N_6832,N_6632,N_6422);
and U6833 (N_6833,N_6602,N_6094);
nor U6834 (N_6834,N_6406,N_6219);
xor U6835 (N_6835,N_6078,N_6303);
nand U6836 (N_6836,N_6008,N_6477);
nor U6837 (N_6837,N_6179,N_6047);
or U6838 (N_6838,N_6441,N_6016);
or U6839 (N_6839,N_6262,N_6054);
nor U6840 (N_6840,N_6587,N_6376);
nor U6841 (N_6841,N_6229,N_6140);
and U6842 (N_6842,N_6524,N_6704);
and U6843 (N_6843,N_6645,N_6199);
xnor U6844 (N_6844,N_6377,N_6416);
xnor U6845 (N_6845,N_6252,N_6384);
nor U6846 (N_6846,N_6226,N_6318);
xnor U6847 (N_6847,N_6528,N_6513);
and U6848 (N_6848,N_6359,N_6488);
nor U6849 (N_6849,N_6481,N_6247);
or U6850 (N_6850,N_6414,N_6652);
and U6851 (N_6851,N_6392,N_6741);
and U6852 (N_6852,N_6677,N_6204);
or U6853 (N_6853,N_6748,N_6216);
xor U6854 (N_6854,N_6511,N_6427);
and U6855 (N_6855,N_6742,N_6669);
nand U6856 (N_6856,N_6139,N_6462);
nor U6857 (N_6857,N_6161,N_6697);
nor U6858 (N_6858,N_6507,N_6128);
nor U6859 (N_6859,N_6604,N_6703);
nand U6860 (N_6860,N_6020,N_6136);
or U6861 (N_6861,N_6418,N_6553);
nor U6862 (N_6862,N_6467,N_6440);
and U6863 (N_6863,N_6284,N_6684);
nand U6864 (N_6864,N_6729,N_6638);
xor U6865 (N_6865,N_6028,N_6598);
and U6866 (N_6866,N_6201,N_6449);
or U6867 (N_6867,N_6182,N_6155);
nand U6868 (N_6868,N_6105,N_6202);
or U6869 (N_6869,N_6048,N_6413);
xnor U6870 (N_6870,N_6230,N_6739);
xor U6871 (N_6871,N_6662,N_6085);
xnor U6872 (N_6872,N_6114,N_6306);
or U6873 (N_6873,N_6334,N_6514);
nand U6874 (N_6874,N_6080,N_6523);
xor U6875 (N_6875,N_6367,N_6269);
and U6876 (N_6876,N_6336,N_6126);
nand U6877 (N_6877,N_6730,N_6738);
nand U6878 (N_6878,N_6231,N_6152);
or U6879 (N_6879,N_6501,N_6393);
and U6880 (N_6880,N_6196,N_6460);
and U6881 (N_6881,N_6244,N_6656);
xnor U6882 (N_6882,N_6211,N_6387);
nand U6883 (N_6883,N_6133,N_6055);
nand U6884 (N_6884,N_6208,N_6205);
nor U6885 (N_6885,N_6256,N_6718);
nor U6886 (N_6886,N_6546,N_6003);
and U6887 (N_6887,N_6264,N_6265);
or U6888 (N_6888,N_6287,N_6436);
or U6889 (N_6889,N_6484,N_6063);
nor U6890 (N_6890,N_6743,N_6675);
nor U6891 (N_6891,N_6509,N_6745);
nor U6892 (N_6892,N_6308,N_6319);
or U6893 (N_6893,N_6578,N_6559);
nor U6894 (N_6894,N_6341,N_6423);
or U6895 (N_6895,N_6640,N_6443);
and U6896 (N_6896,N_6574,N_6371);
xnor U6897 (N_6897,N_6496,N_6668);
and U6898 (N_6898,N_6556,N_6206);
or U6899 (N_6899,N_6615,N_6386);
or U6900 (N_6900,N_6147,N_6213);
nor U6901 (N_6901,N_6679,N_6013);
nand U6902 (N_6902,N_6090,N_6183);
or U6903 (N_6903,N_6554,N_6011);
xor U6904 (N_6904,N_6251,N_6465);
or U6905 (N_6905,N_6576,N_6221);
and U6906 (N_6906,N_6695,N_6451);
or U6907 (N_6907,N_6461,N_6454);
xnor U6908 (N_6908,N_6508,N_6395);
and U6909 (N_6909,N_6163,N_6002);
nand U6910 (N_6910,N_6545,N_6417);
nor U6911 (N_6911,N_6305,N_6603);
or U6912 (N_6912,N_6338,N_6253);
xor U6913 (N_6913,N_6405,N_6599);
nor U6914 (N_6914,N_6722,N_6190);
nand U6915 (N_6915,N_6322,N_6590);
xor U6916 (N_6916,N_6533,N_6001);
nor U6917 (N_6917,N_6606,N_6087);
and U6918 (N_6918,N_6660,N_6498);
nand U6919 (N_6919,N_6701,N_6569);
or U6920 (N_6920,N_6040,N_6240);
nand U6921 (N_6921,N_6271,N_6597);
nor U6922 (N_6922,N_6588,N_6203);
nor U6923 (N_6923,N_6223,N_6685);
or U6924 (N_6924,N_6525,N_6682);
nor U6925 (N_6925,N_6434,N_6382);
or U6926 (N_6926,N_6154,N_6560);
xor U6927 (N_6927,N_6027,N_6447);
or U6928 (N_6928,N_6476,N_6194);
xnor U6929 (N_6929,N_6491,N_6505);
and U6930 (N_6930,N_6014,N_6214);
nand U6931 (N_6931,N_6036,N_6375);
xnor U6932 (N_6932,N_6723,N_6290);
nor U6933 (N_6933,N_6420,N_6734);
and U6934 (N_6934,N_6254,N_6052);
nor U6935 (N_6935,N_6112,N_6641);
nor U6936 (N_6936,N_6479,N_6736);
xor U6937 (N_6937,N_6744,N_6396);
and U6938 (N_6938,N_6289,N_6709);
or U6939 (N_6939,N_6596,N_6153);
and U6940 (N_6940,N_6631,N_6474);
or U6941 (N_6941,N_6307,N_6584);
and U6942 (N_6942,N_6032,N_6493);
or U6943 (N_6943,N_6452,N_6539);
nand U6944 (N_6944,N_6457,N_6728);
nor U6945 (N_6945,N_6132,N_6746);
or U6946 (N_6946,N_6071,N_6268);
xnor U6947 (N_6947,N_6633,N_6589);
and U6948 (N_6948,N_6125,N_6145);
and U6949 (N_6949,N_6494,N_6180);
or U6950 (N_6950,N_6627,N_6165);
nor U6951 (N_6951,N_6100,N_6261);
xor U6952 (N_6952,N_6391,N_6034);
nor U6953 (N_6953,N_6364,N_6162);
and U6954 (N_6954,N_6279,N_6571);
xnor U6955 (N_6955,N_6184,N_6059);
or U6956 (N_6956,N_6459,N_6077);
and U6957 (N_6957,N_6366,N_6532);
and U6958 (N_6958,N_6458,N_6079);
xor U6959 (N_6959,N_6043,N_6121);
nor U6960 (N_6960,N_6072,N_6030);
or U6961 (N_6961,N_6278,N_6402);
nand U6962 (N_6962,N_6655,N_6029);
nor U6963 (N_6963,N_6061,N_6620);
nor U6964 (N_6964,N_6464,N_6239);
or U6965 (N_6965,N_6661,N_6315);
xor U6966 (N_6966,N_6647,N_6169);
or U6967 (N_6967,N_6617,N_6412);
xor U6968 (N_6968,N_6065,N_6410);
and U6969 (N_6969,N_6446,N_6673);
or U6970 (N_6970,N_6358,N_6158);
or U6971 (N_6971,N_6123,N_6717);
nand U6972 (N_6972,N_6593,N_6693);
and U6973 (N_6973,N_6424,N_6678);
nand U6974 (N_6974,N_6686,N_6192);
and U6975 (N_6975,N_6585,N_6594);
nor U6976 (N_6976,N_6073,N_6619);
nor U6977 (N_6977,N_6189,N_6110);
nor U6978 (N_6978,N_6263,N_6168);
nor U6979 (N_6979,N_6033,N_6172);
or U6980 (N_6980,N_6445,N_6705);
or U6981 (N_6981,N_6383,N_6562);
or U6982 (N_6982,N_6657,N_6148);
nand U6983 (N_6983,N_6024,N_6691);
nand U6984 (N_6984,N_6707,N_6159);
and U6985 (N_6985,N_6428,N_6609);
nand U6986 (N_6986,N_6731,N_6694);
and U6987 (N_6987,N_6113,N_6542);
nand U6988 (N_6988,N_6310,N_6512);
nand U6989 (N_6989,N_6176,N_6549);
nor U6990 (N_6990,N_6621,N_6096);
xnor U6991 (N_6991,N_6711,N_6018);
xor U6992 (N_6992,N_6167,N_6053);
nor U6993 (N_6993,N_6634,N_6450);
xnor U6994 (N_6994,N_6463,N_6710);
and U6995 (N_6995,N_6566,N_6555);
nand U6996 (N_6996,N_6667,N_6408);
nand U6997 (N_6997,N_6351,N_6726);
and U6998 (N_6998,N_6050,N_6692);
nor U6999 (N_6999,N_6044,N_6195);
or U7000 (N_7000,N_6236,N_6503);
nor U7001 (N_7001,N_6502,N_6337);
nor U7002 (N_7002,N_6353,N_6051);
xnor U7003 (N_7003,N_6026,N_6345);
nor U7004 (N_7004,N_6623,N_6733);
or U7005 (N_7005,N_6432,N_6389);
and U7006 (N_7006,N_6535,N_6329);
nor U7007 (N_7007,N_6320,N_6374);
or U7008 (N_7008,N_6356,N_6074);
nor U7009 (N_7009,N_6388,N_6489);
and U7010 (N_7010,N_6088,N_6342);
or U7011 (N_7011,N_6312,N_6516);
nand U7012 (N_7012,N_6259,N_6280);
xor U7013 (N_7013,N_6518,N_6538);
nor U7014 (N_7014,N_6644,N_6378);
or U7015 (N_7015,N_6530,N_6004);
xnor U7016 (N_7016,N_6595,N_6057);
nand U7017 (N_7017,N_6309,N_6191);
and U7018 (N_7018,N_6564,N_6702);
nand U7019 (N_7019,N_6098,N_6515);
nor U7020 (N_7020,N_6520,N_6257);
or U7021 (N_7021,N_6651,N_6531);
xnor U7022 (N_7022,N_6225,N_6485);
or U7023 (N_7023,N_6227,N_6706);
xor U7024 (N_7024,N_6671,N_6242);
and U7025 (N_7025,N_6689,N_6699);
or U7026 (N_7026,N_6472,N_6086);
nand U7027 (N_7027,N_6608,N_6688);
xor U7028 (N_7028,N_6437,N_6232);
or U7029 (N_7029,N_6732,N_6012);
nand U7030 (N_7030,N_6298,N_6715);
nand U7031 (N_7031,N_6335,N_6017);
nor U7032 (N_7032,N_6347,N_6212);
nor U7033 (N_7033,N_6558,N_6681);
xnor U7034 (N_7034,N_6005,N_6277);
xnor U7035 (N_7035,N_6069,N_6266);
or U7036 (N_7036,N_6181,N_6720);
nand U7037 (N_7037,N_6586,N_6536);
nor U7038 (N_7038,N_6622,N_6222);
xor U7039 (N_7039,N_6666,N_6327);
and U7040 (N_7040,N_6075,N_6134);
nor U7041 (N_7041,N_6480,N_6111);
or U7042 (N_7042,N_6716,N_6583);
nand U7043 (N_7043,N_6719,N_6089);
nor U7044 (N_7044,N_6325,N_6394);
xor U7045 (N_7045,N_6570,N_6735);
or U7046 (N_7046,N_6646,N_6500);
nand U7047 (N_7047,N_6316,N_6495);
or U7048 (N_7048,N_6350,N_6151);
nor U7049 (N_7049,N_6409,N_6331);
and U7050 (N_7050,N_6698,N_6022);
nand U7051 (N_7051,N_6038,N_6665);
xor U7052 (N_7052,N_6355,N_6295);
xnor U7053 (N_7053,N_6724,N_6529);
xnor U7054 (N_7054,N_6245,N_6360);
nand U7055 (N_7055,N_6178,N_6737);
nand U7056 (N_7056,N_6228,N_6224);
and U7057 (N_7057,N_6565,N_6333);
and U7058 (N_7058,N_6541,N_6200);
or U7059 (N_7059,N_6499,N_6166);
or U7060 (N_7060,N_6064,N_6209);
xnor U7061 (N_7061,N_6234,N_6093);
and U7062 (N_7062,N_6572,N_6400);
nand U7063 (N_7063,N_6015,N_6109);
nor U7064 (N_7064,N_6118,N_6066);
xnor U7065 (N_7065,N_6009,N_6141);
and U7066 (N_7066,N_6272,N_6120);
nand U7067 (N_7067,N_6600,N_6415);
nor U7068 (N_7068,N_6328,N_6135);
nand U7069 (N_7069,N_6547,N_6658);
and U7070 (N_7070,N_6039,N_6713);
nor U7071 (N_7071,N_6398,N_6654);
xnor U7072 (N_7072,N_6116,N_6607);
xor U7073 (N_7073,N_6217,N_6164);
xor U7074 (N_7074,N_6285,N_6614);
and U7075 (N_7075,N_6326,N_6642);
nand U7076 (N_7076,N_6037,N_6317);
xnor U7077 (N_7077,N_6175,N_6276);
nor U7078 (N_7078,N_6149,N_6444);
xnor U7079 (N_7079,N_6399,N_6106);
and U7080 (N_7080,N_6712,N_6700);
and U7081 (N_7081,N_6058,N_6101);
and U7082 (N_7082,N_6000,N_6411);
xnor U7083 (N_7083,N_6468,N_6348);
nand U7084 (N_7084,N_6470,N_6060);
nand U7085 (N_7085,N_6430,N_6250);
and U7086 (N_7086,N_6687,N_6188);
xor U7087 (N_7087,N_6343,N_6273);
nand U7088 (N_7088,N_6124,N_6401);
or U7089 (N_7089,N_6519,N_6321);
and U7090 (N_7090,N_6601,N_6630);
nand U7091 (N_7091,N_6557,N_6103);
or U7092 (N_7092,N_6157,N_6130);
nor U7093 (N_7093,N_6747,N_6429);
and U7094 (N_7094,N_6218,N_6019);
nor U7095 (N_7095,N_6174,N_6592);
xnor U7096 (N_7096,N_6696,N_6007);
and U7097 (N_7097,N_6404,N_6031);
and U7098 (N_7098,N_6439,N_6455);
nand U7099 (N_7099,N_6255,N_6314);
nor U7100 (N_7100,N_6397,N_6357);
or U7101 (N_7101,N_6102,N_6483);
or U7102 (N_7102,N_6193,N_6380);
nand U7103 (N_7103,N_6368,N_6138);
nor U7104 (N_7104,N_6365,N_6352);
nand U7105 (N_7105,N_6177,N_6197);
nand U7106 (N_7106,N_6527,N_6573);
and U7107 (N_7107,N_6369,N_6339);
and U7108 (N_7108,N_6286,N_6083);
nand U7109 (N_7109,N_6249,N_6683);
nand U7110 (N_7110,N_6092,N_6042);
and U7111 (N_7111,N_6067,N_6442);
nand U7112 (N_7112,N_6448,N_6108);
xor U7113 (N_7113,N_6637,N_6049);
nand U7114 (N_7114,N_6370,N_6664);
xor U7115 (N_7115,N_6041,N_6551);
or U7116 (N_7116,N_6363,N_6612);
nor U7117 (N_7117,N_6421,N_6349);
xor U7118 (N_7118,N_6210,N_6611);
nand U7119 (N_7119,N_6475,N_6438);
xor U7120 (N_7120,N_6006,N_6636);
xnor U7121 (N_7121,N_6492,N_6407);
nor U7122 (N_7122,N_6117,N_6143);
xor U7123 (N_7123,N_6068,N_6260);
nor U7124 (N_7124,N_6591,N_6561);
xnor U7125 (N_7125,N_6121,N_6552);
nand U7126 (N_7126,N_6599,N_6704);
xnor U7127 (N_7127,N_6164,N_6081);
and U7128 (N_7128,N_6087,N_6051);
nor U7129 (N_7129,N_6376,N_6022);
and U7130 (N_7130,N_6560,N_6061);
xor U7131 (N_7131,N_6299,N_6657);
nor U7132 (N_7132,N_6653,N_6403);
nor U7133 (N_7133,N_6495,N_6107);
xor U7134 (N_7134,N_6227,N_6327);
or U7135 (N_7135,N_6102,N_6640);
nand U7136 (N_7136,N_6737,N_6463);
xor U7137 (N_7137,N_6533,N_6068);
or U7138 (N_7138,N_6279,N_6315);
or U7139 (N_7139,N_6406,N_6594);
nor U7140 (N_7140,N_6209,N_6048);
nand U7141 (N_7141,N_6416,N_6660);
nor U7142 (N_7142,N_6219,N_6091);
nor U7143 (N_7143,N_6330,N_6325);
xor U7144 (N_7144,N_6470,N_6521);
or U7145 (N_7145,N_6669,N_6399);
nand U7146 (N_7146,N_6264,N_6658);
and U7147 (N_7147,N_6086,N_6229);
nor U7148 (N_7148,N_6094,N_6587);
or U7149 (N_7149,N_6512,N_6087);
xnor U7150 (N_7150,N_6014,N_6583);
nor U7151 (N_7151,N_6280,N_6090);
xnor U7152 (N_7152,N_6373,N_6005);
nand U7153 (N_7153,N_6136,N_6140);
nand U7154 (N_7154,N_6156,N_6148);
or U7155 (N_7155,N_6702,N_6720);
nand U7156 (N_7156,N_6646,N_6692);
or U7157 (N_7157,N_6028,N_6429);
xor U7158 (N_7158,N_6128,N_6682);
xor U7159 (N_7159,N_6422,N_6095);
nor U7160 (N_7160,N_6013,N_6207);
and U7161 (N_7161,N_6305,N_6699);
xor U7162 (N_7162,N_6237,N_6084);
nor U7163 (N_7163,N_6516,N_6477);
nand U7164 (N_7164,N_6440,N_6117);
or U7165 (N_7165,N_6099,N_6316);
xor U7166 (N_7166,N_6010,N_6332);
nand U7167 (N_7167,N_6446,N_6159);
xnor U7168 (N_7168,N_6355,N_6538);
nor U7169 (N_7169,N_6673,N_6187);
nand U7170 (N_7170,N_6739,N_6211);
nor U7171 (N_7171,N_6071,N_6680);
xor U7172 (N_7172,N_6110,N_6023);
or U7173 (N_7173,N_6331,N_6232);
nand U7174 (N_7174,N_6233,N_6173);
nor U7175 (N_7175,N_6234,N_6121);
nor U7176 (N_7176,N_6434,N_6036);
or U7177 (N_7177,N_6055,N_6666);
xnor U7178 (N_7178,N_6570,N_6591);
nand U7179 (N_7179,N_6702,N_6032);
nand U7180 (N_7180,N_6228,N_6645);
and U7181 (N_7181,N_6687,N_6628);
xor U7182 (N_7182,N_6089,N_6360);
nor U7183 (N_7183,N_6020,N_6530);
or U7184 (N_7184,N_6402,N_6593);
or U7185 (N_7185,N_6551,N_6573);
and U7186 (N_7186,N_6162,N_6059);
or U7187 (N_7187,N_6298,N_6290);
xor U7188 (N_7188,N_6542,N_6098);
and U7189 (N_7189,N_6225,N_6533);
xor U7190 (N_7190,N_6335,N_6626);
nor U7191 (N_7191,N_6662,N_6515);
xor U7192 (N_7192,N_6495,N_6678);
and U7193 (N_7193,N_6499,N_6325);
or U7194 (N_7194,N_6210,N_6608);
nand U7195 (N_7195,N_6122,N_6232);
nand U7196 (N_7196,N_6135,N_6026);
nand U7197 (N_7197,N_6002,N_6206);
and U7198 (N_7198,N_6391,N_6551);
xor U7199 (N_7199,N_6019,N_6007);
and U7200 (N_7200,N_6514,N_6622);
xnor U7201 (N_7201,N_6530,N_6367);
and U7202 (N_7202,N_6745,N_6142);
and U7203 (N_7203,N_6295,N_6012);
nand U7204 (N_7204,N_6652,N_6726);
or U7205 (N_7205,N_6362,N_6731);
nand U7206 (N_7206,N_6096,N_6591);
xor U7207 (N_7207,N_6054,N_6605);
and U7208 (N_7208,N_6349,N_6338);
or U7209 (N_7209,N_6060,N_6650);
or U7210 (N_7210,N_6530,N_6090);
nor U7211 (N_7211,N_6740,N_6165);
xor U7212 (N_7212,N_6189,N_6681);
and U7213 (N_7213,N_6629,N_6226);
nand U7214 (N_7214,N_6207,N_6668);
nor U7215 (N_7215,N_6704,N_6228);
nand U7216 (N_7216,N_6029,N_6113);
nor U7217 (N_7217,N_6157,N_6154);
nand U7218 (N_7218,N_6157,N_6026);
xor U7219 (N_7219,N_6160,N_6353);
and U7220 (N_7220,N_6488,N_6442);
nor U7221 (N_7221,N_6359,N_6377);
nor U7222 (N_7222,N_6475,N_6213);
or U7223 (N_7223,N_6579,N_6104);
nor U7224 (N_7224,N_6424,N_6245);
xnor U7225 (N_7225,N_6636,N_6234);
nor U7226 (N_7226,N_6629,N_6698);
nand U7227 (N_7227,N_6597,N_6123);
or U7228 (N_7228,N_6502,N_6710);
and U7229 (N_7229,N_6115,N_6311);
xnor U7230 (N_7230,N_6681,N_6539);
nor U7231 (N_7231,N_6643,N_6121);
nor U7232 (N_7232,N_6321,N_6116);
or U7233 (N_7233,N_6555,N_6410);
xor U7234 (N_7234,N_6318,N_6282);
and U7235 (N_7235,N_6431,N_6586);
xnor U7236 (N_7236,N_6089,N_6283);
nand U7237 (N_7237,N_6030,N_6532);
xnor U7238 (N_7238,N_6449,N_6109);
nand U7239 (N_7239,N_6104,N_6172);
and U7240 (N_7240,N_6475,N_6476);
xnor U7241 (N_7241,N_6225,N_6691);
nand U7242 (N_7242,N_6584,N_6156);
nand U7243 (N_7243,N_6546,N_6443);
and U7244 (N_7244,N_6626,N_6257);
or U7245 (N_7245,N_6725,N_6738);
xor U7246 (N_7246,N_6589,N_6665);
nand U7247 (N_7247,N_6441,N_6715);
nand U7248 (N_7248,N_6127,N_6339);
nand U7249 (N_7249,N_6098,N_6506);
or U7250 (N_7250,N_6344,N_6621);
and U7251 (N_7251,N_6006,N_6292);
nor U7252 (N_7252,N_6023,N_6631);
xnor U7253 (N_7253,N_6614,N_6265);
xnor U7254 (N_7254,N_6406,N_6155);
xor U7255 (N_7255,N_6306,N_6498);
and U7256 (N_7256,N_6196,N_6301);
nand U7257 (N_7257,N_6226,N_6072);
or U7258 (N_7258,N_6099,N_6035);
nor U7259 (N_7259,N_6254,N_6061);
nor U7260 (N_7260,N_6642,N_6737);
nand U7261 (N_7261,N_6505,N_6437);
nand U7262 (N_7262,N_6066,N_6439);
nor U7263 (N_7263,N_6734,N_6095);
and U7264 (N_7264,N_6465,N_6424);
and U7265 (N_7265,N_6168,N_6169);
and U7266 (N_7266,N_6610,N_6053);
xor U7267 (N_7267,N_6173,N_6748);
nand U7268 (N_7268,N_6568,N_6152);
or U7269 (N_7269,N_6114,N_6307);
or U7270 (N_7270,N_6439,N_6743);
nor U7271 (N_7271,N_6645,N_6258);
xor U7272 (N_7272,N_6074,N_6487);
nand U7273 (N_7273,N_6154,N_6074);
nor U7274 (N_7274,N_6335,N_6382);
or U7275 (N_7275,N_6540,N_6488);
xnor U7276 (N_7276,N_6602,N_6721);
or U7277 (N_7277,N_6493,N_6707);
xnor U7278 (N_7278,N_6656,N_6063);
nor U7279 (N_7279,N_6654,N_6621);
nand U7280 (N_7280,N_6039,N_6716);
xor U7281 (N_7281,N_6171,N_6684);
or U7282 (N_7282,N_6007,N_6619);
or U7283 (N_7283,N_6206,N_6231);
and U7284 (N_7284,N_6158,N_6227);
and U7285 (N_7285,N_6014,N_6556);
or U7286 (N_7286,N_6682,N_6048);
and U7287 (N_7287,N_6592,N_6238);
nor U7288 (N_7288,N_6747,N_6374);
and U7289 (N_7289,N_6403,N_6702);
nand U7290 (N_7290,N_6172,N_6601);
xor U7291 (N_7291,N_6259,N_6119);
nor U7292 (N_7292,N_6601,N_6657);
and U7293 (N_7293,N_6683,N_6315);
and U7294 (N_7294,N_6698,N_6200);
or U7295 (N_7295,N_6083,N_6712);
nor U7296 (N_7296,N_6189,N_6697);
nor U7297 (N_7297,N_6073,N_6554);
nor U7298 (N_7298,N_6390,N_6357);
nor U7299 (N_7299,N_6486,N_6186);
and U7300 (N_7300,N_6551,N_6095);
nand U7301 (N_7301,N_6037,N_6435);
xnor U7302 (N_7302,N_6233,N_6552);
and U7303 (N_7303,N_6445,N_6332);
and U7304 (N_7304,N_6487,N_6670);
and U7305 (N_7305,N_6662,N_6331);
nor U7306 (N_7306,N_6387,N_6225);
and U7307 (N_7307,N_6291,N_6621);
and U7308 (N_7308,N_6284,N_6053);
and U7309 (N_7309,N_6433,N_6307);
xnor U7310 (N_7310,N_6237,N_6213);
and U7311 (N_7311,N_6274,N_6084);
or U7312 (N_7312,N_6394,N_6125);
xnor U7313 (N_7313,N_6160,N_6633);
or U7314 (N_7314,N_6418,N_6614);
nor U7315 (N_7315,N_6485,N_6176);
nand U7316 (N_7316,N_6260,N_6119);
and U7317 (N_7317,N_6093,N_6698);
xor U7318 (N_7318,N_6643,N_6088);
or U7319 (N_7319,N_6722,N_6165);
nor U7320 (N_7320,N_6040,N_6306);
nand U7321 (N_7321,N_6646,N_6540);
xnor U7322 (N_7322,N_6487,N_6409);
nor U7323 (N_7323,N_6612,N_6403);
and U7324 (N_7324,N_6227,N_6737);
xor U7325 (N_7325,N_6284,N_6408);
or U7326 (N_7326,N_6398,N_6095);
nand U7327 (N_7327,N_6674,N_6028);
nand U7328 (N_7328,N_6438,N_6636);
nand U7329 (N_7329,N_6475,N_6486);
nand U7330 (N_7330,N_6326,N_6357);
xor U7331 (N_7331,N_6660,N_6085);
or U7332 (N_7332,N_6338,N_6476);
xor U7333 (N_7333,N_6206,N_6485);
and U7334 (N_7334,N_6743,N_6238);
xor U7335 (N_7335,N_6090,N_6527);
and U7336 (N_7336,N_6271,N_6718);
and U7337 (N_7337,N_6259,N_6494);
or U7338 (N_7338,N_6110,N_6477);
nand U7339 (N_7339,N_6529,N_6308);
and U7340 (N_7340,N_6688,N_6419);
xor U7341 (N_7341,N_6511,N_6433);
xor U7342 (N_7342,N_6668,N_6291);
nor U7343 (N_7343,N_6073,N_6468);
nand U7344 (N_7344,N_6270,N_6651);
nand U7345 (N_7345,N_6295,N_6229);
and U7346 (N_7346,N_6144,N_6395);
xor U7347 (N_7347,N_6312,N_6047);
nand U7348 (N_7348,N_6041,N_6109);
or U7349 (N_7349,N_6315,N_6417);
xnor U7350 (N_7350,N_6604,N_6707);
xor U7351 (N_7351,N_6483,N_6632);
nor U7352 (N_7352,N_6074,N_6300);
nand U7353 (N_7353,N_6197,N_6609);
xnor U7354 (N_7354,N_6250,N_6733);
nand U7355 (N_7355,N_6150,N_6505);
and U7356 (N_7356,N_6089,N_6035);
xor U7357 (N_7357,N_6471,N_6090);
and U7358 (N_7358,N_6574,N_6181);
nor U7359 (N_7359,N_6221,N_6081);
or U7360 (N_7360,N_6475,N_6401);
or U7361 (N_7361,N_6060,N_6006);
nand U7362 (N_7362,N_6448,N_6343);
nand U7363 (N_7363,N_6614,N_6713);
nand U7364 (N_7364,N_6221,N_6061);
xnor U7365 (N_7365,N_6073,N_6055);
nand U7366 (N_7366,N_6461,N_6492);
nand U7367 (N_7367,N_6457,N_6015);
xnor U7368 (N_7368,N_6680,N_6032);
nand U7369 (N_7369,N_6338,N_6607);
and U7370 (N_7370,N_6404,N_6193);
xor U7371 (N_7371,N_6607,N_6701);
and U7372 (N_7372,N_6564,N_6650);
nand U7373 (N_7373,N_6340,N_6501);
nand U7374 (N_7374,N_6657,N_6291);
xnor U7375 (N_7375,N_6511,N_6305);
nor U7376 (N_7376,N_6307,N_6024);
xor U7377 (N_7377,N_6493,N_6033);
nand U7378 (N_7378,N_6625,N_6180);
nand U7379 (N_7379,N_6288,N_6330);
or U7380 (N_7380,N_6240,N_6634);
xor U7381 (N_7381,N_6157,N_6345);
nor U7382 (N_7382,N_6222,N_6322);
nand U7383 (N_7383,N_6608,N_6466);
nand U7384 (N_7384,N_6384,N_6724);
or U7385 (N_7385,N_6673,N_6205);
and U7386 (N_7386,N_6298,N_6538);
or U7387 (N_7387,N_6031,N_6565);
xor U7388 (N_7388,N_6244,N_6390);
and U7389 (N_7389,N_6501,N_6099);
and U7390 (N_7390,N_6000,N_6124);
or U7391 (N_7391,N_6090,N_6221);
nand U7392 (N_7392,N_6289,N_6399);
nor U7393 (N_7393,N_6739,N_6420);
nand U7394 (N_7394,N_6387,N_6072);
or U7395 (N_7395,N_6110,N_6217);
and U7396 (N_7396,N_6121,N_6696);
and U7397 (N_7397,N_6093,N_6609);
or U7398 (N_7398,N_6652,N_6579);
xor U7399 (N_7399,N_6265,N_6084);
or U7400 (N_7400,N_6402,N_6706);
or U7401 (N_7401,N_6214,N_6296);
and U7402 (N_7402,N_6120,N_6569);
xnor U7403 (N_7403,N_6669,N_6688);
nor U7404 (N_7404,N_6436,N_6354);
nand U7405 (N_7405,N_6038,N_6025);
nand U7406 (N_7406,N_6058,N_6209);
or U7407 (N_7407,N_6298,N_6056);
or U7408 (N_7408,N_6413,N_6708);
nand U7409 (N_7409,N_6181,N_6235);
and U7410 (N_7410,N_6210,N_6591);
nand U7411 (N_7411,N_6336,N_6499);
or U7412 (N_7412,N_6030,N_6536);
xnor U7413 (N_7413,N_6066,N_6152);
nand U7414 (N_7414,N_6303,N_6345);
xnor U7415 (N_7415,N_6075,N_6216);
nor U7416 (N_7416,N_6000,N_6046);
nor U7417 (N_7417,N_6124,N_6020);
nor U7418 (N_7418,N_6035,N_6350);
or U7419 (N_7419,N_6550,N_6186);
and U7420 (N_7420,N_6542,N_6249);
nand U7421 (N_7421,N_6521,N_6703);
and U7422 (N_7422,N_6002,N_6425);
or U7423 (N_7423,N_6347,N_6070);
and U7424 (N_7424,N_6032,N_6234);
or U7425 (N_7425,N_6427,N_6672);
xor U7426 (N_7426,N_6118,N_6497);
and U7427 (N_7427,N_6424,N_6169);
or U7428 (N_7428,N_6502,N_6643);
nor U7429 (N_7429,N_6500,N_6546);
or U7430 (N_7430,N_6577,N_6103);
xor U7431 (N_7431,N_6405,N_6310);
nor U7432 (N_7432,N_6132,N_6129);
xnor U7433 (N_7433,N_6707,N_6343);
nand U7434 (N_7434,N_6266,N_6290);
xor U7435 (N_7435,N_6402,N_6026);
nand U7436 (N_7436,N_6452,N_6102);
and U7437 (N_7437,N_6748,N_6130);
xor U7438 (N_7438,N_6007,N_6536);
or U7439 (N_7439,N_6671,N_6738);
xnor U7440 (N_7440,N_6550,N_6028);
or U7441 (N_7441,N_6517,N_6009);
or U7442 (N_7442,N_6677,N_6672);
and U7443 (N_7443,N_6461,N_6060);
or U7444 (N_7444,N_6060,N_6715);
xnor U7445 (N_7445,N_6566,N_6048);
nand U7446 (N_7446,N_6166,N_6714);
nor U7447 (N_7447,N_6066,N_6607);
or U7448 (N_7448,N_6677,N_6006);
and U7449 (N_7449,N_6378,N_6562);
nand U7450 (N_7450,N_6268,N_6069);
and U7451 (N_7451,N_6057,N_6388);
and U7452 (N_7452,N_6317,N_6108);
nor U7453 (N_7453,N_6449,N_6145);
nor U7454 (N_7454,N_6464,N_6573);
or U7455 (N_7455,N_6238,N_6090);
and U7456 (N_7456,N_6099,N_6012);
and U7457 (N_7457,N_6314,N_6553);
nand U7458 (N_7458,N_6015,N_6103);
or U7459 (N_7459,N_6735,N_6398);
and U7460 (N_7460,N_6651,N_6386);
nand U7461 (N_7461,N_6469,N_6004);
and U7462 (N_7462,N_6302,N_6590);
xor U7463 (N_7463,N_6070,N_6192);
or U7464 (N_7464,N_6313,N_6006);
nor U7465 (N_7465,N_6598,N_6628);
xnor U7466 (N_7466,N_6537,N_6384);
and U7467 (N_7467,N_6379,N_6277);
or U7468 (N_7468,N_6630,N_6302);
xnor U7469 (N_7469,N_6025,N_6435);
and U7470 (N_7470,N_6201,N_6624);
or U7471 (N_7471,N_6035,N_6637);
xnor U7472 (N_7472,N_6442,N_6456);
xor U7473 (N_7473,N_6158,N_6490);
or U7474 (N_7474,N_6390,N_6310);
nand U7475 (N_7475,N_6172,N_6417);
xor U7476 (N_7476,N_6217,N_6651);
or U7477 (N_7477,N_6360,N_6749);
and U7478 (N_7478,N_6132,N_6126);
xnor U7479 (N_7479,N_6718,N_6374);
or U7480 (N_7480,N_6614,N_6426);
nand U7481 (N_7481,N_6175,N_6598);
or U7482 (N_7482,N_6563,N_6582);
or U7483 (N_7483,N_6153,N_6728);
or U7484 (N_7484,N_6365,N_6141);
or U7485 (N_7485,N_6199,N_6044);
nor U7486 (N_7486,N_6588,N_6422);
nand U7487 (N_7487,N_6553,N_6356);
and U7488 (N_7488,N_6715,N_6088);
xor U7489 (N_7489,N_6292,N_6030);
nand U7490 (N_7490,N_6460,N_6567);
xor U7491 (N_7491,N_6433,N_6217);
nor U7492 (N_7492,N_6133,N_6230);
or U7493 (N_7493,N_6703,N_6479);
or U7494 (N_7494,N_6241,N_6140);
or U7495 (N_7495,N_6281,N_6150);
and U7496 (N_7496,N_6378,N_6299);
xor U7497 (N_7497,N_6273,N_6741);
nor U7498 (N_7498,N_6371,N_6149);
xor U7499 (N_7499,N_6285,N_6437);
nand U7500 (N_7500,N_7020,N_7341);
or U7501 (N_7501,N_6805,N_6841);
and U7502 (N_7502,N_7255,N_7436);
or U7503 (N_7503,N_6764,N_7057);
nor U7504 (N_7504,N_7327,N_6976);
xor U7505 (N_7505,N_7103,N_7395);
nand U7506 (N_7506,N_7035,N_6882);
xor U7507 (N_7507,N_7128,N_7177);
and U7508 (N_7508,N_7046,N_7301);
nand U7509 (N_7509,N_7347,N_7278);
nand U7510 (N_7510,N_7125,N_6955);
xnor U7511 (N_7511,N_6907,N_7424);
nor U7512 (N_7512,N_7201,N_6857);
xnor U7513 (N_7513,N_6799,N_7133);
nor U7514 (N_7514,N_7371,N_6830);
nand U7515 (N_7515,N_6876,N_7446);
xor U7516 (N_7516,N_7202,N_6810);
xnor U7517 (N_7517,N_6944,N_7453);
or U7518 (N_7518,N_7174,N_7153);
xnor U7519 (N_7519,N_6970,N_6793);
and U7520 (N_7520,N_7006,N_7484);
nor U7521 (N_7521,N_7376,N_7088);
nand U7522 (N_7522,N_7498,N_7001);
nor U7523 (N_7523,N_7072,N_6762);
and U7524 (N_7524,N_7486,N_7380);
and U7525 (N_7525,N_7070,N_7195);
and U7526 (N_7526,N_7365,N_7419);
and U7527 (N_7527,N_6833,N_7183);
xnor U7528 (N_7528,N_7363,N_7229);
nand U7529 (N_7529,N_6772,N_6774);
or U7530 (N_7530,N_7404,N_7277);
nand U7531 (N_7531,N_6991,N_7393);
nand U7532 (N_7532,N_7017,N_7156);
nor U7533 (N_7533,N_7176,N_6795);
xor U7534 (N_7534,N_6823,N_7253);
or U7535 (N_7535,N_7318,N_6766);
or U7536 (N_7536,N_7237,N_7242);
and U7537 (N_7537,N_7221,N_6767);
nand U7538 (N_7538,N_6999,N_6779);
nand U7539 (N_7539,N_7455,N_7045);
nand U7540 (N_7540,N_7262,N_7069);
nand U7541 (N_7541,N_7499,N_6753);
nor U7542 (N_7542,N_7286,N_7449);
nand U7543 (N_7543,N_6932,N_6824);
nor U7544 (N_7544,N_6967,N_7215);
and U7545 (N_7545,N_7417,N_7032);
xnor U7546 (N_7546,N_7063,N_7254);
and U7547 (N_7547,N_7245,N_7100);
and U7548 (N_7548,N_7175,N_7367);
or U7549 (N_7549,N_7381,N_7139);
nor U7550 (N_7550,N_6965,N_6820);
nor U7551 (N_7551,N_7060,N_7409);
xor U7552 (N_7552,N_7457,N_7108);
or U7553 (N_7553,N_6868,N_7071);
and U7554 (N_7554,N_7047,N_7299);
and U7555 (N_7555,N_7456,N_6923);
xor U7556 (N_7556,N_6939,N_7137);
nor U7557 (N_7557,N_7192,N_7148);
nand U7558 (N_7558,N_7087,N_7200);
and U7559 (N_7559,N_6780,N_6901);
nand U7560 (N_7560,N_7332,N_7203);
and U7561 (N_7561,N_6849,N_7401);
xor U7562 (N_7562,N_7353,N_7287);
or U7563 (N_7563,N_6804,N_7338);
and U7564 (N_7564,N_6903,N_7317);
and U7565 (N_7565,N_7190,N_7249);
xor U7566 (N_7566,N_7326,N_7468);
nor U7567 (N_7567,N_6773,N_6794);
xnor U7568 (N_7568,N_7225,N_6988);
nand U7569 (N_7569,N_7420,N_7052);
xor U7570 (N_7570,N_6896,N_7272);
xor U7571 (N_7571,N_6872,N_7132);
xor U7572 (N_7572,N_7408,N_7426);
nor U7573 (N_7573,N_7339,N_7012);
and U7574 (N_7574,N_7238,N_7391);
and U7575 (N_7575,N_7403,N_7316);
nand U7576 (N_7576,N_7155,N_7337);
or U7577 (N_7577,N_6775,N_6797);
and U7578 (N_7578,N_7305,N_7102);
and U7579 (N_7579,N_6983,N_7152);
or U7580 (N_7580,N_7437,N_7269);
xnor U7581 (N_7581,N_6898,N_7323);
xnor U7582 (N_7582,N_7368,N_6937);
or U7583 (N_7583,N_6827,N_7230);
xor U7584 (N_7584,N_6812,N_7218);
and U7585 (N_7585,N_7297,N_7000);
nand U7586 (N_7586,N_6931,N_6887);
nor U7587 (N_7587,N_6811,N_6768);
nor U7588 (N_7588,N_6890,N_7370);
and U7589 (N_7589,N_7204,N_7281);
nor U7590 (N_7590,N_7352,N_7092);
nor U7591 (N_7591,N_6886,N_6751);
and U7592 (N_7592,N_6788,N_7428);
nand U7593 (N_7593,N_7488,N_7231);
nor U7594 (N_7594,N_6807,N_7303);
nor U7595 (N_7595,N_7276,N_6935);
nand U7596 (N_7596,N_7232,N_7005);
or U7597 (N_7597,N_7285,N_6835);
nand U7598 (N_7598,N_6761,N_7433);
nor U7599 (N_7599,N_7275,N_7226);
or U7600 (N_7600,N_7270,N_7324);
or U7601 (N_7601,N_7168,N_7350);
and U7602 (N_7602,N_7321,N_6787);
nor U7603 (N_7603,N_7147,N_7165);
nand U7604 (N_7604,N_6997,N_7430);
and U7605 (N_7605,N_7360,N_6836);
and U7606 (N_7606,N_7054,N_7442);
nand U7607 (N_7607,N_6925,N_6930);
or U7608 (N_7608,N_6862,N_6987);
nor U7609 (N_7609,N_7382,N_7173);
xor U7610 (N_7610,N_6879,N_7423);
nor U7611 (N_7611,N_7356,N_7194);
xnor U7612 (N_7612,N_7104,N_6850);
and U7613 (N_7613,N_7333,N_7044);
or U7614 (N_7614,N_6831,N_6863);
or U7615 (N_7615,N_6952,N_6928);
xnor U7616 (N_7616,N_7279,N_7280);
or U7617 (N_7617,N_7043,N_6986);
nand U7618 (N_7618,N_7062,N_7427);
or U7619 (N_7619,N_7157,N_7266);
and U7620 (N_7620,N_7250,N_7127);
and U7621 (N_7621,N_6871,N_7134);
xor U7622 (N_7622,N_7374,N_6782);
and U7623 (N_7623,N_7029,N_7145);
xor U7624 (N_7624,N_6894,N_7079);
nor U7625 (N_7625,N_7251,N_7027);
nor U7626 (N_7626,N_7023,N_7358);
xor U7627 (N_7627,N_6861,N_6984);
and U7628 (N_7628,N_6869,N_7300);
or U7629 (N_7629,N_6834,N_7077);
nor U7630 (N_7630,N_7031,N_7289);
xor U7631 (N_7631,N_7216,N_7246);
nor U7632 (N_7632,N_7328,N_7123);
xnor U7633 (N_7633,N_7463,N_7405);
and U7634 (N_7634,N_6947,N_6927);
nor U7635 (N_7635,N_7078,N_7117);
or U7636 (N_7636,N_6865,N_6832);
xor U7637 (N_7637,N_7344,N_6892);
nand U7638 (N_7638,N_6809,N_7014);
nand U7639 (N_7639,N_7429,N_6956);
and U7640 (N_7640,N_7191,N_7379);
and U7641 (N_7641,N_7091,N_7481);
nor U7642 (N_7642,N_7243,N_7392);
and U7643 (N_7643,N_6874,N_7397);
nand U7644 (N_7644,N_7039,N_6918);
nand U7645 (N_7645,N_6884,N_6900);
or U7646 (N_7646,N_7030,N_6958);
xnor U7647 (N_7647,N_7349,N_7184);
or U7648 (N_7648,N_6974,N_7061);
nor U7649 (N_7649,N_7410,N_7407);
or U7650 (N_7650,N_6888,N_6750);
nand U7651 (N_7651,N_7458,N_7034);
xor U7652 (N_7652,N_7315,N_7329);
nor U7653 (N_7653,N_7056,N_7219);
xnor U7654 (N_7654,N_7386,N_7288);
nand U7655 (N_7655,N_7224,N_7240);
and U7656 (N_7656,N_6929,N_6968);
or U7657 (N_7657,N_6765,N_7434);
xor U7658 (N_7658,N_7389,N_6966);
and U7659 (N_7659,N_6756,N_6808);
nand U7660 (N_7660,N_6770,N_6963);
or U7661 (N_7661,N_6908,N_7460);
xnor U7662 (N_7662,N_6990,N_7252);
nor U7663 (N_7663,N_7473,N_7290);
xor U7664 (N_7664,N_6972,N_7497);
nor U7665 (N_7665,N_7482,N_6798);
nor U7666 (N_7666,N_7098,N_7141);
nand U7667 (N_7667,N_6838,N_7343);
nand U7668 (N_7668,N_7223,N_6942);
and U7669 (N_7669,N_6977,N_7496);
nor U7670 (N_7670,N_6866,N_7009);
xnor U7671 (N_7671,N_7050,N_7115);
or U7672 (N_7672,N_7081,N_7217);
nand U7673 (N_7673,N_7233,N_7443);
or U7674 (N_7674,N_6845,N_7283);
nand U7675 (N_7675,N_6818,N_7049);
nand U7676 (N_7676,N_7227,N_6801);
nand U7677 (N_7677,N_7314,N_7320);
and U7678 (N_7678,N_7161,N_7021);
and U7679 (N_7679,N_6941,N_7065);
or U7680 (N_7680,N_7244,N_7479);
and U7681 (N_7681,N_7179,N_6754);
and U7682 (N_7682,N_6994,N_6904);
and U7683 (N_7683,N_7066,N_7239);
nand U7684 (N_7684,N_7162,N_6895);
nand U7685 (N_7685,N_7263,N_7163);
or U7686 (N_7686,N_7361,N_7124);
or U7687 (N_7687,N_7121,N_7469);
nand U7688 (N_7688,N_6778,N_6909);
or U7689 (N_7689,N_7261,N_7015);
or U7690 (N_7690,N_7222,N_6992);
xor U7691 (N_7691,N_7167,N_6917);
xnor U7692 (N_7692,N_6981,N_6948);
nor U7693 (N_7693,N_7228,N_6945);
xnor U7694 (N_7694,N_6951,N_6755);
and U7695 (N_7695,N_6859,N_7258);
xor U7696 (N_7696,N_6973,N_6971);
xnor U7697 (N_7697,N_6989,N_6791);
nor U7698 (N_7698,N_7051,N_7082);
nand U7699 (N_7699,N_7472,N_6881);
or U7700 (N_7700,N_7490,N_7138);
and U7701 (N_7701,N_7199,N_7189);
and U7702 (N_7702,N_7489,N_6936);
and U7703 (N_7703,N_7094,N_7485);
xor U7704 (N_7704,N_7182,N_7372);
nand U7705 (N_7705,N_6883,N_7295);
or U7706 (N_7706,N_7377,N_7164);
nand U7707 (N_7707,N_7235,N_6960);
and U7708 (N_7708,N_7171,N_7241);
or U7709 (N_7709,N_7055,N_7172);
and U7710 (N_7710,N_7260,N_6950);
nand U7711 (N_7711,N_6852,N_7053);
and U7712 (N_7712,N_6758,N_7435);
nor U7713 (N_7713,N_6815,N_7105);
and U7714 (N_7714,N_6792,N_7418);
xor U7715 (N_7715,N_7438,N_6854);
nand U7716 (N_7716,N_7119,N_7114);
xnor U7717 (N_7717,N_7293,N_6996);
nor U7718 (N_7718,N_7291,N_7159);
nand U7719 (N_7719,N_7096,N_7016);
xor U7720 (N_7720,N_7462,N_7146);
and U7721 (N_7721,N_7450,N_6980);
nor U7722 (N_7722,N_6916,N_7126);
and U7723 (N_7723,N_6906,N_7307);
nand U7724 (N_7724,N_6878,N_7058);
and U7725 (N_7725,N_7467,N_6784);
nand U7726 (N_7726,N_7186,N_6961);
xor U7727 (N_7727,N_7394,N_7109);
xnor U7728 (N_7728,N_7265,N_7267);
and U7729 (N_7729,N_6938,N_7416);
or U7730 (N_7730,N_6949,N_6993);
or U7731 (N_7731,N_7151,N_7169);
and U7732 (N_7732,N_7106,N_6837);
nand U7733 (N_7733,N_7465,N_7075);
or U7734 (N_7734,N_7273,N_7113);
and U7735 (N_7735,N_7441,N_6905);
xnor U7736 (N_7736,N_7256,N_6870);
nand U7737 (N_7737,N_6829,N_7130);
nor U7738 (N_7738,N_6889,N_6803);
nand U7739 (N_7739,N_7129,N_6855);
nor U7740 (N_7740,N_7166,N_7086);
or U7741 (N_7741,N_7451,N_7210);
or U7742 (N_7742,N_7390,N_7154);
or U7743 (N_7743,N_7180,N_7211);
xor U7744 (N_7744,N_7067,N_6821);
nor U7745 (N_7745,N_6819,N_7038);
or U7746 (N_7746,N_7064,N_7214);
xnor U7747 (N_7747,N_7122,N_7111);
and U7748 (N_7748,N_7149,N_6969);
or U7749 (N_7749,N_7493,N_7415);
xor U7750 (N_7750,N_6851,N_7310);
xor U7751 (N_7751,N_7011,N_6919);
xor U7752 (N_7752,N_7306,N_7474);
nand U7753 (N_7753,N_6846,N_7362);
xnor U7754 (N_7754,N_7387,N_6985);
xnor U7755 (N_7755,N_6776,N_7384);
nand U7756 (N_7756,N_7095,N_7355);
nand U7757 (N_7757,N_6840,N_7354);
or U7758 (N_7758,N_7312,N_7158);
and U7759 (N_7759,N_7483,N_6856);
or U7760 (N_7760,N_7010,N_7036);
and U7761 (N_7761,N_7247,N_6806);
xor U7762 (N_7762,N_7447,N_6954);
or U7763 (N_7763,N_7491,N_6897);
xor U7764 (N_7764,N_7383,N_7492);
nor U7765 (N_7765,N_7013,N_6802);
nand U7766 (N_7766,N_7494,N_7378);
xor U7767 (N_7767,N_6825,N_7076);
xor U7768 (N_7768,N_7131,N_6848);
and U7769 (N_7769,N_7298,N_7236);
and U7770 (N_7770,N_7439,N_7110);
xor U7771 (N_7771,N_7373,N_7284);
xnor U7772 (N_7772,N_7425,N_6789);
nand U7773 (N_7773,N_7073,N_7085);
or U7774 (N_7774,N_7059,N_7143);
or U7775 (N_7775,N_7399,N_7282);
or U7776 (N_7776,N_7193,N_7003);
nand U7777 (N_7777,N_7385,N_7406);
xnor U7778 (N_7778,N_7140,N_7336);
nand U7779 (N_7779,N_6864,N_6813);
and U7780 (N_7780,N_7319,N_7388);
and U7781 (N_7781,N_6914,N_6867);
nand U7782 (N_7782,N_6781,N_7431);
xnor U7783 (N_7783,N_6843,N_6785);
nand U7784 (N_7784,N_7413,N_7480);
nand U7785 (N_7785,N_7325,N_7019);
and U7786 (N_7786,N_7364,N_7198);
and U7787 (N_7787,N_7444,N_6964);
or U7788 (N_7788,N_6880,N_7142);
or U7789 (N_7789,N_7432,N_6763);
and U7790 (N_7790,N_7208,N_6899);
or U7791 (N_7791,N_6940,N_7206);
and U7792 (N_7792,N_7268,N_7487);
and U7793 (N_7793,N_7004,N_7026);
or U7794 (N_7794,N_6978,N_6943);
nor U7795 (N_7795,N_6998,N_7335);
or U7796 (N_7796,N_6877,N_6800);
or U7797 (N_7797,N_6995,N_6853);
and U7798 (N_7798,N_7002,N_7340);
and U7799 (N_7799,N_7187,N_7188);
and U7800 (N_7800,N_7178,N_7292);
xnor U7801 (N_7801,N_6911,N_6842);
or U7802 (N_7802,N_6759,N_7099);
nor U7803 (N_7803,N_6822,N_7422);
nor U7804 (N_7804,N_7421,N_7264);
and U7805 (N_7805,N_6962,N_7302);
or U7806 (N_7806,N_6828,N_7037);
and U7807 (N_7807,N_7359,N_6912);
nand U7808 (N_7808,N_6959,N_7478);
and U7809 (N_7809,N_6979,N_7080);
xnor U7810 (N_7810,N_7495,N_7396);
or U7811 (N_7811,N_6816,N_7101);
xnor U7812 (N_7812,N_7093,N_7466);
and U7813 (N_7813,N_7084,N_7322);
nor U7814 (N_7814,N_7118,N_7185);
or U7815 (N_7815,N_7120,N_7028);
nand U7816 (N_7816,N_7346,N_7345);
nor U7817 (N_7817,N_7234,N_7334);
or U7818 (N_7818,N_7411,N_7477);
nor U7819 (N_7819,N_7448,N_7475);
and U7820 (N_7820,N_7083,N_6910);
nand U7821 (N_7821,N_7197,N_7470);
nor U7822 (N_7822,N_7402,N_7311);
xor U7823 (N_7823,N_7412,N_7357);
nand U7824 (N_7824,N_7112,N_7464);
and U7825 (N_7825,N_6926,N_7048);
xnor U7826 (N_7826,N_7342,N_6924);
xnor U7827 (N_7827,N_6826,N_6790);
nor U7828 (N_7828,N_6893,N_7068);
or U7829 (N_7829,N_7207,N_6913);
and U7830 (N_7830,N_7220,N_7271);
nand U7831 (N_7831,N_7040,N_7459);
nor U7832 (N_7832,N_7308,N_7274);
xor U7833 (N_7833,N_7144,N_7471);
nand U7834 (N_7834,N_7351,N_6953);
nand U7835 (N_7835,N_7135,N_6915);
nand U7836 (N_7836,N_6921,N_7476);
nand U7837 (N_7837,N_7018,N_7181);
and U7838 (N_7838,N_7209,N_7022);
nand U7839 (N_7839,N_6760,N_6839);
and U7840 (N_7840,N_7116,N_6858);
xor U7841 (N_7841,N_6769,N_7024);
or U7842 (N_7842,N_7041,N_7454);
or U7843 (N_7843,N_6920,N_6796);
nand U7844 (N_7844,N_7445,N_6891);
nor U7845 (N_7845,N_7150,N_7296);
xnor U7846 (N_7846,N_6982,N_6817);
or U7847 (N_7847,N_6777,N_7348);
nand U7848 (N_7848,N_7400,N_6860);
and U7849 (N_7849,N_6946,N_7414);
and U7850 (N_7850,N_7330,N_6902);
nor U7851 (N_7851,N_7160,N_7090);
nor U7852 (N_7852,N_7196,N_6873);
xnor U7853 (N_7853,N_7309,N_7440);
nand U7854 (N_7854,N_6934,N_7033);
or U7855 (N_7855,N_7366,N_7257);
and U7856 (N_7856,N_7259,N_7248);
nand U7857 (N_7857,N_6771,N_7398);
and U7858 (N_7858,N_6885,N_7025);
nor U7859 (N_7859,N_6847,N_7294);
or U7860 (N_7860,N_7074,N_6875);
nand U7861 (N_7861,N_7331,N_6757);
and U7862 (N_7862,N_7369,N_7461);
or U7863 (N_7863,N_6922,N_7089);
nor U7864 (N_7864,N_7212,N_7107);
xnor U7865 (N_7865,N_7136,N_7205);
nand U7866 (N_7866,N_7042,N_6844);
nor U7867 (N_7867,N_7375,N_6783);
nor U7868 (N_7868,N_6975,N_7213);
nor U7869 (N_7869,N_7452,N_7313);
and U7870 (N_7870,N_7304,N_6786);
and U7871 (N_7871,N_7170,N_6933);
and U7872 (N_7872,N_6814,N_7008);
or U7873 (N_7873,N_7097,N_6957);
xor U7874 (N_7874,N_6752,N_7007);
and U7875 (N_7875,N_7071,N_6931);
nor U7876 (N_7876,N_7308,N_6874);
and U7877 (N_7877,N_7236,N_7246);
or U7878 (N_7878,N_7130,N_7423);
xnor U7879 (N_7879,N_6817,N_6868);
nor U7880 (N_7880,N_6922,N_7170);
and U7881 (N_7881,N_7263,N_7005);
xnor U7882 (N_7882,N_7092,N_6967);
nand U7883 (N_7883,N_7424,N_7385);
and U7884 (N_7884,N_6987,N_7360);
nor U7885 (N_7885,N_6824,N_6865);
xor U7886 (N_7886,N_6957,N_7095);
nor U7887 (N_7887,N_6907,N_7187);
xor U7888 (N_7888,N_6763,N_6835);
xor U7889 (N_7889,N_6894,N_7444);
or U7890 (N_7890,N_6831,N_6767);
nand U7891 (N_7891,N_7134,N_7007);
nand U7892 (N_7892,N_7294,N_6912);
nand U7893 (N_7893,N_6832,N_6913);
nand U7894 (N_7894,N_6900,N_7213);
nor U7895 (N_7895,N_7302,N_6888);
or U7896 (N_7896,N_7182,N_6790);
nor U7897 (N_7897,N_6951,N_7042);
or U7898 (N_7898,N_7243,N_6939);
xor U7899 (N_7899,N_6957,N_7354);
nor U7900 (N_7900,N_7121,N_7448);
or U7901 (N_7901,N_7199,N_7207);
or U7902 (N_7902,N_7108,N_7313);
nand U7903 (N_7903,N_7020,N_6979);
and U7904 (N_7904,N_6876,N_7406);
and U7905 (N_7905,N_7467,N_7441);
nand U7906 (N_7906,N_7458,N_6926);
and U7907 (N_7907,N_7203,N_7426);
and U7908 (N_7908,N_6937,N_7198);
xnor U7909 (N_7909,N_6999,N_7040);
nor U7910 (N_7910,N_6951,N_7301);
or U7911 (N_7911,N_6802,N_7086);
and U7912 (N_7912,N_7336,N_7282);
nand U7913 (N_7913,N_7306,N_7312);
and U7914 (N_7914,N_6844,N_6975);
xor U7915 (N_7915,N_6965,N_7088);
or U7916 (N_7916,N_6780,N_7216);
nand U7917 (N_7917,N_6831,N_6888);
nand U7918 (N_7918,N_6982,N_7236);
nand U7919 (N_7919,N_7419,N_7394);
nor U7920 (N_7920,N_6868,N_6988);
and U7921 (N_7921,N_6964,N_6806);
nand U7922 (N_7922,N_6995,N_7240);
nor U7923 (N_7923,N_7192,N_7325);
nor U7924 (N_7924,N_7046,N_6850);
nand U7925 (N_7925,N_7103,N_7385);
xnor U7926 (N_7926,N_7432,N_7311);
xnor U7927 (N_7927,N_7204,N_7365);
or U7928 (N_7928,N_7062,N_7244);
and U7929 (N_7929,N_7103,N_6807);
or U7930 (N_7930,N_7140,N_7370);
nor U7931 (N_7931,N_6773,N_6893);
xor U7932 (N_7932,N_6753,N_7283);
nand U7933 (N_7933,N_6908,N_7377);
or U7934 (N_7934,N_7480,N_6931);
nor U7935 (N_7935,N_6901,N_7195);
xor U7936 (N_7936,N_7166,N_7152);
xor U7937 (N_7937,N_7420,N_7448);
xnor U7938 (N_7938,N_6798,N_6763);
and U7939 (N_7939,N_7135,N_7020);
and U7940 (N_7940,N_7228,N_7362);
or U7941 (N_7941,N_6935,N_6864);
or U7942 (N_7942,N_7101,N_7452);
and U7943 (N_7943,N_7026,N_7274);
and U7944 (N_7944,N_7484,N_6854);
and U7945 (N_7945,N_7114,N_6893);
xnor U7946 (N_7946,N_6988,N_7181);
nand U7947 (N_7947,N_7316,N_6832);
nor U7948 (N_7948,N_7297,N_7325);
nand U7949 (N_7949,N_7392,N_7263);
nand U7950 (N_7950,N_6984,N_6757);
and U7951 (N_7951,N_7491,N_7440);
nor U7952 (N_7952,N_7039,N_6934);
nand U7953 (N_7953,N_7377,N_7114);
xnor U7954 (N_7954,N_6887,N_6874);
xor U7955 (N_7955,N_7219,N_6793);
nand U7956 (N_7956,N_6839,N_7022);
nand U7957 (N_7957,N_7084,N_6956);
or U7958 (N_7958,N_7439,N_7234);
and U7959 (N_7959,N_7432,N_6839);
or U7960 (N_7960,N_7321,N_6891);
and U7961 (N_7961,N_7446,N_7261);
nand U7962 (N_7962,N_7459,N_7272);
or U7963 (N_7963,N_7079,N_6845);
xor U7964 (N_7964,N_6765,N_7325);
nor U7965 (N_7965,N_7490,N_6801);
or U7966 (N_7966,N_7009,N_6937);
nor U7967 (N_7967,N_6928,N_7121);
and U7968 (N_7968,N_6827,N_7316);
nand U7969 (N_7969,N_6771,N_7432);
nor U7970 (N_7970,N_6774,N_6918);
or U7971 (N_7971,N_7445,N_6818);
or U7972 (N_7972,N_7123,N_6815);
or U7973 (N_7973,N_6923,N_7445);
xnor U7974 (N_7974,N_7199,N_7310);
xnor U7975 (N_7975,N_7221,N_6811);
nand U7976 (N_7976,N_6909,N_7092);
and U7977 (N_7977,N_7057,N_6825);
xnor U7978 (N_7978,N_7204,N_7310);
or U7979 (N_7979,N_7448,N_7308);
and U7980 (N_7980,N_7184,N_7180);
or U7981 (N_7981,N_7062,N_7094);
xnor U7982 (N_7982,N_6953,N_7155);
xnor U7983 (N_7983,N_7057,N_7181);
nand U7984 (N_7984,N_7023,N_6894);
and U7985 (N_7985,N_6815,N_7278);
xor U7986 (N_7986,N_6991,N_6848);
nor U7987 (N_7987,N_7345,N_7381);
nor U7988 (N_7988,N_7370,N_7264);
xnor U7989 (N_7989,N_7413,N_6905);
xor U7990 (N_7990,N_7024,N_7388);
nor U7991 (N_7991,N_7406,N_7140);
xor U7992 (N_7992,N_7209,N_7274);
xnor U7993 (N_7993,N_7290,N_7301);
and U7994 (N_7994,N_7047,N_7391);
or U7995 (N_7995,N_6866,N_7260);
and U7996 (N_7996,N_7436,N_6877);
nor U7997 (N_7997,N_7039,N_6802);
nor U7998 (N_7998,N_7386,N_6832);
xor U7999 (N_7999,N_7477,N_6767);
nor U8000 (N_8000,N_6782,N_6941);
nor U8001 (N_8001,N_6789,N_7107);
or U8002 (N_8002,N_7065,N_6824);
or U8003 (N_8003,N_7297,N_6869);
nand U8004 (N_8004,N_6941,N_7371);
and U8005 (N_8005,N_7148,N_6893);
xor U8006 (N_8006,N_6871,N_6760);
xor U8007 (N_8007,N_7429,N_7124);
and U8008 (N_8008,N_7367,N_6950);
nand U8009 (N_8009,N_7203,N_6907);
xor U8010 (N_8010,N_7336,N_7408);
and U8011 (N_8011,N_6997,N_7381);
nor U8012 (N_8012,N_6831,N_7165);
nor U8013 (N_8013,N_7344,N_7046);
or U8014 (N_8014,N_7279,N_6837);
and U8015 (N_8015,N_7423,N_6809);
and U8016 (N_8016,N_7113,N_7306);
and U8017 (N_8017,N_7430,N_6880);
nor U8018 (N_8018,N_6807,N_7067);
nor U8019 (N_8019,N_7243,N_6813);
xor U8020 (N_8020,N_6790,N_7265);
nor U8021 (N_8021,N_7216,N_7325);
nand U8022 (N_8022,N_6809,N_7294);
nor U8023 (N_8023,N_6804,N_7200);
xor U8024 (N_8024,N_7033,N_7009);
nand U8025 (N_8025,N_7075,N_6965);
xnor U8026 (N_8026,N_6808,N_7442);
nor U8027 (N_8027,N_7479,N_7178);
nor U8028 (N_8028,N_7276,N_6915);
nor U8029 (N_8029,N_7377,N_6820);
xor U8030 (N_8030,N_6917,N_6944);
xnor U8031 (N_8031,N_6823,N_7016);
nor U8032 (N_8032,N_7014,N_7205);
xor U8033 (N_8033,N_7391,N_7057);
or U8034 (N_8034,N_6961,N_6792);
or U8035 (N_8035,N_6815,N_6964);
nor U8036 (N_8036,N_7455,N_6771);
xor U8037 (N_8037,N_6860,N_7430);
xnor U8038 (N_8038,N_6797,N_6853);
nand U8039 (N_8039,N_7425,N_7117);
or U8040 (N_8040,N_6955,N_7372);
and U8041 (N_8041,N_7466,N_7031);
or U8042 (N_8042,N_7136,N_7001);
xnor U8043 (N_8043,N_7259,N_6791);
nor U8044 (N_8044,N_6884,N_7225);
and U8045 (N_8045,N_7409,N_6847);
nand U8046 (N_8046,N_6755,N_7241);
or U8047 (N_8047,N_7409,N_6840);
xor U8048 (N_8048,N_6785,N_6819);
nand U8049 (N_8049,N_7042,N_7179);
nand U8050 (N_8050,N_6852,N_6918);
nor U8051 (N_8051,N_7015,N_7166);
nand U8052 (N_8052,N_7216,N_6933);
or U8053 (N_8053,N_7456,N_7261);
and U8054 (N_8054,N_7275,N_7245);
nor U8055 (N_8055,N_6769,N_7112);
nand U8056 (N_8056,N_6861,N_7386);
or U8057 (N_8057,N_7423,N_7060);
xor U8058 (N_8058,N_7330,N_7159);
or U8059 (N_8059,N_7088,N_7336);
nor U8060 (N_8060,N_7245,N_7376);
or U8061 (N_8061,N_7129,N_7323);
xnor U8062 (N_8062,N_7175,N_6904);
nor U8063 (N_8063,N_7176,N_7285);
nand U8064 (N_8064,N_7414,N_7310);
xor U8065 (N_8065,N_6943,N_7025);
nor U8066 (N_8066,N_7403,N_7175);
nand U8067 (N_8067,N_7161,N_7261);
xor U8068 (N_8068,N_6907,N_7275);
and U8069 (N_8069,N_6773,N_7499);
xnor U8070 (N_8070,N_6952,N_7467);
nor U8071 (N_8071,N_7023,N_7016);
nand U8072 (N_8072,N_7122,N_7461);
xnor U8073 (N_8073,N_6813,N_7337);
nand U8074 (N_8074,N_6862,N_7326);
or U8075 (N_8075,N_7124,N_7043);
nand U8076 (N_8076,N_7319,N_7484);
xor U8077 (N_8077,N_7387,N_6795);
and U8078 (N_8078,N_6917,N_7340);
nor U8079 (N_8079,N_7161,N_6754);
nor U8080 (N_8080,N_7475,N_7442);
or U8081 (N_8081,N_7480,N_7027);
or U8082 (N_8082,N_7281,N_7438);
xor U8083 (N_8083,N_7311,N_7380);
and U8084 (N_8084,N_7150,N_6782);
nand U8085 (N_8085,N_6988,N_7324);
xor U8086 (N_8086,N_7075,N_7254);
xnor U8087 (N_8087,N_7011,N_6890);
nor U8088 (N_8088,N_6915,N_6976);
or U8089 (N_8089,N_7079,N_7343);
and U8090 (N_8090,N_7224,N_7088);
xor U8091 (N_8091,N_7048,N_7495);
nand U8092 (N_8092,N_7362,N_7442);
nand U8093 (N_8093,N_7140,N_7287);
xor U8094 (N_8094,N_7202,N_6931);
xnor U8095 (N_8095,N_6805,N_7474);
and U8096 (N_8096,N_7487,N_7334);
xor U8097 (N_8097,N_6789,N_7208);
nor U8098 (N_8098,N_7246,N_7006);
and U8099 (N_8099,N_7082,N_7288);
xnor U8100 (N_8100,N_7342,N_7367);
nand U8101 (N_8101,N_7481,N_6771);
and U8102 (N_8102,N_7062,N_7363);
or U8103 (N_8103,N_6933,N_7355);
nor U8104 (N_8104,N_7239,N_6878);
nor U8105 (N_8105,N_6911,N_6751);
and U8106 (N_8106,N_7089,N_7018);
nor U8107 (N_8107,N_7231,N_6757);
xor U8108 (N_8108,N_7146,N_7488);
and U8109 (N_8109,N_6842,N_7145);
nand U8110 (N_8110,N_7454,N_7112);
and U8111 (N_8111,N_7132,N_7407);
nand U8112 (N_8112,N_7165,N_7361);
xnor U8113 (N_8113,N_6885,N_7003);
xor U8114 (N_8114,N_6963,N_6814);
and U8115 (N_8115,N_7459,N_7032);
or U8116 (N_8116,N_6773,N_7194);
nand U8117 (N_8117,N_7003,N_6829);
and U8118 (N_8118,N_7347,N_6757);
and U8119 (N_8119,N_7202,N_7007);
or U8120 (N_8120,N_7002,N_7373);
nor U8121 (N_8121,N_7329,N_6969);
or U8122 (N_8122,N_7102,N_6817);
xnor U8123 (N_8123,N_7303,N_7282);
or U8124 (N_8124,N_7332,N_7044);
nor U8125 (N_8125,N_6839,N_6962);
nand U8126 (N_8126,N_7079,N_7027);
xor U8127 (N_8127,N_7387,N_6876);
nor U8128 (N_8128,N_6795,N_6941);
and U8129 (N_8129,N_6777,N_7228);
nand U8130 (N_8130,N_7215,N_7185);
nand U8131 (N_8131,N_6901,N_6872);
nand U8132 (N_8132,N_7376,N_7080);
and U8133 (N_8133,N_7045,N_6768);
and U8134 (N_8134,N_7344,N_7443);
or U8135 (N_8135,N_7331,N_7271);
or U8136 (N_8136,N_7415,N_7212);
and U8137 (N_8137,N_7058,N_7137);
or U8138 (N_8138,N_7020,N_6875);
and U8139 (N_8139,N_6935,N_7491);
nand U8140 (N_8140,N_6802,N_7405);
and U8141 (N_8141,N_6803,N_7011);
nor U8142 (N_8142,N_6948,N_6893);
nand U8143 (N_8143,N_7481,N_7179);
nor U8144 (N_8144,N_7167,N_6983);
nand U8145 (N_8145,N_6826,N_7375);
and U8146 (N_8146,N_6914,N_7363);
nor U8147 (N_8147,N_7304,N_7381);
and U8148 (N_8148,N_7402,N_7473);
or U8149 (N_8149,N_7323,N_7242);
xnor U8150 (N_8150,N_7158,N_7238);
xnor U8151 (N_8151,N_7266,N_7148);
nand U8152 (N_8152,N_7345,N_7207);
nor U8153 (N_8153,N_6905,N_7196);
and U8154 (N_8154,N_7066,N_7289);
and U8155 (N_8155,N_6816,N_7255);
nor U8156 (N_8156,N_7291,N_6817);
xnor U8157 (N_8157,N_7416,N_6817);
nor U8158 (N_8158,N_7193,N_7342);
or U8159 (N_8159,N_6757,N_7100);
xor U8160 (N_8160,N_7212,N_7455);
nand U8161 (N_8161,N_7274,N_6792);
nor U8162 (N_8162,N_7130,N_7450);
xnor U8163 (N_8163,N_7216,N_7039);
nand U8164 (N_8164,N_7034,N_6919);
and U8165 (N_8165,N_6856,N_7360);
or U8166 (N_8166,N_7122,N_7475);
nand U8167 (N_8167,N_6775,N_7354);
nor U8168 (N_8168,N_6788,N_7329);
xnor U8169 (N_8169,N_7380,N_7009);
or U8170 (N_8170,N_7121,N_6782);
and U8171 (N_8171,N_7197,N_7394);
and U8172 (N_8172,N_7212,N_7430);
or U8173 (N_8173,N_6793,N_7139);
xor U8174 (N_8174,N_7430,N_6902);
xor U8175 (N_8175,N_7288,N_7329);
nand U8176 (N_8176,N_7316,N_7063);
nand U8177 (N_8177,N_6802,N_7421);
or U8178 (N_8178,N_7251,N_6982);
xnor U8179 (N_8179,N_7098,N_7382);
nor U8180 (N_8180,N_7077,N_6806);
and U8181 (N_8181,N_7232,N_6997);
or U8182 (N_8182,N_6904,N_7293);
nor U8183 (N_8183,N_7295,N_7074);
xnor U8184 (N_8184,N_7480,N_7067);
and U8185 (N_8185,N_7482,N_7379);
nor U8186 (N_8186,N_6884,N_6930);
xnor U8187 (N_8187,N_6948,N_7049);
nand U8188 (N_8188,N_6914,N_7427);
nand U8189 (N_8189,N_7139,N_7471);
or U8190 (N_8190,N_7174,N_6863);
or U8191 (N_8191,N_7386,N_6941);
and U8192 (N_8192,N_6990,N_7477);
or U8193 (N_8193,N_7069,N_7358);
nand U8194 (N_8194,N_6908,N_6960);
and U8195 (N_8195,N_7444,N_6995);
and U8196 (N_8196,N_7280,N_7257);
or U8197 (N_8197,N_6898,N_7473);
nor U8198 (N_8198,N_6846,N_6943);
nor U8199 (N_8199,N_7017,N_7427);
or U8200 (N_8200,N_7182,N_6962);
xnor U8201 (N_8201,N_6888,N_7462);
xor U8202 (N_8202,N_7458,N_6819);
or U8203 (N_8203,N_7288,N_6950);
nor U8204 (N_8204,N_7003,N_6764);
and U8205 (N_8205,N_6828,N_6783);
nor U8206 (N_8206,N_7454,N_7408);
xor U8207 (N_8207,N_7152,N_7349);
nor U8208 (N_8208,N_7223,N_7018);
or U8209 (N_8209,N_6977,N_6799);
nor U8210 (N_8210,N_6859,N_7048);
nor U8211 (N_8211,N_7025,N_6869);
or U8212 (N_8212,N_7143,N_7094);
or U8213 (N_8213,N_7240,N_7319);
nand U8214 (N_8214,N_7132,N_6808);
and U8215 (N_8215,N_6774,N_7355);
nor U8216 (N_8216,N_7408,N_7455);
or U8217 (N_8217,N_6951,N_6897);
xnor U8218 (N_8218,N_6875,N_6939);
xnor U8219 (N_8219,N_7318,N_7076);
or U8220 (N_8220,N_7022,N_7138);
nor U8221 (N_8221,N_7309,N_7008);
xor U8222 (N_8222,N_6968,N_7403);
nand U8223 (N_8223,N_7097,N_6853);
nor U8224 (N_8224,N_6887,N_7487);
xnor U8225 (N_8225,N_7419,N_6882);
and U8226 (N_8226,N_7203,N_7255);
xnor U8227 (N_8227,N_7087,N_7358);
nand U8228 (N_8228,N_7343,N_7183);
and U8229 (N_8229,N_6953,N_7430);
nor U8230 (N_8230,N_7142,N_6832);
nor U8231 (N_8231,N_7279,N_7270);
or U8232 (N_8232,N_7280,N_7339);
or U8233 (N_8233,N_7161,N_6758);
nand U8234 (N_8234,N_7293,N_7145);
nand U8235 (N_8235,N_6821,N_6795);
xor U8236 (N_8236,N_6775,N_7446);
and U8237 (N_8237,N_7321,N_7333);
and U8238 (N_8238,N_6859,N_6903);
xnor U8239 (N_8239,N_7193,N_6803);
nand U8240 (N_8240,N_6915,N_7399);
nor U8241 (N_8241,N_7334,N_7002);
nor U8242 (N_8242,N_7216,N_7250);
or U8243 (N_8243,N_7199,N_7178);
xnor U8244 (N_8244,N_6948,N_6781);
xnor U8245 (N_8245,N_7023,N_6765);
nand U8246 (N_8246,N_6936,N_7142);
or U8247 (N_8247,N_7109,N_7117);
nor U8248 (N_8248,N_6879,N_7360);
nand U8249 (N_8249,N_6760,N_7448);
nand U8250 (N_8250,N_7571,N_7973);
xnor U8251 (N_8251,N_7603,N_7967);
and U8252 (N_8252,N_7935,N_8126);
or U8253 (N_8253,N_7787,N_8158);
or U8254 (N_8254,N_7535,N_8168);
xor U8255 (N_8255,N_7587,N_7540);
xnor U8256 (N_8256,N_7939,N_7671);
nor U8257 (N_8257,N_7515,N_7864);
nand U8258 (N_8258,N_7969,N_7602);
nor U8259 (N_8259,N_7570,N_8194);
xor U8260 (N_8260,N_7554,N_8098);
nor U8261 (N_8261,N_8161,N_8128);
nand U8262 (N_8262,N_8090,N_7948);
or U8263 (N_8263,N_7985,N_7921);
and U8264 (N_8264,N_7548,N_8046);
or U8265 (N_8265,N_7676,N_7785);
xor U8266 (N_8266,N_7890,N_7522);
xor U8267 (N_8267,N_7523,N_8189);
and U8268 (N_8268,N_7997,N_7803);
xor U8269 (N_8269,N_7632,N_7609);
nor U8270 (N_8270,N_7551,N_7688);
and U8271 (N_8271,N_7937,N_8244);
xor U8272 (N_8272,N_7624,N_7633);
nand U8273 (N_8273,N_7916,N_7812);
nor U8274 (N_8274,N_7516,N_7569);
and U8275 (N_8275,N_7971,N_7737);
and U8276 (N_8276,N_7521,N_7895);
xnor U8277 (N_8277,N_7848,N_8064);
or U8278 (N_8278,N_8080,N_7849);
nand U8279 (N_8279,N_7949,N_7683);
or U8280 (N_8280,N_7684,N_8014);
and U8281 (N_8281,N_7993,N_7505);
or U8282 (N_8282,N_7970,N_8075);
and U8283 (N_8283,N_7865,N_8056);
nor U8284 (N_8284,N_7661,N_7818);
and U8285 (N_8285,N_8035,N_7931);
nor U8286 (N_8286,N_7856,N_8248);
and U8287 (N_8287,N_7835,N_8099);
or U8288 (N_8288,N_7929,N_8155);
or U8289 (N_8289,N_7718,N_8130);
nor U8290 (N_8290,N_7837,N_8204);
nand U8291 (N_8291,N_7513,N_7646);
or U8292 (N_8292,N_8108,N_8234);
nand U8293 (N_8293,N_7964,N_8123);
nor U8294 (N_8294,N_7947,N_7771);
nor U8295 (N_8295,N_7850,N_7592);
or U8296 (N_8296,N_8113,N_7732);
or U8297 (N_8297,N_8227,N_7775);
or U8298 (N_8298,N_7751,N_8079);
nand U8299 (N_8299,N_7976,N_7707);
nand U8300 (N_8300,N_8078,N_7530);
and U8301 (N_8301,N_7582,N_8166);
nor U8302 (N_8302,N_7546,N_7872);
and U8303 (N_8303,N_8029,N_7590);
or U8304 (N_8304,N_8006,N_8001);
xnor U8305 (N_8305,N_8020,N_7839);
nor U8306 (N_8306,N_7857,N_7749);
xnor U8307 (N_8307,N_7722,N_7555);
and U8308 (N_8308,N_7952,N_7902);
nor U8309 (N_8309,N_7754,N_7606);
and U8310 (N_8310,N_7909,N_7504);
nand U8311 (N_8311,N_7574,N_7842);
and U8312 (N_8312,N_7960,N_8096);
and U8313 (N_8313,N_7817,N_7588);
nor U8314 (N_8314,N_7700,N_8135);
xor U8315 (N_8315,N_7901,N_7769);
xnor U8316 (N_8316,N_7752,N_7798);
xnor U8317 (N_8317,N_7730,N_8028);
nor U8318 (N_8318,N_8170,N_7914);
xor U8319 (N_8319,N_8107,N_7987);
xor U8320 (N_8320,N_7986,N_7542);
nand U8321 (N_8321,N_8211,N_7963);
and U8322 (N_8322,N_8110,N_8055);
nand U8323 (N_8323,N_7647,N_7726);
and U8324 (N_8324,N_8171,N_8160);
xor U8325 (N_8325,N_7734,N_7525);
and U8326 (N_8326,N_8019,N_7854);
nand U8327 (N_8327,N_8051,N_7958);
xnor U8328 (N_8328,N_7756,N_7628);
nor U8329 (N_8329,N_7687,N_8238);
nand U8330 (N_8330,N_7644,N_7829);
and U8331 (N_8331,N_7936,N_8149);
or U8332 (N_8332,N_8101,N_7553);
nand U8333 (N_8333,N_7573,N_8232);
xor U8334 (N_8334,N_7673,N_7638);
nor U8335 (N_8335,N_7711,N_7678);
nor U8336 (N_8336,N_7577,N_8216);
and U8337 (N_8337,N_7760,N_7723);
nand U8338 (N_8338,N_7652,N_7799);
or U8339 (N_8339,N_8072,N_7906);
nor U8340 (N_8340,N_7729,N_7928);
xor U8341 (N_8341,N_8132,N_7617);
xnor U8342 (N_8342,N_7637,N_8116);
xor U8343 (N_8343,N_8228,N_8147);
xnor U8344 (N_8344,N_8233,N_7871);
or U8345 (N_8345,N_7648,N_7532);
nor U8346 (N_8346,N_8095,N_8033);
and U8347 (N_8347,N_7873,N_7978);
nand U8348 (N_8348,N_8094,N_7503);
or U8349 (N_8349,N_7630,N_8173);
nor U8350 (N_8350,N_7758,N_8050);
nand U8351 (N_8351,N_7708,N_7656);
xnor U8352 (N_8352,N_7739,N_7717);
and U8353 (N_8353,N_8008,N_7693);
or U8354 (N_8354,N_8102,N_7866);
nand U8355 (N_8355,N_8084,N_7512);
xor U8356 (N_8356,N_8093,N_7537);
and U8357 (N_8357,N_8103,N_8154);
nor U8358 (N_8358,N_7709,N_7980);
or U8359 (N_8359,N_7529,N_7696);
nand U8360 (N_8360,N_7773,N_7955);
or U8361 (N_8361,N_8247,N_7894);
and U8362 (N_8362,N_7520,N_8032);
or U8363 (N_8363,N_7847,N_8097);
xnor U8364 (N_8364,N_7612,N_7927);
and U8365 (N_8365,N_8047,N_8202);
nand U8366 (N_8366,N_7742,N_7932);
nand U8367 (N_8367,N_7527,N_7792);
xnor U8368 (N_8368,N_8203,N_7965);
and U8369 (N_8369,N_8076,N_7740);
and U8370 (N_8370,N_7631,N_7879);
or U8371 (N_8371,N_8212,N_8049);
nor U8372 (N_8372,N_7825,N_8222);
xnor U8373 (N_8373,N_7679,N_8109);
or U8374 (N_8374,N_7579,N_7500);
xnor U8375 (N_8375,N_7713,N_8117);
or U8376 (N_8376,N_7755,N_7618);
nor U8377 (N_8377,N_7727,N_8104);
or U8378 (N_8378,N_7528,N_8140);
nor U8379 (N_8379,N_7905,N_7766);
or U8380 (N_8380,N_7802,N_8010);
nand U8381 (N_8381,N_8119,N_7975);
and U8382 (N_8382,N_7844,N_8125);
xor U8383 (N_8383,N_7580,N_7762);
or U8384 (N_8384,N_7791,N_8086);
nand U8385 (N_8385,N_7922,N_7908);
nor U8386 (N_8386,N_8045,N_7988);
and U8387 (N_8387,N_8068,N_7877);
nor U8388 (N_8388,N_7660,N_8146);
or U8389 (N_8389,N_7822,N_7991);
or U8390 (N_8390,N_7838,N_8036);
and U8391 (N_8391,N_8091,N_7800);
and U8392 (N_8392,N_7820,N_7657);
xor U8393 (N_8393,N_7682,N_8172);
or U8394 (N_8394,N_8180,N_7599);
nand U8395 (N_8395,N_8139,N_7714);
and U8396 (N_8396,N_7852,N_7912);
xnor U8397 (N_8397,N_7999,N_8088);
nand U8398 (N_8398,N_7556,N_7781);
and U8399 (N_8399,N_7998,N_7903);
xnor U8400 (N_8400,N_7809,N_8164);
and U8401 (N_8401,N_7995,N_7990);
or U8402 (N_8402,N_7957,N_8209);
and U8403 (N_8403,N_7539,N_7665);
and U8404 (N_8404,N_7517,N_7886);
nand U8405 (N_8405,N_7526,N_7597);
or U8406 (N_8406,N_7568,N_7830);
nor U8407 (N_8407,N_7904,N_8144);
nand U8408 (N_8408,N_7774,N_7558);
nor U8409 (N_8409,N_7934,N_7804);
nor U8410 (N_8410,N_7744,N_7698);
nand U8411 (N_8411,N_8016,N_7595);
xor U8412 (N_8412,N_8011,N_7600);
nand U8413 (N_8413,N_7941,N_8184);
xnor U8414 (N_8414,N_8214,N_7664);
nor U8415 (N_8415,N_8243,N_7731);
nor U8416 (N_8416,N_7824,N_8200);
or U8417 (N_8417,N_7938,N_7608);
xnor U8418 (N_8418,N_7586,N_7507);
or U8419 (N_8419,N_7946,N_7677);
xnor U8420 (N_8420,N_7757,N_7562);
nor U8421 (N_8421,N_7689,N_7996);
xnor U8422 (N_8422,N_7768,N_7721);
and U8423 (N_8423,N_7510,N_7861);
xor U8424 (N_8424,N_7690,N_8229);
and U8425 (N_8425,N_8137,N_7876);
nand U8426 (N_8426,N_7983,N_7855);
nand U8427 (N_8427,N_8122,N_7736);
xor U8428 (N_8428,N_8159,N_8165);
nor U8429 (N_8429,N_8121,N_7622);
or U8430 (N_8430,N_8039,N_8136);
nand U8431 (N_8431,N_7559,N_7942);
or U8432 (N_8432,N_7669,N_8245);
or U8433 (N_8433,N_8226,N_8213);
nand U8434 (N_8434,N_7702,N_7840);
and U8435 (N_8435,N_7625,N_7794);
nand U8436 (N_8436,N_7668,N_7712);
xor U8437 (N_8437,N_7795,N_7832);
nor U8438 (N_8438,N_7789,N_8151);
and U8439 (N_8439,N_8218,N_7783);
and U8440 (N_8440,N_7953,N_7826);
nand U8441 (N_8441,N_7770,N_7746);
xnor U8442 (N_8442,N_7977,N_7893);
and U8443 (N_8443,N_7544,N_7706);
and U8444 (N_8444,N_8143,N_7549);
or U8445 (N_8445,N_8167,N_7724);
or U8446 (N_8446,N_8174,N_8066);
or U8447 (N_8447,N_7536,N_7979);
nand U8448 (N_8448,N_8013,N_7897);
and U8449 (N_8449,N_7611,N_7870);
nand U8450 (N_8450,N_8067,N_8225);
nand U8451 (N_8451,N_7881,N_7653);
nand U8452 (N_8452,N_7806,N_7959);
xnor U8453 (N_8453,N_8054,N_7649);
nor U8454 (N_8454,N_7620,N_7831);
and U8455 (N_8455,N_7878,N_7502);
and U8456 (N_8456,N_7796,N_7560);
nand U8457 (N_8457,N_7925,N_8092);
or U8458 (N_8458,N_8150,N_7917);
xnor U8459 (N_8459,N_8070,N_8074);
or U8460 (N_8460,N_8007,N_7778);
nor U8461 (N_8461,N_8163,N_7968);
nand U8462 (N_8462,N_8162,N_7508);
or U8463 (N_8463,N_7743,N_7858);
and U8464 (N_8464,N_7810,N_7981);
nand U8465 (N_8465,N_7994,N_7552);
and U8466 (N_8466,N_7930,N_8193);
or U8467 (N_8467,N_8062,N_7918);
and U8468 (N_8468,N_7686,N_7524);
nor U8469 (N_8469,N_8111,N_7889);
xor U8470 (N_8470,N_7843,N_7716);
nor U8471 (N_8471,N_7735,N_8131);
nand U8472 (N_8472,N_8142,N_8105);
or U8473 (N_8473,N_8060,N_8087);
nand U8474 (N_8474,N_7654,N_7626);
nor U8475 (N_8475,N_7641,N_7951);
nor U8476 (N_8476,N_8134,N_8015);
and U8477 (N_8477,N_7915,N_7509);
nor U8478 (N_8478,N_8221,N_8042);
nor U8479 (N_8479,N_7619,N_8053);
nor U8480 (N_8480,N_8187,N_7545);
or U8481 (N_8481,N_8100,N_7614);
nand U8482 (N_8482,N_8156,N_8230);
and U8483 (N_8483,N_7598,N_8148);
nor U8484 (N_8484,N_7884,N_7604);
xnor U8485 (N_8485,N_8195,N_8106);
nand U8486 (N_8486,N_7834,N_7750);
xor U8487 (N_8487,N_7607,N_7761);
xor U8488 (N_8488,N_8120,N_8223);
and U8489 (N_8489,N_7816,N_7629);
xor U8490 (N_8490,N_7704,N_7805);
nand U8491 (N_8491,N_7801,N_8025);
or U8492 (N_8492,N_8157,N_7541);
or U8493 (N_8493,N_7956,N_8215);
xor U8494 (N_8494,N_7610,N_8205);
xnor U8495 (N_8495,N_8127,N_8017);
nand U8496 (N_8496,N_7748,N_7962);
and U8497 (N_8497,N_8040,N_7701);
nor U8498 (N_8498,N_7567,N_8191);
nor U8499 (N_8499,N_8207,N_8038);
nand U8500 (N_8500,N_8175,N_7797);
nand U8501 (N_8501,N_8000,N_7940);
or U8502 (N_8502,N_7883,N_7910);
nand U8503 (N_8503,N_8115,N_7920);
and U8504 (N_8504,N_7911,N_7655);
and U8505 (N_8505,N_7593,N_7880);
nand U8506 (N_8506,N_8192,N_7790);
and U8507 (N_8507,N_7982,N_8188);
and U8508 (N_8508,N_8057,N_7933);
nand U8509 (N_8509,N_7578,N_7591);
and U8510 (N_8510,N_8030,N_7882);
nand U8511 (N_8511,N_8240,N_7788);
and U8512 (N_8512,N_8169,N_7615);
or U8513 (N_8513,N_7601,N_8118);
nor U8514 (N_8514,N_8201,N_8034);
xor U8515 (N_8515,N_7613,N_7720);
xnor U8516 (N_8516,N_7699,N_7945);
nand U8517 (N_8517,N_7819,N_8124);
or U8518 (N_8518,N_7658,N_7913);
and U8519 (N_8519,N_8112,N_7814);
nand U8520 (N_8520,N_7898,N_8089);
and U8521 (N_8521,N_7924,N_7636);
or U8522 (N_8522,N_7859,N_7672);
and U8523 (N_8523,N_8217,N_8018);
nand U8524 (N_8524,N_8241,N_7685);
nor U8525 (N_8525,N_7547,N_8071);
nand U8526 (N_8526,N_7594,N_8182);
nor U8527 (N_8527,N_7900,N_7815);
and U8528 (N_8528,N_7667,N_7896);
nor U8529 (N_8529,N_7623,N_7753);
xnor U8530 (N_8530,N_8178,N_7589);
nand U8531 (N_8531,N_8002,N_7643);
and U8532 (N_8532,N_7862,N_8061);
or U8533 (N_8533,N_7659,N_7892);
and U8534 (N_8534,N_8197,N_7869);
nand U8535 (N_8535,N_7793,N_7585);
xnor U8536 (N_8536,N_8003,N_7888);
and U8537 (N_8537,N_8206,N_8196);
nor U8538 (N_8538,N_7680,N_7845);
or U8539 (N_8539,N_8059,N_7666);
nor U8540 (N_8540,N_7807,N_8249);
nand U8541 (N_8541,N_8183,N_7651);
nor U8542 (N_8542,N_8133,N_8027);
or U8543 (N_8543,N_7944,N_7635);
nor U8544 (N_8544,N_7966,N_7738);
nand U8545 (N_8545,N_7874,N_8186);
nor U8546 (N_8546,N_7823,N_8181);
nor U8547 (N_8547,N_7841,N_7605);
xor U8548 (N_8548,N_7764,N_7674);
xnor U8549 (N_8549,N_7885,N_7972);
nor U8550 (N_8550,N_7782,N_7745);
and U8551 (N_8551,N_7765,N_8129);
nor U8552 (N_8552,N_8041,N_7725);
xnor U8553 (N_8553,N_8153,N_7868);
nand U8554 (N_8554,N_7596,N_8219);
or U8555 (N_8555,N_7645,N_7621);
and U8556 (N_8556,N_8023,N_8236);
and U8557 (N_8557,N_7772,N_7650);
xor U8558 (N_8558,N_7777,N_7784);
and U8559 (N_8559,N_8242,N_7575);
xnor U8560 (N_8560,N_7984,N_8237);
nand U8561 (N_8561,N_7780,N_8026);
and U8562 (N_8562,N_8220,N_8083);
or U8563 (N_8563,N_8179,N_7961);
and U8564 (N_8564,N_7511,N_7808);
and U8565 (N_8565,N_7681,N_7846);
xnor U8566 (N_8566,N_8044,N_7670);
xnor U8567 (N_8567,N_7992,N_7923);
xor U8568 (N_8568,N_8190,N_7950);
and U8569 (N_8569,N_8081,N_8048);
and U8570 (N_8570,N_8073,N_7943);
nor U8571 (N_8571,N_8085,N_8043);
and U8572 (N_8572,N_7827,N_8138);
nand U8573 (N_8573,N_7974,N_8145);
nand U8574 (N_8574,N_7639,N_7583);
and U8575 (N_8575,N_8208,N_7989);
xor U8576 (N_8576,N_7733,N_8235);
or U8577 (N_8577,N_7543,N_8069);
xnor U8578 (N_8578,N_8022,N_8231);
nand U8579 (N_8579,N_7695,N_7703);
and U8580 (N_8580,N_8176,N_7836);
nand U8581 (N_8581,N_7691,N_7581);
nor U8582 (N_8582,N_7747,N_7564);
or U8583 (N_8583,N_8185,N_7710);
nand U8584 (N_8584,N_7811,N_7627);
xnor U8585 (N_8585,N_8114,N_7705);
and U8586 (N_8586,N_8065,N_7875);
and U8587 (N_8587,N_8012,N_7584);
nand U8588 (N_8588,N_7954,N_8198);
or U8589 (N_8589,N_7640,N_7518);
or U8590 (N_8590,N_7692,N_7565);
nand U8591 (N_8591,N_8152,N_7557);
and U8592 (N_8592,N_7642,N_7926);
nor U8593 (N_8593,N_7531,N_7779);
or U8594 (N_8594,N_7561,N_7828);
or U8595 (N_8595,N_7616,N_7694);
xor U8596 (N_8596,N_8239,N_8009);
or U8597 (N_8597,N_7566,N_7514);
nor U8598 (N_8598,N_7728,N_7891);
and U8599 (N_8599,N_8031,N_7741);
or U8600 (N_8600,N_8210,N_8021);
or U8601 (N_8601,N_7662,N_7634);
nor U8602 (N_8602,N_7506,N_7576);
nor U8603 (N_8603,N_7572,N_7851);
nor U8604 (N_8604,N_7538,N_7887);
xnor U8605 (N_8605,N_8037,N_8063);
xor U8606 (N_8606,N_7853,N_8077);
xnor U8607 (N_8607,N_7821,N_8082);
xor U8608 (N_8608,N_8224,N_7534);
nand U8609 (N_8609,N_7776,N_7919);
nor U8610 (N_8610,N_7863,N_7860);
nand U8611 (N_8611,N_7867,N_7697);
and U8612 (N_8612,N_7833,N_8004);
or U8613 (N_8613,N_8024,N_7675);
nand U8614 (N_8614,N_8005,N_7719);
nor U8615 (N_8615,N_7907,N_8246);
xnor U8616 (N_8616,N_8199,N_8141);
and U8617 (N_8617,N_8058,N_7533);
nand U8618 (N_8618,N_8052,N_7663);
nor U8619 (N_8619,N_7519,N_7899);
and U8620 (N_8620,N_7550,N_7767);
or U8621 (N_8621,N_7759,N_7813);
or U8622 (N_8622,N_7501,N_7715);
nor U8623 (N_8623,N_8177,N_7563);
or U8624 (N_8624,N_7763,N_7786);
xor U8625 (N_8625,N_7572,N_7839);
nor U8626 (N_8626,N_7670,N_8102);
xnor U8627 (N_8627,N_7900,N_7832);
or U8628 (N_8628,N_7807,N_8048);
nor U8629 (N_8629,N_7856,N_7510);
or U8630 (N_8630,N_7526,N_7980);
or U8631 (N_8631,N_8204,N_8161);
or U8632 (N_8632,N_8166,N_7592);
and U8633 (N_8633,N_7594,N_8181);
or U8634 (N_8634,N_7670,N_8118);
xnor U8635 (N_8635,N_7632,N_7534);
nand U8636 (N_8636,N_8053,N_8198);
nor U8637 (N_8637,N_7903,N_7965);
xor U8638 (N_8638,N_7977,N_7930);
nor U8639 (N_8639,N_7801,N_7911);
or U8640 (N_8640,N_7980,N_8136);
xor U8641 (N_8641,N_7635,N_7757);
xnor U8642 (N_8642,N_7780,N_7866);
nand U8643 (N_8643,N_7640,N_7765);
nor U8644 (N_8644,N_7739,N_7579);
or U8645 (N_8645,N_8237,N_8211);
and U8646 (N_8646,N_7643,N_8165);
nand U8647 (N_8647,N_7855,N_7836);
nor U8648 (N_8648,N_8032,N_7529);
xor U8649 (N_8649,N_7724,N_7661);
nor U8650 (N_8650,N_8204,N_7756);
and U8651 (N_8651,N_8145,N_7704);
nand U8652 (N_8652,N_7995,N_8166);
and U8653 (N_8653,N_7702,N_8088);
nor U8654 (N_8654,N_8098,N_7538);
xnor U8655 (N_8655,N_8171,N_7601);
or U8656 (N_8656,N_7599,N_8183);
nor U8657 (N_8657,N_8039,N_7703);
nand U8658 (N_8658,N_8182,N_7532);
or U8659 (N_8659,N_8074,N_7532);
nor U8660 (N_8660,N_7911,N_8221);
nor U8661 (N_8661,N_7755,N_8199);
nand U8662 (N_8662,N_7876,N_7913);
xnor U8663 (N_8663,N_7603,N_8109);
xor U8664 (N_8664,N_7672,N_7815);
nor U8665 (N_8665,N_7680,N_7560);
and U8666 (N_8666,N_7937,N_7970);
nand U8667 (N_8667,N_7523,N_7574);
and U8668 (N_8668,N_7937,N_7833);
xor U8669 (N_8669,N_7704,N_7993);
nor U8670 (N_8670,N_8013,N_7710);
nor U8671 (N_8671,N_8198,N_8208);
xor U8672 (N_8672,N_7897,N_7956);
xnor U8673 (N_8673,N_8150,N_7835);
nor U8674 (N_8674,N_8166,N_7620);
and U8675 (N_8675,N_8202,N_7775);
nor U8676 (N_8676,N_8078,N_7952);
nor U8677 (N_8677,N_7799,N_7715);
and U8678 (N_8678,N_7825,N_7901);
and U8679 (N_8679,N_8012,N_8093);
nor U8680 (N_8680,N_8121,N_7923);
nor U8681 (N_8681,N_7826,N_7793);
or U8682 (N_8682,N_7570,N_7625);
xor U8683 (N_8683,N_7854,N_7904);
nor U8684 (N_8684,N_7538,N_8235);
nor U8685 (N_8685,N_7734,N_7770);
or U8686 (N_8686,N_7866,N_7827);
and U8687 (N_8687,N_7840,N_8041);
and U8688 (N_8688,N_7874,N_8144);
nor U8689 (N_8689,N_8119,N_7617);
nor U8690 (N_8690,N_7877,N_8066);
and U8691 (N_8691,N_7534,N_7907);
xor U8692 (N_8692,N_7767,N_7739);
and U8693 (N_8693,N_7970,N_7704);
and U8694 (N_8694,N_7706,N_8073);
and U8695 (N_8695,N_8194,N_7984);
and U8696 (N_8696,N_7985,N_8101);
xnor U8697 (N_8697,N_7685,N_8159);
xnor U8698 (N_8698,N_7575,N_8065);
nor U8699 (N_8699,N_7837,N_8057);
and U8700 (N_8700,N_7683,N_8178);
nor U8701 (N_8701,N_7975,N_8151);
or U8702 (N_8702,N_8048,N_7851);
xor U8703 (N_8703,N_8112,N_7879);
nand U8704 (N_8704,N_7691,N_7657);
or U8705 (N_8705,N_7837,N_7554);
nand U8706 (N_8706,N_7710,N_7997);
nand U8707 (N_8707,N_8044,N_7780);
nor U8708 (N_8708,N_7525,N_7762);
and U8709 (N_8709,N_8037,N_7525);
or U8710 (N_8710,N_7734,N_8234);
nand U8711 (N_8711,N_8123,N_7856);
or U8712 (N_8712,N_7933,N_7912);
xnor U8713 (N_8713,N_7908,N_8071);
xor U8714 (N_8714,N_7692,N_7621);
nor U8715 (N_8715,N_7634,N_8096);
nor U8716 (N_8716,N_7749,N_7836);
nand U8717 (N_8717,N_7756,N_8227);
and U8718 (N_8718,N_8142,N_8029);
xnor U8719 (N_8719,N_7559,N_8096);
nor U8720 (N_8720,N_7525,N_7519);
xor U8721 (N_8721,N_7542,N_8002);
and U8722 (N_8722,N_8020,N_7928);
or U8723 (N_8723,N_8015,N_8086);
xor U8724 (N_8724,N_7888,N_7728);
or U8725 (N_8725,N_8070,N_7819);
and U8726 (N_8726,N_8082,N_7793);
xnor U8727 (N_8727,N_7880,N_7933);
or U8728 (N_8728,N_7734,N_8241);
and U8729 (N_8729,N_7811,N_7941);
nor U8730 (N_8730,N_7542,N_8137);
or U8731 (N_8731,N_7650,N_8138);
and U8732 (N_8732,N_8181,N_7737);
nor U8733 (N_8733,N_8001,N_7760);
or U8734 (N_8734,N_8027,N_7995);
nand U8735 (N_8735,N_8134,N_8135);
nor U8736 (N_8736,N_7808,N_7630);
xnor U8737 (N_8737,N_8218,N_7651);
nand U8738 (N_8738,N_7639,N_7963);
nand U8739 (N_8739,N_7572,N_8165);
and U8740 (N_8740,N_7682,N_7838);
and U8741 (N_8741,N_7985,N_7646);
nand U8742 (N_8742,N_8235,N_7890);
and U8743 (N_8743,N_8094,N_8175);
or U8744 (N_8744,N_8242,N_7792);
xor U8745 (N_8745,N_7747,N_8037);
nor U8746 (N_8746,N_8126,N_7926);
nand U8747 (N_8747,N_8092,N_8180);
xnor U8748 (N_8748,N_8222,N_7802);
nor U8749 (N_8749,N_8140,N_7729);
nand U8750 (N_8750,N_7662,N_7674);
xnor U8751 (N_8751,N_7692,N_7965);
xor U8752 (N_8752,N_8201,N_8162);
nor U8753 (N_8753,N_7954,N_7691);
xnor U8754 (N_8754,N_7564,N_7780);
xnor U8755 (N_8755,N_7515,N_8156);
and U8756 (N_8756,N_8208,N_7502);
xnor U8757 (N_8757,N_7519,N_7943);
xor U8758 (N_8758,N_7987,N_8150);
or U8759 (N_8759,N_7535,N_8098);
xor U8760 (N_8760,N_8170,N_7711);
nor U8761 (N_8761,N_8133,N_7825);
or U8762 (N_8762,N_7589,N_8237);
or U8763 (N_8763,N_7879,N_7860);
xor U8764 (N_8764,N_7916,N_8121);
or U8765 (N_8765,N_8235,N_7571);
and U8766 (N_8766,N_7803,N_8140);
and U8767 (N_8767,N_8171,N_7781);
or U8768 (N_8768,N_8090,N_8026);
and U8769 (N_8769,N_8072,N_7860);
and U8770 (N_8770,N_8134,N_7977);
nor U8771 (N_8771,N_8138,N_8038);
nand U8772 (N_8772,N_7907,N_8028);
or U8773 (N_8773,N_7512,N_7851);
or U8774 (N_8774,N_7887,N_8038);
or U8775 (N_8775,N_8116,N_7928);
xor U8776 (N_8776,N_7842,N_7786);
and U8777 (N_8777,N_8126,N_7874);
nand U8778 (N_8778,N_8037,N_7603);
nor U8779 (N_8779,N_7666,N_7637);
and U8780 (N_8780,N_7962,N_8006);
xnor U8781 (N_8781,N_7725,N_7850);
xnor U8782 (N_8782,N_8124,N_7747);
nand U8783 (N_8783,N_7664,N_7689);
or U8784 (N_8784,N_8186,N_8195);
and U8785 (N_8785,N_7848,N_7855);
xnor U8786 (N_8786,N_8224,N_8049);
or U8787 (N_8787,N_7653,N_7988);
nor U8788 (N_8788,N_7932,N_8165);
nor U8789 (N_8789,N_7871,N_7533);
nor U8790 (N_8790,N_7727,N_8133);
or U8791 (N_8791,N_7639,N_7528);
xor U8792 (N_8792,N_7546,N_7635);
nor U8793 (N_8793,N_7757,N_7993);
nand U8794 (N_8794,N_7629,N_7789);
or U8795 (N_8795,N_7677,N_7661);
nor U8796 (N_8796,N_7567,N_7683);
nor U8797 (N_8797,N_8034,N_7980);
xnor U8798 (N_8798,N_8190,N_7854);
nand U8799 (N_8799,N_8123,N_7548);
nor U8800 (N_8800,N_7668,N_7672);
and U8801 (N_8801,N_7757,N_8244);
nor U8802 (N_8802,N_8088,N_7686);
nand U8803 (N_8803,N_7917,N_7637);
nor U8804 (N_8804,N_7606,N_8040);
nand U8805 (N_8805,N_7620,N_8055);
xor U8806 (N_8806,N_8010,N_8074);
nor U8807 (N_8807,N_8228,N_7772);
xnor U8808 (N_8808,N_7816,N_7630);
xnor U8809 (N_8809,N_7837,N_7663);
xor U8810 (N_8810,N_7551,N_8238);
xnor U8811 (N_8811,N_7505,N_7777);
nor U8812 (N_8812,N_7730,N_7724);
nor U8813 (N_8813,N_8111,N_7994);
xnor U8814 (N_8814,N_8023,N_8161);
nand U8815 (N_8815,N_7569,N_8038);
nor U8816 (N_8816,N_7989,N_7879);
nand U8817 (N_8817,N_7863,N_8155);
or U8818 (N_8818,N_7955,N_8214);
and U8819 (N_8819,N_7768,N_7990);
nor U8820 (N_8820,N_8235,N_8055);
nand U8821 (N_8821,N_7642,N_7869);
and U8822 (N_8822,N_7595,N_7928);
xnor U8823 (N_8823,N_7646,N_7806);
nor U8824 (N_8824,N_8117,N_8171);
nor U8825 (N_8825,N_7902,N_7781);
nand U8826 (N_8826,N_8208,N_8175);
xor U8827 (N_8827,N_7920,N_8026);
and U8828 (N_8828,N_8149,N_7736);
or U8829 (N_8829,N_7564,N_8091);
nand U8830 (N_8830,N_7712,N_7801);
nor U8831 (N_8831,N_7666,N_7654);
nor U8832 (N_8832,N_8092,N_7576);
and U8833 (N_8833,N_8044,N_7633);
and U8834 (N_8834,N_7828,N_7711);
xor U8835 (N_8835,N_7942,N_7806);
nor U8836 (N_8836,N_7518,N_7867);
and U8837 (N_8837,N_7551,N_7946);
xor U8838 (N_8838,N_8002,N_7781);
or U8839 (N_8839,N_7953,N_7510);
and U8840 (N_8840,N_7635,N_7827);
or U8841 (N_8841,N_8194,N_8083);
nor U8842 (N_8842,N_7878,N_7764);
and U8843 (N_8843,N_8231,N_8163);
and U8844 (N_8844,N_8226,N_7637);
xor U8845 (N_8845,N_8110,N_7713);
and U8846 (N_8846,N_8006,N_7728);
nor U8847 (N_8847,N_7672,N_7838);
nand U8848 (N_8848,N_8242,N_8091);
nand U8849 (N_8849,N_8063,N_8160);
nor U8850 (N_8850,N_7668,N_7793);
xor U8851 (N_8851,N_7917,N_7856);
xnor U8852 (N_8852,N_7571,N_7923);
and U8853 (N_8853,N_7607,N_7781);
nor U8854 (N_8854,N_7583,N_8237);
xnor U8855 (N_8855,N_7739,N_7682);
nor U8856 (N_8856,N_8048,N_7671);
or U8857 (N_8857,N_8159,N_7558);
nor U8858 (N_8858,N_7739,N_8219);
or U8859 (N_8859,N_7634,N_7784);
nor U8860 (N_8860,N_7934,N_7924);
nand U8861 (N_8861,N_8150,N_8148);
xor U8862 (N_8862,N_7535,N_8186);
or U8863 (N_8863,N_8163,N_7662);
xnor U8864 (N_8864,N_7806,N_7609);
xor U8865 (N_8865,N_7894,N_7504);
nand U8866 (N_8866,N_7553,N_7525);
nand U8867 (N_8867,N_8075,N_8073);
and U8868 (N_8868,N_7524,N_7908);
nand U8869 (N_8869,N_7881,N_8031);
nand U8870 (N_8870,N_8082,N_7940);
or U8871 (N_8871,N_7949,N_7631);
and U8872 (N_8872,N_7829,N_7655);
xnor U8873 (N_8873,N_7820,N_8001);
xnor U8874 (N_8874,N_7661,N_8096);
xnor U8875 (N_8875,N_7766,N_7755);
nor U8876 (N_8876,N_7709,N_7771);
nand U8877 (N_8877,N_7549,N_8223);
and U8878 (N_8878,N_8218,N_7717);
nand U8879 (N_8879,N_7539,N_7792);
and U8880 (N_8880,N_8139,N_7818);
and U8881 (N_8881,N_7861,N_7760);
and U8882 (N_8882,N_7804,N_8046);
nand U8883 (N_8883,N_7652,N_8157);
xnor U8884 (N_8884,N_7922,N_7819);
nor U8885 (N_8885,N_7929,N_7564);
nand U8886 (N_8886,N_7829,N_7725);
xor U8887 (N_8887,N_7521,N_8112);
xor U8888 (N_8888,N_7786,N_8068);
and U8889 (N_8889,N_8219,N_7636);
nor U8890 (N_8890,N_7662,N_7827);
and U8891 (N_8891,N_7844,N_7927);
and U8892 (N_8892,N_7524,N_7841);
nand U8893 (N_8893,N_7649,N_7909);
or U8894 (N_8894,N_8199,N_7507);
nand U8895 (N_8895,N_7851,N_7527);
nand U8896 (N_8896,N_8214,N_8035);
xnor U8897 (N_8897,N_7718,N_7626);
nand U8898 (N_8898,N_7883,N_8163);
nor U8899 (N_8899,N_7794,N_7547);
or U8900 (N_8900,N_8228,N_7736);
nand U8901 (N_8901,N_7552,N_8104);
and U8902 (N_8902,N_8190,N_7896);
nor U8903 (N_8903,N_8196,N_8130);
nor U8904 (N_8904,N_7794,N_7680);
nor U8905 (N_8905,N_7928,N_7585);
and U8906 (N_8906,N_7615,N_8173);
and U8907 (N_8907,N_8038,N_8170);
xor U8908 (N_8908,N_8175,N_7849);
or U8909 (N_8909,N_7725,N_7791);
or U8910 (N_8910,N_7906,N_7552);
nand U8911 (N_8911,N_8149,N_7770);
and U8912 (N_8912,N_8197,N_7536);
xor U8913 (N_8913,N_7885,N_8174);
and U8914 (N_8914,N_8083,N_7863);
or U8915 (N_8915,N_8218,N_7727);
or U8916 (N_8916,N_7822,N_7716);
nand U8917 (N_8917,N_8177,N_7789);
nor U8918 (N_8918,N_7920,N_7656);
and U8919 (N_8919,N_7655,N_7562);
or U8920 (N_8920,N_7777,N_7736);
nand U8921 (N_8921,N_7901,N_7858);
nand U8922 (N_8922,N_7960,N_7760);
nor U8923 (N_8923,N_7535,N_8190);
and U8924 (N_8924,N_7868,N_7803);
and U8925 (N_8925,N_7754,N_7512);
or U8926 (N_8926,N_8108,N_7895);
or U8927 (N_8927,N_7556,N_7737);
or U8928 (N_8928,N_7836,N_7985);
or U8929 (N_8929,N_8087,N_7705);
nand U8930 (N_8930,N_7805,N_8051);
nor U8931 (N_8931,N_8191,N_7909);
xor U8932 (N_8932,N_7713,N_8044);
or U8933 (N_8933,N_8187,N_7634);
and U8934 (N_8934,N_7634,N_8088);
or U8935 (N_8935,N_8126,N_7695);
xnor U8936 (N_8936,N_7653,N_8089);
or U8937 (N_8937,N_7970,N_8194);
or U8938 (N_8938,N_7655,N_7776);
nor U8939 (N_8939,N_7871,N_7573);
or U8940 (N_8940,N_8119,N_7611);
and U8941 (N_8941,N_7631,N_8093);
or U8942 (N_8942,N_8060,N_8146);
nor U8943 (N_8943,N_7868,N_7648);
or U8944 (N_8944,N_8197,N_7870);
and U8945 (N_8945,N_8202,N_8183);
xnor U8946 (N_8946,N_8111,N_8220);
or U8947 (N_8947,N_8191,N_7835);
xor U8948 (N_8948,N_7725,N_7985);
xor U8949 (N_8949,N_8156,N_7813);
and U8950 (N_8950,N_8175,N_7888);
and U8951 (N_8951,N_7888,N_7551);
and U8952 (N_8952,N_8072,N_8206);
xor U8953 (N_8953,N_7941,N_7836);
and U8954 (N_8954,N_7571,N_7503);
or U8955 (N_8955,N_7904,N_7922);
xnor U8956 (N_8956,N_8147,N_8070);
nand U8957 (N_8957,N_7752,N_8152);
nor U8958 (N_8958,N_7817,N_8233);
xnor U8959 (N_8959,N_7619,N_8067);
nand U8960 (N_8960,N_7903,N_7514);
and U8961 (N_8961,N_8200,N_7631);
or U8962 (N_8962,N_8245,N_7736);
and U8963 (N_8963,N_7526,N_8055);
nand U8964 (N_8964,N_7594,N_7613);
or U8965 (N_8965,N_8086,N_7778);
and U8966 (N_8966,N_7503,N_7988);
xor U8967 (N_8967,N_8077,N_7663);
nand U8968 (N_8968,N_7506,N_7615);
nor U8969 (N_8969,N_7681,N_7530);
xor U8970 (N_8970,N_7748,N_7746);
nand U8971 (N_8971,N_8185,N_7558);
or U8972 (N_8972,N_8103,N_7901);
or U8973 (N_8973,N_8010,N_7969);
nand U8974 (N_8974,N_7713,N_8130);
and U8975 (N_8975,N_7779,N_7683);
and U8976 (N_8976,N_7684,N_7728);
and U8977 (N_8977,N_8013,N_7767);
or U8978 (N_8978,N_7762,N_7832);
or U8979 (N_8979,N_8118,N_8234);
nor U8980 (N_8980,N_8189,N_8181);
nor U8981 (N_8981,N_8074,N_7916);
and U8982 (N_8982,N_7870,N_7705);
xor U8983 (N_8983,N_7907,N_7971);
or U8984 (N_8984,N_7522,N_7856);
or U8985 (N_8985,N_7951,N_8097);
or U8986 (N_8986,N_7997,N_7682);
xor U8987 (N_8987,N_7641,N_8132);
nor U8988 (N_8988,N_7998,N_7787);
nor U8989 (N_8989,N_8121,N_8179);
xor U8990 (N_8990,N_7784,N_8209);
xnor U8991 (N_8991,N_7748,N_7698);
and U8992 (N_8992,N_7775,N_8065);
nor U8993 (N_8993,N_8142,N_7534);
nand U8994 (N_8994,N_7922,N_8082);
nor U8995 (N_8995,N_7648,N_8214);
or U8996 (N_8996,N_7821,N_7833);
nor U8997 (N_8997,N_7783,N_7983);
xnor U8998 (N_8998,N_7651,N_7584);
or U8999 (N_8999,N_8193,N_8153);
and U9000 (N_9000,N_8806,N_8887);
and U9001 (N_9001,N_8713,N_8342);
xor U9002 (N_9002,N_8569,N_8586);
xor U9003 (N_9003,N_8476,N_8423);
and U9004 (N_9004,N_8381,N_8781);
nand U9005 (N_9005,N_8520,N_8572);
nor U9006 (N_9006,N_8928,N_8462);
nor U9007 (N_9007,N_8733,N_8338);
xor U9008 (N_9008,N_8295,N_8922);
nand U9009 (N_9009,N_8517,N_8854);
xor U9010 (N_9010,N_8348,N_8253);
nand U9011 (N_9011,N_8392,N_8876);
nand U9012 (N_9012,N_8536,N_8846);
xor U9013 (N_9013,N_8659,N_8465);
and U9014 (N_9014,N_8848,N_8768);
and U9015 (N_9015,N_8655,N_8608);
nand U9016 (N_9016,N_8672,N_8651);
nor U9017 (N_9017,N_8705,N_8256);
or U9018 (N_9018,N_8686,N_8561);
xnor U9019 (N_9019,N_8716,N_8435);
or U9020 (N_9020,N_8252,N_8552);
or U9021 (N_9021,N_8573,N_8543);
and U9022 (N_9022,N_8680,N_8912);
or U9023 (N_9023,N_8355,N_8653);
or U9024 (N_9024,N_8756,N_8636);
nand U9025 (N_9025,N_8640,N_8769);
or U9026 (N_9026,N_8808,N_8315);
nand U9027 (N_9027,N_8578,N_8766);
nand U9028 (N_9028,N_8558,N_8873);
or U9029 (N_9029,N_8879,N_8981);
nor U9030 (N_9030,N_8683,N_8959);
nand U9031 (N_9031,N_8557,N_8396);
nor U9032 (N_9032,N_8286,N_8376);
and U9033 (N_9033,N_8741,N_8635);
or U9034 (N_9034,N_8383,N_8938);
or U9035 (N_9035,N_8496,N_8633);
nand U9036 (N_9036,N_8772,N_8830);
or U9037 (N_9037,N_8263,N_8298);
xnor U9038 (N_9038,N_8992,N_8625);
nor U9039 (N_9039,N_8841,N_8566);
nor U9040 (N_9040,N_8916,N_8461);
xnor U9041 (N_9041,N_8583,N_8357);
xor U9042 (N_9042,N_8454,N_8626);
xor U9043 (N_9043,N_8388,N_8744);
nand U9044 (N_9044,N_8820,N_8750);
nor U9045 (N_9045,N_8782,N_8731);
xor U9046 (N_9046,N_8466,N_8896);
xnor U9047 (N_9047,N_8732,N_8574);
xor U9048 (N_9048,N_8884,N_8589);
nor U9049 (N_9049,N_8923,N_8949);
and U9050 (N_9050,N_8950,N_8845);
xor U9051 (N_9051,N_8330,N_8762);
xor U9052 (N_9052,N_8765,N_8800);
or U9053 (N_9053,N_8576,N_8620);
nor U9054 (N_9054,N_8555,N_8404);
xnor U9055 (N_9055,N_8260,N_8316);
nor U9056 (N_9056,N_8798,N_8527);
or U9057 (N_9057,N_8774,N_8562);
nor U9058 (N_9058,N_8365,N_8850);
and U9059 (N_9059,N_8508,N_8691);
nand U9060 (N_9060,N_8952,N_8727);
and U9061 (N_9061,N_8832,N_8687);
nor U9062 (N_9062,N_8619,N_8953);
nand U9063 (N_9063,N_8792,N_8825);
and U9064 (N_9064,N_8473,N_8723);
or U9065 (N_9065,N_8585,N_8598);
and U9066 (N_9066,N_8497,N_8826);
nand U9067 (N_9067,N_8682,N_8855);
or U9068 (N_9068,N_8803,N_8936);
nand U9069 (N_9069,N_8991,N_8951);
and U9070 (N_9070,N_8487,N_8307);
or U9071 (N_9071,N_8968,N_8417);
nand U9072 (N_9072,N_8872,N_8665);
and U9073 (N_9073,N_8748,N_8865);
xnor U9074 (N_9074,N_8373,N_8692);
nor U9075 (N_9075,N_8931,N_8455);
and U9076 (N_9076,N_8515,N_8366);
and U9077 (N_9077,N_8451,N_8789);
and U9078 (N_9078,N_8269,N_8394);
nor U9079 (N_9079,N_8804,N_8614);
nand U9080 (N_9080,N_8433,N_8384);
and U9081 (N_9081,N_8697,N_8982);
nor U9082 (N_9082,N_8346,N_8272);
and U9083 (N_9083,N_8282,N_8322);
xnor U9084 (N_9084,N_8324,N_8809);
nand U9085 (N_9085,N_8279,N_8954);
or U9086 (N_9086,N_8314,N_8334);
xor U9087 (N_9087,N_8743,N_8471);
nor U9088 (N_9088,N_8593,N_8823);
nor U9089 (N_9089,N_8345,N_8546);
xor U9090 (N_9090,N_8630,N_8399);
nor U9091 (N_9091,N_8979,N_8746);
nor U9092 (N_9092,N_8313,N_8590);
xnor U9093 (N_9093,N_8507,N_8389);
or U9094 (N_9094,N_8976,N_8791);
or U9095 (N_9095,N_8627,N_8747);
and U9096 (N_9096,N_8988,N_8405);
nor U9097 (N_9097,N_8822,N_8445);
xor U9098 (N_9098,N_8698,N_8251);
nand U9099 (N_9099,N_8980,N_8767);
nor U9100 (N_9100,N_8592,N_8358);
nor U9101 (N_9101,N_8475,N_8450);
or U9102 (N_9102,N_8658,N_8983);
or U9103 (N_9103,N_8693,N_8694);
and U9104 (N_9104,N_8679,N_8479);
or U9105 (N_9105,N_8429,N_8704);
nand U9106 (N_9106,N_8927,N_8641);
nor U9107 (N_9107,N_8901,N_8660);
and U9108 (N_9108,N_8737,N_8439);
xnor U9109 (N_9109,N_8638,N_8794);
nand U9110 (N_9110,N_8735,N_8844);
nand U9111 (N_9111,N_8728,N_8973);
and U9112 (N_9112,N_8637,N_8333);
xor U9113 (N_9113,N_8354,N_8711);
xor U9114 (N_9114,N_8730,N_8814);
and U9115 (N_9115,N_8488,N_8412);
xnor U9116 (N_9116,N_8612,N_8788);
xor U9117 (N_9117,N_8519,N_8472);
and U9118 (N_9118,N_8430,N_8395);
nor U9119 (N_9119,N_8371,N_8734);
nor U9120 (N_9120,N_8784,N_8971);
nand U9121 (N_9121,N_8289,N_8915);
xnor U9122 (N_9122,N_8904,N_8930);
nand U9123 (N_9123,N_8821,N_8288);
nor U9124 (N_9124,N_8828,N_8688);
nand U9125 (N_9125,N_8866,N_8560);
or U9126 (N_9126,N_8761,N_8443);
and U9127 (N_9127,N_8894,N_8646);
nand U9128 (N_9128,N_8382,N_8745);
and U9129 (N_9129,N_8611,N_8531);
nand U9130 (N_9130,N_8588,N_8601);
nand U9131 (N_9131,N_8960,N_8720);
xor U9132 (N_9132,N_8474,N_8427);
or U9133 (N_9133,N_8503,N_8538);
nand U9134 (N_9134,N_8709,N_8287);
nand U9135 (N_9135,N_8993,N_8987);
and U9136 (N_9136,N_8671,N_8736);
or U9137 (N_9137,N_8550,N_8707);
nand U9138 (N_9138,N_8615,N_8575);
xor U9139 (N_9139,N_8401,N_8779);
or U9140 (N_9140,N_8778,N_8514);
nor U9141 (N_9141,N_8926,N_8380);
or U9142 (N_9142,N_8596,N_8512);
or U9143 (N_9143,N_8426,N_8511);
and U9144 (N_9144,N_8858,N_8281);
or U9145 (N_9145,N_8624,N_8668);
nand U9146 (N_9146,N_8403,N_8483);
or U9147 (N_9147,N_8311,N_8363);
xor U9148 (N_9148,N_8861,N_8907);
or U9149 (N_9149,N_8622,N_8852);
or U9150 (N_9150,N_8431,N_8932);
nand U9151 (N_9151,N_8787,N_8890);
nor U9152 (N_9152,N_8262,N_8724);
and U9153 (N_9153,N_8325,N_8336);
nor U9154 (N_9154,N_8886,N_8367);
and U9155 (N_9155,N_8903,N_8347);
or U9156 (N_9156,N_8975,N_8594);
xnor U9157 (N_9157,N_8292,N_8994);
or U9158 (N_9158,N_8948,N_8456);
xnor U9159 (N_9159,N_8621,N_8811);
and U9160 (N_9160,N_8795,N_8463);
and U9161 (N_9161,N_8364,N_8924);
nor U9162 (N_9162,N_8934,N_8917);
nand U9163 (N_9163,N_8985,N_8352);
xnor U9164 (N_9164,N_8967,N_8480);
nor U9165 (N_9165,N_8265,N_8486);
and U9166 (N_9166,N_8397,N_8670);
nand U9167 (N_9167,N_8510,N_8521);
nand U9168 (N_9168,N_8391,N_8437);
and U9169 (N_9169,N_8498,N_8824);
and U9170 (N_9170,N_8673,N_8317);
xnor U9171 (N_9171,N_8897,N_8337);
or U9172 (N_9172,N_8319,N_8742);
xor U9173 (N_9173,N_8356,N_8906);
or U9174 (N_9174,N_8644,N_8947);
and U9175 (N_9175,N_8387,N_8810);
nor U9176 (N_9176,N_8714,N_8564);
nand U9177 (N_9177,N_8977,N_8616);
and U9178 (N_9178,N_8296,N_8489);
nor U9179 (N_9179,N_8604,N_8523);
or U9180 (N_9180,N_8664,N_8532);
nand U9181 (N_9181,N_8999,N_8500);
nor U9182 (N_9182,N_8409,N_8442);
and U9183 (N_9183,N_8819,N_8533);
nor U9184 (N_9184,N_8280,N_8911);
nor U9185 (N_9185,N_8722,N_8448);
or U9186 (N_9186,N_8678,N_8544);
xor U9187 (N_9187,N_8299,N_8353);
nand U9188 (N_9188,N_8413,N_8610);
xor U9189 (N_9189,N_8602,N_8918);
or U9190 (N_9190,N_8955,N_8870);
or U9191 (N_9191,N_8648,N_8470);
and U9192 (N_9192,N_8509,N_8963);
nand U9193 (N_9193,N_8309,N_8266);
xor U9194 (N_9194,N_8502,N_8418);
nand U9195 (N_9195,N_8556,N_8339);
and U9196 (N_9196,N_8888,N_8853);
or U9197 (N_9197,N_8522,N_8343);
nor U9198 (N_9198,N_8892,N_8807);
nor U9199 (N_9199,N_8677,N_8525);
or U9200 (N_9200,N_8283,N_8827);
and U9201 (N_9201,N_8468,N_8940);
or U9202 (N_9202,N_8419,N_8303);
and U9203 (N_9203,N_8817,N_8833);
xnor U9204 (N_9204,N_8494,N_8460);
nand U9205 (N_9205,N_8900,N_8970);
nor U9206 (N_9206,N_8290,N_8889);
xor U9207 (N_9207,N_8681,N_8447);
or U9208 (N_9208,N_8416,N_8554);
nor U9209 (N_9209,N_8293,N_8529);
nor U9210 (N_9210,N_8368,N_8351);
xnor U9211 (N_9211,N_8751,N_8754);
or U9212 (N_9212,N_8831,N_8542);
and U9213 (N_9213,N_8871,N_8607);
nand U9214 (N_9214,N_8905,N_8493);
or U9215 (N_9215,N_8370,N_8689);
xnor U9216 (N_9216,N_8857,N_8440);
xor U9217 (N_9217,N_8882,N_8577);
and U9218 (N_9218,N_8261,N_8535);
nand U9219 (N_9219,N_8268,N_8377);
or U9220 (N_9220,N_8941,N_8258);
xor U9221 (N_9221,N_8643,N_8839);
xor U9222 (N_9222,N_8267,N_8835);
and U9223 (N_9223,N_8801,N_8369);
nor U9224 (N_9224,N_8972,N_8524);
nor U9225 (N_9225,N_8790,N_8320);
xnor U9226 (N_9226,N_8895,N_8652);
xnor U9227 (N_9227,N_8961,N_8410);
xnor U9228 (N_9228,N_8591,N_8957);
xor U9229 (N_9229,N_8250,N_8780);
and U9230 (N_9230,N_8675,N_8402);
xnor U9231 (N_9231,N_8582,N_8937);
nor U9232 (N_9232,N_8703,N_8385);
xor U9233 (N_9233,N_8492,N_8306);
xor U9234 (N_9234,N_8308,N_8793);
nand U9235 (N_9235,N_8829,N_8838);
xnor U9236 (N_9236,N_8818,N_8669);
nor U9237 (N_9237,N_8899,N_8965);
and U9238 (N_9238,N_8883,N_8464);
nand U9239 (N_9239,N_8939,N_8603);
or U9240 (N_9240,N_8541,N_8729);
nor U9241 (N_9241,N_8302,N_8706);
xor U9242 (N_9242,N_8378,N_8432);
and U9243 (N_9243,N_8696,N_8579);
xor U9244 (N_9244,N_8415,N_8327);
xnor U9245 (N_9245,N_8504,N_8540);
xnor U9246 (N_9246,N_8294,N_8700);
xor U9247 (N_9247,N_8919,N_8332);
nand U9248 (N_9248,N_8843,N_8485);
nor U9249 (N_9249,N_8783,N_8860);
or U9250 (N_9250,N_8869,N_8974);
or U9251 (N_9251,N_8946,N_8875);
nand U9252 (N_9252,N_8942,N_8274);
and U9253 (N_9253,N_8548,N_8726);
nor U9254 (N_9254,N_8534,N_8847);
xnor U9255 (N_9255,N_8910,N_8329);
nand U9256 (N_9256,N_8349,N_8717);
or U9257 (N_9257,N_8943,N_8587);
nor U9258 (N_9258,N_8446,N_8702);
and U9259 (N_9259,N_8816,N_8285);
nand U9260 (N_9260,N_8372,N_8914);
or U9261 (N_9261,N_8570,N_8851);
and U9262 (N_9262,N_8701,N_8467);
xor U9263 (N_9263,N_8760,N_8457);
nor U9264 (N_9264,N_8469,N_8259);
nand U9265 (N_9265,N_8537,N_8759);
and U9266 (N_9266,N_8305,N_8318);
or U9267 (N_9267,N_8528,N_8868);
nor U9268 (N_9268,N_8254,N_8300);
and U9269 (N_9269,N_8505,N_8998);
xnor U9270 (N_9270,N_8559,N_8453);
or U9271 (N_9271,N_8849,N_8933);
and U9272 (N_9272,N_8859,N_8813);
or U9273 (N_9273,N_8618,N_8490);
or U9274 (N_9274,N_8962,N_8597);
or U9275 (N_9275,N_8571,N_8799);
nor U9276 (N_9276,N_8506,N_8771);
and U9277 (N_9277,N_8609,N_8770);
nand U9278 (N_9278,N_8374,N_8877);
nand U9279 (N_9279,N_8725,N_8501);
or U9280 (N_9280,N_8921,N_8545);
nor U9281 (N_9281,N_8639,N_8301);
and U9282 (N_9282,N_8721,N_8495);
or U9283 (N_9283,N_8909,N_8398);
xor U9284 (N_9284,N_8478,N_8777);
nor U9285 (N_9285,N_8264,N_8328);
or U9286 (N_9286,N_8805,N_8277);
or U9287 (N_9287,N_8708,N_8898);
xnor U9288 (N_9288,N_8599,N_8323);
nand U9289 (N_9289,N_8499,N_8902);
and U9290 (N_9290,N_8891,N_8856);
nand U9291 (N_9291,N_8815,N_8386);
and U9292 (N_9292,N_8913,N_8321);
or U9293 (N_9293,N_8441,N_8996);
and U9294 (N_9294,N_8629,N_8749);
nor U9295 (N_9295,N_8958,N_8656);
and U9296 (N_9296,N_8458,N_8436);
nor U9297 (N_9297,N_8565,N_8553);
xor U9298 (N_9298,N_8617,N_8925);
and U9299 (N_9299,N_8796,N_8956);
nor U9300 (N_9300,N_8567,N_8812);
and U9301 (N_9301,N_8874,N_8929);
nand U9302 (N_9302,N_8802,N_8428);
nor U9303 (N_9303,N_8797,N_8563);
nand U9304 (N_9304,N_8667,N_8491);
xnor U9305 (N_9305,N_8908,N_8526);
nand U9306 (N_9306,N_8775,N_8840);
nor U9307 (N_9307,N_8752,N_8864);
and U9308 (N_9308,N_8642,N_8530);
nor U9309 (N_9309,N_8863,N_8628);
nor U9310 (N_9310,N_8271,N_8758);
nand U9311 (N_9311,N_8710,N_8676);
nor U9312 (N_9312,N_8657,N_8757);
nand U9313 (N_9313,N_8390,N_8661);
nand U9314 (N_9314,N_8695,N_8837);
nor U9315 (N_9315,N_8477,N_8362);
or U9316 (N_9316,N_8513,N_8878);
nor U9317 (N_9317,N_8284,N_8674);
or U9318 (N_9318,N_8966,N_8989);
or U9319 (N_9319,N_8393,N_8920);
or U9320 (N_9320,N_8880,N_8885);
nor U9321 (N_9321,N_8278,N_8763);
and U9322 (N_9322,N_8663,N_8964);
xor U9323 (N_9323,N_8862,N_8684);
and U9324 (N_9324,N_8740,N_8690);
and U9325 (N_9325,N_8990,N_8755);
nand U9326 (N_9326,N_8407,N_8595);
nand U9327 (N_9327,N_8379,N_8547);
xnor U9328 (N_9328,N_8411,N_8580);
and U9329 (N_9329,N_8685,N_8786);
or U9330 (N_9330,N_8312,N_8275);
nand U9331 (N_9331,N_8484,N_8945);
nand U9332 (N_9332,N_8834,N_8360);
xor U9333 (N_9333,N_8406,N_8986);
nand U9334 (N_9334,N_8935,N_8631);
and U9335 (N_9335,N_8449,N_8273);
and U9336 (N_9336,N_8341,N_8632);
and U9337 (N_9337,N_8257,N_8424);
or U9338 (N_9338,N_8359,N_8785);
and U9339 (N_9339,N_8568,N_8984);
or U9340 (N_9340,N_8662,N_8764);
nor U9341 (N_9341,N_8944,N_8422);
nor U9342 (N_9342,N_8421,N_8481);
nand U9343 (N_9343,N_8276,N_8350);
nor U9344 (N_9344,N_8623,N_8438);
or U9345 (N_9345,N_8995,N_8400);
or U9346 (N_9346,N_8715,N_8255);
nand U9347 (N_9347,N_8344,N_8739);
xnor U9348 (N_9348,N_8634,N_8551);
nor U9349 (N_9349,N_8650,N_8335);
nand U9350 (N_9350,N_8753,N_8654);
or U9351 (N_9351,N_8997,N_8605);
nand U9352 (N_9352,N_8270,N_8539);
nand U9353 (N_9353,N_8776,N_8581);
nor U9354 (N_9354,N_8375,N_8452);
nor U9355 (N_9355,N_8414,N_8645);
xor U9356 (N_9356,N_8978,N_8647);
xnor U9357 (N_9357,N_8304,N_8600);
and U9358 (N_9358,N_8420,N_8459);
xnor U9359 (N_9359,N_8893,N_8606);
and U9360 (N_9360,N_8340,N_8326);
and U9361 (N_9361,N_8613,N_8549);
xnor U9362 (N_9362,N_8773,N_8712);
xnor U9363 (N_9363,N_8310,N_8518);
and U9364 (N_9364,N_8738,N_8649);
nand U9365 (N_9365,N_8291,N_8434);
nand U9366 (N_9366,N_8719,N_8297);
or U9367 (N_9367,N_8718,N_8666);
or U9368 (N_9368,N_8867,N_8842);
and U9369 (N_9369,N_8482,N_8331);
xor U9370 (N_9370,N_8584,N_8969);
and U9371 (N_9371,N_8836,N_8444);
xnor U9372 (N_9372,N_8408,N_8881);
or U9373 (N_9373,N_8425,N_8361);
nand U9374 (N_9374,N_8699,N_8516);
or U9375 (N_9375,N_8298,N_8333);
and U9376 (N_9376,N_8755,N_8824);
nand U9377 (N_9377,N_8344,N_8734);
xor U9378 (N_9378,N_8331,N_8776);
and U9379 (N_9379,N_8545,N_8341);
xor U9380 (N_9380,N_8375,N_8457);
or U9381 (N_9381,N_8846,N_8374);
nor U9382 (N_9382,N_8887,N_8975);
or U9383 (N_9383,N_8826,N_8784);
nand U9384 (N_9384,N_8585,N_8793);
xnor U9385 (N_9385,N_8327,N_8450);
or U9386 (N_9386,N_8364,N_8680);
nand U9387 (N_9387,N_8950,N_8876);
and U9388 (N_9388,N_8886,N_8494);
or U9389 (N_9389,N_8964,N_8458);
or U9390 (N_9390,N_8761,N_8300);
xnor U9391 (N_9391,N_8532,N_8547);
and U9392 (N_9392,N_8283,N_8256);
and U9393 (N_9393,N_8558,N_8751);
or U9394 (N_9394,N_8468,N_8319);
xor U9395 (N_9395,N_8846,N_8336);
or U9396 (N_9396,N_8970,N_8649);
nor U9397 (N_9397,N_8580,N_8786);
nor U9398 (N_9398,N_8476,N_8467);
xor U9399 (N_9399,N_8671,N_8517);
or U9400 (N_9400,N_8391,N_8456);
nand U9401 (N_9401,N_8295,N_8431);
or U9402 (N_9402,N_8813,N_8321);
and U9403 (N_9403,N_8974,N_8814);
nor U9404 (N_9404,N_8896,N_8424);
xor U9405 (N_9405,N_8410,N_8914);
and U9406 (N_9406,N_8593,N_8951);
nor U9407 (N_9407,N_8592,N_8551);
or U9408 (N_9408,N_8525,N_8397);
nand U9409 (N_9409,N_8851,N_8555);
nand U9410 (N_9410,N_8923,N_8580);
nand U9411 (N_9411,N_8838,N_8503);
nand U9412 (N_9412,N_8467,N_8915);
nor U9413 (N_9413,N_8326,N_8632);
or U9414 (N_9414,N_8596,N_8714);
or U9415 (N_9415,N_8512,N_8430);
xor U9416 (N_9416,N_8644,N_8949);
nor U9417 (N_9417,N_8458,N_8685);
nand U9418 (N_9418,N_8440,N_8334);
xor U9419 (N_9419,N_8504,N_8622);
and U9420 (N_9420,N_8854,N_8495);
or U9421 (N_9421,N_8392,N_8840);
or U9422 (N_9422,N_8573,N_8991);
and U9423 (N_9423,N_8522,N_8709);
or U9424 (N_9424,N_8934,N_8957);
or U9425 (N_9425,N_8894,N_8716);
and U9426 (N_9426,N_8882,N_8646);
nand U9427 (N_9427,N_8488,N_8388);
or U9428 (N_9428,N_8653,N_8785);
nand U9429 (N_9429,N_8437,N_8723);
xnor U9430 (N_9430,N_8337,N_8718);
and U9431 (N_9431,N_8624,N_8671);
nand U9432 (N_9432,N_8358,N_8481);
nor U9433 (N_9433,N_8908,N_8701);
nand U9434 (N_9434,N_8342,N_8546);
nand U9435 (N_9435,N_8360,N_8784);
and U9436 (N_9436,N_8986,N_8271);
nor U9437 (N_9437,N_8923,N_8779);
nand U9438 (N_9438,N_8785,N_8784);
xnor U9439 (N_9439,N_8802,N_8553);
and U9440 (N_9440,N_8888,N_8609);
xnor U9441 (N_9441,N_8446,N_8609);
nand U9442 (N_9442,N_8576,N_8548);
nand U9443 (N_9443,N_8588,N_8554);
xnor U9444 (N_9444,N_8974,N_8413);
and U9445 (N_9445,N_8330,N_8258);
nor U9446 (N_9446,N_8525,N_8709);
and U9447 (N_9447,N_8517,N_8430);
and U9448 (N_9448,N_8633,N_8449);
and U9449 (N_9449,N_8278,N_8873);
or U9450 (N_9450,N_8280,N_8393);
nor U9451 (N_9451,N_8828,N_8398);
or U9452 (N_9452,N_8871,N_8527);
and U9453 (N_9453,N_8350,N_8498);
xor U9454 (N_9454,N_8555,N_8333);
nor U9455 (N_9455,N_8729,N_8673);
or U9456 (N_9456,N_8438,N_8906);
nor U9457 (N_9457,N_8913,N_8710);
xor U9458 (N_9458,N_8475,N_8519);
xnor U9459 (N_9459,N_8300,N_8797);
xnor U9460 (N_9460,N_8809,N_8658);
nor U9461 (N_9461,N_8395,N_8802);
nor U9462 (N_9462,N_8487,N_8330);
or U9463 (N_9463,N_8946,N_8255);
nor U9464 (N_9464,N_8646,N_8462);
nand U9465 (N_9465,N_8665,N_8703);
nand U9466 (N_9466,N_8760,N_8260);
nand U9467 (N_9467,N_8251,N_8381);
and U9468 (N_9468,N_8739,N_8336);
nor U9469 (N_9469,N_8638,N_8634);
nor U9470 (N_9470,N_8990,N_8758);
nand U9471 (N_9471,N_8428,N_8920);
or U9472 (N_9472,N_8549,N_8985);
and U9473 (N_9473,N_8852,N_8832);
nand U9474 (N_9474,N_8985,N_8271);
xnor U9475 (N_9475,N_8837,N_8653);
xnor U9476 (N_9476,N_8389,N_8917);
and U9477 (N_9477,N_8955,N_8741);
xnor U9478 (N_9478,N_8766,N_8988);
xnor U9479 (N_9479,N_8844,N_8451);
nand U9480 (N_9480,N_8854,N_8520);
and U9481 (N_9481,N_8882,N_8617);
and U9482 (N_9482,N_8803,N_8741);
xnor U9483 (N_9483,N_8867,N_8632);
nor U9484 (N_9484,N_8849,N_8344);
nand U9485 (N_9485,N_8874,N_8812);
or U9486 (N_9486,N_8278,N_8495);
xnor U9487 (N_9487,N_8386,N_8943);
xor U9488 (N_9488,N_8751,N_8927);
nor U9489 (N_9489,N_8467,N_8755);
xor U9490 (N_9490,N_8560,N_8961);
or U9491 (N_9491,N_8719,N_8943);
or U9492 (N_9492,N_8503,N_8528);
or U9493 (N_9493,N_8641,N_8766);
nand U9494 (N_9494,N_8935,N_8975);
nand U9495 (N_9495,N_8278,N_8877);
nor U9496 (N_9496,N_8715,N_8644);
nand U9497 (N_9497,N_8944,N_8459);
and U9498 (N_9498,N_8820,N_8892);
or U9499 (N_9499,N_8412,N_8433);
xor U9500 (N_9500,N_8719,N_8784);
nand U9501 (N_9501,N_8496,N_8368);
xor U9502 (N_9502,N_8608,N_8252);
xnor U9503 (N_9503,N_8584,N_8929);
nor U9504 (N_9504,N_8507,N_8713);
nand U9505 (N_9505,N_8689,N_8546);
or U9506 (N_9506,N_8582,N_8977);
xnor U9507 (N_9507,N_8386,N_8276);
xnor U9508 (N_9508,N_8278,N_8795);
nor U9509 (N_9509,N_8594,N_8292);
and U9510 (N_9510,N_8788,N_8420);
and U9511 (N_9511,N_8476,N_8386);
xnor U9512 (N_9512,N_8937,N_8547);
and U9513 (N_9513,N_8326,N_8618);
xor U9514 (N_9514,N_8701,N_8706);
nor U9515 (N_9515,N_8490,N_8648);
or U9516 (N_9516,N_8910,N_8490);
or U9517 (N_9517,N_8366,N_8955);
xnor U9518 (N_9518,N_8851,N_8930);
or U9519 (N_9519,N_8964,N_8919);
and U9520 (N_9520,N_8412,N_8341);
nor U9521 (N_9521,N_8420,N_8769);
and U9522 (N_9522,N_8390,N_8727);
or U9523 (N_9523,N_8632,N_8840);
xor U9524 (N_9524,N_8437,N_8778);
nand U9525 (N_9525,N_8702,N_8721);
nor U9526 (N_9526,N_8981,N_8969);
nand U9527 (N_9527,N_8717,N_8670);
xnor U9528 (N_9528,N_8444,N_8902);
and U9529 (N_9529,N_8436,N_8979);
nand U9530 (N_9530,N_8560,N_8693);
xnor U9531 (N_9531,N_8790,N_8914);
nand U9532 (N_9532,N_8898,N_8368);
xor U9533 (N_9533,N_8552,N_8603);
or U9534 (N_9534,N_8674,N_8542);
xor U9535 (N_9535,N_8442,N_8401);
nor U9536 (N_9536,N_8932,N_8601);
and U9537 (N_9537,N_8776,N_8436);
or U9538 (N_9538,N_8291,N_8991);
xnor U9539 (N_9539,N_8269,N_8842);
nand U9540 (N_9540,N_8353,N_8697);
nand U9541 (N_9541,N_8411,N_8524);
xor U9542 (N_9542,N_8798,N_8559);
nand U9543 (N_9543,N_8267,N_8882);
nand U9544 (N_9544,N_8958,N_8716);
xor U9545 (N_9545,N_8692,N_8909);
nor U9546 (N_9546,N_8298,N_8671);
nand U9547 (N_9547,N_8862,N_8568);
xnor U9548 (N_9548,N_8343,N_8607);
or U9549 (N_9549,N_8684,N_8886);
nor U9550 (N_9550,N_8676,N_8975);
or U9551 (N_9551,N_8491,N_8664);
and U9552 (N_9552,N_8268,N_8471);
or U9553 (N_9553,N_8416,N_8567);
or U9554 (N_9554,N_8887,N_8587);
or U9555 (N_9555,N_8802,N_8290);
nor U9556 (N_9556,N_8628,N_8531);
and U9557 (N_9557,N_8588,N_8463);
and U9558 (N_9558,N_8430,N_8504);
or U9559 (N_9559,N_8674,N_8920);
xor U9560 (N_9560,N_8436,N_8919);
nor U9561 (N_9561,N_8684,N_8873);
xnor U9562 (N_9562,N_8360,N_8622);
nand U9563 (N_9563,N_8339,N_8572);
or U9564 (N_9564,N_8803,N_8975);
or U9565 (N_9565,N_8366,N_8800);
or U9566 (N_9566,N_8477,N_8301);
xor U9567 (N_9567,N_8777,N_8421);
xor U9568 (N_9568,N_8255,N_8672);
or U9569 (N_9569,N_8727,N_8558);
nor U9570 (N_9570,N_8973,N_8912);
xnor U9571 (N_9571,N_8796,N_8743);
and U9572 (N_9572,N_8570,N_8544);
xor U9573 (N_9573,N_8268,N_8408);
nor U9574 (N_9574,N_8390,N_8376);
nor U9575 (N_9575,N_8722,N_8584);
or U9576 (N_9576,N_8273,N_8690);
or U9577 (N_9577,N_8512,N_8403);
nor U9578 (N_9578,N_8552,N_8451);
nor U9579 (N_9579,N_8649,N_8252);
nand U9580 (N_9580,N_8414,N_8660);
nor U9581 (N_9581,N_8793,N_8410);
and U9582 (N_9582,N_8642,N_8753);
or U9583 (N_9583,N_8930,N_8605);
and U9584 (N_9584,N_8799,N_8365);
nand U9585 (N_9585,N_8495,N_8891);
and U9586 (N_9586,N_8722,N_8924);
and U9587 (N_9587,N_8356,N_8980);
nand U9588 (N_9588,N_8668,N_8455);
and U9589 (N_9589,N_8938,N_8369);
nor U9590 (N_9590,N_8369,N_8446);
nand U9591 (N_9591,N_8962,N_8584);
nor U9592 (N_9592,N_8491,N_8943);
nor U9593 (N_9593,N_8674,N_8724);
nand U9594 (N_9594,N_8409,N_8854);
nand U9595 (N_9595,N_8417,N_8843);
or U9596 (N_9596,N_8525,N_8568);
nor U9597 (N_9597,N_8535,N_8265);
and U9598 (N_9598,N_8720,N_8747);
and U9599 (N_9599,N_8580,N_8911);
xnor U9600 (N_9600,N_8535,N_8459);
nor U9601 (N_9601,N_8648,N_8843);
or U9602 (N_9602,N_8326,N_8522);
nand U9603 (N_9603,N_8912,N_8637);
and U9604 (N_9604,N_8857,N_8782);
nor U9605 (N_9605,N_8632,N_8580);
nand U9606 (N_9606,N_8748,N_8949);
nor U9607 (N_9607,N_8539,N_8784);
xnor U9608 (N_9608,N_8993,N_8454);
nand U9609 (N_9609,N_8625,N_8485);
or U9610 (N_9610,N_8769,N_8622);
xnor U9611 (N_9611,N_8549,N_8744);
nor U9612 (N_9612,N_8716,N_8402);
xor U9613 (N_9613,N_8919,N_8834);
xor U9614 (N_9614,N_8364,N_8602);
xor U9615 (N_9615,N_8877,N_8862);
or U9616 (N_9616,N_8968,N_8701);
or U9617 (N_9617,N_8509,N_8567);
nor U9618 (N_9618,N_8262,N_8833);
or U9619 (N_9619,N_8684,N_8440);
xor U9620 (N_9620,N_8347,N_8411);
or U9621 (N_9621,N_8878,N_8778);
and U9622 (N_9622,N_8668,N_8446);
nor U9623 (N_9623,N_8453,N_8936);
xor U9624 (N_9624,N_8595,N_8417);
nor U9625 (N_9625,N_8253,N_8953);
nor U9626 (N_9626,N_8471,N_8983);
and U9627 (N_9627,N_8899,N_8947);
xnor U9628 (N_9628,N_8716,N_8979);
or U9629 (N_9629,N_8854,N_8719);
xnor U9630 (N_9630,N_8660,N_8574);
xor U9631 (N_9631,N_8638,N_8678);
xnor U9632 (N_9632,N_8547,N_8858);
nor U9633 (N_9633,N_8492,N_8846);
nor U9634 (N_9634,N_8788,N_8510);
or U9635 (N_9635,N_8796,N_8327);
nand U9636 (N_9636,N_8467,N_8493);
nor U9637 (N_9637,N_8717,N_8820);
xnor U9638 (N_9638,N_8666,N_8739);
nor U9639 (N_9639,N_8785,N_8689);
and U9640 (N_9640,N_8534,N_8356);
and U9641 (N_9641,N_8267,N_8948);
xor U9642 (N_9642,N_8598,N_8949);
or U9643 (N_9643,N_8639,N_8946);
xnor U9644 (N_9644,N_8336,N_8661);
and U9645 (N_9645,N_8280,N_8864);
xor U9646 (N_9646,N_8444,N_8856);
or U9647 (N_9647,N_8784,N_8289);
or U9648 (N_9648,N_8688,N_8883);
or U9649 (N_9649,N_8435,N_8955);
nand U9650 (N_9650,N_8745,N_8814);
xor U9651 (N_9651,N_8507,N_8328);
nand U9652 (N_9652,N_8699,N_8309);
and U9653 (N_9653,N_8509,N_8873);
nand U9654 (N_9654,N_8926,N_8961);
and U9655 (N_9655,N_8724,N_8737);
nand U9656 (N_9656,N_8383,N_8766);
and U9657 (N_9657,N_8690,N_8374);
xor U9658 (N_9658,N_8505,N_8859);
nand U9659 (N_9659,N_8790,N_8370);
nand U9660 (N_9660,N_8679,N_8633);
or U9661 (N_9661,N_8325,N_8693);
and U9662 (N_9662,N_8551,N_8271);
or U9663 (N_9663,N_8751,N_8886);
nand U9664 (N_9664,N_8687,N_8799);
nor U9665 (N_9665,N_8767,N_8755);
xor U9666 (N_9666,N_8492,N_8382);
xor U9667 (N_9667,N_8681,N_8409);
and U9668 (N_9668,N_8294,N_8506);
nand U9669 (N_9669,N_8602,N_8550);
or U9670 (N_9670,N_8716,N_8882);
nor U9671 (N_9671,N_8685,N_8582);
xnor U9672 (N_9672,N_8338,N_8360);
and U9673 (N_9673,N_8705,N_8410);
nor U9674 (N_9674,N_8460,N_8522);
nor U9675 (N_9675,N_8877,N_8976);
or U9676 (N_9676,N_8688,N_8845);
and U9677 (N_9677,N_8546,N_8616);
nand U9678 (N_9678,N_8440,N_8450);
nor U9679 (N_9679,N_8528,N_8740);
xnor U9680 (N_9680,N_8393,N_8370);
nor U9681 (N_9681,N_8522,N_8520);
xnor U9682 (N_9682,N_8956,N_8268);
and U9683 (N_9683,N_8871,N_8316);
or U9684 (N_9684,N_8269,N_8918);
or U9685 (N_9685,N_8406,N_8771);
or U9686 (N_9686,N_8532,N_8731);
and U9687 (N_9687,N_8876,N_8722);
and U9688 (N_9688,N_8498,N_8310);
or U9689 (N_9689,N_8440,N_8904);
xor U9690 (N_9690,N_8720,N_8712);
nor U9691 (N_9691,N_8654,N_8468);
nand U9692 (N_9692,N_8619,N_8590);
or U9693 (N_9693,N_8769,N_8491);
and U9694 (N_9694,N_8573,N_8796);
nor U9695 (N_9695,N_8618,N_8610);
xnor U9696 (N_9696,N_8628,N_8416);
or U9697 (N_9697,N_8634,N_8421);
nand U9698 (N_9698,N_8579,N_8733);
and U9699 (N_9699,N_8339,N_8346);
and U9700 (N_9700,N_8745,N_8860);
nor U9701 (N_9701,N_8926,N_8291);
nand U9702 (N_9702,N_8403,N_8556);
or U9703 (N_9703,N_8449,N_8702);
nor U9704 (N_9704,N_8552,N_8806);
xor U9705 (N_9705,N_8288,N_8555);
nor U9706 (N_9706,N_8628,N_8849);
or U9707 (N_9707,N_8956,N_8314);
or U9708 (N_9708,N_8431,N_8827);
nand U9709 (N_9709,N_8664,N_8496);
or U9710 (N_9710,N_8635,N_8640);
or U9711 (N_9711,N_8966,N_8819);
or U9712 (N_9712,N_8653,N_8595);
nor U9713 (N_9713,N_8931,N_8629);
xor U9714 (N_9714,N_8710,N_8780);
xor U9715 (N_9715,N_8339,N_8333);
xnor U9716 (N_9716,N_8440,N_8323);
xor U9717 (N_9717,N_8855,N_8451);
and U9718 (N_9718,N_8895,N_8763);
and U9719 (N_9719,N_8477,N_8268);
xor U9720 (N_9720,N_8772,N_8902);
nand U9721 (N_9721,N_8698,N_8672);
nand U9722 (N_9722,N_8653,N_8322);
or U9723 (N_9723,N_8533,N_8268);
and U9724 (N_9724,N_8521,N_8736);
nor U9725 (N_9725,N_8912,N_8250);
nand U9726 (N_9726,N_8965,N_8840);
or U9727 (N_9727,N_8442,N_8934);
and U9728 (N_9728,N_8464,N_8988);
nor U9729 (N_9729,N_8594,N_8442);
nand U9730 (N_9730,N_8818,N_8881);
nor U9731 (N_9731,N_8613,N_8401);
nor U9732 (N_9732,N_8482,N_8511);
xor U9733 (N_9733,N_8780,N_8784);
nand U9734 (N_9734,N_8799,N_8363);
nor U9735 (N_9735,N_8852,N_8772);
nor U9736 (N_9736,N_8562,N_8422);
nand U9737 (N_9737,N_8799,N_8372);
nor U9738 (N_9738,N_8483,N_8266);
nand U9739 (N_9739,N_8636,N_8392);
nand U9740 (N_9740,N_8293,N_8629);
nor U9741 (N_9741,N_8713,N_8561);
xor U9742 (N_9742,N_8590,N_8758);
nor U9743 (N_9743,N_8709,N_8981);
xor U9744 (N_9744,N_8688,N_8600);
and U9745 (N_9745,N_8755,N_8570);
and U9746 (N_9746,N_8782,N_8361);
nand U9747 (N_9747,N_8457,N_8627);
nor U9748 (N_9748,N_8698,N_8762);
or U9749 (N_9749,N_8768,N_8775);
nor U9750 (N_9750,N_9532,N_9159);
nand U9751 (N_9751,N_9102,N_9723);
or U9752 (N_9752,N_9058,N_9016);
xor U9753 (N_9753,N_9247,N_9418);
nand U9754 (N_9754,N_9089,N_9316);
and U9755 (N_9755,N_9365,N_9455);
and U9756 (N_9756,N_9632,N_9651);
and U9757 (N_9757,N_9174,N_9691);
and U9758 (N_9758,N_9330,N_9127);
or U9759 (N_9759,N_9409,N_9588);
nor U9760 (N_9760,N_9508,N_9457);
or U9761 (N_9761,N_9347,N_9630);
nor U9762 (N_9762,N_9494,N_9150);
nor U9763 (N_9763,N_9042,N_9272);
and U9764 (N_9764,N_9211,N_9143);
and U9765 (N_9765,N_9487,N_9614);
nand U9766 (N_9766,N_9379,N_9022);
or U9767 (N_9767,N_9542,N_9729);
xor U9768 (N_9768,N_9038,N_9524);
nor U9769 (N_9769,N_9196,N_9587);
and U9770 (N_9770,N_9141,N_9543);
nand U9771 (N_9771,N_9334,N_9177);
and U9772 (N_9772,N_9721,N_9615);
or U9773 (N_9773,N_9315,N_9286);
nor U9774 (N_9774,N_9660,N_9373);
nor U9775 (N_9775,N_9342,N_9185);
or U9776 (N_9776,N_9064,N_9546);
nor U9777 (N_9777,N_9206,N_9402);
nor U9778 (N_9778,N_9311,N_9000);
and U9779 (N_9779,N_9426,N_9120);
xnor U9780 (N_9780,N_9167,N_9152);
or U9781 (N_9781,N_9259,N_9564);
nor U9782 (N_9782,N_9221,N_9730);
and U9783 (N_9783,N_9212,N_9095);
and U9784 (N_9784,N_9656,N_9571);
xnor U9785 (N_9785,N_9121,N_9345);
and U9786 (N_9786,N_9434,N_9018);
or U9787 (N_9787,N_9733,N_9085);
xor U9788 (N_9788,N_9153,N_9555);
and U9789 (N_9789,N_9623,N_9386);
or U9790 (N_9790,N_9551,N_9190);
nand U9791 (N_9791,N_9662,N_9428);
nand U9792 (N_9792,N_9617,N_9215);
nor U9793 (N_9793,N_9590,N_9126);
xnor U9794 (N_9794,N_9154,N_9696);
nor U9795 (N_9795,N_9222,N_9682);
xnor U9796 (N_9796,N_9366,N_9318);
or U9797 (N_9797,N_9357,N_9319);
xor U9798 (N_9798,N_9395,N_9351);
or U9799 (N_9799,N_9341,N_9383);
nor U9800 (N_9800,N_9541,N_9568);
nor U9801 (N_9801,N_9622,N_9589);
xnor U9802 (N_9802,N_9640,N_9059);
or U9803 (N_9803,N_9021,N_9111);
nor U9804 (N_9804,N_9382,N_9145);
or U9805 (N_9805,N_9529,N_9056);
and U9806 (N_9806,N_9332,N_9453);
or U9807 (N_9807,N_9037,N_9236);
nand U9808 (N_9808,N_9425,N_9181);
or U9809 (N_9809,N_9531,N_9253);
nor U9810 (N_9810,N_9399,N_9192);
nor U9811 (N_9811,N_9636,N_9336);
or U9812 (N_9812,N_9262,N_9309);
nand U9813 (N_9813,N_9256,N_9470);
and U9814 (N_9814,N_9371,N_9681);
or U9815 (N_9815,N_9579,N_9234);
xnor U9816 (N_9816,N_9337,N_9398);
nor U9817 (N_9817,N_9155,N_9563);
xnor U9818 (N_9818,N_9747,N_9575);
and U9819 (N_9819,N_9308,N_9360);
or U9820 (N_9820,N_9675,N_9420);
or U9821 (N_9821,N_9702,N_9739);
xor U9822 (N_9822,N_9294,N_9549);
or U9823 (N_9823,N_9157,N_9556);
nor U9824 (N_9824,N_9736,N_9732);
or U9825 (N_9825,N_9668,N_9118);
nand U9826 (N_9826,N_9582,N_9025);
xnor U9827 (N_9827,N_9458,N_9176);
nand U9828 (N_9828,N_9014,N_9197);
and U9829 (N_9829,N_9325,N_9381);
nand U9830 (N_9830,N_9741,N_9481);
nand U9831 (N_9831,N_9217,N_9209);
nor U9832 (N_9832,N_9602,N_9231);
nor U9833 (N_9833,N_9686,N_9519);
nor U9834 (N_9834,N_9712,N_9094);
nand U9835 (N_9835,N_9082,N_9639);
nand U9836 (N_9836,N_9628,N_9725);
or U9837 (N_9837,N_9214,N_9722);
nand U9838 (N_9838,N_9535,N_9044);
xor U9839 (N_9839,N_9719,N_9260);
xnor U9840 (N_9840,N_9727,N_9296);
or U9841 (N_9841,N_9377,N_9201);
xnor U9842 (N_9842,N_9241,N_9497);
nor U9843 (N_9843,N_9720,N_9665);
nand U9844 (N_9844,N_9269,N_9258);
and U9845 (N_9845,N_9243,N_9103);
nor U9846 (N_9846,N_9117,N_9306);
and U9847 (N_9847,N_9005,N_9276);
and U9848 (N_9848,N_9084,N_9271);
nor U9849 (N_9849,N_9653,N_9267);
xnor U9850 (N_9850,N_9580,N_9449);
and U9851 (N_9851,N_9637,N_9616);
nand U9852 (N_9852,N_9384,N_9548);
and U9853 (N_9853,N_9061,N_9188);
and U9854 (N_9854,N_9518,N_9277);
and U9855 (N_9855,N_9027,N_9048);
nand U9856 (N_9856,N_9068,N_9255);
xnor U9857 (N_9857,N_9677,N_9525);
xor U9858 (N_9858,N_9700,N_9592);
nand U9859 (N_9859,N_9020,N_9164);
nand U9860 (N_9860,N_9456,N_9716);
or U9861 (N_9861,N_9029,N_9685);
xor U9862 (N_9862,N_9179,N_9421);
xnor U9863 (N_9863,N_9718,N_9092);
xor U9864 (N_9864,N_9075,N_9431);
and U9865 (N_9865,N_9045,N_9060);
or U9866 (N_9866,N_9292,N_9112);
xnor U9867 (N_9867,N_9125,N_9432);
xnor U9868 (N_9868,N_9631,N_9607);
or U9869 (N_9869,N_9430,N_9172);
nand U9870 (N_9870,N_9328,N_9046);
nand U9871 (N_9871,N_9080,N_9654);
nor U9872 (N_9872,N_9410,N_9105);
nor U9873 (N_9873,N_9039,N_9119);
nor U9874 (N_9874,N_9239,N_9063);
nand U9875 (N_9875,N_9626,N_9444);
nand U9876 (N_9876,N_9363,N_9545);
and U9877 (N_9877,N_9687,N_9326);
or U9878 (N_9878,N_9405,N_9619);
nor U9879 (N_9879,N_9570,N_9202);
xor U9880 (N_9880,N_9069,N_9087);
xor U9881 (N_9881,N_9144,N_9472);
xor U9882 (N_9882,N_9643,N_9099);
nand U9883 (N_9883,N_9704,N_9109);
and U9884 (N_9884,N_9408,N_9690);
or U9885 (N_9885,N_9055,N_9062);
and U9886 (N_9886,N_9140,N_9376);
or U9887 (N_9887,N_9728,N_9744);
nor U9888 (N_9888,N_9367,N_9265);
or U9889 (N_9889,N_9633,N_9354);
and U9890 (N_9890,N_9527,N_9439);
xor U9891 (N_9891,N_9635,N_9599);
nor U9892 (N_9892,N_9344,N_9358);
nand U9893 (N_9893,N_9163,N_9011);
nor U9894 (N_9894,N_9715,N_9275);
or U9895 (N_9895,N_9013,N_9473);
nor U9896 (N_9896,N_9469,N_9650);
and U9897 (N_9897,N_9618,N_9544);
nor U9898 (N_9898,N_9624,N_9684);
or U9899 (N_9899,N_9506,N_9605);
and U9900 (N_9900,N_9339,N_9520);
nand U9901 (N_9901,N_9165,N_9248);
or U9902 (N_9902,N_9178,N_9244);
and U9903 (N_9903,N_9693,N_9323);
and U9904 (N_9904,N_9407,N_9225);
nand U9905 (N_9905,N_9284,N_9368);
or U9906 (N_9906,N_9051,N_9268);
nand U9907 (N_9907,N_9394,N_9695);
or U9908 (N_9908,N_9437,N_9249);
or U9909 (N_9909,N_9310,N_9133);
nand U9910 (N_9910,N_9151,N_9043);
and U9911 (N_9911,N_9200,N_9370);
xor U9912 (N_9912,N_9134,N_9303);
and U9913 (N_9913,N_9385,N_9440);
nor U9914 (N_9914,N_9499,N_9521);
nand U9915 (N_9915,N_9387,N_9419);
nor U9916 (N_9916,N_9738,N_9740);
nand U9917 (N_9917,N_9040,N_9565);
and U9918 (N_9918,N_9187,N_9389);
nand U9919 (N_9919,N_9475,N_9698);
or U9920 (N_9920,N_9466,N_9227);
nand U9921 (N_9921,N_9608,N_9638);
or U9922 (N_9922,N_9581,N_9516);
or U9923 (N_9923,N_9658,N_9547);
and U9924 (N_9924,N_9246,N_9742);
and U9925 (N_9925,N_9476,N_9274);
nand U9926 (N_9926,N_9572,N_9707);
nor U9927 (N_9927,N_9604,N_9024);
nand U9928 (N_9928,N_9297,N_9735);
nor U9929 (N_9929,N_9203,N_9372);
xor U9930 (N_9930,N_9071,N_9380);
xnor U9931 (N_9931,N_9350,N_9603);
or U9932 (N_9932,N_9673,N_9442);
xor U9933 (N_9933,N_9083,N_9184);
or U9934 (N_9934,N_9158,N_9004);
xor U9935 (N_9935,N_9705,N_9595);
nand U9936 (N_9936,N_9574,N_9355);
nand U9937 (N_9937,N_9500,N_9391);
and U9938 (N_9938,N_9173,N_9593);
nand U9939 (N_9939,N_9321,N_9406);
nor U9940 (N_9940,N_9417,N_9034);
xor U9941 (N_9941,N_9359,N_9454);
and U9942 (N_9942,N_9411,N_9671);
and U9943 (N_9943,N_9030,N_9288);
nand U9944 (N_9944,N_9135,N_9436);
nor U9945 (N_9945,N_9403,N_9511);
xor U9946 (N_9946,N_9509,N_9186);
and U9947 (N_9947,N_9213,N_9647);
and U9948 (N_9948,N_9642,N_9329);
and U9949 (N_9949,N_9289,N_9017);
nor U9950 (N_9950,N_9412,N_9077);
nor U9951 (N_9951,N_9333,N_9703);
xnor U9952 (N_9952,N_9540,N_9210);
or U9953 (N_9953,N_9191,N_9467);
or U9954 (N_9954,N_9287,N_9193);
nor U9955 (N_9955,N_9375,N_9072);
and U9956 (N_9956,N_9734,N_9007);
and U9957 (N_9957,N_9218,N_9404);
xnor U9958 (N_9958,N_9232,N_9010);
or U9959 (N_9959,N_9086,N_9460);
and U9960 (N_9960,N_9422,N_9317);
and U9961 (N_9961,N_9504,N_9313);
or U9962 (N_9962,N_9251,N_9298);
and U9963 (N_9963,N_9331,N_9114);
nand U9964 (N_9964,N_9629,N_9340);
xnor U9965 (N_9965,N_9204,N_9220);
nor U9966 (N_9966,N_9674,N_9012);
nor U9967 (N_9967,N_9512,N_9362);
nor U9968 (N_9968,N_9139,N_9346);
xor U9969 (N_9969,N_9584,N_9283);
and U9970 (N_9970,N_9503,N_9250);
xnor U9971 (N_9971,N_9001,N_9464);
nand U9972 (N_9972,N_9076,N_9352);
nor U9973 (N_9973,N_9433,N_9672);
and U9974 (N_9974,N_9560,N_9388);
nand U9975 (N_9975,N_9706,N_9445);
xnor U9976 (N_9976,N_9280,N_9136);
nand U9977 (N_9977,N_9229,N_9390);
xor U9978 (N_9978,N_9353,N_9414);
or U9979 (N_9979,N_9237,N_9663);
or U9980 (N_9980,N_9281,N_9567);
or U9981 (N_9981,N_9447,N_9216);
nor U9982 (N_9982,N_9116,N_9067);
or U9983 (N_9983,N_9528,N_9462);
nand U9984 (N_9984,N_9392,N_9160);
nand U9985 (N_9985,N_9393,N_9659);
or U9986 (N_9986,N_9149,N_9429);
or U9987 (N_9987,N_9664,N_9356);
or U9988 (N_9988,N_9463,N_9110);
nand U9989 (N_9989,N_9226,N_9378);
nand U9990 (N_9990,N_9245,N_9031);
or U9991 (N_9991,N_9609,N_9261);
nor U9992 (N_9992,N_9423,N_9486);
xor U9993 (N_9993,N_9492,N_9523);
nand U9994 (N_9994,N_9238,N_9746);
nand U9995 (N_9995,N_9290,N_9307);
xor U9996 (N_9996,N_9070,N_9537);
xor U9997 (N_9997,N_9557,N_9198);
nand U9998 (N_9998,N_9015,N_9745);
and U9999 (N_9999,N_9107,N_9676);
nor U10000 (N_10000,N_9416,N_9634);
nand U10001 (N_10001,N_9611,N_9219);
xor U10002 (N_10002,N_9270,N_9097);
or U10003 (N_10003,N_9396,N_9263);
and U10004 (N_10004,N_9559,N_9468);
nand U10005 (N_10005,N_9301,N_9279);
nand U10006 (N_10006,N_9074,N_9726);
nor U10007 (N_10007,N_9438,N_9285);
and U10008 (N_10008,N_9131,N_9023);
nand U10009 (N_10009,N_9090,N_9471);
or U10010 (N_10010,N_9312,N_9553);
nand U10011 (N_10011,N_9566,N_9724);
xnor U10012 (N_10012,N_9036,N_9533);
xnor U10013 (N_10013,N_9562,N_9148);
and U10014 (N_10014,N_9098,N_9495);
or U10015 (N_10015,N_9714,N_9088);
nor U10016 (N_10016,N_9169,N_9006);
and U10017 (N_10017,N_9295,N_9578);
xnor U10018 (N_10018,N_9465,N_9199);
nand U10019 (N_10019,N_9709,N_9057);
xnor U10020 (N_10020,N_9490,N_9510);
nand U10021 (N_10021,N_9079,N_9073);
xor U10022 (N_10022,N_9670,N_9669);
nor U10023 (N_10023,N_9485,N_9147);
nor U10024 (N_10024,N_9601,N_9450);
xor U10025 (N_10025,N_9257,N_9701);
nand U10026 (N_10026,N_9240,N_9101);
xnor U10027 (N_10027,N_9343,N_9517);
or U10028 (N_10028,N_9302,N_9620);
and U10029 (N_10029,N_9327,N_9550);
or U10030 (N_10030,N_9266,N_9539);
nor U10031 (N_10031,N_9349,N_9482);
or U10032 (N_10032,N_9171,N_9597);
nand U10033 (N_10033,N_9132,N_9708);
and U10034 (N_10034,N_9513,N_9596);
or U10035 (N_10035,N_9166,N_9451);
nand U10036 (N_10036,N_9019,N_9606);
or U10037 (N_10037,N_9003,N_9106);
nand U10038 (N_10038,N_9711,N_9026);
nor U10039 (N_10039,N_9522,N_9415);
nor U10040 (N_10040,N_9583,N_9273);
xnor U10041 (N_10041,N_9452,N_9731);
and U10042 (N_10042,N_9032,N_9479);
and U10043 (N_10043,N_9401,N_9293);
xnor U10044 (N_10044,N_9304,N_9554);
and U10045 (N_10045,N_9613,N_9480);
nor U10046 (N_10046,N_9113,N_9666);
and U10047 (N_10047,N_9137,N_9223);
nand U10048 (N_10048,N_9054,N_9282);
nand U10049 (N_10049,N_9096,N_9502);
nand U10050 (N_10050,N_9493,N_9322);
nor U10051 (N_10051,N_9124,N_9577);
and U10052 (N_10052,N_9717,N_9129);
or U10053 (N_10053,N_9644,N_9498);
and U10054 (N_10054,N_9461,N_9641);
nand U10055 (N_10055,N_9252,N_9175);
or U10056 (N_10056,N_9530,N_9162);
and U10057 (N_10057,N_9514,N_9364);
nand U10058 (N_10058,N_9443,N_9002);
or U10059 (N_10059,N_9678,N_9627);
xor U10060 (N_10060,N_9008,N_9123);
nor U10061 (N_10061,N_9081,N_9091);
and U10062 (N_10062,N_9320,N_9335);
and U10063 (N_10063,N_9361,N_9491);
nand U10064 (N_10064,N_9652,N_9488);
and U10065 (N_10065,N_9183,N_9348);
and U10066 (N_10066,N_9424,N_9299);
nand U10067 (N_10067,N_9400,N_9576);
nor U10068 (N_10068,N_9625,N_9585);
nor U10069 (N_10069,N_9066,N_9697);
or U10070 (N_10070,N_9446,N_9168);
nand U10071 (N_10071,N_9427,N_9305);
xnor U10072 (N_10072,N_9489,N_9561);
xor U10073 (N_10073,N_9435,N_9536);
or U10074 (N_10074,N_9600,N_9009);
and U10075 (N_10075,N_9254,N_9594);
xnor U10076 (N_10076,N_9680,N_9041);
xnor U10077 (N_10077,N_9161,N_9093);
or U10078 (N_10078,N_9689,N_9646);
or U10079 (N_10079,N_9737,N_9078);
nor U10080 (N_10080,N_9208,N_9477);
nand U10081 (N_10081,N_9156,N_9526);
and U10082 (N_10082,N_9291,N_9338);
nand U10083 (N_10083,N_9028,N_9748);
nand U10084 (N_10084,N_9235,N_9515);
nor U10085 (N_10085,N_9047,N_9122);
nor U10086 (N_10086,N_9692,N_9586);
nor U10087 (N_10087,N_9128,N_9374);
nor U10088 (N_10088,N_9448,N_9195);
or U10089 (N_10089,N_9033,N_9035);
xor U10090 (N_10090,N_9694,N_9052);
nor U10091 (N_10091,N_9242,N_9710);
xnor U10092 (N_10092,N_9507,N_9228);
or U10093 (N_10093,N_9648,N_9534);
nor U10094 (N_10094,N_9170,N_9699);
xor U10095 (N_10095,N_9612,N_9324);
xnor U10096 (N_10096,N_9189,N_9538);
and U10097 (N_10097,N_9050,N_9104);
and U10098 (N_10098,N_9552,N_9108);
and U10099 (N_10099,N_9369,N_9474);
and U10100 (N_10100,N_9621,N_9496);
nor U10101 (N_10101,N_9713,N_9314);
and U10102 (N_10102,N_9478,N_9130);
or U10103 (N_10103,N_9207,N_9138);
or U10104 (N_10104,N_9413,N_9441);
nand U10105 (N_10105,N_9459,N_9610);
and U10106 (N_10106,N_9142,N_9278);
xnor U10107 (N_10107,N_9053,N_9655);
or U10108 (N_10108,N_9146,N_9749);
and U10109 (N_10109,N_9591,N_9224);
xor U10110 (N_10110,N_9688,N_9501);
or U10111 (N_10111,N_9679,N_9115);
nand U10112 (N_10112,N_9649,N_9049);
nor U10113 (N_10113,N_9194,N_9065);
nand U10114 (N_10114,N_9661,N_9645);
nor U10115 (N_10115,N_9233,N_9397);
or U10116 (N_10116,N_9743,N_9598);
and U10117 (N_10117,N_9573,N_9484);
and U10118 (N_10118,N_9683,N_9667);
or U10119 (N_10119,N_9483,N_9569);
or U10120 (N_10120,N_9264,N_9505);
xnor U10121 (N_10121,N_9657,N_9300);
xor U10122 (N_10122,N_9182,N_9180);
nand U10123 (N_10123,N_9100,N_9230);
xor U10124 (N_10124,N_9205,N_9558);
xnor U10125 (N_10125,N_9412,N_9384);
nor U10126 (N_10126,N_9132,N_9144);
nand U10127 (N_10127,N_9664,N_9259);
xor U10128 (N_10128,N_9665,N_9729);
and U10129 (N_10129,N_9566,N_9484);
nor U10130 (N_10130,N_9664,N_9684);
xnor U10131 (N_10131,N_9545,N_9403);
nor U10132 (N_10132,N_9410,N_9529);
xnor U10133 (N_10133,N_9384,N_9145);
nand U10134 (N_10134,N_9260,N_9276);
xnor U10135 (N_10135,N_9008,N_9251);
or U10136 (N_10136,N_9114,N_9034);
or U10137 (N_10137,N_9596,N_9522);
and U10138 (N_10138,N_9202,N_9260);
and U10139 (N_10139,N_9418,N_9184);
and U10140 (N_10140,N_9578,N_9645);
and U10141 (N_10141,N_9064,N_9075);
and U10142 (N_10142,N_9463,N_9426);
xor U10143 (N_10143,N_9189,N_9726);
nand U10144 (N_10144,N_9098,N_9207);
nand U10145 (N_10145,N_9532,N_9304);
nand U10146 (N_10146,N_9522,N_9429);
nor U10147 (N_10147,N_9425,N_9182);
nor U10148 (N_10148,N_9272,N_9043);
or U10149 (N_10149,N_9168,N_9411);
and U10150 (N_10150,N_9471,N_9322);
nand U10151 (N_10151,N_9387,N_9619);
nor U10152 (N_10152,N_9080,N_9652);
nor U10153 (N_10153,N_9433,N_9064);
nor U10154 (N_10154,N_9645,N_9431);
or U10155 (N_10155,N_9719,N_9221);
nor U10156 (N_10156,N_9621,N_9733);
nor U10157 (N_10157,N_9388,N_9518);
xnor U10158 (N_10158,N_9337,N_9089);
nor U10159 (N_10159,N_9260,N_9319);
or U10160 (N_10160,N_9191,N_9168);
or U10161 (N_10161,N_9284,N_9319);
and U10162 (N_10162,N_9614,N_9267);
and U10163 (N_10163,N_9057,N_9728);
or U10164 (N_10164,N_9618,N_9189);
and U10165 (N_10165,N_9319,N_9164);
nor U10166 (N_10166,N_9085,N_9086);
nand U10167 (N_10167,N_9749,N_9086);
or U10168 (N_10168,N_9446,N_9397);
and U10169 (N_10169,N_9532,N_9568);
and U10170 (N_10170,N_9234,N_9015);
nor U10171 (N_10171,N_9624,N_9659);
nand U10172 (N_10172,N_9050,N_9299);
xor U10173 (N_10173,N_9036,N_9514);
or U10174 (N_10174,N_9190,N_9307);
xor U10175 (N_10175,N_9044,N_9137);
xnor U10176 (N_10176,N_9455,N_9662);
or U10177 (N_10177,N_9692,N_9694);
and U10178 (N_10178,N_9369,N_9327);
nand U10179 (N_10179,N_9312,N_9429);
and U10180 (N_10180,N_9268,N_9495);
and U10181 (N_10181,N_9708,N_9730);
nor U10182 (N_10182,N_9412,N_9416);
nor U10183 (N_10183,N_9422,N_9522);
and U10184 (N_10184,N_9572,N_9303);
nand U10185 (N_10185,N_9092,N_9429);
or U10186 (N_10186,N_9682,N_9689);
or U10187 (N_10187,N_9546,N_9297);
nor U10188 (N_10188,N_9224,N_9341);
xnor U10189 (N_10189,N_9464,N_9518);
or U10190 (N_10190,N_9539,N_9501);
and U10191 (N_10191,N_9607,N_9275);
xor U10192 (N_10192,N_9384,N_9572);
and U10193 (N_10193,N_9111,N_9417);
or U10194 (N_10194,N_9190,N_9471);
xor U10195 (N_10195,N_9080,N_9665);
xnor U10196 (N_10196,N_9523,N_9590);
nor U10197 (N_10197,N_9542,N_9168);
nor U10198 (N_10198,N_9745,N_9283);
nor U10199 (N_10199,N_9537,N_9668);
nor U10200 (N_10200,N_9034,N_9612);
or U10201 (N_10201,N_9097,N_9105);
nor U10202 (N_10202,N_9625,N_9012);
xnor U10203 (N_10203,N_9214,N_9090);
nor U10204 (N_10204,N_9345,N_9168);
xnor U10205 (N_10205,N_9684,N_9626);
and U10206 (N_10206,N_9347,N_9568);
nor U10207 (N_10207,N_9329,N_9504);
and U10208 (N_10208,N_9129,N_9449);
nor U10209 (N_10209,N_9188,N_9527);
or U10210 (N_10210,N_9740,N_9442);
nand U10211 (N_10211,N_9262,N_9192);
and U10212 (N_10212,N_9522,N_9044);
nand U10213 (N_10213,N_9262,N_9127);
nor U10214 (N_10214,N_9230,N_9461);
nand U10215 (N_10215,N_9518,N_9076);
xnor U10216 (N_10216,N_9623,N_9019);
nor U10217 (N_10217,N_9721,N_9452);
or U10218 (N_10218,N_9406,N_9228);
or U10219 (N_10219,N_9668,N_9368);
xnor U10220 (N_10220,N_9158,N_9567);
or U10221 (N_10221,N_9022,N_9043);
or U10222 (N_10222,N_9473,N_9087);
nor U10223 (N_10223,N_9341,N_9256);
or U10224 (N_10224,N_9037,N_9313);
and U10225 (N_10225,N_9282,N_9641);
and U10226 (N_10226,N_9204,N_9039);
xor U10227 (N_10227,N_9472,N_9332);
xor U10228 (N_10228,N_9568,N_9491);
xnor U10229 (N_10229,N_9426,N_9025);
nor U10230 (N_10230,N_9747,N_9643);
or U10231 (N_10231,N_9175,N_9059);
xor U10232 (N_10232,N_9023,N_9357);
or U10233 (N_10233,N_9641,N_9227);
nand U10234 (N_10234,N_9627,N_9573);
xor U10235 (N_10235,N_9663,N_9610);
and U10236 (N_10236,N_9090,N_9525);
or U10237 (N_10237,N_9623,N_9568);
nand U10238 (N_10238,N_9111,N_9601);
and U10239 (N_10239,N_9540,N_9537);
nand U10240 (N_10240,N_9411,N_9290);
nand U10241 (N_10241,N_9700,N_9314);
xnor U10242 (N_10242,N_9272,N_9274);
nand U10243 (N_10243,N_9607,N_9427);
nor U10244 (N_10244,N_9287,N_9047);
nor U10245 (N_10245,N_9661,N_9441);
or U10246 (N_10246,N_9115,N_9617);
nor U10247 (N_10247,N_9457,N_9470);
xnor U10248 (N_10248,N_9708,N_9100);
xnor U10249 (N_10249,N_9658,N_9006);
xnor U10250 (N_10250,N_9216,N_9275);
xnor U10251 (N_10251,N_9385,N_9606);
or U10252 (N_10252,N_9713,N_9708);
or U10253 (N_10253,N_9215,N_9434);
nand U10254 (N_10254,N_9674,N_9712);
nor U10255 (N_10255,N_9349,N_9232);
nor U10256 (N_10256,N_9074,N_9399);
xor U10257 (N_10257,N_9698,N_9674);
nand U10258 (N_10258,N_9351,N_9191);
and U10259 (N_10259,N_9505,N_9533);
nand U10260 (N_10260,N_9041,N_9042);
and U10261 (N_10261,N_9525,N_9244);
and U10262 (N_10262,N_9159,N_9080);
and U10263 (N_10263,N_9045,N_9378);
and U10264 (N_10264,N_9465,N_9572);
nand U10265 (N_10265,N_9323,N_9342);
nand U10266 (N_10266,N_9619,N_9510);
nand U10267 (N_10267,N_9621,N_9611);
and U10268 (N_10268,N_9007,N_9747);
or U10269 (N_10269,N_9568,N_9368);
nor U10270 (N_10270,N_9686,N_9111);
or U10271 (N_10271,N_9460,N_9541);
xor U10272 (N_10272,N_9609,N_9348);
nor U10273 (N_10273,N_9065,N_9650);
nand U10274 (N_10274,N_9655,N_9518);
nand U10275 (N_10275,N_9048,N_9256);
nand U10276 (N_10276,N_9015,N_9030);
or U10277 (N_10277,N_9550,N_9351);
xnor U10278 (N_10278,N_9318,N_9138);
nand U10279 (N_10279,N_9415,N_9010);
nand U10280 (N_10280,N_9430,N_9626);
or U10281 (N_10281,N_9337,N_9016);
nor U10282 (N_10282,N_9712,N_9222);
and U10283 (N_10283,N_9030,N_9092);
nand U10284 (N_10284,N_9103,N_9032);
nand U10285 (N_10285,N_9622,N_9270);
and U10286 (N_10286,N_9065,N_9251);
or U10287 (N_10287,N_9507,N_9660);
nor U10288 (N_10288,N_9500,N_9680);
nor U10289 (N_10289,N_9100,N_9095);
nor U10290 (N_10290,N_9372,N_9699);
nand U10291 (N_10291,N_9671,N_9394);
xor U10292 (N_10292,N_9216,N_9603);
or U10293 (N_10293,N_9555,N_9308);
nor U10294 (N_10294,N_9356,N_9612);
and U10295 (N_10295,N_9064,N_9468);
or U10296 (N_10296,N_9556,N_9266);
xnor U10297 (N_10297,N_9441,N_9678);
nor U10298 (N_10298,N_9563,N_9747);
nand U10299 (N_10299,N_9227,N_9438);
nor U10300 (N_10300,N_9224,N_9606);
nand U10301 (N_10301,N_9208,N_9218);
and U10302 (N_10302,N_9470,N_9300);
nand U10303 (N_10303,N_9563,N_9169);
xor U10304 (N_10304,N_9248,N_9132);
nor U10305 (N_10305,N_9743,N_9379);
nand U10306 (N_10306,N_9114,N_9104);
nand U10307 (N_10307,N_9276,N_9594);
nor U10308 (N_10308,N_9738,N_9589);
nor U10309 (N_10309,N_9028,N_9107);
xor U10310 (N_10310,N_9518,N_9218);
nand U10311 (N_10311,N_9666,N_9005);
or U10312 (N_10312,N_9175,N_9458);
or U10313 (N_10313,N_9038,N_9263);
nand U10314 (N_10314,N_9498,N_9233);
nor U10315 (N_10315,N_9400,N_9374);
xor U10316 (N_10316,N_9306,N_9378);
and U10317 (N_10317,N_9385,N_9384);
xnor U10318 (N_10318,N_9168,N_9351);
and U10319 (N_10319,N_9709,N_9274);
nor U10320 (N_10320,N_9299,N_9370);
nand U10321 (N_10321,N_9282,N_9182);
and U10322 (N_10322,N_9470,N_9290);
or U10323 (N_10323,N_9476,N_9645);
xnor U10324 (N_10324,N_9147,N_9550);
nand U10325 (N_10325,N_9122,N_9278);
nand U10326 (N_10326,N_9342,N_9365);
nand U10327 (N_10327,N_9712,N_9175);
xnor U10328 (N_10328,N_9084,N_9286);
xnor U10329 (N_10329,N_9078,N_9457);
nand U10330 (N_10330,N_9645,N_9022);
and U10331 (N_10331,N_9390,N_9426);
and U10332 (N_10332,N_9100,N_9031);
or U10333 (N_10333,N_9579,N_9625);
or U10334 (N_10334,N_9215,N_9528);
nand U10335 (N_10335,N_9271,N_9107);
or U10336 (N_10336,N_9571,N_9562);
xnor U10337 (N_10337,N_9369,N_9333);
nand U10338 (N_10338,N_9601,N_9492);
nand U10339 (N_10339,N_9021,N_9344);
nor U10340 (N_10340,N_9482,N_9578);
nand U10341 (N_10341,N_9473,N_9230);
or U10342 (N_10342,N_9186,N_9665);
nor U10343 (N_10343,N_9063,N_9116);
nor U10344 (N_10344,N_9196,N_9642);
or U10345 (N_10345,N_9227,N_9418);
and U10346 (N_10346,N_9140,N_9338);
nand U10347 (N_10347,N_9208,N_9037);
and U10348 (N_10348,N_9662,N_9288);
nor U10349 (N_10349,N_9037,N_9411);
xnor U10350 (N_10350,N_9139,N_9214);
and U10351 (N_10351,N_9468,N_9230);
nand U10352 (N_10352,N_9082,N_9698);
nor U10353 (N_10353,N_9447,N_9256);
and U10354 (N_10354,N_9111,N_9165);
xnor U10355 (N_10355,N_9434,N_9038);
xnor U10356 (N_10356,N_9088,N_9601);
and U10357 (N_10357,N_9033,N_9252);
and U10358 (N_10358,N_9417,N_9065);
xor U10359 (N_10359,N_9739,N_9232);
nor U10360 (N_10360,N_9049,N_9620);
nand U10361 (N_10361,N_9200,N_9578);
and U10362 (N_10362,N_9060,N_9279);
or U10363 (N_10363,N_9065,N_9346);
or U10364 (N_10364,N_9059,N_9613);
nand U10365 (N_10365,N_9056,N_9390);
and U10366 (N_10366,N_9645,N_9544);
xnor U10367 (N_10367,N_9647,N_9549);
nand U10368 (N_10368,N_9221,N_9635);
or U10369 (N_10369,N_9615,N_9572);
and U10370 (N_10370,N_9275,N_9203);
and U10371 (N_10371,N_9632,N_9307);
nor U10372 (N_10372,N_9032,N_9417);
xor U10373 (N_10373,N_9069,N_9363);
nand U10374 (N_10374,N_9155,N_9317);
or U10375 (N_10375,N_9128,N_9707);
and U10376 (N_10376,N_9102,N_9516);
nand U10377 (N_10377,N_9034,N_9385);
or U10378 (N_10378,N_9729,N_9410);
and U10379 (N_10379,N_9540,N_9193);
and U10380 (N_10380,N_9246,N_9014);
nor U10381 (N_10381,N_9512,N_9716);
or U10382 (N_10382,N_9740,N_9369);
nor U10383 (N_10383,N_9580,N_9336);
or U10384 (N_10384,N_9147,N_9351);
or U10385 (N_10385,N_9297,N_9167);
xnor U10386 (N_10386,N_9651,N_9560);
xor U10387 (N_10387,N_9130,N_9409);
and U10388 (N_10388,N_9060,N_9030);
nor U10389 (N_10389,N_9284,N_9536);
xnor U10390 (N_10390,N_9461,N_9748);
or U10391 (N_10391,N_9104,N_9570);
and U10392 (N_10392,N_9115,N_9234);
and U10393 (N_10393,N_9730,N_9028);
or U10394 (N_10394,N_9277,N_9506);
nand U10395 (N_10395,N_9283,N_9057);
nand U10396 (N_10396,N_9246,N_9361);
or U10397 (N_10397,N_9166,N_9613);
and U10398 (N_10398,N_9266,N_9414);
and U10399 (N_10399,N_9280,N_9307);
nand U10400 (N_10400,N_9016,N_9579);
nor U10401 (N_10401,N_9193,N_9743);
and U10402 (N_10402,N_9615,N_9604);
or U10403 (N_10403,N_9173,N_9567);
xor U10404 (N_10404,N_9478,N_9372);
nor U10405 (N_10405,N_9444,N_9543);
nor U10406 (N_10406,N_9483,N_9653);
nor U10407 (N_10407,N_9164,N_9162);
or U10408 (N_10408,N_9479,N_9313);
nor U10409 (N_10409,N_9208,N_9012);
xnor U10410 (N_10410,N_9144,N_9692);
and U10411 (N_10411,N_9303,N_9428);
nand U10412 (N_10412,N_9401,N_9505);
and U10413 (N_10413,N_9063,N_9398);
nor U10414 (N_10414,N_9560,N_9509);
or U10415 (N_10415,N_9689,N_9737);
or U10416 (N_10416,N_9108,N_9720);
or U10417 (N_10417,N_9358,N_9650);
nand U10418 (N_10418,N_9647,N_9005);
xnor U10419 (N_10419,N_9607,N_9205);
or U10420 (N_10420,N_9647,N_9069);
and U10421 (N_10421,N_9254,N_9455);
and U10422 (N_10422,N_9423,N_9158);
xnor U10423 (N_10423,N_9308,N_9655);
nand U10424 (N_10424,N_9518,N_9661);
or U10425 (N_10425,N_9109,N_9122);
and U10426 (N_10426,N_9740,N_9662);
and U10427 (N_10427,N_9331,N_9321);
nand U10428 (N_10428,N_9093,N_9128);
nand U10429 (N_10429,N_9056,N_9179);
or U10430 (N_10430,N_9400,N_9353);
nand U10431 (N_10431,N_9004,N_9701);
or U10432 (N_10432,N_9318,N_9434);
xnor U10433 (N_10433,N_9157,N_9020);
xor U10434 (N_10434,N_9441,N_9575);
nor U10435 (N_10435,N_9067,N_9398);
nand U10436 (N_10436,N_9180,N_9435);
nand U10437 (N_10437,N_9223,N_9018);
nand U10438 (N_10438,N_9171,N_9001);
xnor U10439 (N_10439,N_9470,N_9555);
nor U10440 (N_10440,N_9576,N_9580);
xnor U10441 (N_10441,N_9418,N_9037);
and U10442 (N_10442,N_9124,N_9312);
and U10443 (N_10443,N_9598,N_9117);
or U10444 (N_10444,N_9050,N_9538);
nand U10445 (N_10445,N_9515,N_9527);
xor U10446 (N_10446,N_9249,N_9006);
xnor U10447 (N_10447,N_9479,N_9485);
xor U10448 (N_10448,N_9609,N_9273);
xnor U10449 (N_10449,N_9098,N_9340);
or U10450 (N_10450,N_9097,N_9195);
xor U10451 (N_10451,N_9699,N_9275);
or U10452 (N_10452,N_9424,N_9501);
and U10453 (N_10453,N_9637,N_9142);
xnor U10454 (N_10454,N_9479,N_9224);
nor U10455 (N_10455,N_9274,N_9004);
nand U10456 (N_10456,N_9414,N_9725);
or U10457 (N_10457,N_9059,N_9623);
xor U10458 (N_10458,N_9686,N_9401);
or U10459 (N_10459,N_9100,N_9082);
nand U10460 (N_10460,N_9710,N_9085);
or U10461 (N_10461,N_9398,N_9295);
or U10462 (N_10462,N_9226,N_9228);
or U10463 (N_10463,N_9246,N_9420);
and U10464 (N_10464,N_9155,N_9161);
and U10465 (N_10465,N_9711,N_9730);
or U10466 (N_10466,N_9743,N_9668);
nor U10467 (N_10467,N_9588,N_9466);
xnor U10468 (N_10468,N_9050,N_9566);
xor U10469 (N_10469,N_9330,N_9570);
and U10470 (N_10470,N_9145,N_9699);
nor U10471 (N_10471,N_9498,N_9048);
nand U10472 (N_10472,N_9697,N_9327);
or U10473 (N_10473,N_9098,N_9260);
or U10474 (N_10474,N_9029,N_9009);
or U10475 (N_10475,N_9097,N_9449);
or U10476 (N_10476,N_9611,N_9178);
and U10477 (N_10477,N_9678,N_9324);
and U10478 (N_10478,N_9192,N_9073);
nand U10479 (N_10479,N_9549,N_9628);
xor U10480 (N_10480,N_9624,N_9394);
nand U10481 (N_10481,N_9288,N_9183);
or U10482 (N_10482,N_9298,N_9435);
or U10483 (N_10483,N_9173,N_9107);
or U10484 (N_10484,N_9665,N_9626);
nand U10485 (N_10485,N_9171,N_9058);
and U10486 (N_10486,N_9092,N_9728);
and U10487 (N_10487,N_9452,N_9287);
xnor U10488 (N_10488,N_9395,N_9163);
xnor U10489 (N_10489,N_9384,N_9488);
nor U10490 (N_10490,N_9534,N_9587);
or U10491 (N_10491,N_9507,N_9459);
or U10492 (N_10492,N_9528,N_9747);
and U10493 (N_10493,N_9247,N_9645);
xor U10494 (N_10494,N_9068,N_9090);
nor U10495 (N_10495,N_9131,N_9414);
and U10496 (N_10496,N_9492,N_9350);
nor U10497 (N_10497,N_9331,N_9542);
xnor U10498 (N_10498,N_9205,N_9499);
or U10499 (N_10499,N_9498,N_9507);
nand U10500 (N_10500,N_10048,N_10027);
nand U10501 (N_10501,N_10179,N_10317);
nand U10502 (N_10502,N_10059,N_9794);
nor U10503 (N_10503,N_9861,N_9813);
xor U10504 (N_10504,N_10396,N_10232);
or U10505 (N_10505,N_10283,N_10119);
or U10506 (N_10506,N_10345,N_10056);
xnor U10507 (N_10507,N_10407,N_10094);
xor U10508 (N_10508,N_9761,N_10159);
or U10509 (N_10509,N_10450,N_9974);
nand U10510 (N_10510,N_10004,N_9903);
nor U10511 (N_10511,N_10164,N_9826);
nor U10512 (N_10512,N_10281,N_10052);
or U10513 (N_10513,N_10416,N_9940);
and U10514 (N_10514,N_10168,N_9853);
nand U10515 (N_10515,N_9783,N_9837);
and U10516 (N_10516,N_9816,N_10028);
and U10517 (N_10517,N_9988,N_10008);
nor U10518 (N_10518,N_9867,N_10394);
nand U10519 (N_10519,N_10270,N_10492);
nor U10520 (N_10520,N_9991,N_10442);
or U10521 (N_10521,N_9948,N_10477);
and U10522 (N_10522,N_10136,N_10334);
nor U10523 (N_10523,N_9963,N_10252);
and U10524 (N_10524,N_10458,N_10221);
nor U10525 (N_10525,N_10390,N_10089);
nand U10526 (N_10526,N_10378,N_10403);
xnor U10527 (N_10527,N_10397,N_10393);
nor U10528 (N_10528,N_10014,N_10034);
nor U10529 (N_10529,N_9844,N_10408);
or U10530 (N_10530,N_9842,N_9845);
nor U10531 (N_10531,N_10031,N_10101);
xnor U10532 (N_10532,N_10349,N_10006);
or U10533 (N_10533,N_9777,N_9976);
nand U10534 (N_10534,N_10488,N_10234);
and U10535 (N_10535,N_10333,N_10395);
or U10536 (N_10536,N_10124,N_10447);
xnor U10537 (N_10537,N_10026,N_9788);
xnor U10538 (N_10538,N_10371,N_10466);
and U10539 (N_10539,N_9793,N_9970);
and U10540 (N_10540,N_10181,N_10023);
nand U10541 (N_10541,N_10385,N_10263);
xnor U10542 (N_10542,N_10370,N_10498);
nor U10543 (N_10543,N_9756,N_9967);
xnor U10544 (N_10544,N_9764,N_10248);
nor U10545 (N_10545,N_10173,N_10314);
and U10546 (N_10546,N_10228,N_9854);
nand U10547 (N_10547,N_10068,N_10104);
or U10548 (N_10548,N_10233,N_9901);
and U10549 (N_10549,N_9921,N_10446);
xor U10550 (N_10550,N_10099,N_10236);
nand U10551 (N_10551,N_10318,N_9876);
or U10552 (N_10552,N_9910,N_10042);
xnor U10553 (N_10553,N_10142,N_10432);
or U10554 (N_10554,N_9857,N_10376);
xor U10555 (N_10555,N_10086,N_10231);
nor U10556 (N_10556,N_10463,N_10346);
nor U10557 (N_10557,N_10344,N_10340);
or U10558 (N_10558,N_9997,N_10046);
and U10559 (N_10559,N_9993,N_10058);
nand U10560 (N_10560,N_10037,N_10342);
nor U10561 (N_10561,N_10377,N_10448);
or U10562 (N_10562,N_10276,N_10194);
and U10563 (N_10563,N_10067,N_10215);
or U10564 (N_10564,N_9961,N_9886);
nor U10565 (N_10565,N_10125,N_9787);
or U10566 (N_10566,N_10130,N_9980);
nand U10567 (N_10567,N_10241,N_10325);
and U10568 (N_10568,N_10435,N_10108);
nand U10569 (N_10569,N_10444,N_10080);
and U10570 (N_10570,N_9949,N_9931);
xnor U10571 (N_10571,N_10409,N_9850);
or U10572 (N_10572,N_10404,N_9778);
nand U10573 (N_10573,N_10122,N_10485);
nor U10574 (N_10574,N_9800,N_10392);
nand U10575 (N_10575,N_10123,N_10030);
or U10576 (N_10576,N_10296,N_10003);
or U10577 (N_10577,N_9965,N_10284);
or U10578 (N_10578,N_10041,N_10206);
and U10579 (N_10579,N_9899,N_9977);
and U10580 (N_10580,N_9798,N_10106);
xor U10581 (N_10581,N_10480,N_10468);
nor U10582 (N_10582,N_9913,N_10256);
nor U10583 (N_10583,N_10237,N_10309);
and U10584 (N_10584,N_9916,N_10338);
xnor U10585 (N_10585,N_10029,N_10322);
or U10586 (N_10586,N_10210,N_9807);
xor U10587 (N_10587,N_9972,N_10483);
nor U10588 (N_10588,N_10065,N_10077);
xor U10589 (N_10589,N_9796,N_9932);
and U10590 (N_10590,N_10329,N_10151);
xnor U10591 (N_10591,N_9797,N_10311);
or U10592 (N_10592,N_10272,N_10487);
xnor U10593 (N_10593,N_9811,N_10091);
nor U10594 (N_10594,N_9862,N_10182);
and U10595 (N_10595,N_10096,N_10118);
nand U10596 (N_10596,N_10440,N_9926);
nand U10597 (N_10597,N_9960,N_9866);
nand U10598 (N_10598,N_10022,N_9819);
nor U10599 (N_10599,N_10259,N_9964);
nand U10600 (N_10600,N_9814,N_10481);
or U10601 (N_10601,N_10454,N_10001);
nand U10602 (N_10602,N_9776,N_10304);
and U10603 (N_10603,N_9873,N_10364);
nor U10604 (N_10604,N_9839,N_10083);
and U10605 (N_10605,N_9896,N_10465);
and U10606 (N_10606,N_10245,N_10285);
nor U10607 (N_10607,N_10074,N_10307);
or U10608 (N_10608,N_10093,N_9922);
nor U10609 (N_10609,N_10290,N_9805);
xor U10610 (N_10610,N_10105,N_9894);
and U10611 (N_10611,N_10191,N_9933);
xnor U10612 (N_10612,N_10186,N_10484);
nand U10613 (N_10613,N_10464,N_10359);
nand U10614 (N_10614,N_9898,N_9834);
xor U10615 (N_10615,N_10145,N_9982);
or U10616 (N_10616,N_10043,N_10354);
nor U10617 (N_10617,N_9950,N_10266);
nand U10618 (N_10618,N_10461,N_10439);
xor U10619 (N_10619,N_10496,N_10475);
nor U10620 (N_10620,N_10121,N_10131);
and U10621 (N_10621,N_9944,N_9841);
xnor U10622 (N_10622,N_9752,N_9897);
and U10623 (N_10623,N_10459,N_10032);
or U10624 (N_10624,N_9835,N_10147);
xor U10625 (N_10625,N_9846,N_10391);
nand U10626 (N_10626,N_10189,N_10295);
and U10627 (N_10627,N_9979,N_10209);
or U10628 (N_10628,N_9924,N_9969);
nand U10629 (N_10629,N_10117,N_9840);
or U10630 (N_10630,N_10286,N_10177);
or U10631 (N_10631,N_10453,N_10471);
nor U10632 (N_10632,N_9789,N_9986);
and U10633 (N_10633,N_10375,N_9773);
xnor U10634 (N_10634,N_10313,N_9824);
xor U10635 (N_10635,N_10161,N_10187);
xnor U10636 (N_10636,N_9851,N_10462);
nand U10637 (N_10637,N_10347,N_10335);
nor U10638 (N_10638,N_9829,N_9911);
or U10639 (N_10639,N_10456,N_9904);
nand U10640 (N_10640,N_9860,N_9781);
nor U10641 (N_10641,N_10428,N_10102);
nor U10642 (N_10642,N_10415,N_10425);
nand U10643 (N_10643,N_10064,N_10242);
nor U10644 (N_10644,N_9930,N_10353);
nand U10645 (N_10645,N_10024,N_10383);
or U10646 (N_10646,N_10156,N_10040);
nand U10647 (N_10647,N_9989,N_9992);
nor U10648 (N_10648,N_10146,N_9808);
xnor U10649 (N_10649,N_10305,N_10414);
nor U10650 (N_10650,N_9996,N_10293);
xor U10651 (N_10651,N_10424,N_9848);
nand U10652 (N_10652,N_10257,N_10380);
and U10653 (N_10653,N_9772,N_9920);
xor U10654 (N_10654,N_9809,N_9919);
or U10655 (N_10655,N_10116,N_10054);
or U10656 (N_10656,N_10264,N_10036);
nand U10657 (N_10657,N_9943,N_9833);
nand U10658 (N_10658,N_10160,N_10298);
nand U10659 (N_10659,N_10114,N_10148);
and U10660 (N_10660,N_10216,N_10417);
or U10661 (N_10661,N_10207,N_10012);
xor U10662 (N_10662,N_10129,N_10153);
nand U10663 (N_10663,N_9875,N_9954);
and U10664 (N_10664,N_10184,N_9900);
and U10665 (N_10665,N_10165,N_10192);
xor U10666 (N_10666,N_10111,N_9892);
xor U10667 (N_10667,N_10332,N_9768);
nand U10668 (N_10668,N_9951,N_10324);
nand U10669 (N_10669,N_9975,N_10323);
or U10670 (N_10670,N_10127,N_10306);
xnor U10671 (N_10671,N_9971,N_10490);
xnor U10672 (N_10672,N_10388,N_10002);
nand U10673 (N_10673,N_10015,N_9831);
xnor U10674 (N_10674,N_10204,N_9874);
nand U10675 (N_10675,N_10066,N_10382);
nor U10676 (N_10676,N_10467,N_10398);
or U10677 (N_10677,N_10261,N_10365);
nand U10678 (N_10678,N_10198,N_10292);
nand U10679 (N_10679,N_10452,N_9865);
nand U10680 (N_10680,N_10087,N_9935);
nor U10681 (N_10681,N_10132,N_10282);
and U10682 (N_10682,N_10235,N_10433);
xor U10683 (N_10683,N_9998,N_10300);
nand U10684 (N_10684,N_10482,N_10355);
xor U10685 (N_10685,N_10260,N_9864);
xor U10686 (N_10686,N_10202,N_10176);
xnor U10687 (N_10687,N_10128,N_10339);
or U10688 (N_10688,N_10497,N_10138);
and U10689 (N_10689,N_10076,N_10188);
or U10690 (N_10690,N_9959,N_9812);
and U10691 (N_10691,N_10197,N_9906);
nor U10692 (N_10692,N_10288,N_10410);
or U10693 (N_10693,N_10273,N_10294);
nor U10694 (N_10694,N_10268,N_9871);
nor U10695 (N_10695,N_10357,N_9868);
nor U10696 (N_10696,N_10170,N_9784);
xnor U10697 (N_10697,N_9891,N_10211);
and U10698 (N_10698,N_9966,N_10438);
nand U10699 (N_10699,N_10049,N_10372);
and U10700 (N_10700,N_10443,N_10238);
or U10701 (N_10701,N_10071,N_9804);
xor U10702 (N_10702,N_10251,N_9887);
xnor U10703 (N_10703,N_10180,N_9942);
xor U10704 (N_10704,N_9877,N_10280);
or U10705 (N_10705,N_9858,N_9987);
xnor U10706 (N_10706,N_9774,N_10254);
xnor U10707 (N_10707,N_10402,N_10472);
and U10708 (N_10708,N_9879,N_9782);
nand U10709 (N_10709,N_10045,N_10301);
nor U10710 (N_10710,N_10149,N_10038);
nand U10711 (N_10711,N_9762,N_10434);
nor U10712 (N_10712,N_10474,N_10449);
nand U10713 (N_10713,N_9936,N_10223);
nand U10714 (N_10714,N_9759,N_9999);
xor U10715 (N_10715,N_10203,N_9770);
nor U10716 (N_10716,N_10360,N_10208);
and U10717 (N_10717,N_10158,N_10494);
xor U10718 (N_10718,N_10374,N_9817);
nor U10719 (N_10719,N_10411,N_9792);
and U10720 (N_10720,N_10356,N_10229);
xnor U10721 (N_10721,N_10009,N_9983);
xnor U10722 (N_10722,N_10381,N_10244);
nand U10723 (N_10723,N_9820,N_10423);
nand U10724 (N_10724,N_10098,N_10451);
nor U10725 (N_10725,N_9908,N_10315);
nand U10726 (N_10726,N_9815,N_9823);
xnor U10727 (N_10727,N_10057,N_10139);
or U10728 (N_10728,N_10289,N_9765);
and U10729 (N_10729,N_9863,N_9849);
xnor U10730 (N_10730,N_10088,N_10469);
nand U10731 (N_10731,N_10412,N_9767);
xor U10732 (N_10732,N_10476,N_10169);
nand U10733 (N_10733,N_10219,N_9890);
nand U10734 (N_10734,N_10312,N_10175);
xnor U10735 (N_10735,N_10150,N_10455);
xnor U10736 (N_10736,N_9843,N_10362);
or U10737 (N_10737,N_9918,N_10007);
nor U10738 (N_10738,N_10016,N_10230);
nor U10739 (N_10739,N_10072,N_10269);
and U10740 (N_10740,N_10274,N_10051);
nor U10741 (N_10741,N_9995,N_10431);
xnor U10742 (N_10742,N_10092,N_10243);
or U10743 (N_10743,N_10299,N_10155);
xnor U10744 (N_10744,N_9914,N_10060);
or U10745 (N_10745,N_10140,N_10427);
and U10746 (N_10746,N_9779,N_10271);
xor U10747 (N_10747,N_9907,N_9895);
and U10748 (N_10748,N_9880,N_10025);
xnor U10749 (N_10749,N_10011,N_10120);
xnor U10750 (N_10750,N_10258,N_10134);
nand U10751 (N_10751,N_9818,N_10033);
nand U10752 (N_10752,N_10419,N_10070);
and U10753 (N_10753,N_10073,N_10321);
and U10754 (N_10754,N_10133,N_10441);
nand U10755 (N_10755,N_10010,N_9881);
and U10756 (N_10756,N_9923,N_10328);
and U10757 (N_10757,N_10316,N_10174);
or U10758 (N_10758,N_9821,N_9828);
xnor U10759 (N_10759,N_10199,N_10069);
xnor U10760 (N_10760,N_10250,N_9937);
and U10761 (N_10761,N_10200,N_10302);
nor U10762 (N_10762,N_10291,N_9915);
xor U10763 (N_10763,N_10227,N_10361);
or U10764 (N_10764,N_9822,N_10095);
or U10765 (N_10765,N_10220,N_10247);
nand U10766 (N_10766,N_10386,N_9855);
and U10767 (N_10767,N_9754,N_9925);
or U10768 (N_10768,N_10255,N_10367);
and U10769 (N_10769,N_10107,N_10308);
or U10770 (N_10770,N_10172,N_10141);
xnor U10771 (N_10771,N_10368,N_9763);
nor U10772 (N_10772,N_9909,N_10167);
or U10773 (N_10773,N_9938,N_10144);
or U10774 (N_10774,N_10422,N_10115);
or U10775 (N_10775,N_9984,N_10152);
and U10776 (N_10776,N_9775,N_9827);
nor U10777 (N_10777,N_10429,N_10000);
xor U10778 (N_10778,N_10278,N_9780);
and U10779 (N_10779,N_9978,N_10479);
nor U10780 (N_10780,N_9883,N_9994);
or U10781 (N_10781,N_9803,N_10097);
xor U10782 (N_10782,N_9847,N_9990);
or U10783 (N_10783,N_10082,N_9928);
nand U10784 (N_10784,N_9795,N_10436);
nand U10785 (N_10785,N_10019,N_10062);
and U10786 (N_10786,N_9889,N_9927);
nor U10787 (N_10787,N_10413,N_10326);
or U10788 (N_10788,N_10226,N_10470);
nor U10789 (N_10789,N_9791,N_9882);
and U10790 (N_10790,N_9902,N_9878);
and U10791 (N_10791,N_10103,N_10491);
nand U10792 (N_10792,N_10421,N_9755);
xor U10793 (N_10793,N_10075,N_10253);
xnor U10794 (N_10794,N_10337,N_10426);
nor U10795 (N_10795,N_9750,N_10499);
nor U10796 (N_10796,N_10166,N_10135);
or U10797 (N_10797,N_10320,N_9859);
or U10798 (N_10798,N_10478,N_9825);
nand U10799 (N_10799,N_9893,N_9766);
xor U10800 (N_10800,N_10400,N_10217);
xor U10801 (N_10801,N_9786,N_9957);
nor U10802 (N_10802,N_10369,N_10239);
nor U10803 (N_10803,N_10109,N_9832);
and U10804 (N_10804,N_9872,N_9985);
and U10805 (N_10805,N_10017,N_10489);
xor U10806 (N_10806,N_9758,N_10420);
xnor U10807 (N_10807,N_9929,N_10373);
or U10808 (N_10808,N_10044,N_10418);
nor U10809 (N_10809,N_10039,N_10113);
and U10810 (N_10810,N_10085,N_10047);
nor U10811 (N_10811,N_10240,N_10350);
and U10812 (N_10812,N_9802,N_9941);
nor U10813 (N_10813,N_10021,N_9806);
nor U10814 (N_10814,N_9956,N_10279);
and U10815 (N_10815,N_9785,N_10212);
and U10816 (N_10816,N_10437,N_10084);
xor U10817 (N_10817,N_10343,N_10366);
or U10818 (N_10818,N_10265,N_10100);
xor U10819 (N_10819,N_9945,N_10363);
or U10820 (N_10820,N_9934,N_10020);
nor U10821 (N_10821,N_10157,N_10050);
or U10822 (N_10822,N_10225,N_10389);
or U10823 (N_10823,N_10310,N_10195);
or U10824 (N_10824,N_10384,N_9905);
xnor U10825 (N_10825,N_9757,N_10473);
or U10826 (N_10826,N_10185,N_10224);
or U10827 (N_10827,N_9939,N_9856);
or U10828 (N_10828,N_10336,N_10331);
xnor U10829 (N_10829,N_9760,N_9947);
nor U10830 (N_10830,N_10406,N_10348);
xnor U10831 (N_10831,N_9973,N_9946);
or U10832 (N_10832,N_10078,N_10277);
nor U10833 (N_10833,N_9751,N_10399);
nor U10834 (N_10834,N_10081,N_9958);
nor U10835 (N_10835,N_10162,N_10457);
nor U10836 (N_10836,N_9838,N_10183);
nand U10837 (N_10837,N_10246,N_9830);
or U10838 (N_10838,N_9912,N_10287);
nand U10839 (N_10839,N_10090,N_10445);
xnor U10840 (N_10840,N_10112,N_9852);
and U10841 (N_10841,N_10387,N_10327);
nor U10842 (N_10842,N_10196,N_10143);
and U10843 (N_10843,N_10275,N_10079);
and U10844 (N_10844,N_10262,N_10201);
nor U10845 (N_10845,N_9953,N_9955);
xnor U10846 (N_10846,N_10495,N_10297);
nand U10847 (N_10847,N_10137,N_10205);
xor U10848 (N_10848,N_10218,N_10126);
and U10849 (N_10849,N_10055,N_10053);
and U10850 (N_10850,N_10222,N_10341);
nand U10851 (N_10851,N_10267,N_9917);
nand U10852 (N_10852,N_10460,N_10035);
nor U10853 (N_10853,N_9870,N_10154);
nor U10854 (N_10854,N_10486,N_10249);
or U10855 (N_10855,N_9836,N_10171);
nor U10856 (N_10856,N_9810,N_10358);
or U10857 (N_10857,N_9790,N_10401);
xnor U10858 (N_10858,N_9981,N_10319);
or U10859 (N_10859,N_9884,N_10178);
nor U10860 (N_10860,N_10214,N_10110);
or U10861 (N_10861,N_9769,N_10405);
xnor U10862 (N_10862,N_10330,N_10061);
or U10863 (N_10863,N_10018,N_9771);
xnor U10864 (N_10864,N_9952,N_10430);
nand U10865 (N_10865,N_9888,N_10193);
nor U10866 (N_10866,N_9968,N_9885);
and U10867 (N_10867,N_10063,N_10005);
and U10868 (N_10868,N_10352,N_10351);
or U10869 (N_10869,N_9869,N_10493);
and U10870 (N_10870,N_10213,N_10163);
nand U10871 (N_10871,N_10190,N_10303);
nor U10872 (N_10872,N_9962,N_9801);
and U10873 (N_10873,N_9753,N_9799);
nand U10874 (N_10874,N_10379,N_10013);
and U10875 (N_10875,N_9910,N_10493);
nand U10876 (N_10876,N_9837,N_9847);
nor U10877 (N_10877,N_9764,N_10296);
nor U10878 (N_10878,N_10085,N_10149);
or U10879 (N_10879,N_9881,N_10360);
nor U10880 (N_10880,N_10147,N_9795);
nand U10881 (N_10881,N_9857,N_9792);
xnor U10882 (N_10882,N_10303,N_10231);
nand U10883 (N_10883,N_9972,N_10312);
or U10884 (N_10884,N_9916,N_10154);
nand U10885 (N_10885,N_10434,N_10110);
and U10886 (N_10886,N_10409,N_10280);
and U10887 (N_10887,N_9966,N_9789);
nand U10888 (N_10888,N_10163,N_10054);
and U10889 (N_10889,N_10029,N_10464);
nand U10890 (N_10890,N_9987,N_10405);
xnor U10891 (N_10891,N_9974,N_9897);
xnor U10892 (N_10892,N_9993,N_10436);
nand U10893 (N_10893,N_10007,N_10147);
nor U10894 (N_10894,N_10378,N_10167);
nor U10895 (N_10895,N_10352,N_9968);
xor U10896 (N_10896,N_9836,N_9929);
xnor U10897 (N_10897,N_10453,N_9843);
nor U10898 (N_10898,N_10243,N_9867);
nor U10899 (N_10899,N_9831,N_10140);
or U10900 (N_10900,N_9933,N_9955);
nand U10901 (N_10901,N_10472,N_10440);
nor U10902 (N_10902,N_10059,N_10275);
and U10903 (N_10903,N_9896,N_9873);
nor U10904 (N_10904,N_10421,N_9861);
and U10905 (N_10905,N_9826,N_9898);
and U10906 (N_10906,N_10453,N_10263);
nor U10907 (N_10907,N_10297,N_9835);
nor U10908 (N_10908,N_9885,N_10213);
and U10909 (N_10909,N_9894,N_10412);
or U10910 (N_10910,N_10189,N_9959);
and U10911 (N_10911,N_10239,N_10317);
xor U10912 (N_10912,N_10376,N_10151);
and U10913 (N_10913,N_10042,N_10273);
or U10914 (N_10914,N_10260,N_9955);
and U10915 (N_10915,N_9916,N_10435);
nor U10916 (N_10916,N_9842,N_10224);
nor U10917 (N_10917,N_10011,N_10113);
or U10918 (N_10918,N_9946,N_10292);
nand U10919 (N_10919,N_10465,N_10337);
nor U10920 (N_10920,N_9922,N_10342);
and U10921 (N_10921,N_10347,N_10314);
nand U10922 (N_10922,N_10066,N_9944);
and U10923 (N_10923,N_10090,N_9808);
or U10924 (N_10924,N_10350,N_10100);
or U10925 (N_10925,N_10035,N_9780);
nand U10926 (N_10926,N_9886,N_10360);
nor U10927 (N_10927,N_10411,N_10239);
nand U10928 (N_10928,N_10359,N_10494);
and U10929 (N_10929,N_9765,N_10102);
nor U10930 (N_10930,N_9831,N_10122);
nor U10931 (N_10931,N_9771,N_10029);
xnor U10932 (N_10932,N_10339,N_10358);
xnor U10933 (N_10933,N_10493,N_10319);
and U10934 (N_10934,N_10442,N_9976);
nor U10935 (N_10935,N_9754,N_9769);
xor U10936 (N_10936,N_10291,N_10470);
xnor U10937 (N_10937,N_10110,N_9836);
nor U10938 (N_10938,N_10082,N_9978);
or U10939 (N_10939,N_9997,N_9773);
xnor U10940 (N_10940,N_9820,N_10135);
nor U10941 (N_10941,N_10466,N_9753);
or U10942 (N_10942,N_10031,N_9963);
nand U10943 (N_10943,N_10409,N_10249);
and U10944 (N_10944,N_9915,N_10192);
and U10945 (N_10945,N_10106,N_10080);
nand U10946 (N_10946,N_10012,N_10411);
or U10947 (N_10947,N_10065,N_10218);
nor U10948 (N_10948,N_10355,N_10372);
and U10949 (N_10949,N_10428,N_10338);
or U10950 (N_10950,N_10296,N_10223);
nor U10951 (N_10951,N_9924,N_10303);
xor U10952 (N_10952,N_10261,N_10413);
and U10953 (N_10953,N_9943,N_10226);
and U10954 (N_10954,N_10325,N_9924);
nand U10955 (N_10955,N_10162,N_9979);
nand U10956 (N_10956,N_10393,N_10278);
nand U10957 (N_10957,N_10469,N_10266);
nor U10958 (N_10958,N_10408,N_10454);
and U10959 (N_10959,N_10071,N_9962);
and U10960 (N_10960,N_10161,N_10406);
xnor U10961 (N_10961,N_9807,N_10158);
and U10962 (N_10962,N_10471,N_10143);
nor U10963 (N_10963,N_10211,N_10339);
or U10964 (N_10964,N_9771,N_10325);
nor U10965 (N_10965,N_10313,N_9799);
or U10966 (N_10966,N_10260,N_10238);
or U10967 (N_10967,N_10084,N_10264);
and U10968 (N_10968,N_10083,N_10403);
and U10969 (N_10969,N_10241,N_10284);
nand U10970 (N_10970,N_10465,N_10167);
nand U10971 (N_10971,N_10030,N_10308);
nor U10972 (N_10972,N_10308,N_9755);
nor U10973 (N_10973,N_9861,N_10447);
nand U10974 (N_10974,N_9789,N_10086);
and U10975 (N_10975,N_9979,N_10488);
or U10976 (N_10976,N_10101,N_10164);
xnor U10977 (N_10977,N_10320,N_10214);
nand U10978 (N_10978,N_9884,N_10099);
nand U10979 (N_10979,N_10239,N_9918);
or U10980 (N_10980,N_10343,N_10244);
nor U10981 (N_10981,N_9951,N_9754);
xnor U10982 (N_10982,N_10161,N_10261);
and U10983 (N_10983,N_10188,N_9884);
and U10984 (N_10984,N_10344,N_10466);
nor U10985 (N_10985,N_10294,N_10416);
or U10986 (N_10986,N_10171,N_10231);
nor U10987 (N_10987,N_10242,N_10306);
nor U10988 (N_10988,N_9852,N_10021);
nor U10989 (N_10989,N_10489,N_10429);
or U10990 (N_10990,N_10251,N_10452);
xor U10991 (N_10991,N_10011,N_10396);
nand U10992 (N_10992,N_10143,N_10013);
or U10993 (N_10993,N_9908,N_10434);
or U10994 (N_10994,N_9980,N_10001);
or U10995 (N_10995,N_10271,N_9880);
nor U10996 (N_10996,N_9774,N_9800);
nor U10997 (N_10997,N_10100,N_10407);
or U10998 (N_10998,N_9829,N_10168);
nor U10999 (N_10999,N_9823,N_9959);
nand U11000 (N_11000,N_9784,N_10017);
and U11001 (N_11001,N_9772,N_10225);
xnor U11002 (N_11002,N_9960,N_10046);
and U11003 (N_11003,N_9876,N_10204);
nor U11004 (N_11004,N_9931,N_10054);
nor U11005 (N_11005,N_9936,N_10444);
or U11006 (N_11006,N_10061,N_9972);
or U11007 (N_11007,N_10277,N_9994);
and U11008 (N_11008,N_10121,N_10374);
nor U11009 (N_11009,N_10005,N_10067);
nor U11010 (N_11010,N_10443,N_9869);
xnor U11011 (N_11011,N_10041,N_10264);
xor U11012 (N_11012,N_10173,N_10066);
and U11013 (N_11013,N_10485,N_10133);
and U11014 (N_11014,N_9798,N_10369);
or U11015 (N_11015,N_10252,N_10216);
nor U11016 (N_11016,N_10168,N_9794);
or U11017 (N_11017,N_9961,N_10421);
nand U11018 (N_11018,N_9949,N_9821);
or U11019 (N_11019,N_10339,N_10219);
nor U11020 (N_11020,N_10318,N_10081);
and U11021 (N_11021,N_9975,N_10064);
xnor U11022 (N_11022,N_9878,N_10197);
or U11023 (N_11023,N_10467,N_10243);
and U11024 (N_11024,N_10141,N_10358);
and U11025 (N_11025,N_10392,N_10408);
xnor U11026 (N_11026,N_10201,N_10061);
nor U11027 (N_11027,N_10330,N_10315);
nand U11028 (N_11028,N_10405,N_9816);
nand U11029 (N_11029,N_9982,N_9763);
xnor U11030 (N_11030,N_9942,N_9754);
nand U11031 (N_11031,N_10195,N_9990);
and U11032 (N_11032,N_10281,N_10497);
or U11033 (N_11033,N_9899,N_10412);
xnor U11034 (N_11034,N_9932,N_10082);
xor U11035 (N_11035,N_10413,N_10291);
xor U11036 (N_11036,N_10388,N_10399);
and U11037 (N_11037,N_9933,N_9805);
xor U11038 (N_11038,N_10172,N_10461);
xnor U11039 (N_11039,N_10424,N_10318);
or U11040 (N_11040,N_9907,N_9804);
nor U11041 (N_11041,N_9854,N_9774);
nor U11042 (N_11042,N_9789,N_9756);
nor U11043 (N_11043,N_10138,N_10349);
xnor U11044 (N_11044,N_9886,N_10178);
and U11045 (N_11045,N_10264,N_10464);
or U11046 (N_11046,N_9942,N_10362);
and U11047 (N_11047,N_9877,N_10176);
nor U11048 (N_11048,N_10042,N_10023);
xor U11049 (N_11049,N_10195,N_9757);
or U11050 (N_11050,N_10423,N_9772);
or U11051 (N_11051,N_10044,N_9950);
nand U11052 (N_11052,N_10390,N_9966);
and U11053 (N_11053,N_10086,N_10292);
or U11054 (N_11054,N_9847,N_9994);
xor U11055 (N_11055,N_10290,N_10155);
xor U11056 (N_11056,N_10381,N_9843);
and U11057 (N_11057,N_10380,N_10106);
or U11058 (N_11058,N_10387,N_9844);
nor U11059 (N_11059,N_9763,N_9852);
or U11060 (N_11060,N_10171,N_10304);
and U11061 (N_11061,N_9907,N_10038);
nand U11062 (N_11062,N_9959,N_10039);
nor U11063 (N_11063,N_10422,N_9932);
nand U11064 (N_11064,N_10491,N_10183);
or U11065 (N_11065,N_9994,N_9767);
and U11066 (N_11066,N_9859,N_10171);
xor U11067 (N_11067,N_9832,N_10383);
and U11068 (N_11068,N_10062,N_9825);
nor U11069 (N_11069,N_10078,N_10235);
nor U11070 (N_11070,N_10497,N_10229);
or U11071 (N_11071,N_9810,N_10124);
nor U11072 (N_11072,N_9976,N_10197);
or U11073 (N_11073,N_10374,N_9845);
and U11074 (N_11074,N_9856,N_9919);
or U11075 (N_11075,N_10215,N_9832);
or U11076 (N_11076,N_10351,N_10470);
xor U11077 (N_11077,N_10264,N_10403);
and U11078 (N_11078,N_10170,N_10426);
or U11079 (N_11079,N_10002,N_10268);
xor U11080 (N_11080,N_10063,N_9916);
or U11081 (N_11081,N_10000,N_9900);
xnor U11082 (N_11082,N_9926,N_10157);
and U11083 (N_11083,N_9784,N_9816);
or U11084 (N_11084,N_10290,N_10394);
xor U11085 (N_11085,N_10346,N_10248);
and U11086 (N_11086,N_10067,N_9980);
nand U11087 (N_11087,N_10032,N_10061);
nor U11088 (N_11088,N_10060,N_9832);
nor U11089 (N_11089,N_9946,N_9951);
and U11090 (N_11090,N_10429,N_10245);
nor U11091 (N_11091,N_9974,N_10471);
nor U11092 (N_11092,N_9975,N_9795);
nor U11093 (N_11093,N_10022,N_9789);
nand U11094 (N_11094,N_10047,N_10192);
xnor U11095 (N_11095,N_10346,N_10094);
xor U11096 (N_11096,N_9956,N_10443);
nand U11097 (N_11097,N_10297,N_9760);
or U11098 (N_11098,N_9869,N_10145);
xnor U11099 (N_11099,N_10041,N_9965);
nor U11100 (N_11100,N_10313,N_9932);
xnor U11101 (N_11101,N_9971,N_9789);
or U11102 (N_11102,N_10140,N_10100);
xor U11103 (N_11103,N_10060,N_10059);
nor U11104 (N_11104,N_10088,N_9935);
nor U11105 (N_11105,N_9827,N_10102);
nor U11106 (N_11106,N_9806,N_10144);
or U11107 (N_11107,N_9826,N_10228);
nand U11108 (N_11108,N_10382,N_10354);
and U11109 (N_11109,N_9970,N_10011);
and U11110 (N_11110,N_9982,N_10069);
and U11111 (N_11111,N_9754,N_10243);
nand U11112 (N_11112,N_10043,N_10179);
nor U11113 (N_11113,N_9953,N_10488);
nand U11114 (N_11114,N_10323,N_10040);
nor U11115 (N_11115,N_10001,N_10047);
and U11116 (N_11116,N_9777,N_9847);
xor U11117 (N_11117,N_10057,N_9966);
or U11118 (N_11118,N_10096,N_9817);
and U11119 (N_11119,N_10277,N_10407);
nand U11120 (N_11120,N_10112,N_10230);
xnor U11121 (N_11121,N_9972,N_9943);
nor U11122 (N_11122,N_9906,N_10234);
xor U11123 (N_11123,N_9920,N_10387);
or U11124 (N_11124,N_9977,N_10411);
and U11125 (N_11125,N_9791,N_9880);
xor U11126 (N_11126,N_10410,N_9870);
nor U11127 (N_11127,N_9917,N_10178);
or U11128 (N_11128,N_10186,N_10376);
and U11129 (N_11129,N_9857,N_10224);
or U11130 (N_11130,N_10431,N_10164);
and U11131 (N_11131,N_10275,N_10237);
xor U11132 (N_11132,N_9895,N_10453);
nor U11133 (N_11133,N_10431,N_9970);
nor U11134 (N_11134,N_10010,N_10334);
xnor U11135 (N_11135,N_10051,N_9804);
nor U11136 (N_11136,N_9802,N_10133);
nand U11137 (N_11137,N_10343,N_10039);
nor U11138 (N_11138,N_9994,N_10492);
nor U11139 (N_11139,N_10163,N_10010);
or U11140 (N_11140,N_9962,N_10110);
xor U11141 (N_11141,N_9785,N_9954);
xor U11142 (N_11142,N_10424,N_9757);
xnor U11143 (N_11143,N_10203,N_10112);
and U11144 (N_11144,N_10207,N_9809);
nand U11145 (N_11145,N_9883,N_10016);
nand U11146 (N_11146,N_10410,N_10222);
xor U11147 (N_11147,N_9999,N_10400);
xor U11148 (N_11148,N_9949,N_9987);
or U11149 (N_11149,N_9751,N_9942);
xor U11150 (N_11150,N_10492,N_10109);
or U11151 (N_11151,N_10020,N_9915);
and U11152 (N_11152,N_10130,N_9869);
or U11153 (N_11153,N_10101,N_10341);
xnor U11154 (N_11154,N_10189,N_10378);
xor U11155 (N_11155,N_10057,N_10162);
or U11156 (N_11156,N_9950,N_9761);
or U11157 (N_11157,N_10230,N_9770);
xor U11158 (N_11158,N_10180,N_10438);
nor U11159 (N_11159,N_10074,N_9867);
nor U11160 (N_11160,N_9941,N_10445);
or U11161 (N_11161,N_10358,N_9877);
nand U11162 (N_11162,N_10365,N_10201);
xor U11163 (N_11163,N_10352,N_10175);
or U11164 (N_11164,N_10477,N_10120);
xor U11165 (N_11165,N_9824,N_9772);
and U11166 (N_11166,N_10408,N_10422);
xnor U11167 (N_11167,N_10048,N_9909);
nor U11168 (N_11168,N_9987,N_9846);
nor U11169 (N_11169,N_10131,N_9959);
xnor U11170 (N_11170,N_10205,N_10209);
nor U11171 (N_11171,N_10000,N_10430);
or U11172 (N_11172,N_10194,N_10079);
nor U11173 (N_11173,N_9771,N_10279);
nand U11174 (N_11174,N_9812,N_10125);
nand U11175 (N_11175,N_10413,N_10001);
and U11176 (N_11176,N_10148,N_10117);
xnor U11177 (N_11177,N_9849,N_10031);
or U11178 (N_11178,N_10030,N_9894);
nand U11179 (N_11179,N_9785,N_10368);
nor U11180 (N_11180,N_10033,N_9997);
nand U11181 (N_11181,N_10046,N_10466);
and U11182 (N_11182,N_10360,N_10103);
or U11183 (N_11183,N_10193,N_10326);
nor U11184 (N_11184,N_9935,N_10168);
and U11185 (N_11185,N_10467,N_9925);
nor U11186 (N_11186,N_10409,N_9966);
nor U11187 (N_11187,N_9887,N_9938);
nand U11188 (N_11188,N_10079,N_10443);
nand U11189 (N_11189,N_10133,N_9816);
nor U11190 (N_11190,N_10165,N_10482);
or U11191 (N_11191,N_10253,N_9894);
nor U11192 (N_11192,N_10256,N_10202);
or U11193 (N_11193,N_9861,N_9953);
nor U11194 (N_11194,N_9773,N_10492);
or U11195 (N_11195,N_10053,N_10059);
nor U11196 (N_11196,N_10044,N_10293);
xor U11197 (N_11197,N_10189,N_10418);
nor U11198 (N_11198,N_10082,N_10441);
nor U11199 (N_11199,N_9858,N_10044);
nor U11200 (N_11200,N_9898,N_10392);
xor U11201 (N_11201,N_9890,N_10091);
or U11202 (N_11202,N_10200,N_9786);
xnor U11203 (N_11203,N_10106,N_9805);
or U11204 (N_11204,N_9858,N_10472);
and U11205 (N_11205,N_9773,N_9826);
nor U11206 (N_11206,N_10376,N_10374);
xor U11207 (N_11207,N_9906,N_10340);
xnor U11208 (N_11208,N_10389,N_9857);
or U11209 (N_11209,N_10317,N_10120);
nand U11210 (N_11210,N_9900,N_10049);
nand U11211 (N_11211,N_10023,N_10196);
nand U11212 (N_11212,N_10298,N_10222);
nand U11213 (N_11213,N_9800,N_10049);
and U11214 (N_11214,N_10272,N_10415);
and U11215 (N_11215,N_10470,N_10215);
and U11216 (N_11216,N_10006,N_10038);
or U11217 (N_11217,N_10395,N_10069);
nand U11218 (N_11218,N_10224,N_10380);
nor U11219 (N_11219,N_10455,N_9984);
and U11220 (N_11220,N_10442,N_9962);
nand U11221 (N_11221,N_10189,N_10260);
and U11222 (N_11222,N_10076,N_10323);
nor U11223 (N_11223,N_10128,N_9967);
nand U11224 (N_11224,N_10399,N_9930);
nand U11225 (N_11225,N_10244,N_10370);
nor U11226 (N_11226,N_10317,N_10178);
xor U11227 (N_11227,N_10319,N_9908);
xor U11228 (N_11228,N_10014,N_10038);
nor U11229 (N_11229,N_9753,N_9925);
nand U11230 (N_11230,N_10424,N_9858);
or U11231 (N_11231,N_10226,N_10031);
and U11232 (N_11232,N_10418,N_9801);
or U11233 (N_11233,N_9904,N_9844);
nor U11234 (N_11234,N_10288,N_9769);
nand U11235 (N_11235,N_9984,N_10329);
nor U11236 (N_11236,N_10120,N_10461);
and U11237 (N_11237,N_10080,N_10126);
nor U11238 (N_11238,N_10141,N_10227);
nand U11239 (N_11239,N_9802,N_10002);
nor U11240 (N_11240,N_9871,N_10398);
and U11241 (N_11241,N_10307,N_10139);
and U11242 (N_11242,N_10457,N_10310);
and U11243 (N_11243,N_10396,N_10268);
or U11244 (N_11244,N_10320,N_9880);
nor U11245 (N_11245,N_10015,N_9756);
nand U11246 (N_11246,N_10141,N_9788);
nand U11247 (N_11247,N_10314,N_10082);
nor U11248 (N_11248,N_9786,N_10442);
nor U11249 (N_11249,N_10017,N_9908);
nor U11250 (N_11250,N_10665,N_11083);
and U11251 (N_11251,N_10944,N_11114);
or U11252 (N_11252,N_10997,N_10788);
or U11253 (N_11253,N_10830,N_10890);
or U11254 (N_11254,N_10948,N_11118);
xor U11255 (N_11255,N_10821,N_10990);
or U11256 (N_11256,N_10770,N_10529);
and U11257 (N_11257,N_10612,N_10886);
or U11258 (N_11258,N_10701,N_10561);
nand U11259 (N_11259,N_10909,N_10924);
nand U11260 (N_11260,N_10978,N_10740);
or U11261 (N_11261,N_10777,N_11033);
xor U11262 (N_11262,N_10863,N_10992);
and U11263 (N_11263,N_10522,N_10689);
nor U11264 (N_11264,N_11106,N_10707);
or U11265 (N_11265,N_11010,N_11075);
and U11266 (N_11266,N_10706,N_10817);
nor U11267 (N_11267,N_11037,N_10624);
or U11268 (N_11268,N_10808,N_10754);
and U11269 (N_11269,N_10648,N_10938);
or U11270 (N_11270,N_11188,N_10858);
or U11271 (N_11271,N_10542,N_10799);
and U11272 (N_11272,N_10585,N_11042);
xnor U11273 (N_11273,N_11204,N_11101);
nand U11274 (N_11274,N_10703,N_10669);
and U11275 (N_11275,N_11052,N_11142);
nor U11276 (N_11276,N_10818,N_10537);
and U11277 (N_11277,N_11121,N_10608);
xor U11278 (N_11278,N_10932,N_11243);
xor U11279 (N_11279,N_10991,N_10575);
nand U11280 (N_11280,N_10719,N_10599);
nor U11281 (N_11281,N_10763,N_11181);
nor U11282 (N_11282,N_10896,N_10828);
or U11283 (N_11283,N_10617,N_11191);
xnor U11284 (N_11284,N_10778,N_10766);
and U11285 (N_11285,N_11081,N_11129);
or U11286 (N_11286,N_10792,N_11195);
or U11287 (N_11287,N_10743,N_10979);
nor U11288 (N_11288,N_10996,N_10839);
xor U11289 (N_11289,N_11066,N_11143);
nand U11290 (N_11290,N_10520,N_10903);
xnor U11291 (N_11291,N_10510,N_11125);
nor U11292 (N_11292,N_10543,N_10810);
nor U11293 (N_11293,N_10524,N_11079);
xnor U11294 (N_11294,N_10551,N_10836);
nand U11295 (N_11295,N_10637,N_11094);
nor U11296 (N_11296,N_11110,N_10692);
and U11297 (N_11297,N_10729,N_11043);
nand U11298 (N_11298,N_11124,N_11225);
xor U11299 (N_11299,N_11161,N_10962);
nor U11300 (N_11300,N_11002,N_10586);
nor U11301 (N_11301,N_10718,N_10774);
nor U11302 (N_11302,N_10658,N_10872);
nor U11303 (N_11303,N_10564,N_11004);
xnor U11304 (N_11304,N_10732,N_11148);
or U11305 (N_11305,N_11227,N_10627);
and U11306 (N_11306,N_10713,N_11202);
or U11307 (N_11307,N_10697,N_10682);
nor U11308 (N_11308,N_10712,N_11230);
or U11309 (N_11309,N_11153,N_10504);
xor U11310 (N_11310,N_11147,N_11130);
and U11311 (N_11311,N_10717,N_10789);
and U11312 (N_11312,N_10931,N_11067);
and U11313 (N_11313,N_11242,N_10755);
or U11314 (N_11314,N_10936,N_10738);
nand U11315 (N_11315,N_10734,N_10653);
and U11316 (N_11316,N_10654,N_11017);
xor U11317 (N_11317,N_10640,N_11011);
nand U11318 (N_11318,N_10906,N_11013);
or U11319 (N_11319,N_10593,N_10678);
nand U11320 (N_11320,N_10780,N_10993);
nand U11321 (N_11321,N_10860,N_10984);
or U11322 (N_11322,N_11201,N_10814);
nor U11323 (N_11323,N_11208,N_11123);
and U11324 (N_11324,N_10735,N_10911);
nand U11325 (N_11325,N_10570,N_11203);
xor U11326 (N_11326,N_11064,N_10843);
and U11327 (N_11327,N_10917,N_11117);
or U11328 (N_11328,N_10771,N_10609);
and U11329 (N_11329,N_11175,N_11174);
nand U11330 (N_11330,N_11077,N_10667);
and U11331 (N_11331,N_11249,N_11172);
xnor U11332 (N_11332,N_11109,N_11169);
or U11333 (N_11333,N_10753,N_10871);
or U11334 (N_11334,N_11080,N_10604);
and U11335 (N_11335,N_10832,N_11107);
and U11336 (N_11336,N_10711,N_10968);
xnor U11337 (N_11337,N_10566,N_10567);
xor U11338 (N_11338,N_10534,N_11054);
and U11339 (N_11339,N_11116,N_10927);
nand U11340 (N_11340,N_10518,N_10698);
nor U11341 (N_11341,N_10869,N_11163);
xnor U11342 (N_11342,N_10574,N_10532);
nand U11343 (N_11343,N_10602,N_11138);
xnor U11344 (N_11344,N_10904,N_10730);
or U11345 (N_11345,N_11089,N_10633);
or U11346 (N_11346,N_10824,N_10761);
xnor U11347 (N_11347,N_11157,N_10866);
nand U11348 (N_11348,N_10555,N_10623);
and U11349 (N_11349,N_11196,N_10864);
nor U11350 (N_11350,N_11218,N_10922);
nand U11351 (N_11351,N_11132,N_10807);
and U11352 (N_11352,N_11084,N_10894);
or U11353 (N_11353,N_10538,N_10556);
nand U11354 (N_11354,N_11005,N_10893);
and U11355 (N_11355,N_10842,N_11165);
nor U11356 (N_11356,N_10680,N_11194);
xor U11357 (N_11357,N_11020,N_11179);
and U11358 (N_11358,N_11028,N_10649);
xnor U11359 (N_11359,N_10949,N_10723);
nor U11360 (N_11360,N_10583,N_11187);
nor U11361 (N_11361,N_10549,N_10565);
xnor U11362 (N_11362,N_10523,N_11058);
nand U11363 (N_11363,N_11168,N_11183);
or U11364 (N_11364,N_11093,N_10702);
xnor U11365 (N_11365,N_10796,N_10739);
nand U11366 (N_11366,N_11237,N_10884);
or U11367 (N_11367,N_10643,N_10577);
or U11368 (N_11368,N_11244,N_10889);
and U11369 (N_11369,N_10539,N_11245);
or U11370 (N_11370,N_10946,N_11222);
xor U11371 (N_11371,N_10600,N_10631);
xnor U11372 (N_11372,N_11087,N_10744);
and U11373 (N_11373,N_11006,N_10512);
or U11374 (N_11374,N_10785,N_10625);
nand U11375 (N_11375,N_10541,N_10913);
and U11376 (N_11376,N_10554,N_10614);
nor U11377 (N_11377,N_10562,N_10786);
xor U11378 (N_11378,N_10501,N_10651);
xor U11379 (N_11379,N_10725,N_10929);
nand U11380 (N_11380,N_11158,N_11149);
and U11381 (N_11381,N_10919,N_11205);
nand U11382 (N_11382,N_10868,N_11078);
and U11383 (N_11383,N_10550,N_11055);
and U11384 (N_11384,N_11247,N_10960);
xor U11385 (N_11385,N_10528,N_10705);
or U11386 (N_11386,N_10751,N_10772);
nor U11387 (N_11387,N_10581,N_10989);
nand U11388 (N_11388,N_11217,N_10519);
nor U11389 (N_11389,N_11056,N_10629);
and U11390 (N_11390,N_10969,N_10974);
and U11391 (N_11391,N_10937,N_11051);
xor U11392 (N_11392,N_10910,N_10831);
xnor U11393 (N_11393,N_10632,N_10745);
xor U11394 (N_11394,N_10662,N_11214);
or U11395 (N_11395,N_10742,N_11088);
nor U11396 (N_11396,N_10521,N_11212);
nor U11397 (N_11397,N_10673,N_11145);
nor U11398 (N_11398,N_10835,N_11224);
or U11399 (N_11399,N_10659,N_10731);
and U11400 (N_11400,N_11009,N_10657);
xnor U11401 (N_11401,N_10797,N_11103);
nor U11402 (N_11402,N_10897,N_10964);
and U11403 (N_11403,N_11197,N_10722);
and U11404 (N_11404,N_11238,N_10784);
xnor U11405 (N_11405,N_10597,N_11156);
nor U11406 (N_11406,N_10582,N_10876);
or U11407 (N_11407,N_10620,N_10900);
nand U11408 (N_11408,N_11008,N_10694);
nor U11409 (N_11409,N_11039,N_10733);
xor U11410 (N_11410,N_10656,N_10918);
nor U11411 (N_11411,N_10502,N_11029);
xor U11412 (N_11412,N_10768,N_10601);
nand U11413 (N_11413,N_11231,N_10645);
and U11414 (N_11414,N_10916,N_10857);
and U11415 (N_11415,N_10811,N_11131);
and U11416 (N_11416,N_10973,N_11198);
and U11417 (N_11417,N_10795,N_11108);
or U11418 (N_11418,N_10802,N_10957);
xnor U11419 (N_11419,N_11137,N_10880);
nor U11420 (N_11420,N_11085,N_11105);
or U11421 (N_11421,N_10700,N_10563);
or U11422 (N_11422,N_10813,N_10545);
and U11423 (N_11423,N_10767,N_11233);
xor U11424 (N_11424,N_10558,N_10812);
nor U11425 (N_11425,N_11022,N_11192);
nor U11426 (N_11426,N_11032,N_10675);
or U11427 (N_11427,N_10681,N_10741);
and U11428 (N_11428,N_10677,N_11152);
and U11429 (N_11429,N_10513,N_10769);
nor U11430 (N_11430,N_11026,N_10588);
nand U11431 (N_11431,N_10580,N_10547);
or U11432 (N_11432,N_10695,N_10639);
nor U11433 (N_11433,N_10605,N_10569);
or U11434 (N_11434,N_10888,N_10899);
nor U11435 (N_11435,N_10652,N_11049);
nor U11436 (N_11436,N_10848,N_10995);
xor U11437 (N_11437,N_10686,N_10933);
nand U11438 (N_11438,N_11070,N_10934);
nand U11439 (N_11439,N_11047,N_10972);
nand U11440 (N_11440,N_11090,N_10572);
and U11441 (N_11441,N_10816,N_10533);
or U11442 (N_11442,N_11035,N_10947);
or U11443 (N_11443,N_11021,N_10939);
nand U11444 (N_11444,N_11061,N_10553);
nor U11445 (N_11445,N_10514,N_11228);
nor U11446 (N_11446,N_10970,N_10619);
and U11447 (N_11447,N_11177,N_10829);
or U11448 (N_11448,N_10750,N_10596);
and U11449 (N_11449,N_10925,N_10546);
nand U11450 (N_11450,N_10515,N_10994);
and U11451 (N_11451,N_11193,N_10980);
nand U11452 (N_11452,N_10950,N_10966);
nor U11453 (N_11453,N_10663,N_11031);
xnor U11454 (N_11454,N_11003,N_10676);
xnor U11455 (N_11455,N_11189,N_10881);
or U11456 (N_11456,N_10636,N_11007);
nand U11457 (N_11457,N_10806,N_10887);
or U11458 (N_11458,N_10591,N_11164);
or U11459 (N_11459,N_10527,N_10958);
and U11460 (N_11460,N_11068,N_10727);
xnor U11461 (N_11461,N_11232,N_10650);
or U11462 (N_11462,N_10794,N_10775);
nor U11463 (N_11463,N_10671,N_10668);
and U11464 (N_11464,N_10940,N_11014);
or U11465 (N_11465,N_10737,N_10613);
nand U11466 (N_11466,N_10759,N_10517);
or U11467 (N_11467,N_10781,N_10862);
xnor U11468 (N_11468,N_10757,N_10954);
nand U11469 (N_11469,N_10846,N_11016);
or U11470 (N_11470,N_10891,N_11234);
or U11471 (N_11471,N_10809,N_10976);
or U11472 (N_11472,N_11173,N_11122);
and U11473 (N_11473,N_11045,N_10660);
and U11474 (N_11474,N_10760,N_10559);
or U11475 (N_11475,N_10756,N_11166);
or U11476 (N_11476,N_10953,N_10883);
nor U11477 (N_11477,N_11178,N_10672);
and U11478 (N_11478,N_11199,N_11119);
xnor U11479 (N_11479,N_11115,N_10699);
nand U11480 (N_11480,N_10815,N_10849);
and U11481 (N_11481,N_10710,N_10837);
and U11482 (N_11482,N_10595,N_10762);
nor U11483 (N_11483,N_10961,N_10507);
nand U11484 (N_11484,N_10803,N_11159);
nand U11485 (N_11485,N_10838,N_11040);
xnor U11486 (N_11486,N_11057,N_10622);
nand U11487 (N_11487,N_11112,N_10804);
nand U11488 (N_11488,N_11113,N_11018);
and U11489 (N_11489,N_10854,N_10509);
or U11490 (N_11490,N_10721,N_11207);
nand U11491 (N_11491,N_10847,N_10870);
or U11492 (N_11492,N_11099,N_11190);
xor U11493 (N_11493,N_11133,N_10758);
and U11494 (N_11494,N_10536,N_10877);
nand U11495 (N_11495,N_10915,N_10967);
nand U11496 (N_11496,N_10661,N_11160);
nor U11497 (N_11497,N_11001,N_10971);
nor U11498 (N_11498,N_10747,N_10607);
nor U11499 (N_11499,N_11206,N_10644);
or U11500 (N_11500,N_11226,N_10670);
xnor U11501 (N_11501,N_10749,N_10791);
xor U11502 (N_11502,N_10875,N_11030);
nand U11503 (N_11503,N_10895,N_11102);
or U11504 (N_11504,N_11211,N_10867);
and U11505 (N_11505,N_11246,N_10603);
xnor U11506 (N_11506,N_10798,N_10959);
xor U11507 (N_11507,N_11139,N_10505);
and U11508 (N_11508,N_11072,N_11210);
xor U11509 (N_11509,N_10560,N_11098);
and U11510 (N_11510,N_10679,N_10861);
nor U11511 (N_11511,N_10674,N_10827);
xor U11512 (N_11512,N_10845,N_10764);
or U11513 (N_11513,N_11126,N_10859);
xnor U11514 (N_11514,N_11053,N_11036);
and U11515 (N_11515,N_10982,N_10691);
nand U11516 (N_11516,N_10865,N_10508);
nand U11517 (N_11517,N_10610,N_10986);
nor U11518 (N_11518,N_10885,N_10587);
xor U11519 (N_11519,N_10882,N_10683);
nand U11520 (N_11520,N_11135,N_10955);
or U11521 (N_11521,N_10800,N_11136);
or U11522 (N_11522,N_10998,N_11182);
and U11523 (N_11523,N_11044,N_10664);
or U11524 (N_11524,N_10878,N_10557);
xor U11525 (N_11525,N_10655,N_10914);
nor U11526 (N_11526,N_10855,N_10535);
nand U11527 (N_11527,N_10942,N_11151);
xnor U11528 (N_11528,N_11091,N_11180);
or U11529 (N_11529,N_10898,N_10983);
or U11530 (N_11530,N_10590,N_10779);
or U11531 (N_11531,N_11041,N_11074);
or U11532 (N_11532,N_10615,N_11027);
nor U11533 (N_11533,N_10500,N_10526);
xnor U11534 (N_11534,N_10975,N_10988);
and U11535 (N_11535,N_10641,N_10840);
xor U11536 (N_11536,N_11071,N_11176);
xnor U11537 (N_11537,N_10684,N_10685);
or U11538 (N_11538,N_11241,N_10908);
nor U11539 (N_11539,N_11186,N_10985);
nor U11540 (N_11540,N_10726,N_11162);
nor U11541 (N_11541,N_11063,N_10920);
nor U11542 (N_11542,N_10856,N_10576);
nand U11543 (N_11543,N_10606,N_10621);
or U11544 (N_11544,N_11097,N_10912);
nand U11545 (N_11545,N_11248,N_11155);
and U11546 (N_11546,N_10787,N_11086);
nand U11547 (N_11547,N_10571,N_10724);
nand U11548 (N_11548,N_10977,N_10822);
nor U11549 (N_11549,N_10635,N_11216);
xnor U11550 (N_11550,N_11171,N_10573);
nand U11551 (N_11551,N_11034,N_10965);
nor U11552 (N_11552,N_10951,N_10765);
and U11553 (N_11553,N_10584,N_11069);
or U11554 (N_11554,N_11000,N_11221);
and U11555 (N_11555,N_11185,N_10525);
nor U11556 (N_11556,N_10752,N_11048);
nor U11557 (N_11557,N_11170,N_11120);
xor U11558 (N_11558,N_10708,N_10943);
or U11559 (N_11559,N_10825,N_10928);
nand U11560 (N_11560,N_10935,N_10999);
xnor U11561 (N_11561,N_11060,N_10793);
and U11562 (N_11562,N_11015,N_10823);
and U11563 (N_11563,N_10592,N_10696);
and U11564 (N_11564,N_10892,N_11236);
or U11565 (N_11565,N_10941,N_10850);
xnor U11566 (N_11566,N_10748,N_10981);
nor U11567 (N_11567,N_11046,N_10626);
nand U11568 (N_11568,N_10544,N_10568);
nor U11569 (N_11569,N_10851,N_10616);
nor U11570 (N_11570,N_11023,N_11140);
and U11571 (N_11571,N_10618,N_11141);
nand U11572 (N_11572,N_10782,N_11100);
or U11573 (N_11573,N_11082,N_11220);
nand U11574 (N_11574,N_10728,N_10776);
and U11575 (N_11575,N_10819,N_10902);
xor U11576 (N_11576,N_10901,N_10714);
or U11577 (N_11577,N_10987,N_10746);
nor U11578 (N_11578,N_11229,N_10905);
nand U11579 (N_11579,N_10921,N_10790);
and U11580 (N_11580,N_11050,N_10853);
or U11581 (N_11581,N_10716,N_11127);
or U11582 (N_11582,N_10945,N_11213);
nor U11583 (N_11583,N_11184,N_10963);
or U11584 (N_11584,N_11134,N_10628);
nor U11585 (N_11585,N_11111,N_10956);
nand U11586 (N_11586,N_10548,N_10611);
or U11587 (N_11587,N_11062,N_10688);
and U11588 (N_11588,N_11025,N_10923);
xnor U11589 (N_11589,N_10736,N_11092);
nand U11590 (N_11590,N_11235,N_10834);
nand U11591 (N_11591,N_10634,N_10666);
and U11592 (N_11592,N_11012,N_10506);
or U11593 (N_11593,N_11095,N_10530);
nand U11594 (N_11594,N_10930,N_11019);
and U11595 (N_11595,N_11209,N_11065);
xor U11596 (N_11596,N_11239,N_11200);
or U11597 (N_11597,N_10579,N_11076);
and U11598 (N_11598,N_11073,N_11038);
xor U11599 (N_11599,N_10646,N_11059);
nor U11600 (N_11600,N_10704,N_10720);
or U11601 (N_11601,N_10594,N_10690);
and U11602 (N_11602,N_10826,N_10952);
or U11603 (N_11603,N_11024,N_10874);
nor U11604 (N_11604,N_10873,N_10578);
xor U11605 (N_11605,N_11240,N_10844);
nand U11606 (N_11606,N_10511,N_10820);
xor U11607 (N_11607,N_10805,N_10503);
nor U11608 (N_11608,N_10540,N_10589);
xnor U11609 (N_11609,N_10516,N_10841);
nor U11610 (N_11610,N_10642,N_10693);
xnor U11611 (N_11611,N_11096,N_11167);
nor U11612 (N_11612,N_11215,N_10531);
nand U11613 (N_11613,N_10687,N_11128);
nand U11614 (N_11614,N_10801,N_11154);
nor U11615 (N_11615,N_10715,N_10552);
nand U11616 (N_11616,N_10630,N_10907);
and U11617 (N_11617,N_10879,N_10833);
xor U11618 (N_11618,N_11146,N_10852);
and U11619 (N_11619,N_10638,N_10647);
and U11620 (N_11620,N_11219,N_10598);
and U11621 (N_11621,N_11144,N_10783);
xor U11622 (N_11622,N_11150,N_10709);
and U11623 (N_11623,N_10926,N_11223);
xor U11624 (N_11624,N_11104,N_10773);
and U11625 (N_11625,N_10831,N_11110);
nor U11626 (N_11626,N_10508,N_10628);
nand U11627 (N_11627,N_10790,N_10930);
xnor U11628 (N_11628,N_10506,N_11000);
or U11629 (N_11629,N_10764,N_11173);
nor U11630 (N_11630,N_10897,N_10672);
xor U11631 (N_11631,N_10678,N_10500);
nand U11632 (N_11632,N_10939,N_11006);
nand U11633 (N_11633,N_10535,N_11040);
and U11634 (N_11634,N_10959,N_11247);
nand U11635 (N_11635,N_10968,N_11121);
or U11636 (N_11636,N_10955,N_11083);
and U11637 (N_11637,N_11180,N_10978);
nand U11638 (N_11638,N_10809,N_11138);
nand U11639 (N_11639,N_10958,N_11110);
nor U11640 (N_11640,N_11197,N_10782);
nor U11641 (N_11641,N_11124,N_10720);
or U11642 (N_11642,N_10543,N_10741);
or U11643 (N_11643,N_10752,N_11116);
xnor U11644 (N_11644,N_10568,N_10832);
or U11645 (N_11645,N_10625,N_11204);
nor U11646 (N_11646,N_10937,N_10962);
or U11647 (N_11647,N_10788,N_10619);
and U11648 (N_11648,N_10593,N_10799);
and U11649 (N_11649,N_10896,N_10626);
and U11650 (N_11650,N_11125,N_10767);
nand U11651 (N_11651,N_10725,N_10894);
and U11652 (N_11652,N_10983,N_11002);
xnor U11653 (N_11653,N_10698,N_10545);
xor U11654 (N_11654,N_10520,N_10701);
nor U11655 (N_11655,N_10698,N_10759);
nand U11656 (N_11656,N_10752,N_11221);
nor U11657 (N_11657,N_11160,N_10767);
nor U11658 (N_11658,N_11172,N_10717);
nand U11659 (N_11659,N_10772,N_10824);
xor U11660 (N_11660,N_10931,N_10614);
nor U11661 (N_11661,N_11036,N_10508);
and U11662 (N_11662,N_11196,N_10588);
nor U11663 (N_11663,N_10543,N_11104);
nand U11664 (N_11664,N_10525,N_11177);
nor U11665 (N_11665,N_10839,N_10830);
or U11666 (N_11666,N_11161,N_10790);
nand U11667 (N_11667,N_10984,N_10818);
or U11668 (N_11668,N_10597,N_11226);
nand U11669 (N_11669,N_10950,N_10731);
nor U11670 (N_11670,N_10833,N_10664);
nand U11671 (N_11671,N_11028,N_10938);
nor U11672 (N_11672,N_11186,N_10833);
xor U11673 (N_11673,N_10504,N_10537);
xor U11674 (N_11674,N_10852,N_10685);
nand U11675 (N_11675,N_10592,N_10947);
nand U11676 (N_11676,N_11238,N_10985);
nor U11677 (N_11677,N_10804,N_10818);
xnor U11678 (N_11678,N_10663,N_10515);
or U11679 (N_11679,N_11100,N_10590);
xnor U11680 (N_11680,N_10692,N_10525);
and U11681 (N_11681,N_10548,N_10707);
nor U11682 (N_11682,N_10961,N_10524);
and U11683 (N_11683,N_10641,N_10697);
or U11684 (N_11684,N_11245,N_11188);
xnor U11685 (N_11685,N_11091,N_10630);
and U11686 (N_11686,N_10849,N_11022);
nor U11687 (N_11687,N_10570,N_10507);
or U11688 (N_11688,N_10812,N_11211);
or U11689 (N_11689,N_10615,N_11084);
nand U11690 (N_11690,N_10616,N_10994);
and U11691 (N_11691,N_11107,N_10683);
or U11692 (N_11692,N_10837,N_10972);
nor U11693 (N_11693,N_10618,N_10699);
and U11694 (N_11694,N_10738,N_10837);
and U11695 (N_11695,N_11061,N_10688);
and U11696 (N_11696,N_10925,N_10574);
nand U11697 (N_11697,N_11218,N_10587);
xnor U11698 (N_11698,N_11226,N_10842);
xnor U11699 (N_11699,N_10680,N_11165);
or U11700 (N_11700,N_11192,N_11054);
nand U11701 (N_11701,N_10924,N_11147);
or U11702 (N_11702,N_10780,N_11034);
and U11703 (N_11703,N_10691,N_10658);
and U11704 (N_11704,N_10881,N_11119);
nand U11705 (N_11705,N_11180,N_10827);
nor U11706 (N_11706,N_10924,N_11073);
xor U11707 (N_11707,N_11185,N_10825);
and U11708 (N_11708,N_10628,N_11177);
xnor U11709 (N_11709,N_11021,N_10569);
and U11710 (N_11710,N_11149,N_10500);
nor U11711 (N_11711,N_10594,N_10936);
xor U11712 (N_11712,N_10816,N_11149);
xor U11713 (N_11713,N_11120,N_10628);
nor U11714 (N_11714,N_10855,N_11150);
and U11715 (N_11715,N_10870,N_10814);
or U11716 (N_11716,N_11189,N_10877);
nand U11717 (N_11717,N_11014,N_11035);
nor U11718 (N_11718,N_10606,N_11050);
xor U11719 (N_11719,N_10965,N_11243);
nand U11720 (N_11720,N_10576,N_11053);
or U11721 (N_11721,N_11057,N_11065);
and U11722 (N_11722,N_10945,N_11022);
nor U11723 (N_11723,N_10885,N_10620);
and U11724 (N_11724,N_10591,N_10513);
nor U11725 (N_11725,N_10950,N_10573);
or U11726 (N_11726,N_10707,N_11241);
nor U11727 (N_11727,N_10867,N_11109);
or U11728 (N_11728,N_10596,N_10969);
and U11729 (N_11729,N_10732,N_11000);
or U11730 (N_11730,N_10889,N_10931);
nand U11731 (N_11731,N_10809,N_10624);
nand U11732 (N_11732,N_10831,N_11119);
and U11733 (N_11733,N_10935,N_11246);
or U11734 (N_11734,N_11133,N_10719);
nand U11735 (N_11735,N_11221,N_10787);
xnor U11736 (N_11736,N_10512,N_10528);
xnor U11737 (N_11737,N_10605,N_10774);
and U11738 (N_11738,N_10615,N_11152);
xnor U11739 (N_11739,N_11110,N_10641);
nand U11740 (N_11740,N_10503,N_10615);
or U11741 (N_11741,N_11017,N_10752);
or U11742 (N_11742,N_11124,N_10740);
nor U11743 (N_11743,N_10838,N_10998);
xor U11744 (N_11744,N_10660,N_11036);
xor U11745 (N_11745,N_10746,N_11154);
or U11746 (N_11746,N_10762,N_10574);
xnor U11747 (N_11747,N_10587,N_10941);
nor U11748 (N_11748,N_11227,N_10947);
or U11749 (N_11749,N_10756,N_10699);
xor U11750 (N_11750,N_10957,N_10547);
or U11751 (N_11751,N_10539,N_10603);
nor U11752 (N_11752,N_11199,N_10650);
and U11753 (N_11753,N_10705,N_10697);
or U11754 (N_11754,N_10879,N_10986);
or U11755 (N_11755,N_10611,N_10927);
xor U11756 (N_11756,N_11249,N_10804);
and U11757 (N_11757,N_11245,N_10994);
nor U11758 (N_11758,N_10726,N_11088);
nand U11759 (N_11759,N_11145,N_10762);
or U11760 (N_11760,N_10920,N_10657);
and U11761 (N_11761,N_10925,N_10650);
or U11762 (N_11762,N_11047,N_11131);
xor U11763 (N_11763,N_10709,N_11106);
nor U11764 (N_11764,N_11033,N_11245);
xor U11765 (N_11765,N_10696,N_10889);
nor U11766 (N_11766,N_10877,N_10823);
nor U11767 (N_11767,N_10958,N_10956);
or U11768 (N_11768,N_10918,N_10779);
and U11769 (N_11769,N_11101,N_10704);
and U11770 (N_11770,N_10880,N_11190);
nor U11771 (N_11771,N_11056,N_10622);
nor U11772 (N_11772,N_10945,N_10959);
xor U11773 (N_11773,N_10507,N_10721);
or U11774 (N_11774,N_10569,N_10650);
nand U11775 (N_11775,N_11149,N_10525);
and U11776 (N_11776,N_11097,N_10610);
nor U11777 (N_11777,N_10601,N_10559);
or U11778 (N_11778,N_10673,N_10506);
xnor U11779 (N_11779,N_10666,N_10607);
nand U11780 (N_11780,N_10940,N_10732);
nand U11781 (N_11781,N_10667,N_10567);
or U11782 (N_11782,N_11055,N_10726);
xnor U11783 (N_11783,N_10826,N_11237);
xnor U11784 (N_11784,N_11239,N_11220);
and U11785 (N_11785,N_11204,N_11214);
nand U11786 (N_11786,N_10735,N_11136);
nand U11787 (N_11787,N_11144,N_10640);
xor U11788 (N_11788,N_11039,N_11160);
or U11789 (N_11789,N_11044,N_10672);
or U11790 (N_11790,N_10573,N_10616);
and U11791 (N_11791,N_10539,N_10622);
or U11792 (N_11792,N_10756,N_10988);
or U11793 (N_11793,N_11224,N_10998);
or U11794 (N_11794,N_10744,N_10710);
nand U11795 (N_11795,N_11190,N_10700);
nand U11796 (N_11796,N_10540,N_11232);
and U11797 (N_11797,N_10767,N_10544);
xor U11798 (N_11798,N_10835,N_11247);
xnor U11799 (N_11799,N_11033,N_10840);
nand U11800 (N_11800,N_10680,N_10515);
nor U11801 (N_11801,N_10878,N_10815);
or U11802 (N_11802,N_10644,N_11073);
and U11803 (N_11803,N_11018,N_10803);
nand U11804 (N_11804,N_10572,N_11062);
xnor U11805 (N_11805,N_10851,N_10725);
and U11806 (N_11806,N_10750,N_11015);
and U11807 (N_11807,N_10707,N_10794);
xor U11808 (N_11808,N_10659,N_10831);
nand U11809 (N_11809,N_10650,N_11007);
and U11810 (N_11810,N_10964,N_11032);
nor U11811 (N_11811,N_11168,N_11167);
or U11812 (N_11812,N_10780,N_10679);
or U11813 (N_11813,N_10534,N_10853);
xor U11814 (N_11814,N_11013,N_10669);
and U11815 (N_11815,N_10555,N_11191);
xor U11816 (N_11816,N_10630,N_10993);
nand U11817 (N_11817,N_10914,N_10636);
or U11818 (N_11818,N_11229,N_11205);
and U11819 (N_11819,N_10993,N_10582);
xnor U11820 (N_11820,N_11009,N_10559);
or U11821 (N_11821,N_11197,N_10512);
nor U11822 (N_11822,N_11069,N_10712);
xnor U11823 (N_11823,N_10514,N_10839);
or U11824 (N_11824,N_10688,N_10880);
nand U11825 (N_11825,N_11009,N_11231);
nand U11826 (N_11826,N_10524,N_10762);
xnor U11827 (N_11827,N_10601,N_10850);
xnor U11828 (N_11828,N_11235,N_11177);
or U11829 (N_11829,N_10610,N_10867);
xnor U11830 (N_11830,N_10692,N_10978);
and U11831 (N_11831,N_11017,N_10540);
and U11832 (N_11832,N_11242,N_11186);
or U11833 (N_11833,N_11201,N_11224);
nand U11834 (N_11834,N_10878,N_10802);
nor U11835 (N_11835,N_11005,N_11021);
and U11836 (N_11836,N_11008,N_10502);
and U11837 (N_11837,N_10793,N_11127);
and U11838 (N_11838,N_10595,N_10635);
and U11839 (N_11839,N_10856,N_10757);
nor U11840 (N_11840,N_10618,N_10714);
or U11841 (N_11841,N_10585,N_11090);
nand U11842 (N_11842,N_10541,N_10530);
or U11843 (N_11843,N_10564,N_11168);
and U11844 (N_11844,N_11070,N_10703);
xnor U11845 (N_11845,N_10818,N_10827);
and U11846 (N_11846,N_10608,N_10653);
and U11847 (N_11847,N_10676,N_11193);
nand U11848 (N_11848,N_10841,N_11139);
nand U11849 (N_11849,N_10908,N_11188);
and U11850 (N_11850,N_10891,N_10717);
or U11851 (N_11851,N_10618,N_11097);
nand U11852 (N_11852,N_11072,N_11171);
or U11853 (N_11853,N_11169,N_10558);
xnor U11854 (N_11854,N_10911,N_10847);
nor U11855 (N_11855,N_11048,N_11231);
or U11856 (N_11856,N_11103,N_10737);
nor U11857 (N_11857,N_11142,N_11134);
nand U11858 (N_11858,N_10622,N_10559);
nand U11859 (N_11859,N_10666,N_11123);
or U11860 (N_11860,N_10571,N_11099);
nand U11861 (N_11861,N_11188,N_11189);
or U11862 (N_11862,N_11131,N_10661);
xnor U11863 (N_11863,N_10781,N_11159);
xor U11864 (N_11864,N_11081,N_10862);
nand U11865 (N_11865,N_10623,N_11228);
or U11866 (N_11866,N_11226,N_10736);
xnor U11867 (N_11867,N_10847,N_11043);
nand U11868 (N_11868,N_10972,N_10676);
nand U11869 (N_11869,N_10582,N_10855);
nand U11870 (N_11870,N_10764,N_10716);
or U11871 (N_11871,N_10822,N_10928);
nor U11872 (N_11872,N_10674,N_10939);
and U11873 (N_11873,N_10548,N_10688);
and U11874 (N_11874,N_10989,N_11154);
and U11875 (N_11875,N_10593,N_10748);
nand U11876 (N_11876,N_11087,N_11115);
nor U11877 (N_11877,N_11236,N_10977);
nand U11878 (N_11878,N_10781,N_11095);
nand U11879 (N_11879,N_10984,N_10853);
and U11880 (N_11880,N_10514,N_11211);
and U11881 (N_11881,N_10550,N_10772);
nor U11882 (N_11882,N_11038,N_11223);
xor U11883 (N_11883,N_10851,N_11095);
nand U11884 (N_11884,N_10837,N_11096);
and U11885 (N_11885,N_10699,N_10585);
nor U11886 (N_11886,N_10856,N_10514);
nor U11887 (N_11887,N_10605,N_11236);
xor U11888 (N_11888,N_10556,N_10666);
and U11889 (N_11889,N_10777,N_10965);
and U11890 (N_11890,N_10838,N_11191);
xor U11891 (N_11891,N_10803,N_10947);
or U11892 (N_11892,N_11234,N_10801);
nand U11893 (N_11893,N_10969,N_11215);
nor U11894 (N_11894,N_10616,N_10662);
and U11895 (N_11895,N_11021,N_10627);
nand U11896 (N_11896,N_10959,N_11166);
nor U11897 (N_11897,N_10924,N_10803);
and U11898 (N_11898,N_10507,N_10541);
or U11899 (N_11899,N_11091,N_10922);
nand U11900 (N_11900,N_10644,N_10508);
nand U11901 (N_11901,N_11224,N_11016);
and U11902 (N_11902,N_11108,N_10687);
and U11903 (N_11903,N_10540,N_10787);
and U11904 (N_11904,N_10503,N_10600);
nand U11905 (N_11905,N_10637,N_10772);
nand U11906 (N_11906,N_11203,N_11035);
nor U11907 (N_11907,N_10922,N_10668);
or U11908 (N_11908,N_10981,N_11144);
nor U11909 (N_11909,N_10957,N_10988);
or U11910 (N_11910,N_10825,N_10773);
and U11911 (N_11911,N_11081,N_10570);
nor U11912 (N_11912,N_11019,N_10829);
xor U11913 (N_11913,N_10610,N_10692);
or U11914 (N_11914,N_10739,N_10763);
xor U11915 (N_11915,N_10798,N_10840);
nand U11916 (N_11916,N_10535,N_11174);
and U11917 (N_11917,N_11204,N_10748);
or U11918 (N_11918,N_11058,N_11126);
or U11919 (N_11919,N_10989,N_10803);
nand U11920 (N_11920,N_11122,N_10802);
nor U11921 (N_11921,N_10935,N_10885);
and U11922 (N_11922,N_11014,N_10648);
nand U11923 (N_11923,N_11078,N_10771);
xor U11924 (N_11924,N_10932,N_11118);
nand U11925 (N_11925,N_10715,N_10821);
or U11926 (N_11926,N_10599,N_10530);
xor U11927 (N_11927,N_10876,N_11077);
or U11928 (N_11928,N_10808,N_10936);
xor U11929 (N_11929,N_11180,N_10527);
nand U11930 (N_11930,N_10905,N_10954);
xor U11931 (N_11931,N_10871,N_10954);
and U11932 (N_11932,N_10863,N_10647);
or U11933 (N_11933,N_10662,N_10657);
xor U11934 (N_11934,N_10719,N_10660);
xor U11935 (N_11935,N_10550,N_10500);
and U11936 (N_11936,N_10709,N_11129);
or U11937 (N_11937,N_10734,N_10708);
xor U11938 (N_11938,N_10633,N_11050);
and U11939 (N_11939,N_11057,N_10998);
xnor U11940 (N_11940,N_10509,N_11183);
and U11941 (N_11941,N_10901,N_10786);
nor U11942 (N_11942,N_11012,N_11205);
or U11943 (N_11943,N_11127,N_10566);
xnor U11944 (N_11944,N_10993,N_10569);
and U11945 (N_11945,N_10624,N_10813);
xor U11946 (N_11946,N_11021,N_10584);
xor U11947 (N_11947,N_11196,N_10685);
nor U11948 (N_11948,N_11235,N_10985);
xnor U11949 (N_11949,N_10680,N_10813);
nor U11950 (N_11950,N_11170,N_11223);
xor U11951 (N_11951,N_10618,N_10599);
nor U11952 (N_11952,N_11011,N_10826);
nor U11953 (N_11953,N_10620,N_11105);
xor U11954 (N_11954,N_10511,N_10966);
and U11955 (N_11955,N_10688,N_11100);
nor U11956 (N_11956,N_11162,N_11155);
nand U11957 (N_11957,N_10610,N_11247);
or U11958 (N_11958,N_10561,N_10853);
nor U11959 (N_11959,N_10828,N_10542);
nand U11960 (N_11960,N_10730,N_10691);
nor U11961 (N_11961,N_10949,N_10558);
xnor U11962 (N_11962,N_11225,N_10720);
xnor U11963 (N_11963,N_11030,N_10810);
nand U11964 (N_11964,N_10885,N_10729);
and U11965 (N_11965,N_11078,N_10999);
and U11966 (N_11966,N_10745,N_10811);
nand U11967 (N_11967,N_10671,N_10819);
and U11968 (N_11968,N_11090,N_11055);
and U11969 (N_11969,N_11138,N_10594);
nand U11970 (N_11970,N_10527,N_11214);
and U11971 (N_11971,N_11084,N_10994);
or U11972 (N_11972,N_10956,N_10533);
or U11973 (N_11973,N_11000,N_11060);
nor U11974 (N_11974,N_10799,N_10556);
or U11975 (N_11975,N_10678,N_10914);
and U11976 (N_11976,N_10913,N_10887);
nand U11977 (N_11977,N_10778,N_11062);
xnor U11978 (N_11978,N_10630,N_11014);
or U11979 (N_11979,N_11056,N_10799);
or U11980 (N_11980,N_11051,N_10811);
or U11981 (N_11981,N_10911,N_10577);
nand U11982 (N_11982,N_10731,N_11020);
nand U11983 (N_11983,N_10987,N_11208);
and U11984 (N_11984,N_10771,N_10637);
or U11985 (N_11985,N_10531,N_11001);
xor U11986 (N_11986,N_11236,N_10830);
xor U11987 (N_11987,N_11167,N_10699);
nand U11988 (N_11988,N_11111,N_10841);
nor U11989 (N_11989,N_10567,N_10984);
and U11990 (N_11990,N_10808,N_11232);
or U11991 (N_11991,N_10871,N_10818);
nor U11992 (N_11992,N_10739,N_10734);
or U11993 (N_11993,N_11222,N_10680);
or U11994 (N_11994,N_11082,N_10643);
nand U11995 (N_11995,N_10904,N_10737);
nor U11996 (N_11996,N_11114,N_11100);
or U11997 (N_11997,N_11098,N_11046);
and U11998 (N_11998,N_10717,N_11024);
and U11999 (N_11999,N_10537,N_11151);
nand U12000 (N_12000,N_11397,N_11371);
or U12001 (N_12001,N_11434,N_11395);
and U12002 (N_12002,N_11714,N_11711);
xor U12003 (N_12003,N_11413,N_11912);
and U12004 (N_12004,N_11270,N_11406);
xor U12005 (N_12005,N_11688,N_11463);
nor U12006 (N_12006,N_11330,N_11704);
and U12007 (N_12007,N_11307,N_11416);
or U12008 (N_12008,N_11781,N_11755);
or U12009 (N_12009,N_11503,N_11545);
or U12010 (N_12010,N_11532,N_11908);
nand U12011 (N_12011,N_11658,N_11581);
and U12012 (N_12012,N_11424,N_11309);
and U12013 (N_12013,N_11622,N_11932);
nor U12014 (N_12014,N_11647,N_11967);
and U12015 (N_12015,N_11611,N_11841);
or U12016 (N_12016,N_11756,N_11376);
or U12017 (N_12017,N_11881,N_11517);
nand U12018 (N_12018,N_11619,N_11883);
nor U12019 (N_12019,N_11402,N_11437);
nand U12020 (N_12020,N_11701,N_11880);
and U12021 (N_12021,N_11775,N_11316);
xnor U12022 (N_12022,N_11964,N_11389);
and U12023 (N_12023,N_11925,N_11926);
and U12024 (N_12024,N_11420,N_11540);
or U12025 (N_12025,N_11329,N_11610);
nand U12026 (N_12026,N_11910,N_11885);
nand U12027 (N_12027,N_11888,N_11591);
and U12028 (N_12028,N_11509,N_11414);
nor U12029 (N_12029,N_11620,N_11957);
and U12030 (N_12030,N_11575,N_11914);
nand U12031 (N_12031,N_11853,N_11308);
or U12032 (N_12032,N_11296,N_11454);
xor U12033 (N_12033,N_11977,N_11810);
nand U12034 (N_12034,N_11823,N_11537);
or U12035 (N_12035,N_11806,N_11678);
nand U12036 (N_12036,N_11900,N_11455);
or U12037 (N_12037,N_11822,N_11483);
nor U12038 (N_12038,N_11663,N_11759);
nor U12039 (N_12039,N_11572,N_11699);
or U12040 (N_12040,N_11857,N_11854);
nand U12041 (N_12041,N_11727,N_11758);
nand U12042 (N_12042,N_11562,N_11916);
and U12043 (N_12043,N_11733,N_11868);
nor U12044 (N_12044,N_11673,N_11605);
xor U12045 (N_12045,N_11835,N_11478);
nor U12046 (N_12046,N_11825,N_11828);
or U12047 (N_12047,N_11633,N_11544);
and U12048 (N_12048,N_11263,N_11566);
nand U12049 (N_12049,N_11936,N_11335);
nand U12050 (N_12050,N_11837,N_11726);
and U12051 (N_12051,N_11831,N_11506);
nand U12052 (N_12052,N_11675,N_11617);
xor U12053 (N_12053,N_11363,N_11482);
nor U12054 (N_12054,N_11426,N_11978);
nor U12055 (N_12055,N_11418,N_11584);
nor U12056 (N_12056,N_11366,N_11290);
nand U12057 (N_12057,N_11762,N_11312);
or U12058 (N_12058,N_11576,N_11808);
and U12059 (N_12059,N_11928,N_11834);
and U12060 (N_12060,N_11452,N_11267);
and U12061 (N_12061,N_11535,N_11986);
or U12062 (N_12062,N_11346,N_11842);
nor U12063 (N_12063,N_11486,N_11404);
xor U12064 (N_12064,N_11720,N_11310);
nand U12065 (N_12065,N_11660,N_11930);
nor U12066 (N_12066,N_11466,N_11253);
nand U12067 (N_12067,N_11268,N_11898);
xnor U12068 (N_12068,N_11737,N_11798);
nand U12069 (N_12069,N_11645,N_11909);
nand U12070 (N_12070,N_11878,N_11777);
xor U12071 (N_12071,N_11281,N_11636);
and U12072 (N_12072,N_11951,N_11311);
or U12073 (N_12073,N_11264,N_11332);
nor U12074 (N_12074,N_11648,N_11696);
and U12075 (N_12075,N_11796,N_11919);
and U12076 (N_12076,N_11355,N_11628);
xor U12077 (N_12077,N_11856,N_11554);
nand U12078 (N_12078,N_11342,N_11784);
and U12079 (N_12079,N_11833,N_11860);
or U12080 (N_12080,N_11724,N_11456);
and U12081 (N_12081,N_11412,N_11975);
xor U12082 (N_12082,N_11565,N_11937);
and U12083 (N_12083,N_11642,N_11892);
or U12084 (N_12084,N_11300,N_11322);
xor U12085 (N_12085,N_11783,N_11971);
nand U12086 (N_12086,N_11470,N_11719);
nor U12087 (N_12087,N_11985,N_11644);
nand U12088 (N_12088,N_11713,N_11879);
xnor U12089 (N_12089,N_11973,N_11315);
nand U12090 (N_12090,N_11543,N_11379);
and U12091 (N_12091,N_11508,N_11811);
and U12092 (N_12092,N_11741,N_11336);
nor U12093 (N_12093,N_11408,N_11561);
xnor U12094 (N_12094,N_11409,N_11702);
nor U12095 (N_12095,N_11996,N_11255);
xnor U12096 (N_12096,N_11867,N_11390);
and U12097 (N_12097,N_11694,N_11326);
nand U12098 (N_12098,N_11260,N_11616);
nor U12099 (N_12099,N_11657,N_11443);
nor U12100 (N_12100,N_11305,N_11906);
nand U12101 (N_12101,N_11374,N_11933);
xnor U12102 (N_12102,N_11794,N_11638);
and U12103 (N_12103,N_11415,N_11552);
nor U12104 (N_12104,N_11349,N_11417);
and U12105 (N_12105,N_11556,N_11635);
nor U12106 (N_12106,N_11323,N_11907);
nor U12107 (N_12107,N_11585,N_11604);
or U12108 (N_12108,N_11449,N_11624);
or U12109 (N_12109,N_11457,N_11380);
nor U12110 (N_12110,N_11812,N_11966);
or U12111 (N_12111,N_11634,N_11943);
nor U12112 (N_12112,N_11364,N_11493);
nand U12113 (N_12113,N_11788,N_11952);
nand U12114 (N_12114,N_11448,N_11266);
nor U12115 (N_12115,N_11829,N_11498);
xnor U12116 (N_12116,N_11859,N_11570);
xnor U12117 (N_12117,N_11950,N_11496);
and U12118 (N_12118,N_11827,N_11304);
or U12119 (N_12119,N_11958,N_11563);
xor U12120 (N_12120,N_11525,N_11626);
nand U12121 (N_12121,N_11725,N_11601);
nor U12122 (N_12122,N_11684,N_11887);
nor U12123 (N_12123,N_11350,N_11385);
nand U12124 (N_12124,N_11671,N_11301);
and U12125 (N_12125,N_11716,N_11394);
nor U12126 (N_12126,N_11499,N_11836);
or U12127 (N_12127,N_11941,N_11847);
nand U12128 (N_12128,N_11459,N_11718);
nor U12129 (N_12129,N_11286,N_11484);
nor U12130 (N_12130,N_11472,N_11793);
nand U12131 (N_12131,N_11344,N_11410);
nor U12132 (N_12132,N_11770,N_11513);
xor U12133 (N_12133,N_11766,N_11785);
or U12134 (N_12134,N_11608,N_11451);
or U12135 (N_12135,N_11567,N_11970);
xor U12136 (N_12136,N_11993,N_11803);
and U12137 (N_12137,N_11365,N_11747);
and U12138 (N_12138,N_11594,N_11757);
nand U12139 (N_12139,N_11961,N_11817);
or U12140 (N_12140,N_11297,N_11539);
or U12141 (N_12141,N_11999,N_11795);
xor U12142 (N_12142,N_11786,N_11516);
or U12143 (N_12143,N_11272,N_11818);
nor U12144 (N_12144,N_11771,N_11987);
nor U12145 (N_12145,N_11627,N_11816);
xnor U12146 (N_12146,N_11918,N_11685);
and U12147 (N_12147,N_11790,N_11754);
or U12148 (N_12148,N_11615,N_11676);
nor U12149 (N_12149,N_11614,N_11686);
nand U12150 (N_12150,N_11821,N_11799);
xnor U12151 (N_12151,N_11938,N_11369);
xnor U12152 (N_12152,N_11876,N_11613);
or U12153 (N_12153,N_11949,N_11820);
nor U12154 (N_12154,N_11843,N_11729);
and U12155 (N_12155,N_11889,N_11935);
and U12156 (N_12156,N_11924,N_11846);
or U12157 (N_12157,N_11431,N_11998);
and U12158 (N_12158,N_11292,N_11683);
or U12159 (N_12159,N_11929,N_11893);
xnor U12160 (N_12160,N_11746,N_11809);
or U12161 (N_12161,N_11579,N_11564);
xor U12162 (N_12162,N_11273,N_11862);
and U12163 (N_12163,N_11728,N_11722);
and U12164 (N_12164,N_11779,N_11712);
nor U12165 (N_12165,N_11618,N_11805);
and U12166 (N_12166,N_11444,N_11460);
xor U12167 (N_12167,N_11595,N_11739);
or U12168 (N_12168,N_11400,N_11709);
xnor U12169 (N_12169,N_11652,N_11681);
nand U12170 (N_12170,N_11661,N_11436);
xnor U12171 (N_12171,N_11874,N_11972);
or U12172 (N_12172,N_11801,N_11774);
xnor U12173 (N_12173,N_11715,N_11778);
or U12174 (N_12174,N_11468,N_11844);
nand U12175 (N_12175,N_11959,N_11873);
or U12176 (N_12176,N_11501,N_11599);
or U12177 (N_12177,N_11473,N_11692);
nand U12178 (N_12178,N_11597,N_11407);
and U12179 (N_12179,N_11515,N_11465);
nor U12180 (N_12180,N_11639,N_11334);
nor U12181 (N_12181,N_11851,N_11587);
nand U12182 (N_12182,N_11863,N_11979);
nand U12183 (N_12183,N_11668,N_11531);
nand U12184 (N_12184,N_11588,N_11769);
nor U12185 (N_12185,N_11871,N_11477);
and U12186 (N_12186,N_11962,N_11838);
xnor U12187 (N_12187,N_11954,N_11441);
xor U12188 (N_12188,N_11621,N_11682);
and U12189 (N_12189,N_11403,N_11432);
nor U12190 (N_12190,N_11731,N_11491);
and U12191 (N_12191,N_11352,N_11705);
and U12192 (N_12192,N_11849,N_11523);
nor U12193 (N_12193,N_11277,N_11845);
or U12194 (N_12194,N_11283,N_11596);
or U12195 (N_12195,N_11401,N_11446);
nand U12196 (N_12196,N_11666,N_11734);
nor U12197 (N_12197,N_11373,N_11419);
or U12198 (N_12198,N_11697,N_11299);
nor U12199 (N_12199,N_11869,N_11968);
nand U12200 (N_12200,N_11679,N_11398);
xnor U12201 (N_12201,N_11589,N_11505);
nor U12202 (N_12202,N_11861,N_11953);
xor U12203 (N_12203,N_11302,N_11631);
xnor U12204 (N_12204,N_11577,N_11314);
xnor U12205 (N_12205,N_11956,N_11677);
or U12206 (N_12206,N_11745,N_11367);
xnor U12207 (N_12207,N_11573,N_11280);
nor U12208 (N_12208,N_11659,N_11359);
or U12209 (N_12209,N_11667,N_11534);
xnor U12210 (N_12210,N_11687,N_11982);
xnor U12211 (N_12211,N_11288,N_11522);
nand U12212 (N_12212,N_11378,N_11640);
nand U12213 (N_12213,N_11923,N_11442);
nand U12214 (N_12214,N_11293,N_11422);
and U12215 (N_12215,N_11824,N_11467);
or U12216 (N_12216,N_11259,N_11538);
nand U12217 (N_12217,N_11607,N_11313);
xnor U12218 (N_12218,N_11768,N_11333);
or U12219 (N_12219,N_11665,N_11319);
xnor U12220 (N_12220,N_11751,N_11995);
nor U12221 (N_12221,N_11934,N_11511);
nand U12222 (N_12222,N_11852,N_11598);
xor U12223 (N_12223,N_11875,N_11603);
xor U12224 (N_12224,N_11984,N_11429);
and U12225 (N_12225,N_11551,N_11946);
and U12226 (N_12226,N_11568,N_11902);
and U12227 (N_12227,N_11753,N_11730);
and U12228 (N_12228,N_11490,N_11555);
nand U12229 (N_12229,N_11289,N_11592);
nand U12230 (N_12230,N_11340,N_11927);
or U12231 (N_12231,N_11435,N_11760);
or U12232 (N_12232,N_11370,N_11362);
nor U12233 (N_12233,N_11321,N_11976);
xnor U12234 (N_12234,N_11502,N_11317);
and U12235 (N_12235,N_11519,N_11947);
nand U12236 (N_12236,N_11942,N_11530);
xnor U12237 (N_12237,N_11433,N_11580);
nor U12238 (N_12238,N_11328,N_11285);
or U12239 (N_12239,N_11269,N_11558);
nor U12240 (N_12240,N_11480,N_11318);
and U12241 (N_12241,N_11262,N_11695);
or U12242 (N_12242,N_11690,N_11251);
or U12243 (N_12243,N_11858,N_11654);
xor U12244 (N_12244,N_11680,N_11629);
nand U12245 (N_12245,N_11423,N_11710);
xnor U12246 (N_12246,N_11440,N_11819);
nand U12247 (N_12247,N_11495,N_11903);
xnor U12248 (N_12248,N_11578,N_11476);
xnor U12249 (N_12249,N_11399,N_11430);
and U12250 (N_12250,N_11913,N_11593);
nor U12251 (N_12251,N_11797,N_11643);
and U12252 (N_12252,N_11960,N_11388);
nand U12253 (N_12253,N_11717,N_11981);
and U12254 (N_12254,N_11361,N_11965);
xnor U12255 (N_12255,N_11662,N_11773);
nor U12256 (N_12256,N_11814,N_11276);
and U12257 (N_12257,N_11649,N_11877);
nor U12258 (N_12258,N_11750,N_11707);
and U12259 (N_12259,N_11391,N_11890);
nand U12260 (N_12260,N_11469,N_11375);
xnor U12261 (N_12261,N_11765,N_11529);
nand U12262 (N_12262,N_11396,N_11504);
or U12263 (N_12263,N_11325,N_11761);
xor U12264 (N_12264,N_11895,N_11736);
and U12265 (N_12265,N_11904,N_11347);
or U12266 (N_12266,N_11655,N_11708);
or U12267 (N_12267,N_11298,N_11343);
and U12268 (N_12268,N_11899,N_11815);
nand U12269 (N_12269,N_11339,N_11945);
or U12270 (N_12270,N_11291,N_11258);
xnor U12271 (N_12271,N_11991,N_11732);
xnor U12272 (N_12272,N_11358,N_11533);
nand U12273 (N_12273,N_11915,N_11354);
and U12274 (N_12274,N_11590,N_11360);
nor U12275 (N_12275,N_11743,N_11421);
nand U12276 (N_12276,N_11439,N_11782);
nand U12277 (N_12277,N_11341,N_11921);
xnor U12278 (N_12278,N_11274,N_11650);
or U12279 (N_12279,N_11691,N_11632);
or U12280 (N_12280,N_11911,N_11672);
nand U12281 (N_12281,N_11527,N_11284);
xor U12282 (N_12282,N_11461,N_11521);
nor U12283 (N_12283,N_11997,N_11646);
nor U12284 (N_12284,N_11494,N_11475);
nand U12285 (N_12285,N_11948,N_11536);
or U12286 (N_12286,N_11252,N_11485);
nor U12287 (N_12287,N_11520,N_11767);
xnor U12288 (N_12288,N_11807,N_11275);
and U12289 (N_12289,N_11507,N_11586);
nand U12290 (N_12290,N_11602,N_11377);
and U12291 (N_12291,N_11392,N_11693);
or U12292 (N_12292,N_11653,N_11939);
xnor U12293 (N_12293,N_11748,N_11353);
or U12294 (N_12294,N_11487,N_11337);
xor U12295 (N_12295,N_11901,N_11582);
xnor U12296 (N_12296,N_11866,N_11839);
nor U12297 (N_12297,N_11357,N_11600);
and U12298 (N_12298,N_11891,N_11800);
or U12299 (N_12299,N_11630,N_11489);
and U12300 (N_12300,N_11792,N_11855);
xor U12301 (N_12301,N_11327,N_11453);
xnor U12302 (N_12302,N_11664,N_11992);
or U12303 (N_12303,N_11850,N_11872);
nor U12304 (N_12304,N_11983,N_11787);
and U12305 (N_12305,N_11546,N_11387);
nor U12306 (N_12306,N_11382,N_11703);
or U12307 (N_12307,N_11752,N_11848);
or U12308 (N_12308,N_11381,N_11669);
nand U12309 (N_12309,N_11742,N_11338);
and U12310 (N_12310,N_11479,N_11514);
xnor U12311 (N_12311,N_11560,N_11840);
and U12312 (N_12312,N_11922,N_11279);
xor U12313 (N_12313,N_11882,N_11512);
nor U12314 (N_12314,N_11813,N_11955);
nor U12315 (N_12315,N_11791,N_11550);
and U12316 (N_12316,N_11306,N_11612);
nor U12317 (N_12317,N_11278,N_11524);
nand U12318 (N_12318,N_11492,N_11651);
nand U12319 (N_12319,N_11749,N_11896);
nor U12320 (N_12320,N_11721,N_11569);
nor U12321 (N_12321,N_11884,N_11763);
nand U12322 (N_12322,N_11510,N_11674);
or U12323 (N_12323,N_11351,N_11303);
nand U12324 (N_12324,N_11497,N_11700);
and U12325 (N_12325,N_11518,N_11723);
nor U12326 (N_12326,N_11804,N_11557);
nand U12327 (N_12327,N_11989,N_11864);
nor U12328 (N_12328,N_11789,N_11894);
or U12329 (N_12329,N_11427,N_11331);
nor U12330 (N_12330,N_11356,N_11706);
nand U12331 (N_12331,N_11294,N_11559);
nor U12332 (N_12332,N_11780,N_11897);
nand U12333 (N_12333,N_11656,N_11944);
xnor U12334 (N_12334,N_11637,N_11772);
nor U12335 (N_12335,N_11571,N_11990);
or U12336 (N_12336,N_11740,N_11865);
nand U12337 (N_12337,N_11384,N_11553);
and U12338 (N_12338,N_11261,N_11282);
nand U12339 (N_12339,N_11542,N_11257);
or U12340 (N_12340,N_11428,N_11474);
or U12341 (N_12341,N_11411,N_11287);
nor U12342 (N_12342,N_11393,N_11905);
and U12343 (N_12343,N_11764,N_11368);
nand U12344 (N_12344,N_11802,N_11445);
nor U12345 (N_12345,N_11623,N_11980);
nand U12346 (N_12346,N_11826,N_11547);
nor U12347 (N_12347,N_11583,N_11458);
or U12348 (N_12348,N_11548,N_11549);
nand U12349 (N_12349,N_11609,N_11250);
nand U12350 (N_12350,N_11886,N_11735);
or U12351 (N_12351,N_11450,N_11974);
or U12352 (N_12352,N_11526,N_11940);
xor U12353 (N_12353,N_11462,N_11625);
xnor U12354 (N_12354,N_11744,N_11698);
xnor U12355 (N_12355,N_11670,N_11372);
xor U12356 (N_12356,N_11830,N_11541);
and U12357 (N_12357,N_11738,N_11254);
or U12358 (N_12358,N_11641,N_11447);
and U12359 (N_12359,N_11574,N_11464);
xnor U12360 (N_12360,N_11386,N_11471);
nand U12361 (N_12361,N_11606,N_11265);
xor U12362 (N_12362,N_11320,N_11383);
and U12363 (N_12363,N_11776,N_11425);
nor U12364 (N_12364,N_11994,N_11438);
nand U12365 (N_12365,N_11528,N_11271);
xnor U12366 (N_12366,N_11348,N_11832);
nand U12367 (N_12367,N_11345,N_11295);
and U12368 (N_12368,N_11481,N_11405);
nor U12369 (N_12369,N_11920,N_11969);
xnor U12370 (N_12370,N_11917,N_11870);
or U12371 (N_12371,N_11324,N_11689);
nand U12372 (N_12372,N_11988,N_11500);
and U12373 (N_12373,N_11488,N_11256);
or U12374 (N_12374,N_11931,N_11963);
xnor U12375 (N_12375,N_11426,N_11563);
and U12376 (N_12376,N_11672,N_11540);
and U12377 (N_12377,N_11621,N_11343);
xnor U12378 (N_12378,N_11317,N_11905);
nor U12379 (N_12379,N_11428,N_11642);
and U12380 (N_12380,N_11362,N_11739);
nor U12381 (N_12381,N_11953,N_11258);
nand U12382 (N_12382,N_11819,N_11532);
nor U12383 (N_12383,N_11251,N_11930);
xor U12384 (N_12384,N_11541,N_11746);
xnor U12385 (N_12385,N_11655,N_11768);
and U12386 (N_12386,N_11584,N_11937);
nor U12387 (N_12387,N_11695,N_11918);
nor U12388 (N_12388,N_11420,N_11594);
xnor U12389 (N_12389,N_11340,N_11929);
xor U12390 (N_12390,N_11981,N_11562);
or U12391 (N_12391,N_11496,N_11610);
nand U12392 (N_12392,N_11746,N_11389);
or U12393 (N_12393,N_11400,N_11688);
or U12394 (N_12394,N_11591,N_11543);
and U12395 (N_12395,N_11402,N_11524);
or U12396 (N_12396,N_11592,N_11966);
nor U12397 (N_12397,N_11525,N_11537);
and U12398 (N_12398,N_11969,N_11650);
nand U12399 (N_12399,N_11457,N_11256);
and U12400 (N_12400,N_11549,N_11421);
xnor U12401 (N_12401,N_11982,N_11913);
nor U12402 (N_12402,N_11868,N_11831);
xnor U12403 (N_12403,N_11753,N_11292);
xnor U12404 (N_12404,N_11325,N_11923);
nor U12405 (N_12405,N_11310,N_11619);
xor U12406 (N_12406,N_11426,N_11979);
or U12407 (N_12407,N_11728,N_11778);
xor U12408 (N_12408,N_11814,N_11907);
or U12409 (N_12409,N_11677,N_11647);
nand U12410 (N_12410,N_11934,N_11641);
and U12411 (N_12411,N_11485,N_11638);
xor U12412 (N_12412,N_11478,N_11523);
nor U12413 (N_12413,N_11603,N_11999);
nor U12414 (N_12414,N_11580,N_11747);
or U12415 (N_12415,N_11532,N_11708);
nand U12416 (N_12416,N_11292,N_11771);
nand U12417 (N_12417,N_11403,N_11491);
xnor U12418 (N_12418,N_11671,N_11368);
nor U12419 (N_12419,N_11669,N_11731);
or U12420 (N_12420,N_11315,N_11481);
nor U12421 (N_12421,N_11914,N_11890);
nor U12422 (N_12422,N_11374,N_11757);
or U12423 (N_12423,N_11642,N_11684);
and U12424 (N_12424,N_11725,N_11303);
xnor U12425 (N_12425,N_11813,N_11568);
xnor U12426 (N_12426,N_11280,N_11719);
nor U12427 (N_12427,N_11677,N_11987);
xnor U12428 (N_12428,N_11426,N_11704);
or U12429 (N_12429,N_11567,N_11806);
and U12430 (N_12430,N_11675,N_11792);
or U12431 (N_12431,N_11786,N_11254);
and U12432 (N_12432,N_11849,N_11559);
nor U12433 (N_12433,N_11775,N_11607);
and U12434 (N_12434,N_11303,N_11313);
nor U12435 (N_12435,N_11787,N_11710);
or U12436 (N_12436,N_11288,N_11425);
or U12437 (N_12437,N_11373,N_11980);
xor U12438 (N_12438,N_11841,N_11504);
nor U12439 (N_12439,N_11864,N_11651);
nand U12440 (N_12440,N_11725,N_11513);
xor U12441 (N_12441,N_11970,N_11873);
or U12442 (N_12442,N_11773,N_11652);
or U12443 (N_12443,N_11391,N_11994);
and U12444 (N_12444,N_11308,N_11293);
or U12445 (N_12445,N_11489,N_11876);
xnor U12446 (N_12446,N_11962,N_11850);
nand U12447 (N_12447,N_11780,N_11519);
nor U12448 (N_12448,N_11487,N_11866);
nor U12449 (N_12449,N_11533,N_11364);
or U12450 (N_12450,N_11338,N_11661);
nand U12451 (N_12451,N_11376,N_11686);
and U12452 (N_12452,N_11741,N_11993);
nor U12453 (N_12453,N_11550,N_11893);
and U12454 (N_12454,N_11360,N_11387);
nand U12455 (N_12455,N_11727,N_11368);
nand U12456 (N_12456,N_11265,N_11383);
and U12457 (N_12457,N_11565,N_11551);
xnor U12458 (N_12458,N_11408,N_11690);
xor U12459 (N_12459,N_11644,N_11814);
nor U12460 (N_12460,N_11262,N_11871);
xnor U12461 (N_12461,N_11719,N_11558);
xor U12462 (N_12462,N_11601,N_11363);
or U12463 (N_12463,N_11821,N_11500);
xor U12464 (N_12464,N_11759,N_11653);
nor U12465 (N_12465,N_11942,N_11776);
and U12466 (N_12466,N_11822,N_11288);
or U12467 (N_12467,N_11559,N_11416);
or U12468 (N_12468,N_11909,N_11876);
and U12469 (N_12469,N_11765,N_11285);
nand U12470 (N_12470,N_11649,N_11317);
xor U12471 (N_12471,N_11695,N_11542);
xnor U12472 (N_12472,N_11499,N_11766);
or U12473 (N_12473,N_11981,N_11992);
or U12474 (N_12474,N_11946,N_11586);
nor U12475 (N_12475,N_11555,N_11314);
or U12476 (N_12476,N_11528,N_11647);
nor U12477 (N_12477,N_11972,N_11626);
or U12478 (N_12478,N_11470,N_11883);
nor U12479 (N_12479,N_11254,N_11657);
xnor U12480 (N_12480,N_11568,N_11680);
xor U12481 (N_12481,N_11932,N_11311);
xor U12482 (N_12482,N_11871,N_11393);
xor U12483 (N_12483,N_11450,N_11555);
and U12484 (N_12484,N_11980,N_11429);
nor U12485 (N_12485,N_11537,N_11723);
or U12486 (N_12486,N_11793,N_11737);
or U12487 (N_12487,N_11935,N_11565);
xnor U12488 (N_12488,N_11666,N_11735);
nand U12489 (N_12489,N_11437,N_11611);
xor U12490 (N_12490,N_11970,N_11767);
xnor U12491 (N_12491,N_11574,N_11671);
and U12492 (N_12492,N_11871,N_11602);
nor U12493 (N_12493,N_11979,N_11441);
and U12494 (N_12494,N_11264,N_11560);
nand U12495 (N_12495,N_11805,N_11386);
nor U12496 (N_12496,N_11601,N_11748);
nand U12497 (N_12497,N_11667,N_11776);
xnor U12498 (N_12498,N_11373,N_11589);
xor U12499 (N_12499,N_11999,N_11695);
nor U12500 (N_12500,N_11326,N_11876);
xor U12501 (N_12501,N_11776,N_11699);
or U12502 (N_12502,N_11695,N_11470);
or U12503 (N_12503,N_11727,N_11769);
xor U12504 (N_12504,N_11388,N_11512);
nand U12505 (N_12505,N_11271,N_11884);
or U12506 (N_12506,N_11797,N_11464);
or U12507 (N_12507,N_11786,N_11416);
and U12508 (N_12508,N_11828,N_11550);
xor U12509 (N_12509,N_11902,N_11539);
nor U12510 (N_12510,N_11545,N_11659);
nand U12511 (N_12511,N_11884,N_11659);
or U12512 (N_12512,N_11407,N_11543);
and U12513 (N_12513,N_11460,N_11421);
and U12514 (N_12514,N_11393,N_11830);
or U12515 (N_12515,N_11811,N_11587);
or U12516 (N_12516,N_11420,N_11560);
nor U12517 (N_12517,N_11757,N_11568);
or U12518 (N_12518,N_11967,N_11574);
and U12519 (N_12519,N_11972,N_11411);
nand U12520 (N_12520,N_11319,N_11686);
nand U12521 (N_12521,N_11545,N_11372);
nor U12522 (N_12522,N_11692,N_11501);
or U12523 (N_12523,N_11689,N_11494);
nor U12524 (N_12524,N_11951,N_11828);
or U12525 (N_12525,N_11929,N_11252);
or U12526 (N_12526,N_11723,N_11803);
nand U12527 (N_12527,N_11428,N_11666);
xnor U12528 (N_12528,N_11518,N_11940);
nand U12529 (N_12529,N_11996,N_11772);
or U12530 (N_12530,N_11877,N_11300);
nor U12531 (N_12531,N_11649,N_11871);
xnor U12532 (N_12532,N_11587,N_11889);
or U12533 (N_12533,N_11622,N_11406);
nor U12534 (N_12534,N_11431,N_11301);
nand U12535 (N_12535,N_11381,N_11503);
and U12536 (N_12536,N_11643,N_11831);
nand U12537 (N_12537,N_11273,N_11416);
nor U12538 (N_12538,N_11713,N_11485);
nand U12539 (N_12539,N_11672,N_11265);
nor U12540 (N_12540,N_11719,N_11258);
xor U12541 (N_12541,N_11622,N_11404);
nand U12542 (N_12542,N_11566,N_11607);
xor U12543 (N_12543,N_11698,N_11416);
or U12544 (N_12544,N_11911,N_11499);
or U12545 (N_12545,N_11897,N_11399);
nor U12546 (N_12546,N_11482,N_11832);
and U12547 (N_12547,N_11487,N_11445);
or U12548 (N_12548,N_11441,N_11317);
nor U12549 (N_12549,N_11435,N_11855);
or U12550 (N_12550,N_11565,N_11270);
xnor U12551 (N_12551,N_11481,N_11586);
or U12552 (N_12552,N_11347,N_11935);
and U12553 (N_12553,N_11837,N_11709);
and U12554 (N_12554,N_11946,N_11255);
or U12555 (N_12555,N_11489,N_11844);
or U12556 (N_12556,N_11905,N_11800);
and U12557 (N_12557,N_11800,N_11991);
and U12558 (N_12558,N_11814,N_11402);
and U12559 (N_12559,N_11910,N_11653);
and U12560 (N_12560,N_11298,N_11447);
nand U12561 (N_12561,N_11858,N_11673);
or U12562 (N_12562,N_11744,N_11471);
and U12563 (N_12563,N_11936,N_11670);
and U12564 (N_12564,N_11659,N_11308);
and U12565 (N_12565,N_11316,N_11656);
nor U12566 (N_12566,N_11904,N_11688);
nand U12567 (N_12567,N_11910,N_11958);
nor U12568 (N_12568,N_11287,N_11485);
or U12569 (N_12569,N_11725,N_11550);
and U12570 (N_12570,N_11823,N_11630);
nand U12571 (N_12571,N_11881,N_11786);
and U12572 (N_12572,N_11948,N_11837);
nor U12573 (N_12573,N_11651,N_11868);
or U12574 (N_12574,N_11750,N_11756);
xor U12575 (N_12575,N_11738,N_11507);
nand U12576 (N_12576,N_11947,N_11772);
nor U12577 (N_12577,N_11781,N_11825);
xor U12578 (N_12578,N_11380,N_11687);
nand U12579 (N_12579,N_11742,N_11522);
nand U12580 (N_12580,N_11710,N_11625);
nor U12581 (N_12581,N_11897,N_11546);
nand U12582 (N_12582,N_11950,N_11619);
nand U12583 (N_12583,N_11523,N_11579);
xnor U12584 (N_12584,N_11830,N_11305);
and U12585 (N_12585,N_11605,N_11647);
xor U12586 (N_12586,N_11276,N_11846);
xnor U12587 (N_12587,N_11559,N_11532);
nor U12588 (N_12588,N_11271,N_11300);
nand U12589 (N_12589,N_11897,N_11665);
and U12590 (N_12590,N_11408,N_11751);
or U12591 (N_12591,N_11970,N_11294);
nand U12592 (N_12592,N_11925,N_11989);
xor U12593 (N_12593,N_11561,N_11692);
xor U12594 (N_12594,N_11418,N_11813);
and U12595 (N_12595,N_11701,N_11516);
nor U12596 (N_12596,N_11654,N_11584);
nor U12597 (N_12597,N_11746,N_11526);
nand U12598 (N_12598,N_11256,N_11499);
or U12599 (N_12599,N_11497,N_11840);
and U12600 (N_12600,N_11334,N_11272);
nor U12601 (N_12601,N_11428,N_11718);
and U12602 (N_12602,N_11835,N_11969);
and U12603 (N_12603,N_11799,N_11961);
and U12604 (N_12604,N_11600,N_11622);
nand U12605 (N_12605,N_11735,N_11442);
xnor U12606 (N_12606,N_11358,N_11676);
and U12607 (N_12607,N_11764,N_11445);
or U12608 (N_12608,N_11483,N_11832);
nand U12609 (N_12609,N_11618,N_11823);
xnor U12610 (N_12610,N_11563,N_11921);
xor U12611 (N_12611,N_11906,N_11397);
xor U12612 (N_12612,N_11738,N_11898);
or U12613 (N_12613,N_11936,N_11904);
or U12614 (N_12614,N_11688,N_11780);
or U12615 (N_12615,N_11694,N_11954);
xor U12616 (N_12616,N_11490,N_11659);
nor U12617 (N_12617,N_11692,N_11312);
and U12618 (N_12618,N_11531,N_11526);
nand U12619 (N_12619,N_11935,N_11650);
nand U12620 (N_12620,N_11628,N_11953);
nand U12621 (N_12621,N_11350,N_11365);
nor U12622 (N_12622,N_11429,N_11875);
nand U12623 (N_12623,N_11544,N_11447);
and U12624 (N_12624,N_11295,N_11590);
xnor U12625 (N_12625,N_11881,N_11305);
nand U12626 (N_12626,N_11554,N_11267);
nand U12627 (N_12627,N_11508,N_11660);
nand U12628 (N_12628,N_11578,N_11254);
or U12629 (N_12629,N_11318,N_11420);
nor U12630 (N_12630,N_11523,N_11296);
or U12631 (N_12631,N_11488,N_11325);
nand U12632 (N_12632,N_11957,N_11910);
xor U12633 (N_12633,N_11280,N_11736);
xnor U12634 (N_12634,N_11793,N_11476);
or U12635 (N_12635,N_11695,N_11507);
or U12636 (N_12636,N_11398,N_11623);
nor U12637 (N_12637,N_11470,N_11834);
nor U12638 (N_12638,N_11495,N_11921);
or U12639 (N_12639,N_11250,N_11300);
nor U12640 (N_12640,N_11753,N_11418);
nand U12641 (N_12641,N_11253,N_11283);
xor U12642 (N_12642,N_11647,N_11643);
nand U12643 (N_12643,N_11994,N_11635);
and U12644 (N_12644,N_11832,N_11484);
or U12645 (N_12645,N_11392,N_11663);
xor U12646 (N_12646,N_11908,N_11829);
nand U12647 (N_12647,N_11387,N_11420);
nand U12648 (N_12648,N_11822,N_11302);
xnor U12649 (N_12649,N_11379,N_11481);
or U12650 (N_12650,N_11716,N_11585);
nand U12651 (N_12651,N_11544,N_11820);
nand U12652 (N_12652,N_11853,N_11512);
nand U12653 (N_12653,N_11786,N_11388);
nor U12654 (N_12654,N_11725,N_11713);
or U12655 (N_12655,N_11514,N_11658);
and U12656 (N_12656,N_11284,N_11903);
nand U12657 (N_12657,N_11364,N_11719);
nand U12658 (N_12658,N_11736,N_11847);
nor U12659 (N_12659,N_11446,N_11434);
nor U12660 (N_12660,N_11576,N_11840);
or U12661 (N_12661,N_11464,N_11269);
and U12662 (N_12662,N_11329,N_11874);
nand U12663 (N_12663,N_11491,N_11904);
nand U12664 (N_12664,N_11856,N_11911);
and U12665 (N_12665,N_11867,N_11387);
xor U12666 (N_12666,N_11704,N_11701);
and U12667 (N_12667,N_11785,N_11824);
xnor U12668 (N_12668,N_11384,N_11952);
or U12669 (N_12669,N_11573,N_11769);
nor U12670 (N_12670,N_11677,N_11379);
or U12671 (N_12671,N_11705,N_11269);
nor U12672 (N_12672,N_11868,N_11818);
nand U12673 (N_12673,N_11665,N_11697);
xor U12674 (N_12674,N_11527,N_11711);
and U12675 (N_12675,N_11473,N_11480);
nor U12676 (N_12676,N_11454,N_11452);
nor U12677 (N_12677,N_11454,N_11260);
and U12678 (N_12678,N_11871,N_11735);
nand U12679 (N_12679,N_11939,N_11690);
nand U12680 (N_12680,N_11909,N_11519);
and U12681 (N_12681,N_11886,N_11524);
nand U12682 (N_12682,N_11691,N_11284);
nand U12683 (N_12683,N_11697,N_11429);
nand U12684 (N_12684,N_11386,N_11514);
or U12685 (N_12685,N_11798,N_11627);
nor U12686 (N_12686,N_11310,N_11478);
xnor U12687 (N_12687,N_11981,N_11734);
or U12688 (N_12688,N_11668,N_11384);
and U12689 (N_12689,N_11370,N_11810);
nor U12690 (N_12690,N_11460,N_11989);
nand U12691 (N_12691,N_11976,N_11795);
nand U12692 (N_12692,N_11637,N_11936);
nor U12693 (N_12693,N_11620,N_11723);
or U12694 (N_12694,N_11329,N_11616);
xor U12695 (N_12695,N_11307,N_11313);
nand U12696 (N_12696,N_11339,N_11657);
xnor U12697 (N_12697,N_11704,N_11716);
xnor U12698 (N_12698,N_11359,N_11335);
xor U12699 (N_12699,N_11630,N_11313);
xnor U12700 (N_12700,N_11927,N_11296);
or U12701 (N_12701,N_11911,N_11832);
nor U12702 (N_12702,N_11458,N_11814);
nand U12703 (N_12703,N_11942,N_11700);
or U12704 (N_12704,N_11510,N_11485);
nand U12705 (N_12705,N_11791,N_11315);
and U12706 (N_12706,N_11588,N_11898);
nand U12707 (N_12707,N_11473,N_11582);
or U12708 (N_12708,N_11447,N_11554);
nor U12709 (N_12709,N_11646,N_11543);
or U12710 (N_12710,N_11314,N_11280);
nor U12711 (N_12711,N_11509,N_11521);
nand U12712 (N_12712,N_11536,N_11907);
or U12713 (N_12713,N_11666,N_11958);
or U12714 (N_12714,N_11566,N_11892);
and U12715 (N_12715,N_11482,N_11852);
xor U12716 (N_12716,N_11478,N_11626);
and U12717 (N_12717,N_11606,N_11782);
nor U12718 (N_12718,N_11382,N_11481);
and U12719 (N_12719,N_11922,N_11982);
and U12720 (N_12720,N_11570,N_11577);
nor U12721 (N_12721,N_11403,N_11764);
nor U12722 (N_12722,N_11443,N_11695);
nor U12723 (N_12723,N_11624,N_11832);
nor U12724 (N_12724,N_11986,N_11362);
xnor U12725 (N_12725,N_11317,N_11267);
or U12726 (N_12726,N_11667,N_11708);
xor U12727 (N_12727,N_11408,N_11403);
xnor U12728 (N_12728,N_11660,N_11986);
nor U12729 (N_12729,N_11451,N_11886);
nand U12730 (N_12730,N_11989,N_11733);
or U12731 (N_12731,N_11324,N_11614);
nand U12732 (N_12732,N_11672,N_11684);
nand U12733 (N_12733,N_11340,N_11373);
nor U12734 (N_12734,N_11455,N_11662);
or U12735 (N_12735,N_11921,N_11926);
nor U12736 (N_12736,N_11537,N_11440);
or U12737 (N_12737,N_11459,N_11450);
xnor U12738 (N_12738,N_11816,N_11812);
and U12739 (N_12739,N_11525,N_11361);
xnor U12740 (N_12740,N_11832,N_11945);
and U12741 (N_12741,N_11878,N_11488);
and U12742 (N_12742,N_11296,N_11478);
or U12743 (N_12743,N_11387,N_11627);
nor U12744 (N_12744,N_11733,N_11985);
nor U12745 (N_12745,N_11644,N_11745);
xor U12746 (N_12746,N_11777,N_11469);
nand U12747 (N_12747,N_11912,N_11351);
and U12748 (N_12748,N_11773,N_11548);
or U12749 (N_12749,N_11822,N_11812);
xnor U12750 (N_12750,N_12010,N_12019);
or U12751 (N_12751,N_12582,N_12489);
xnor U12752 (N_12752,N_12468,N_12435);
or U12753 (N_12753,N_12202,N_12702);
xor U12754 (N_12754,N_12369,N_12555);
or U12755 (N_12755,N_12340,N_12673);
or U12756 (N_12756,N_12033,N_12532);
or U12757 (N_12757,N_12520,N_12235);
and U12758 (N_12758,N_12306,N_12691);
or U12759 (N_12759,N_12545,N_12635);
and U12760 (N_12760,N_12368,N_12497);
nand U12761 (N_12761,N_12571,N_12097);
or U12762 (N_12762,N_12357,N_12240);
or U12763 (N_12763,N_12507,N_12102);
nor U12764 (N_12764,N_12709,N_12644);
nor U12765 (N_12765,N_12243,N_12004);
and U12766 (N_12766,N_12650,N_12111);
and U12767 (N_12767,N_12136,N_12621);
nand U12768 (N_12768,N_12364,N_12351);
and U12769 (N_12769,N_12182,N_12190);
nor U12770 (N_12770,N_12050,N_12409);
nand U12771 (N_12771,N_12261,N_12365);
xor U12772 (N_12772,N_12639,N_12200);
or U12773 (N_12773,N_12230,N_12397);
nor U12774 (N_12774,N_12001,N_12616);
nor U12775 (N_12775,N_12177,N_12407);
nor U12776 (N_12776,N_12228,N_12653);
and U12777 (N_12777,N_12484,N_12331);
nor U12778 (N_12778,N_12370,N_12375);
and U12779 (N_12779,N_12557,N_12374);
or U12780 (N_12780,N_12419,N_12104);
or U12781 (N_12781,N_12335,N_12494);
and U12782 (N_12782,N_12637,N_12056);
and U12783 (N_12783,N_12605,N_12062);
and U12784 (N_12784,N_12137,N_12508);
nand U12785 (N_12785,N_12721,N_12444);
nand U12786 (N_12786,N_12147,N_12543);
and U12787 (N_12787,N_12611,N_12420);
and U12788 (N_12788,N_12149,N_12451);
or U12789 (N_12789,N_12246,N_12713);
nand U12790 (N_12790,N_12126,N_12201);
or U12791 (N_12791,N_12674,N_12633);
nor U12792 (N_12792,N_12417,N_12712);
nor U12793 (N_12793,N_12334,N_12135);
and U12794 (N_12794,N_12423,N_12130);
xor U12795 (N_12795,N_12692,N_12167);
nor U12796 (N_12796,N_12474,N_12382);
nor U12797 (N_12797,N_12502,N_12552);
and U12798 (N_12798,N_12366,N_12522);
xor U12799 (N_12799,N_12092,N_12448);
and U12800 (N_12800,N_12666,N_12481);
nor U12801 (N_12801,N_12677,N_12400);
xor U12802 (N_12802,N_12363,N_12421);
and U12803 (N_12803,N_12378,N_12689);
nand U12804 (N_12804,N_12372,N_12734);
or U12805 (N_12805,N_12081,N_12008);
or U12806 (N_12806,N_12082,N_12337);
xnor U12807 (N_12807,N_12745,N_12128);
xnor U12808 (N_12808,N_12730,N_12003);
xor U12809 (N_12809,N_12184,N_12722);
nand U12810 (N_12810,N_12453,N_12452);
or U12811 (N_12811,N_12257,N_12185);
nor U12812 (N_12812,N_12509,N_12120);
nand U12813 (N_12813,N_12096,N_12477);
or U12814 (N_12814,N_12099,N_12029);
nand U12815 (N_12815,N_12274,N_12353);
and U12816 (N_12816,N_12410,N_12226);
or U12817 (N_12817,N_12715,N_12112);
or U12818 (N_12818,N_12500,N_12179);
xnor U12819 (N_12819,N_12017,N_12704);
and U12820 (N_12820,N_12441,N_12401);
and U12821 (N_12821,N_12160,N_12627);
or U12822 (N_12822,N_12040,N_12649);
nand U12823 (N_12823,N_12744,N_12558);
nand U12824 (N_12824,N_12073,N_12089);
nand U12825 (N_12825,N_12381,N_12586);
nor U12826 (N_12826,N_12476,N_12269);
or U12827 (N_12827,N_12318,N_12594);
nand U12828 (N_12828,N_12101,N_12483);
xor U12829 (N_12829,N_12268,N_12422);
and U12830 (N_12830,N_12525,N_12169);
nor U12831 (N_12831,N_12032,N_12161);
xor U12832 (N_12832,N_12542,N_12654);
and U12833 (N_12833,N_12630,N_12186);
or U12834 (N_12834,N_12678,N_12292);
xnor U12835 (N_12835,N_12675,N_12533);
nand U12836 (N_12836,N_12220,N_12505);
xor U12837 (N_12837,N_12232,N_12071);
nand U12838 (N_12838,N_12205,N_12206);
xnor U12839 (N_12839,N_12255,N_12242);
and U12840 (N_12840,N_12562,N_12597);
nor U12841 (N_12841,N_12224,N_12581);
nor U12842 (N_12842,N_12229,N_12035);
nand U12843 (N_12843,N_12356,N_12253);
nand U12844 (N_12844,N_12325,N_12203);
nor U12845 (N_12845,N_12574,N_12227);
nor U12846 (N_12846,N_12643,N_12113);
nor U12847 (N_12847,N_12701,N_12090);
xnor U12848 (N_12848,N_12563,N_12659);
xor U12849 (N_12849,N_12194,N_12516);
and U12850 (N_12850,N_12345,N_12125);
nor U12851 (N_12851,N_12188,N_12303);
and U12852 (N_12852,N_12640,N_12736);
or U12853 (N_12853,N_12433,N_12030);
and U12854 (N_12854,N_12593,N_12168);
nand U12855 (N_12855,N_12540,N_12612);
and U12856 (N_12856,N_12214,N_12121);
and U12857 (N_12857,N_12454,N_12068);
nand U12858 (N_12858,N_12725,N_12287);
nor U12859 (N_12859,N_12462,N_12596);
or U12860 (N_12860,N_12283,N_12385);
xor U12861 (N_12861,N_12060,N_12549);
or U12862 (N_12862,N_12459,N_12642);
nor U12863 (N_12863,N_12355,N_12157);
and U12864 (N_12864,N_12426,N_12587);
xnor U12865 (N_12865,N_12607,N_12100);
xor U12866 (N_12866,N_12084,N_12564);
or U12867 (N_12867,N_12732,N_12519);
nor U12868 (N_12868,N_12020,N_12670);
nor U12869 (N_12869,N_12580,N_12150);
nand U12870 (N_12870,N_12265,N_12272);
nand U12871 (N_12871,N_12387,N_12620);
nor U12872 (N_12872,N_12350,N_12626);
and U12873 (N_12873,N_12535,N_12195);
nand U12874 (N_12874,N_12389,N_12648);
and U12875 (N_12875,N_12687,N_12493);
nand U12876 (N_12876,N_12395,N_12191);
xnor U12877 (N_12877,N_12314,N_12298);
and U12878 (N_12878,N_12538,N_12039);
or U12879 (N_12879,N_12609,N_12601);
or U12880 (N_12880,N_12207,N_12221);
nor U12881 (N_12881,N_12367,N_12339);
nand U12882 (N_12882,N_12002,N_12405);
nor U12883 (N_12883,N_12399,N_12492);
nand U12884 (N_12884,N_12480,N_12568);
or U12885 (N_12885,N_12037,N_12553);
and U12886 (N_12886,N_12437,N_12748);
nor U12887 (N_12887,N_12544,N_12313);
nor U12888 (N_12888,N_12290,N_12438);
and U12889 (N_12889,N_12731,N_12264);
and U12890 (N_12890,N_12210,N_12672);
nor U12891 (N_12891,N_12067,N_12436);
nand U12892 (N_12892,N_12212,N_12371);
and U12893 (N_12893,N_12280,N_12373);
nor U12894 (N_12894,N_12153,N_12131);
xor U12895 (N_12895,N_12647,N_12416);
nor U12896 (N_12896,N_12000,N_12254);
and U12897 (N_12897,N_12527,N_12077);
nor U12898 (N_12898,N_12315,N_12379);
and U12899 (N_12899,N_12565,N_12457);
or U12900 (N_12900,N_12536,N_12295);
or U12901 (N_12901,N_12575,N_12349);
and U12902 (N_12902,N_12384,N_12139);
or U12903 (N_12903,N_12718,N_12332);
xor U12904 (N_12904,N_12170,N_12576);
nor U12905 (N_12905,N_12348,N_12152);
and U12906 (N_12906,N_12663,N_12259);
nand U12907 (N_12907,N_12324,N_12471);
or U12908 (N_12908,N_12705,N_12510);
nor U12909 (N_12909,N_12110,N_12703);
or U12910 (N_12910,N_12107,N_12052);
xnor U12911 (N_12911,N_12219,N_12260);
or U12912 (N_12912,N_12258,N_12078);
or U12913 (N_12913,N_12218,N_12708);
or U12914 (N_12914,N_12682,N_12386);
and U12915 (N_12915,N_12449,N_12285);
and U12916 (N_12916,N_12693,N_12178);
nor U12917 (N_12917,N_12733,N_12487);
or U12918 (N_12918,N_12662,N_12541);
and U12919 (N_12919,N_12415,N_12531);
or U12920 (N_12920,N_12529,N_12144);
nor U12921 (N_12921,N_12720,N_12430);
xor U12922 (N_12922,N_12041,N_12236);
or U12923 (N_12923,N_12684,N_12685);
nor U12924 (N_12924,N_12589,N_12171);
xnor U12925 (N_12925,N_12636,N_12512);
nand U12926 (N_12926,N_12239,N_12700);
nor U12927 (N_12927,N_12223,N_12641);
nand U12928 (N_12928,N_12049,N_12667);
or U12929 (N_12929,N_12276,N_12294);
nor U12930 (N_12930,N_12479,N_12045);
and U12931 (N_12931,N_12517,N_12180);
nor U12932 (N_12932,N_12284,N_12066);
and U12933 (N_12933,N_12572,N_12461);
nand U12934 (N_12934,N_12727,N_12076);
xnor U12935 (N_12935,N_12263,N_12183);
xnor U12936 (N_12936,N_12065,N_12646);
and U12937 (N_12937,N_12679,N_12117);
nand U12938 (N_12938,N_12301,N_12598);
and U12939 (N_12939,N_12523,N_12455);
and U12940 (N_12940,N_12322,N_12070);
and U12941 (N_12941,N_12083,N_12015);
nor U12942 (N_12942,N_12310,N_12606);
xor U12943 (N_12943,N_12312,N_12323);
and U12944 (N_12944,N_12726,N_12442);
nand U12945 (N_12945,N_12034,N_12025);
nand U12946 (N_12946,N_12634,N_12600);
and U12947 (N_12947,N_12012,N_12539);
nand U12948 (N_12948,N_12446,N_12354);
nand U12949 (N_12949,N_12059,N_12584);
or U12950 (N_12950,N_12680,N_12450);
nor U12951 (N_12951,N_12087,N_12380);
and U12952 (N_12952,N_12724,N_12208);
and U12953 (N_12953,N_12173,N_12159);
nor U12954 (N_12954,N_12316,N_12164);
or U12955 (N_12955,N_12115,N_12391);
or U12956 (N_12956,N_12463,N_12573);
and U12957 (N_12957,N_12628,N_12602);
or U12958 (N_12958,N_12683,N_12638);
nor U12959 (N_12959,N_12028,N_12105);
nor U12960 (N_12960,N_12749,N_12222);
xor U12961 (N_12961,N_12114,N_12281);
and U12962 (N_12962,N_12559,N_12016);
nor U12963 (N_12963,N_12618,N_12515);
nor U12964 (N_12964,N_12664,N_12406);
or U12965 (N_12965,N_12554,N_12155);
nor U12966 (N_12966,N_12362,N_12590);
nand U12967 (N_12967,N_12005,N_12079);
and U12968 (N_12968,N_12530,N_12022);
or U12969 (N_12969,N_12342,N_12352);
and U12970 (N_12970,N_12176,N_12424);
or U12971 (N_12971,N_12319,N_12737);
and U12972 (N_12972,N_12645,N_12622);
or U12973 (N_12973,N_12490,N_12696);
nand U12974 (N_12974,N_12439,N_12109);
xnor U12975 (N_12975,N_12729,N_12361);
or U12976 (N_12976,N_12244,N_12192);
xnor U12977 (N_12977,N_12690,N_12418);
nor U12978 (N_12978,N_12311,N_12278);
or U12979 (N_12979,N_12556,N_12506);
xnor U12980 (N_12980,N_12328,N_12098);
and U12981 (N_12981,N_12093,N_12614);
and U12982 (N_12982,N_12140,N_12069);
nand U12983 (N_12983,N_12181,N_12617);
xor U12984 (N_12984,N_12163,N_12404);
nand U12985 (N_12985,N_12695,N_12009);
nor U12986 (N_12986,N_12583,N_12247);
xor U12987 (N_12987,N_12534,N_12036);
nand U12988 (N_12988,N_12706,N_12688);
xnor U12989 (N_12989,N_12566,N_12347);
and U12990 (N_12990,N_12189,N_12528);
xor U12991 (N_12991,N_12570,N_12716);
nor U12992 (N_12992,N_12495,N_12046);
nor U12993 (N_12993,N_12344,N_12445);
nor U12994 (N_12994,N_12658,N_12055);
or U12995 (N_12995,N_12469,N_12127);
and U12996 (N_12996,N_12482,N_12216);
nor U12997 (N_12997,N_12669,N_12403);
or U12998 (N_12998,N_12699,N_12485);
and U12999 (N_12999,N_12146,N_12498);
nor U13000 (N_13000,N_12021,N_12051);
nor U13001 (N_13001,N_12333,N_12151);
xor U13002 (N_13002,N_12320,N_12133);
nor U13003 (N_13003,N_12376,N_12198);
nand U13004 (N_13004,N_12251,N_12063);
nor U13005 (N_13005,N_12624,N_12383);
nor U13006 (N_13006,N_12546,N_12697);
nand U13007 (N_13007,N_12359,N_12388);
or U13008 (N_13008,N_12657,N_12631);
nand U13009 (N_13009,N_12511,N_12377);
xor U13010 (N_13010,N_12560,N_12158);
and U13011 (N_13011,N_12739,N_12300);
nand U13012 (N_13012,N_12698,N_12478);
nor U13013 (N_13013,N_12141,N_12307);
nor U13014 (N_13014,N_12551,N_12209);
or U13015 (N_13015,N_12156,N_12547);
nor U13016 (N_13016,N_12148,N_12393);
nor U13017 (N_13017,N_12488,N_12305);
or U13018 (N_13018,N_12579,N_12585);
xor U13019 (N_13019,N_12526,N_12486);
and U13020 (N_13020,N_12231,N_12327);
nand U13021 (N_13021,N_12175,N_12714);
nor U13022 (N_13022,N_12042,N_12217);
xor U13023 (N_13023,N_12738,N_12668);
nor U13024 (N_13024,N_12123,N_12094);
nand U13025 (N_13025,N_12743,N_12694);
or U13026 (N_13026,N_12431,N_12047);
xor U13027 (N_13027,N_12610,N_12129);
nor U13028 (N_13028,N_12427,N_12719);
nor U13029 (N_13029,N_12432,N_12723);
nor U13030 (N_13030,N_12475,N_12711);
xor U13031 (N_13031,N_12023,N_12308);
xor U13032 (N_13032,N_12599,N_12728);
nor U13033 (N_13033,N_12262,N_12499);
nand U13034 (N_13034,N_12007,N_12613);
or U13035 (N_13035,N_12241,N_12443);
nand U13036 (N_13036,N_12414,N_12116);
nor U13037 (N_13037,N_12011,N_12304);
nor U13038 (N_13038,N_12501,N_12248);
or U13039 (N_13039,N_12425,N_12266);
and U13040 (N_13040,N_12317,N_12142);
and U13041 (N_13041,N_12548,N_12103);
xnor U13042 (N_13042,N_12465,N_12651);
and U13043 (N_13043,N_12595,N_12473);
and U13044 (N_13044,N_12604,N_12740);
and U13045 (N_13045,N_12245,N_12411);
or U13046 (N_13046,N_12686,N_12119);
nand U13047 (N_13047,N_12394,N_12237);
nor U13048 (N_13048,N_12271,N_12434);
and U13049 (N_13049,N_12655,N_12013);
or U13050 (N_13050,N_12398,N_12024);
nor U13051 (N_13051,N_12085,N_12429);
nand U13052 (N_13052,N_12326,N_12681);
nand U13053 (N_13053,N_12569,N_12741);
xnor U13054 (N_13054,N_12252,N_12336);
and U13055 (N_13055,N_12632,N_12591);
and U13056 (N_13056,N_12309,N_12625);
nand U13057 (N_13057,N_12145,N_12249);
and U13058 (N_13058,N_12166,N_12619);
nor U13059 (N_13059,N_12256,N_12118);
nor U13060 (N_13060,N_12031,N_12286);
xnor U13061 (N_13061,N_12018,N_12456);
nor U13062 (N_13062,N_12057,N_12058);
or U13063 (N_13063,N_12006,N_12088);
nor U13064 (N_13064,N_12472,N_12134);
and U13065 (N_13065,N_12282,N_12108);
nor U13066 (N_13066,N_12338,N_12291);
or U13067 (N_13067,N_12615,N_12124);
nand U13068 (N_13068,N_12233,N_12289);
and U13069 (N_13069,N_12661,N_12106);
nor U13070 (N_13070,N_12048,N_12402);
xnor U13071 (N_13071,N_12143,N_12458);
nand U13072 (N_13072,N_12464,N_12080);
or U13073 (N_13073,N_12747,N_12413);
and U13074 (N_13074,N_12054,N_12196);
nor U13075 (N_13075,N_12267,N_12428);
or U13076 (N_13076,N_12710,N_12504);
nand U13077 (N_13077,N_12717,N_12038);
nor U13078 (N_13078,N_12392,N_12341);
nor U13079 (N_13079,N_12250,N_12652);
xnor U13080 (N_13080,N_12412,N_12296);
and U13081 (N_13081,N_12225,N_12466);
or U13082 (N_13082,N_12467,N_12578);
or U13083 (N_13083,N_12470,N_12238);
nor U13084 (N_13084,N_12321,N_12293);
and U13085 (N_13085,N_12358,N_12608);
or U13086 (N_13086,N_12279,N_12091);
nor U13087 (N_13087,N_12288,N_12676);
nand U13088 (N_13088,N_12302,N_12027);
and U13089 (N_13089,N_12656,N_12273);
xor U13090 (N_13090,N_12588,N_12270);
or U13091 (N_13091,N_12199,N_12440);
or U13092 (N_13092,N_12213,N_12174);
nand U13093 (N_13093,N_12074,N_12053);
or U13094 (N_13094,N_12577,N_12043);
xor U13095 (N_13095,N_12197,N_12396);
xor U13096 (N_13096,N_12521,N_12503);
nor U13097 (N_13097,N_12044,N_12561);
nor U13098 (N_13098,N_12603,N_12162);
nor U13099 (N_13099,N_12095,N_12447);
or U13100 (N_13100,N_12623,N_12707);
nor U13101 (N_13101,N_12026,N_12204);
xnor U13102 (N_13102,N_12660,N_12671);
or U13103 (N_13103,N_12215,N_12343);
or U13104 (N_13104,N_12408,N_12496);
nor U13105 (N_13105,N_12132,N_12172);
and U13106 (N_13106,N_12346,N_12187);
nand U13107 (N_13107,N_12742,N_12360);
and U13108 (N_13108,N_12629,N_12138);
nand U13109 (N_13109,N_12211,N_12275);
and U13110 (N_13110,N_12329,N_12075);
nor U13111 (N_13111,N_12014,N_12537);
or U13112 (N_13112,N_12299,N_12061);
or U13113 (N_13113,N_12330,N_12234);
or U13114 (N_13114,N_12514,N_12064);
or U13115 (N_13115,N_12524,N_12072);
nor U13116 (N_13116,N_12154,N_12277);
xor U13117 (N_13117,N_12491,N_12122);
xor U13118 (N_13118,N_12735,N_12567);
xor U13119 (N_13119,N_12665,N_12513);
or U13120 (N_13120,N_12550,N_12165);
nand U13121 (N_13121,N_12297,N_12746);
and U13122 (N_13122,N_12390,N_12086);
nand U13123 (N_13123,N_12193,N_12518);
or U13124 (N_13124,N_12592,N_12460);
nand U13125 (N_13125,N_12446,N_12312);
or U13126 (N_13126,N_12240,N_12461);
and U13127 (N_13127,N_12609,N_12160);
xor U13128 (N_13128,N_12116,N_12172);
and U13129 (N_13129,N_12165,N_12612);
or U13130 (N_13130,N_12194,N_12665);
nand U13131 (N_13131,N_12467,N_12618);
nor U13132 (N_13132,N_12662,N_12394);
nor U13133 (N_13133,N_12005,N_12481);
and U13134 (N_13134,N_12504,N_12002);
nand U13135 (N_13135,N_12650,N_12542);
or U13136 (N_13136,N_12479,N_12650);
nand U13137 (N_13137,N_12008,N_12438);
or U13138 (N_13138,N_12631,N_12362);
and U13139 (N_13139,N_12342,N_12188);
nor U13140 (N_13140,N_12128,N_12606);
and U13141 (N_13141,N_12193,N_12066);
xor U13142 (N_13142,N_12730,N_12421);
xnor U13143 (N_13143,N_12315,N_12414);
and U13144 (N_13144,N_12412,N_12432);
and U13145 (N_13145,N_12248,N_12227);
and U13146 (N_13146,N_12096,N_12217);
xnor U13147 (N_13147,N_12356,N_12437);
nand U13148 (N_13148,N_12131,N_12147);
and U13149 (N_13149,N_12155,N_12419);
nand U13150 (N_13150,N_12072,N_12405);
and U13151 (N_13151,N_12210,N_12700);
nor U13152 (N_13152,N_12556,N_12587);
xnor U13153 (N_13153,N_12457,N_12550);
or U13154 (N_13154,N_12162,N_12215);
and U13155 (N_13155,N_12201,N_12268);
and U13156 (N_13156,N_12342,N_12451);
nand U13157 (N_13157,N_12722,N_12077);
nand U13158 (N_13158,N_12617,N_12488);
xnor U13159 (N_13159,N_12096,N_12049);
and U13160 (N_13160,N_12233,N_12484);
nand U13161 (N_13161,N_12608,N_12260);
nor U13162 (N_13162,N_12433,N_12517);
and U13163 (N_13163,N_12645,N_12589);
nor U13164 (N_13164,N_12432,N_12138);
xnor U13165 (N_13165,N_12658,N_12031);
and U13166 (N_13166,N_12412,N_12670);
or U13167 (N_13167,N_12380,N_12326);
xnor U13168 (N_13168,N_12677,N_12512);
and U13169 (N_13169,N_12044,N_12265);
nand U13170 (N_13170,N_12704,N_12063);
nand U13171 (N_13171,N_12047,N_12244);
nand U13172 (N_13172,N_12562,N_12063);
or U13173 (N_13173,N_12510,N_12695);
or U13174 (N_13174,N_12473,N_12532);
xor U13175 (N_13175,N_12337,N_12735);
xnor U13176 (N_13176,N_12175,N_12651);
nor U13177 (N_13177,N_12671,N_12728);
and U13178 (N_13178,N_12136,N_12422);
nand U13179 (N_13179,N_12447,N_12348);
nand U13180 (N_13180,N_12431,N_12093);
nand U13181 (N_13181,N_12499,N_12613);
xnor U13182 (N_13182,N_12695,N_12574);
nand U13183 (N_13183,N_12172,N_12642);
and U13184 (N_13184,N_12336,N_12259);
or U13185 (N_13185,N_12331,N_12536);
and U13186 (N_13186,N_12644,N_12364);
and U13187 (N_13187,N_12185,N_12123);
xnor U13188 (N_13188,N_12007,N_12093);
xor U13189 (N_13189,N_12517,N_12355);
nor U13190 (N_13190,N_12039,N_12329);
and U13191 (N_13191,N_12162,N_12322);
nor U13192 (N_13192,N_12633,N_12560);
nor U13193 (N_13193,N_12175,N_12426);
and U13194 (N_13194,N_12224,N_12497);
nor U13195 (N_13195,N_12643,N_12693);
xnor U13196 (N_13196,N_12215,N_12210);
or U13197 (N_13197,N_12330,N_12389);
nor U13198 (N_13198,N_12468,N_12270);
xnor U13199 (N_13199,N_12029,N_12476);
nor U13200 (N_13200,N_12373,N_12377);
or U13201 (N_13201,N_12332,N_12317);
or U13202 (N_13202,N_12083,N_12624);
or U13203 (N_13203,N_12455,N_12203);
xnor U13204 (N_13204,N_12403,N_12124);
nand U13205 (N_13205,N_12088,N_12278);
nand U13206 (N_13206,N_12723,N_12550);
nand U13207 (N_13207,N_12377,N_12157);
xor U13208 (N_13208,N_12428,N_12623);
xnor U13209 (N_13209,N_12049,N_12214);
nor U13210 (N_13210,N_12379,N_12288);
nand U13211 (N_13211,N_12139,N_12719);
nor U13212 (N_13212,N_12207,N_12687);
nor U13213 (N_13213,N_12545,N_12114);
or U13214 (N_13214,N_12348,N_12419);
nand U13215 (N_13215,N_12545,N_12484);
nor U13216 (N_13216,N_12724,N_12386);
and U13217 (N_13217,N_12338,N_12433);
nor U13218 (N_13218,N_12526,N_12718);
xor U13219 (N_13219,N_12155,N_12584);
xnor U13220 (N_13220,N_12732,N_12462);
xnor U13221 (N_13221,N_12158,N_12371);
nor U13222 (N_13222,N_12278,N_12353);
nand U13223 (N_13223,N_12144,N_12679);
nand U13224 (N_13224,N_12421,N_12731);
xnor U13225 (N_13225,N_12663,N_12695);
or U13226 (N_13226,N_12543,N_12010);
xor U13227 (N_13227,N_12527,N_12154);
nand U13228 (N_13228,N_12142,N_12390);
or U13229 (N_13229,N_12610,N_12439);
nand U13230 (N_13230,N_12294,N_12307);
xnor U13231 (N_13231,N_12051,N_12134);
and U13232 (N_13232,N_12484,N_12063);
and U13233 (N_13233,N_12444,N_12104);
and U13234 (N_13234,N_12172,N_12559);
nor U13235 (N_13235,N_12456,N_12550);
xnor U13236 (N_13236,N_12479,N_12513);
or U13237 (N_13237,N_12148,N_12240);
or U13238 (N_13238,N_12496,N_12132);
and U13239 (N_13239,N_12002,N_12725);
xnor U13240 (N_13240,N_12310,N_12053);
and U13241 (N_13241,N_12472,N_12169);
nor U13242 (N_13242,N_12400,N_12454);
and U13243 (N_13243,N_12334,N_12575);
and U13244 (N_13244,N_12122,N_12195);
nor U13245 (N_13245,N_12436,N_12221);
nand U13246 (N_13246,N_12672,N_12584);
xnor U13247 (N_13247,N_12625,N_12387);
and U13248 (N_13248,N_12533,N_12725);
and U13249 (N_13249,N_12333,N_12069);
and U13250 (N_13250,N_12031,N_12293);
xnor U13251 (N_13251,N_12538,N_12730);
xnor U13252 (N_13252,N_12709,N_12134);
nor U13253 (N_13253,N_12044,N_12477);
or U13254 (N_13254,N_12736,N_12697);
nor U13255 (N_13255,N_12010,N_12395);
and U13256 (N_13256,N_12429,N_12384);
or U13257 (N_13257,N_12697,N_12039);
nor U13258 (N_13258,N_12119,N_12571);
or U13259 (N_13259,N_12303,N_12557);
and U13260 (N_13260,N_12686,N_12307);
and U13261 (N_13261,N_12468,N_12410);
and U13262 (N_13262,N_12632,N_12354);
and U13263 (N_13263,N_12327,N_12246);
nand U13264 (N_13264,N_12362,N_12661);
xnor U13265 (N_13265,N_12163,N_12443);
xnor U13266 (N_13266,N_12375,N_12705);
nand U13267 (N_13267,N_12174,N_12357);
and U13268 (N_13268,N_12251,N_12312);
nand U13269 (N_13269,N_12005,N_12389);
or U13270 (N_13270,N_12359,N_12512);
and U13271 (N_13271,N_12013,N_12642);
and U13272 (N_13272,N_12088,N_12276);
nand U13273 (N_13273,N_12718,N_12625);
or U13274 (N_13274,N_12449,N_12453);
xor U13275 (N_13275,N_12676,N_12307);
nor U13276 (N_13276,N_12649,N_12227);
and U13277 (N_13277,N_12676,N_12265);
nor U13278 (N_13278,N_12223,N_12474);
nand U13279 (N_13279,N_12326,N_12530);
and U13280 (N_13280,N_12318,N_12474);
nor U13281 (N_13281,N_12721,N_12294);
xnor U13282 (N_13282,N_12352,N_12524);
xnor U13283 (N_13283,N_12052,N_12262);
xnor U13284 (N_13284,N_12625,N_12481);
nand U13285 (N_13285,N_12259,N_12664);
xnor U13286 (N_13286,N_12313,N_12695);
nand U13287 (N_13287,N_12647,N_12106);
and U13288 (N_13288,N_12451,N_12416);
or U13289 (N_13289,N_12704,N_12567);
and U13290 (N_13290,N_12082,N_12175);
and U13291 (N_13291,N_12304,N_12710);
nor U13292 (N_13292,N_12698,N_12534);
nand U13293 (N_13293,N_12583,N_12286);
or U13294 (N_13294,N_12400,N_12197);
and U13295 (N_13295,N_12577,N_12178);
nor U13296 (N_13296,N_12411,N_12026);
and U13297 (N_13297,N_12572,N_12348);
nand U13298 (N_13298,N_12133,N_12435);
or U13299 (N_13299,N_12659,N_12749);
nor U13300 (N_13300,N_12528,N_12561);
nand U13301 (N_13301,N_12665,N_12454);
xor U13302 (N_13302,N_12309,N_12253);
and U13303 (N_13303,N_12471,N_12299);
nor U13304 (N_13304,N_12563,N_12452);
or U13305 (N_13305,N_12529,N_12173);
xor U13306 (N_13306,N_12550,N_12070);
or U13307 (N_13307,N_12708,N_12199);
or U13308 (N_13308,N_12666,N_12733);
nand U13309 (N_13309,N_12273,N_12124);
or U13310 (N_13310,N_12620,N_12316);
nand U13311 (N_13311,N_12629,N_12331);
xor U13312 (N_13312,N_12189,N_12675);
xor U13313 (N_13313,N_12075,N_12551);
and U13314 (N_13314,N_12541,N_12202);
nand U13315 (N_13315,N_12046,N_12269);
and U13316 (N_13316,N_12657,N_12155);
nor U13317 (N_13317,N_12334,N_12140);
xnor U13318 (N_13318,N_12337,N_12169);
nand U13319 (N_13319,N_12073,N_12653);
or U13320 (N_13320,N_12688,N_12321);
nand U13321 (N_13321,N_12579,N_12023);
or U13322 (N_13322,N_12614,N_12256);
and U13323 (N_13323,N_12668,N_12496);
or U13324 (N_13324,N_12445,N_12266);
or U13325 (N_13325,N_12588,N_12272);
or U13326 (N_13326,N_12290,N_12689);
and U13327 (N_13327,N_12470,N_12411);
xnor U13328 (N_13328,N_12570,N_12089);
nand U13329 (N_13329,N_12675,N_12551);
and U13330 (N_13330,N_12594,N_12348);
nor U13331 (N_13331,N_12259,N_12567);
or U13332 (N_13332,N_12236,N_12639);
nor U13333 (N_13333,N_12139,N_12009);
xor U13334 (N_13334,N_12078,N_12350);
or U13335 (N_13335,N_12228,N_12196);
xor U13336 (N_13336,N_12711,N_12388);
or U13337 (N_13337,N_12428,N_12090);
and U13338 (N_13338,N_12030,N_12256);
and U13339 (N_13339,N_12191,N_12676);
or U13340 (N_13340,N_12239,N_12631);
and U13341 (N_13341,N_12462,N_12414);
nand U13342 (N_13342,N_12360,N_12217);
and U13343 (N_13343,N_12627,N_12093);
and U13344 (N_13344,N_12701,N_12389);
nand U13345 (N_13345,N_12675,N_12116);
nand U13346 (N_13346,N_12728,N_12144);
xor U13347 (N_13347,N_12316,N_12704);
nand U13348 (N_13348,N_12324,N_12598);
or U13349 (N_13349,N_12631,N_12178);
or U13350 (N_13350,N_12245,N_12051);
nor U13351 (N_13351,N_12431,N_12168);
or U13352 (N_13352,N_12725,N_12239);
and U13353 (N_13353,N_12077,N_12719);
and U13354 (N_13354,N_12259,N_12337);
nand U13355 (N_13355,N_12615,N_12237);
xnor U13356 (N_13356,N_12541,N_12322);
nand U13357 (N_13357,N_12634,N_12063);
and U13358 (N_13358,N_12671,N_12323);
xnor U13359 (N_13359,N_12618,N_12367);
nor U13360 (N_13360,N_12595,N_12104);
and U13361 (N_13361,N_12074,N_12226);
and U13362 (N_13362,N_12467,N_12044);
nor U13363 (N_13363,N_12115,N_12074);
nand U13364 (N_13364,N_12073,N_12122);
xnor U13365 (N_13365,N_12085,N_12114);
nor U13366 (N_13366,N_12734,N_12015);
nor U13367 (N_13367,N_12339,N_12615);
xnor U13368 (N_13368,N_12701,N_12017);
or U13369 (N_13369,N_12027,N_12047);
nor U13370 (N_13370,N_12556,N_12694);
nand U13371 (N_13371,N_12334,N_12114);
nor U13372 (N_13372,N_12148,N_12314);
nand U13373 (N_13373,N_12234,N_12298);
and U13374 (N_13374,N_12535,N_12001);
or U13375 (N_13375,N_12618,N_12478);
and U13376 (N_13376,N_12677,N_12207);
nand U13377 (N_13377,N_12452,N_12241);
nor U13378 (N_13378,N_12144,N_12498);
nand U13379 (N_13379,N_12106,N_12214);
nor U13380 (N_13380,N_12062,N_12259);
and U13381 (N_13381,N_12748,N_12269);
xor U13382 (N_13382,N_12128,N_12018);
nand U13383 (N_13383,N_12641,N_12362);
nand U13384 (N_13384,N_12355,N_12573);
nand U13385 (N_13385,N_12328,N_12307);
nor U13386 (N_13386,N_12004,N_12143);
xor U13387 (N_13387,N_12230,N_12702);
or U13388 (N_13388,N_12122,N_12582);
xor U13389 (N_13389,N_12345,N_12746);
and U13390 (N_13390,N_12584,N_12081);
nand U13391 (N_13391,N_12482,N_12045);
nor U13392 (N_13392,N_12636,N_12418);
nor U13393 (N_13393,N_12741,N_12598);
xnor U13394 (N_13394,N_12536,N_12491);
or U13395 (N_13395,N_12536,N_12459);
and U13396 (N_13396,N_12353,N_12707);
xor U13397 (N_13397,N_12553,N_12401);
nor U13398 (N_13398,N_12303,N_12209);
nor U13399 (N_13399,N_12203,N_12041);
and U13400 (N_13400,N_12367,N_12727);
nand U13401 (N_13401,N_12390,N_12353);
nand U13402 (N_13402,N_12131,N_12517);
nand U13403 (N_13403,N_12438,N_12539);
xor U13404 (N_13404,N_12552,N_12586);
nor U13405 (N_13405,N_12576,N_12595);
xnor U13406 (N_13406,N_12076,N_12534);
nor U13407 (N_13407,N_12636,N_12619);
nor U13408 (N_13408,N_12656,N_12489);
nor U13409 (N_13409,N_12468,N_12351);
and U13410 (N_13410,N_12481,N_12418);
nand U13411 (N_13411,N_12198,N_12596);
or U13412 (N_13412,N_12297,N_12098);
or U13413 (N_13413,N_12618,N_12504);
and U13414 (N_13414,N_12514,N_12362);
nand U13415 (N_13415,N_12531,N_12704);
or U13416 (N_13416,N_12705,N_12081);
and U13417 (N_13417,N_12564,N_12519);
nand U13418 (N_13418,N_12613,N_12070);
nor U13419 (N_13419,N_12391,N_12412);
and U13420 (N_13420,N_12715,N_12681);
xor U13421 (N_13421,N_12705,N_12147);
nor U13422 (N_13422,N_12114,N_12686);
nand U13423 (N_13423,N_12418,N_12584);
or U13424 (N_13424,N_12247,N_12236);
or U13425 (N_13425,N_12646,N_12434);
nor U13426 (N_13426,N_12201,N_12108);
or U13427 (N_13427,N_12728,N_12294);
or U13428 (N_13428,N_12290,N_12375);
nand U13429 (N_13429,N_12050,N_12544);
nand U13430 (N_13430,N_12129,N_12502);
or U13431 (N_13431,N_12486,N_12650);
nor U13432 (N_13432,N_12690,N_12653);
or U13433 (N_13433,N_12287,N_12081);
or U13434 (N_13434,N_12221,N_12346);
nand U13435 (N_13435,N_12274,N_12519);
nand U13436 (N_13436,N_12621,N_12715);
nand U13437 (N_13437,N_12462,N_12513);
or U13438 (N_13438,N_12316,N_12510);
and U13439 (N_13439,N_12228,N_12188);
xnor U13440 (N_13440,N_12169,N_12282);
nor U13441 (N_13441,N_12620,N_12708);
nor U13442 (N_13442,N_12167,N_12087);
or U13443 (N_13443,N_12084,N_12037);
nand U13444 (N_13444,N_12246,N_12594);
and U13445 (N_13445,N_12542,N_12254);
or U13446 (N_13446,N_12500,N_12541);
nor U13447 (N_13447,N_12162,N_12721);
nand U13448 (N_13448,N_12479,N_12030);
nand U13449 (N_13449,N_12487,N_12636);
nand U13450 (N_13450,N_12674,N_12133);
xor U13451 (N_13451,N_12229,N_12360);
nor U13452 (N_13452,N_12135,N_12046);
or U13453 (N_13453,N_12349,N_12425);
nor U13454 (N_13454,N_12547,N_12649);
nand U13455 (N_13455,N_12368,N_12462);
and U13456 (N_13456,N_12665,N_12634);
and U13457 (N_13457,N_12520,N_12339);
nand U13458 (N_13458,N_12103,N_12175);
xor U13459 (N_13459,N_12316,N_12467);
nor U13460 (N_13460,N_12230,N_12663);
or U13461 (N_13461,N_12453,N_12631);
or U13462 (N_13462,N_12059,N_12498);
xnor U13463 (N_13463,N_12169,N_12674);
or U13464 (N_13464,N_12328,N_12573);
xor U13465 (N_13465,N_12238,N_12609);
and U13466 (N_13466,N_12144,N_12028);
nor U13467 (N_13467,N_12677,N_12605);
xor U13468 (N_13468,N_12558,N_12049);
xnor U13469 (N_13469,N_12380,N_12249);
and U13470 (N_13470,N_12280,N_12622);
xor U13471 (N_13471,N_12220,N_12487);
nand U13472 (N_13472,N_12336,N_12067);
or U13473 (N_13473,N_12580,N_12032);
nor U13474 (N_13474,N_12357,N_12053);
nor U13475 (N_13475,N_12384,N_12012);
xor U13476 (N_13476,N_12462,N_12243);
nand U13477 (N_13477,N_12069,N_12437);
or U13478 (N_13478,N_12380,N_12491);
nor U13479 (N_13479,N_12726,N_12559);
nand U13480 (N_13480,N_12356,N_12357);
or U13481 (N_13481,N_12141,N_12722);
or U13482 (N_13482,N_12037,N_12167);
nor U13483 (N_13483,N_12086,N_12459);
and U13484 (N_13484,N_12011,N_12143);
and U13485 (N_13485,N_12681,N_12639);
xnor U13486 (N_13486,N_12047,N_12432);
or U13487 (N_13487,N_12340,N_12699);
nor U13488 (N_13488,N_12217,N_12187);
nand U13489 (N_13489,N_12096,N_12399);
nand U13490 (N_13490,N_12364,N_12336);
xor U13491 (N_13491,N_12226,N_12042);
and U13492 (N_13492,N_12195,N_12425);
nor U13493 (N_13493,N_12205,N_12615);
nor U13494 (N_13494,N_12336,N_12140);
or U13495 (N_13495,N_12516,N_12274);
xor U13496 (N_13496,N_12349,N_12717);
nand U13497 (N_13497,N_12083,N_12547);
or U13498 (N_13498,N_12161,N_12477);
or U13499 (N_13499,N_12102,N_12099);
nor U13500 (N_13500,N_13043,N_13289);
nand U13501 (N_13501,N_12786,N_13339);
xnor U13502 (N_13502,N_12782,N_12957);
or U13503 (N_13503,N_12986,N_13297);
or U13504 (N_13504,N_13257,N_13458);
and U13505 (N_13505,N_13016,N_13116);
xnor U13506 (N_13506,N_13120,N_12959);
nor U13507 (N_13507,N_13060,N_13171);
or U13508 (N_13508,N_12921,N_12886);
xnor U13509 (N_13509,N_12754,N_13184);
nand U13510 (N_13510,N_13360,N_13266);
xor U13511 (N_13511,N_13051,N_13274);
xnor U13512 (N_13512,N_13209,N_12814);
nand U13513 (N_13513,N_13306,N_13372);
xor U13514 (N_13514,N_13149,N_13211);
nand U13515 (N_13515,N_13197,N_13110);
nor U13516 (N_13516,N_12811,N_13026);
xor U13517 (N_13517,N_13053,N_13041);
nor U13518 (N_13518,N_13292,N_13454);
nor U13519 (N_13519,N_12777,N_13222);
or U13520 (N_13520,N_13400,N_13334);
and U13521 (N_13521,N_13245,N_13300);
and U13522 (N_13522,N_13384,N_12845);
or U13523 (N_13523,N_13188,N_13073);
and U13524 (N_13524,N_13457,N_13336);
or U13525 (N_13525,N_13392,N_12912);
and U13526 (N_13526,N_13276,N_13240);
xor U13527 (N_13527,N_12828,N_12996);
nor U13528 (N_13528,N_13479,N_13040);
xor U13529 (N_13529,N_13082,N_13196);
nor U13530 (N_13530,N_13439,N_12929);
nor U13531 (N_13531,N_12830,N_13282);
nand U13532 (N_13532,N_12968,N_13452);
or U13533 (N_13533,N_12893,N_13168);
or U13534 (N_13534,N_12881,N_13448);
nor U13535 (N_13535,N_13288,N_12988);
xor U13536 (N_13536,N_12859,N_13337);
xor U13537 (N_13537,N_12755,N_13150);
and U13538 (N_13538,N_13286,N_13258);
nand U13539 (N_13539,N_12823,N_13461);
and U13540 (N_13540,N_13230,N_12948);
nand U13541 (N_13541,N_12846,N_13017);
or U13542 (N_13542,N_12788,N_13371);
xnor U13543 (N_13543,N_13355,N_12756);
xor U13544 (N_13544,N_13162,N_12961);
or U13545 (N_13545,N_12888,N_12861);
nand U13546 (N_13546,N_12834,N_12910);
nand U13547 (N_13547,N_13233,N_12764);
nand U13548 (N_13548,N_13363,N_12776);
and U13549 (N_13549,N_12971,N_13054);
nand U13550 (N_13550,N_13343,N_13381);
and U13551 (N_13551,N_13057,N_13158);
nand U13552 (N_13552,N_12796,N_13025);
or U13553 (N_13553,N_12994,N_12752);
and U13554 (N_13554,N_13156,N_13304);
or U13555 (N_13555,N_13335,N_12839);
xnor U13556 (N_13556,N_12938,N_13011);
xnor U13557 (N_13557,N_13079,N_13242);
nor U13558 (N_13558,N_13291,N_12915);
nand U13559 (N_13559,N_12805,N_12891);
nor U13560 (N_13560,N_12867,N_12821);
and U13561 (N_13561,N_13071,N_13200);
or U13562 (N_13562,N_13256,N_13208);
xor U13563 (N_13563,N_13191,N_12972);
or U13564 (N_13564,N_13166,N_12887);
nand U13565 (N_13565,N_12779,N_13278);
nor U13566 (N_13566,N_13409,N_13492);
and U13567 (N_13567,N_13103,N_12781);
xnor U13568 (N_13568,N_12880,N_13024);
nand U13569 (N_13569,N_12984,N_12843);
or U13570 (N_13570,N_13033,N_13391);
nor U13571 (N_13571,N_12815,N_13421);
nand U13572 (N_13572,N_12758,N_12765);
nand U13573 (N_13573,N_13499,N_13124);
xnor U13574 (N_13574,N_12790,N_12901);
or U13575 (N_13575,N_12979,N_12899);
xnor U13576 (N_13576,N_13248,N_13204);
and U13577 (N_13577,N_13497,N_13189);
nand U13578 (N_13578,N_13318,N_12847);
xor U13579 (N_13579,N_12759,N_13126);
xor U13580 (N_13580,N_13213,N_13219);
nor U13581 (N_13581,N_12851,N_13078);
or U13582 (N_13582,N_12930,N_13093);
xor U13583 (N_13583,N_13022,N_13013);
nand U13584 (N_13584,N_12762,N_12939);
nand U13585 (N_13585,N_13021,N_13344);
and U13586 (N_13586,N_13405,N_13307);
and U13587 (N_13587,N_13161,N_12772);
xnor U13588 (N_13588,N_12833,N_13345);
nand U13589 (N_13589,N_12985,N_13328);
xor U13590 (N_13590,N_13244,N_13128);
and U13591 (N_13591,N_13473,N_13032);
nand U13592 (N_13592,N_12974,N_13396);
xor U13593 (N_13593,N_13246,N_13359);
and U13594 (N_13594,N_13046,N_13069);
and U13595 (N_13595,N_12991,N_12773);
or U13596 (N_13596,N_13283,N_13450);
and U13597 (N_13597,N_12969,N_13305);
xnor U13598 (N_13598,N_12956,N_13481);
xor U13599 (N_13599,N_13420,N_12873);
xor U13600 (N_13600,N_12935,N_12826);
and U13601 (N_13601,N_13068,N_13349);
and U13602 (N_13602,N_12941,N_13401);
nor U13603 (N_13603,N_13379,N_12934);
and U13604 (N_13604,N_12866,N_13139);
and U13605 (N_13605,N_13399,N_12852);
xor U13606 (N_13606,N_13098,N_12778);
and U13607 (N_13607,N_12923,N_12835);
xnor U13608 (N_13608,N_13027,N_12952);
and U13609 (N_13609,N_13395,N_13111);
nand U13610 (N_13610,N_12919,N_13152);
nand U13611 (N_13611,N_13247,N_13353);
and U13612 (N_13612,N_13301,N_13085);
xor U13613 (N_13613,N_13309,N_13169);
xnor U13614 (N_13614,N_12962,N_13470);
nor U13615 (N_13615,N_13218,N_12883);
or U13616 (N_13616,N_13472,N_13020);
or U13617 (N_13617,N_13327,N_12937);
nor U13618 (N_13618,N_13004,N_12989);
xnor U13619 (N_13619,N_13005,N_13207);
xor U13620 (N_13620,N_13322,N_13142);
or U13621 (N_13621,N_12854,N_13319);
xor U13622 (N_13622,N_13469,N_13096);
or U13623 (N_13623,N_13066,N_12841);
nand U13624 (N_13624,N_13237,N_13133);
nand U13625 (N_13625,N_12768,N_12973);
nor U13626 (N_13626,N_12848,N_13403);
nand U13627 (N_13627,N_12897,N_12884);
or U13628 (N_13628,N_12797,N_12920);
xor U13629 (N_13629,N_13329,N_12840);
xnor U13630 (N_13630,N_13100,N_13270);
and U13631 (N_13631,N_13157,N_12760);
xor U13632 (N_13632,N_13127,N_13195);
and U13633 (N_13633,N_13387,N_13351);
xnor U13634 (N_13634,N_13170,N_13296);
nand U13635 (N_13635,N_13368,N_12949);
and U13636 (N_13636,N_12855,N_13357);
or U13637 (N_13637,N_12770,N_12983);
nand U13638 (N_13638,N_13007,N_12990);
xnor U13639 (N_13639,N_12872,N_13455);
or U13640 (N_13640,N_13378,N_13178);
nand U13641 (N_13641,N_12791,N_13147);
and U13642 (N_13642,N_13003,N_12998);
and U13643 (N_13643,N_13036,N_12947);
and U13644 (N_13644,N_12864,N_12799);
nor U13645 (N_13645,N_13284,N_13431);
xnor U13646 (N_13646,N_13084,N_12775);
nand U13647 (N_13647,N_13061,N_13348);
nand U13648 (N_13648,N_13221,N_12785);
xor U13649 (N_13649,N_13143,N_13261);
xnor U13650 (N_13650,N_12812,N_13125);
and U13651 (N_13651,N_13201,N_12900);
nor U13652 (N_13652,N_12806,N_13310);
xor U13653 (N_13653,N_13228,N_13052);
nor U13654 (N_13654,N_13251,N_13480);
or U13655 (N_13655,N_13267,N_12964);
xor U13656 (N_13656,N_13364,N_12831);
nand U13657 (N_13657,N_12824,N_13373);
and U13658 (N_13658,N_12896,N_12829);
nand U13659 (N_13659,N_13000,N_13441);
nand U13660 (N_13660,N_13175,N_13308);
nand U13661 (N_13661,N_12951,N_13179);
nor U13662 (N_13662,N_12783,N_12774);
xor U13663 (N_13663,N_12955,N_12943);
xor U13664 (N_13664,N_13253,N_13148);
xor U13665 (N_13665,N_12795,N_12810);
and U13666 (N_13666,N_13214,N_13451);
nor U13667 (N_13667,N_12763,N_13031);
or U13668 (N_13668,N_12863,N_13056);
xnor U13669 (N_13669,N_13092,N_12794);
nand U13670 (N_13670,N_13101,N_13440);
nor U13671 (N_13671,N_13366,N_13141);
nand U13672 (N_13672,N_13490,N_13476);
nand U13673 (N_13673,N_13235,N_13465);
or U13674 (N_13674,N_12885,N_13122);
xnor U13675 (N_13675,N_13065,N_13239);
and U13676 (N_13676,N_13315,N_13193);
xor U13677 (N_13677,N_13462,N_13155);
xor U13678 (N_13678,N_13427,N_12928);
nor U13679 (N_13679,N_13483,N_13097);
or U13680 (N_13680,N_13159,N_13181);
and U13681 (N_13681,N_12789,N_13134);
xor U13682 (N_13682,N_13446,N_13443);
and U13683 (N_13683,N_13397,N_13482);
nand U13684 (N_13684,N_13095,N_13123);
nor U13685 (N_13685,N_12987,N_13419);
nor U13686 (N_13686,N_13486,N_13418);
nor U13687 (N_13687,N_13252,N_13114);
and U13688 (N_13688,N_13295,N_13478);
or U13689 (N_13689,N_12967,N_13434);
and U13690 (N_13690,N_12903,N_12879);
or U13691 (N_13691,N_13338,N_13199);
nor U13692 (N_13692,N_13394,N_13416);
nor U13693 (N_13693,N_13254,N_13102);
and U13694 (N_13694,N_13393,N_12818);
or U13695 (N_13695,N_13493,N_13165);
or U13696 (N_13696,N_13390,N_13176);
or U13697 (N_13697,N_12849,N_12932);
or U13698 (N_13698,N_12793,N_12958);
and U13699 (N_13699,N_12890,N_13186);
nor U13700 (N_13700,N_12960,N_13112);
and U13701 (N_13701,N_13090,N_13070);
nor U13702 (N_13702,N_13019,N_13398);
nor U13703 (N_13703,N_13311,N_13108);
nor U13704 (N_13704,N_13280,N_12917);
and U13705 (N_13705,N_12945,N_12808);
xor U13706 (N_13706,N_12819,N_12942);
and U13707 (N_13707,N_13049,N_13410);
or U13708 (N_13708,N_13365,N_13350);
or U13709 (N_13709,N_13340,N_12950);
and U13710 (N_13710,N_13081,N_13389);
nor U13711 (N_13711,N_13263,N_13223);
nand U13712 (N_13712,N_13272,N_13277);
nand U13713 (N_13713,N_13456,N_13488);
or U13714 (N_13714,N_13382,N_13487);
nand U13715 (N_13715,N_13153,N_13083);
nand U13716 (N_13716,N_13442,N_12817);
xor U13717 (N_13717,N_13411,N_13109);
or U13718 (N_13718,N_12944,N_12980);
nand U13719 (N_13719,N_12902,N_12875);
xnor U13720 (N_13720,N_13225,N_13113);
xor U13721 (N_13721,N_13136,N_13015);
xor U13722 (N_13722,N_12853,N_12822);
nand U13723 (N_13723,N_13323,N_13055);
xor U13724 (N_13724,N_13231,N_13459);
nand U13725 (N_13725,N_13115,N_13206);
or U13726 (N_13726,N_13002,N_13279);
or U13727 (N_13727,N_13494,N_13063);
xnor U13728 (N_13728,N_12933,N_13467);
nor U13729 (N_13729,N_13135,N_13151);
xnor U13730 (N_13730,N_13466,N_13173);
nor U13731 (N_13731,N_13058,N_13062);
xnor U13732 (N_13732,N_13485,N_12892);
or U13733 (N_13733,N_13273,N_13413);
nand U13734 (N_13734,N_12865,N_13265);
and U13735 (N_13735,N_13302,N_13435);
and U13736 (N_13736,N_12750,N_12911);
xnor U13737 (N_13737,N_12757,N_12850);
nor U13738 (N_13738,N_13331,N_13038);
nand U13739 (N_13739,N_13006,N_13474);
and U13740 (N_13740,N_13077,N_13080);
nor U13741 (N_13741,N_13496,N_13298);
nand U13742 (N_13742,N_13034,N_12769);
nor U13743 (N_13743,N_12992,N_13106);
nor U13744 (N_13744,N_13180,N_12954);
nand U13745 (N_13745,N_12981,N_12807);
and U13746 (N_13746,N_12842,N_12771);
nor U13747 (N_13747,N_13330,N_13243);
nand U13748 (N_13748,N_12792,N_13138);
or U13749 (N_13749,N_13172,N_13198);
or U13750 (N_13750,N_13075,N_13464);
xor U13751 (N_13751,N_13259,N_12976);
or U13752 (N_13752,N_13471,N_12836);
nor U13753 (N_13753,N_13121,N_13119);
or U13754 (N_13754,N_12925,N_13453);
and U13755 (N_13755,N_13303,N_13447);
or U13756 (N_13756,N_12860,N_12761);
xnor U13757 (N_13757,N_13491,N_13424);
nand U13758 (N_13758,N_12978,N_12918);
or U13759 (N_13759,N_13341,N_13160);
nor U13760 (N_13760,N_12993,N_12907);
and U13761 (N_13761,N_12837,N_13285);
nor U13762 (N_13762,N_12898,N_13324);
xor U13763 (N_13763,N_13294,N_13406);
or U13764 (N_13764,N_13129,N_12787);
nor U13765 (N_13765,N_13187,N_12926);
or U13766 (N_13766,N_13087,N_13347);
and U13767 (N_13767,N_13316,N_13463);
and U13768 (N_13768,N_13037,N_13313);
xnor U13769 (N_13769,N_12904,N_13354);
nand U13770 (N_13770,N_12905,N_13192);
nand U13771 (N_13771,N_13249,N_13074);
xnor U13772 (N_13772,N_13131,N_12780);
or U13773 (N_13773,N_13388,N_12946);
and U13774 (N_13774,N_12800,N_13072);
nor U13775 (N_13775,N_12827,N_13226);
nor U13776 (N_13776,N_12868,N_13414);
and U13777 (N_13777,N_12894,N_12965);
nor U13778 (N_13778,N_13203,N_13432);
nor U13779 (N_13779,N_13210,N_13383);
nand U13780 (N_13780,N_13099,N_13408);
and U13781 (N_13781,N_13425,N_13234);
nor U13782 (N_13782,N_13346,N_12816);
xor U13783 (N_13783,N_13012,N_13132);
and U13784 (N_13784,N_12832,N_13437);
nand U13785 (N_13785,N_13029,N_13352);
and U13786 (N_13786,N_13385,N_12895);
nand U13787 (N_13787,N_13023,N_13404);
nand U13788 (N_13788,N_12982,N_13001);
nor U13789 (N_13789,N_12878,N_13386);
and U13790 (N_13790,N_13264,N_13047);
or U13791 (N_13791,N_12809,N_12995);
nand U13792 (N_13792,N_13140,N_13216);
xor U13793 (N_13793,N_13380,N_12999);
and U13794 (N_13794,N_13118,N_13255);
and U13795 (N_13795,N_13361,N_13444);
or U13796 (N_13796,N_12963,N_13104);
or U13797 (N_13797,N_13164,N_12876);
nand U13798 (N_13798,N_12767,N_13039);
xnor U13799 (N_13799,N_13333,N_13402);
nand U13800 (N_13800,N_13215,N_13174);
nor U13801 (N_13801,N_12820,N_13250);
or U13802 (N_13802,N_13362,N_13241);
nor U13803 (N_13803,N_13375,N_12862);
xnor U13804 (N_13804,N_12825,N_13048);
and U13805 (N_13805,N_13317,N_13287);
or U13806 (N_13806,N_13194,N_13426);
and U13807 (N_13807,N_12977,N_12844);
nor U13808 (N_13808,N_13144,N_13460);
and U13809 (N_13809,N_13260,N_13088);
nor U13810 (N_13810,N_12813,N_12856);
nor U13811 (N_13811,N_13202,N_13167);
xnor U13812 (N_13812,N_12751,N_13227);
xnor U13813 (N_13813,N_12924,N_13275);
nor U13814 (N_13814,N_13477,N_13436);
and U13815 (N_13815,N_12975,N_12857);
and U13816 (N_13816,N_12922,N_13212);
or U13817 (N_13817,N_13137,N_12906);
and U13818 (N_13818,N_13367,N_13177);
nor U13819 (N_13819,N_13205,N_12798);
nand U13820 (N_13820,N_12801,N_13190);
nor U13821 (N_13821,N_13429,N_13091);
and U13822 (N_13822,N_12909,N_13089);
or U13823 (N_13823,N_12908,N_13430);
nand U13824 (N_13824,N_13008,N_13030);
xor U13825 (N_13825,N_13484,N_13018);
xor U13826 (N_13826,N_13045,N_13094);
or U13827 (N_13827,N_13183,N_13042);
or U13828 (N_13828,N_12874,N_13224);
nor U13829 (N_13829,N_13417,N_13332);
and U13830 (N_13830,N_13412,N_13236);
xnor U13831 (N_13831,N_13064,N_12803);
nand U13832 (N_13832,N_12914,N_13154);
nand U13833 (N_13833,N_13067,N_13076);
nor U13834 (N_13834,N_13369,N_13445);
nand U13835 (N_13835,N_12940,N_13238);
xor U13836 (N_13836,N_13314,N_12871);
or U13837 (N_13837,N_13423,N_13107);
xor U13838 (N_13838,N_13358,N_13342);
or U13839 (N_13839,N_12953,N_13105);
nor U13840 (N_13840,N_13312,N_13325);
and U13841 (N_13841,N_13262,N_13009);
or U13842 (N_13842,N_13182,N_13290);
nor U13843 (N_13843,N_12838,N_13415);
and U13844 (N_13844,N_13163,N_13229);
xnor U13845 (N_13845,N_13146,N_12916);
nand U13846 (N_13846,N_13468,N_13326);
xor U13847 (N_13847,N_13475,N_13374);
or U13848 (N_13848,N_12870,N_13281);
or U13849 (N_13849,N_12766,N_13428);
and U13850 (N_13850,N_12913,N_12877);
and U13851 (N_13851,N_13044,N_13271);
xor U13852 (N_13852,N_13498,N_12997);
or U13853 (N_13853,N_13422,N_13299);
nand U13854 (N_13854,N_13035,N_12804);
nor U13855 (N_13855,N_13117,N_12753);
nand U13856 (N_13856,N_12927,N_13449);
nand U13857 (N_13857,N_13433,N_13028);
nor U13858 (N_13858,N_12802,N_13268);
or U13859 (N_13859,N_12931,N_13320);
xnor U13860 (N_13860,N_13407,N_13014);
nor U13861 (N_13861,N_12966,N_12869);
or U13862 (N_13862,N_13370,N_12970);
nor U13863 (N_13863,N_13232,N_12882);
nor U13864 (N_13864,N_13185,N_13376);
and U13865 (N_13865,N_12784,N_13356);
nor U13866 (N_13866,N_13377,N_13293);
xor U13867 (N_13867,N_13220,N_13059);
nand U13868 (N_13868,N_13050,N_13086);
nand U13869 (N_13869,N_13438,N_12936);
nor U13870 (N_13870,N_13130,N_13495);
nor U13871 (N_13871,N_13321,N_13010);
and U13872 (N_13872,N_12858,N_13217);
or U13873 (N_13873,N_13269,N_13145);
and U13874 (N_13874,N_12889,N_13489);
nand U13875 (N_13875,N_13290,N_13201);
nand U13876 (N_13876,N_13087,N_13071);
nand U13877 (N_13877,N_13210,N_13248);
nand U13878 (N_13878,N_12818,N_13047);
or U13879 (N_13879,N_13416,N_13468);
or U13880 (N_13880,N_12953,N_12904);
nor U13881 (N_13881,N_13155,N_13055);
xor U13882 (N_13882,N_12890,N_13105);
nor U13883 (N_13883,N_12934,N_13221);
or U13884 (N_13884,N_13070,N_13301);
xnor U13885 (N_13885,N_12750,N_12882);
nor U13886 (N_13886,N_12884,N_13415);
and U13887 (N_13887,N_13198,N_13279);
or U13888 (N_13888,N_13454,N_12941);
xor U13889 (N_13889,N_13323,N_12922);
or U13890 (N_13890,N_13282,N_12819);
nor U13891 (N_13891,N_13081,N_12784);
and U13892 (N_13892,N_12760,N_13305);
xnor U13893 (N_13893,N_13196,N_13091);
nand U13894 (N_13894,N_12766,N_12925);
nor U13895 (N_13895,N_13443,N_13362);
or U13896 (N_13896,N_13229,N_13271);
and U13897 (N_13897,N_13348,N_13403);
nor U13898 (N_13898,N_12987,N_13168);
nand U13899 (N_13899,N_13183,N_12863);
or U13900 (N_13900,N_12826,N_13073);
xor U13901 (N_13901,N_12987,N_12871);
nand U13902 (N_13902,N_13459,N_13114);
and U13903 (N_13903,N_13467,N_13144);
nor U13904 (N_13904,N_13406,N_13278);
nor U13905 (N_13905,N_13050,N_13401);
xnor U13906 (N_13906,N_12985,N_13139);
nand U13907 (N_13907,N_12807,N_13082);
or U13908 (N_13908,N_12750,N_13080);
nor U13909 (N_13909,N_13278,N_13334);
xor U13910 (N_13910,N_13454,N_13436);
nor U13911 (N_13911,N_13254,N_13004);
or U13912 (N_13912,N_13094,N_12980);
xnor U13913 (N_13913,N_13005,N_13464);
xnor U13914 (N_13914,N_13059,N_13362);
or U13915 (N_13915,N_13324,N_13143);
nand U13916 (N_13916,N_13314,N_13469);
nand U13917 (N_13917,N_13487,N_13388);
and U13918 (N_13918,N_13165,N_12775);
and U13919 (N_13919,N_12820,N_13020);
nand U13920 (N_13920,N_13427,N_12961);
and U13921 (N_13921,N_13017,N_13349);
nand U13922 (N_13922,N_13233,N_13135);
nand U13923 (N_13923,N_13045,N_13258);
xnor U13924 (N_13924,N_13291,N_12890);
or U13925 (N_13925,N_12787,N_12798);
and U13926 (N_13926,N_13450,N_12891);
xnor U13927 (N_13927,N_12855,N_13335);
nand U13928 (N_13928,N_13398,N_13357);
nor U13929 (N_13929,N_13029,N_13051);
and U13930 (N_13930,N_12896,N_13013);
nor U13931 (N_13931,N_12918,N_13003);
nor U13932 (N_13932,N_12893,N_12959);
nand U13933 (N_13933,N_12982,N_12782);
or U13934 (N_13934,N_12897,N_13063);
nand U13935 (N_13935,N_13191,N_13384);
xor U13936 (N_13936,N_13454,N_13217);
nand U13937 (N_13937,N_13375,N_13312);
nor U13938 (N_13938,N_13058,N_13265);
nand U13939 (N_13939,N_13344,N_13271);
xnor U13940 (N_13940,N_13492,N_12983);
nor U13941 (N_13941,N_13311,N_13478);
and U13942 (N_13942,N_13285,N_12861);
xor U13943 (N_13943,N_13431,N_12750);
and U13944 (N_13944,N_13074,N_12931);
xor U13945 (N_13945,N_13485,N_13060);
and U13946 (N_13946,N_13272,N_13322);
and U13947 (N_13947,N_12958,N_12972);
or U13948 (N_13948,N_12947,N_13333);
or U13949 (N_13949,N_12765,N_13165);
nor U13950 (N_13950,N_13169,N_13490);
xnor U13951 (N_13951,N_12817,N_13008);
nand U13952 (N_13952,N_13374,N_13122);
and U13953 (N_13953,N_13147,N_13310);
xor U13954 (N_13954,N_13110,N_12991);
or U13955 (N_13955,N_12795,N_13051);
and U13956 (N_13956,N_12874,N_13368);
and U13957 (N_13957,N_13190,N_12988);
and U13958 (N_13958,N_12976,N_12914);
nor U13959 (N_13959,N_12931,N_12871);
nand U13960 (N_13960,N_12763,N_13486);
and U13961 (N_13961,N_13139,N_12803);
xnor U13962 (N_13962,N_12957,N_13424);
or U13963 (N_13963,N_12979,N_13398);
xnor U13964 (N_13964,N_12818,N_13332);
or U13965 (N_13965,N_13262,N_13136);
nor U13966 (N_13966,N_12787,N_13246);
and U13967 (N_13967,N_12802,N_13301);
or U13968 (N_13968,N_13167,N_13070);
xor U13969 (N_13969,N_13266,N_13480);
nand U13970 (N_13970,N_13133,N_13058);
xnor U13971 (N_13971,N_13039,N_13196);
xnor U13972 (N_13972,N_12921,N_13352);
nand U13973 (N_13973,N_13496,N_13499);
nand U13974 (N_13974,N_12856,N_12919);
or U13975 (N_13975,N_13076,N_13025);
nor U13976 (N_13976,N_13158,N_13440);
nand U13977 (N_13977,N_13034,N_13495);
xnor U13978 (N_13978,N_13335,N_12841);
nand U13979 (N_13979,N_13347,N_13061);
or U13980 (N_13980,N_13016,N_13469);
and U13981 (N_13981,N_13001,N_13430);
or U13982 (N_13982,N_13314,N_13234);
nor U13983 (N_13983,N_13347,N_13364);
nand U13984 (N_13984,N_13469,N_13437);
xor U13985 (N_13985,N_12783,N_13033);
and U13986 (N_13986,N_12809,N_12988);
or U13987 (N_13987,N_13133,N_13449);
xor U13988 (N_13988,N_12823,N_13138);
xnor U13989 (N_13989,N_12755,N_13431);
nand U13990 (N_13990,N_12945,N_13022);
nor U13991 (N_13991,N_12874,N_13357);
nand U13992 (N_13992,N_13085,N_13479);
or U13993 (N_13993,N_12824,N_12989);
and U13994 (N_13994,N_13057,N_13135);
and U13995 (N_13995,N_13481,N_13010);
or U13996 (N_13996,N_12830,N_13372);
and U13997 (N_13997,N_12936,N_12859);
or U13998 (N_13998,N_13266,N_12966);
or U13999 (N_13999,N_13398,N_12976);
nand U14000 (N_14000,N_12828,N_13316);
nor U14001 (N_14001,N_13041,N_13428);
xor U14002 (N_14002,N_13209,N_13018);
nor U14003 (N_14003,N_13437,N_13174);
or U14004 (N_14004,N_13478,N_13373);
nor U14005 (N_14005,N_13303,N_12786);
nand U14006 (N_14006,N_13161,N_13198);
nor U14007 (N_14007,N_13190,N_13055);
nand U14008 (N_14008,N_12951,N_12788);
or U14009 (N_14009,N_12896,N_12810);
xor U14010 (N_14010,N_12953,N_13043);
nand U14011 (N_14011,N_13402,N_13454);
and U14012 (N_14012,N_13233,N_13126);
or U14013 (N_14013,N_12836,N_12762);
and U14014 (N_14014,N_12999,N_12845);
xor U14015 (N_14015,N_13225,N_13473);
or U14016 (N_14016,N_12954,N_12869);
nor U14017 (N_14017,N_13342,N_12939);
nand U14018 (N_14018,N_13118,N_12782);
or U14019 (N_14019,N_12818,N_12877);
xnor U14020 (N_14020,N_12930,N_13230);
or U14021 (N_14021,N_12803,N_12848);
or U14022 (N_14022,N_12960,N_13461);
xnor U14023 (N_14023,N_13002,N_13063);
xnor U14024 (N_14024,N_13226,N_12909);
xnor U14025 (N_14025,N_13137,N_13110);
or U14026 (N_14026,N_13073,N_13055);
and U14027 (N_14027,N_13379,N_12757);
and U14028 (N_14028,N_13137,N_13028);
xnor U14029 (N_14029,N_13228,N_13477);
xor U14030 (N_14030,N_13248,N_13008);
nor U14031 (N_14031,N_13474,N_13015);
nand U14032 (N_14032,N_12884,N_13173);
xnor U14033 (N_14033,N_13379,N_13048);
xor U14034 (N_14034,N_13386,N_13140);
xor U14035 (N_14035,N_13153,N_13315);
nor U14036 (N_14036,N_13479,N_13174);
xnor U14037 (N_14037,N_12849,N_13107);
xnor U14038 (N_14038,N_12945,N_13013);
and U14039 (N_14039,N_13241,N_13413);
or U14040 (N_14040,N_13084,N_13040);
and U14041 (N_14041,N_13357,N_13458);
nor U14042 (N_14042,N_12992,N_13208);
or U14043 (N_14043,N_13017,N_13174);
xnor U14044 (N_14044,N_13028,N_13284);
xnor U14045 (N_14045,N_13333,N_12800);
nor U14046 (N_14046,N_13471,N_13243);
xor U14047 (N_14047,N_12934,N_12918);
or U14048 (N_14048,N_12953,N_13005);
and U14049 (N_14049,N_12975,N_12995);
or U14050 (N_14050,N_12900,N_13225);
and U14051 (N_14051,N_13077,N_12755);
nor U14052 (N_14052,N_13175,N_13440);
and U14053 (N_14053,N_12915,N_13403);
nor U14054 (N_14054,N_13062,N_12977);
nand U14055 (N_14055,N_12877,N_13277);
or U14056 (N_14056,N_13157,N_12850);
xnor U14057 (N_14057,N_13264,N_13386);
or U14058 (N_14058,N_12868,N_13498);
and U14059 (N_14059,N_13143,N_13292);
xor U14060 (N_14060,N_13422,N_13343);
or U14061 (N_14061,N_13139,N_13263);
xnor U14062 (N_14062,N_12945,N_12846);
xnor U14063 (N_14063,N_12912,N_12781);
and U14064 (N_14064,N_13022,N_13473);
or U14065 (N_14065,N_13002,N_13439);
nor U14066 (N_14066,N_13240,N_13039);
nand U14067 (N_14067,N_13489,N_13456);
or U14068 (N_14068,N_12803,N_13268);
and U14069 (N_14069,N_12884,N_12933);
nand U14070 (N_14070,N_12844,N_13000);
and U14071 (N_14071,N_13315,N_13102);
nand U14072 (N_14072,N_13070,N_12815);
xnor U14073 (N_14073,N_13410,N_13421);
xor U14074 (N_14074,N_13460,N_13275);
nand U14075 (N_14075,N_13442,N_12792);
xnor U14076 (N_14076,N_12947,N_13390);
or U14077 (N_14077,N_13019,N_13165);
xor U14078 (N_14078,N_12937,N_12877);
or U14079 (N_14079,N_13054,N_13198);
xnor U14080 (N_14080,N_13334,N_13199);
nand U14081 (N_14081,N_13006,N_12762);
or U14082 (N_14082,N_12780,N_12888);
nand U14083 (N_14083,N_13111,N_13176);
or U14084 (N_14084,N_12909,N_13122);
and U14085 (N_14085,N_13291,N_12763);
xnor U14086 (N_14086,N_13298,N_12986);
xor U14087 (N_14087,N_13392,N_13295);
xor U14088 (N_14088,N_13335,N_13201);
nor U14089 (N_14089,N_13060,N_13362);
or U14090 (N_14090,N_13081,N_13040);
and U14091 (N_14091,N_12763,N_13044);
and U14092 (N_14092,N_13205,N_13332);
xor U14093 (N_14093,N_12919,N_13250);
and U14094 (N_14094,N_13313,N_12932);
or U14095 (N_14095,N_12872,N_13481);
nand U14096 (N_14096,N_12806,N_12907);
or U14097 (N_14097,N_13011,N_13071);
nor U14098 (N_14098,N_13115,N_13065);
nor U14099 (N_14099,N_13178,N_13409);
xor U14100 (N_14100,N_13206,N_12901);
xnor U14101 (N_14101,N_13426,N_12970);
nor U14102 (N_14102,N_12900,N_13068);
or U14103 (N_14103,N_13008,N_12786);
xor U14104 (N_14104,N_13077,N_12880);
xnor U14105 (N_14105,N_13004,N_12895);
xnor U14106 (N_14106,N_13184,N_12975);
nor U14107 (N_14107,N_13350,N_13088);
and U14108 (N_14108,N_12771,N_13145);
or U14109 (N_14109,N_12946,N_13119);
nor U14110 (N_14110,N_13306,N_12837);
xnor U14111 (N_14111,N_13142,N_13000);
nor U14112 (N_14112,N_13218,N_13168);
nor U14113 (N_14113,N_13481,N_12841);
nor U14114 (N_14114,N_13366,N_13099);
xor U14115 (N_14115,N_12865,N_12885);
and U14116 (N_14116,N_13074,N_12862);
xnor U14117 (N_14117,N_12893,N_12888);
nor U14118 (N_14118,N_13498,N_12895);
nand U14119 (N_14119,N_12788,N_13062);
xor U14120 (N_14120,N_13289,N_13072);
nor U14121 (N_14121,N_13391,N_13343);
and U14122 (N_14122,N_12976,N_13456);
xnor U14123 (N_14123,N_13172,N_12752);
nand U14124 (N_14124,N_13234,N_13033);
nand U14125 (N_14125,N_13188,N_12913);
nor U14126 (N_14126,N_13046,N_12848);
xnor U14127 (N_14127,N_13093,N_12818);
and U14128 (N_14128,N_13318,N_12876);
nand U14129 (N_14129,N_13465,N_13163);
or U14130 (N_14130,N_13193,N_13076);
xor U14131 (N_14131,N_13076,N_13368);
xnor U14132 (N_14132,N_12869,N_12947);
nand U14133 (N_14133,N_13127,N_13212);
and U14134 (N_14134,N_13104,N_13169);
and U14135 (N_14135,N_13256,N_13447);
or U14136 (N_14136,N_12785,N_12857);
xor U14137 (N_14137,N_13042,N_12994);
xnor U14138 (N_14138,N_13357,N_12966);
xor U14139 (N_14139,N_13230,N_12892);
and U14140 (N_14140,N_12989,N_13368);
nor U14141 (N_14141,N_13423,N_13492);
or U14142 (N_14142,N_12877,N_13390);
nand U14143 (N_14143,N_13086,N_13410);
nand U14144 (N_14144,N_13286,N_13070);
nand U14145 (N_14145,N_13116,N_12755);
nand U14146 (N_14146,N_13232,N_13263);
nand U14147 (N_14147,N_12936,N_12750);
or U14148 (N_14148,N_13211,N_13289);
and U14149 (N_14149,N_13013,N_12890);
nor U14150 (N_14150,N_13434,N_13235);
and U14151 (N_14151,N_13235,N_13075);
xnor U14152 (N_14152,N_13311,N_12963);
nor U14153 (N_14153,N_13253,N_13325);
or U14154 (N_14154,N_13197,N_13454);
nor U14155 (N_14155,N_12814,N_13174);
and U14156 (N_14156,N_13302,N_13240);
nor U14157 (N_14157,N_13447,N_13446);
nor U14158 (N_14158,N_12857,N_13125);
nor U14159 (N_14159,N_13411,N_12801);
and U14160 (N_14160,N_13414,N_12787);
xor U14161 (N_14161,N_13256,N_13244);
and U14162 (N_14162,N_12866,N_13315);
xnor U14163 (N_14163,N_12782,N_13424);
or U14164 (N_14164,N_13027,N_13190);
nand U14165 (N_14165,N_13474,N_13185);
nor U14166 (N_14166,N_13424,N_13066);
and U14167 (N_14167,N_12922,N_12943);
nand U14168 (N_14168,N_12822,N_12995);
and U14169 (N_14169,N_13397,N_13306);
or U14170 (N_14170,N_12960,N_12999);
nor U14171 (N_14171,N_13222,N_13361);
nand U14172 (N_14172,N_12833,N_12813);
nor U14173 (N_14173,N_13155,N_13321);
and U14174 (N_14174,N_12947,N_12881);
and U14175 (N_14175,N_13083,N_13009);
and U14176 (N_14176,N_13149,N_13304);
xor U14177 (N_14177,N_13473,N_13330);
xnor U14178 (N_14178,N_13495,N_12759);
nor U14179 (N_14179,N_12960,N_13297);
xnor U14180 (N_14180,N_12797,N_13151);
nor U14181 (N_14181,N_12825,N_12863);
nand U14182 (N_14182,N_13139,N_12975);
xnor U14183 (N_14183,N_13047,N_13243);
xnor U14184 (N_14184,N_12961,N_12946);
nor U14185 (N_14185,N_13010,N_13371);
xor U14186 (N_14186,N_13102,N_13060);
xor U14187 (N_14187,N_13094,N_13059);
or U14188 (N_14188,N_13028,N_13206);
xor U14189 (N_14189,N_13400,N_13190);
and U14190 (N_14190,N_13286,N_12785);
nand U14191 (N_14191,N_12972,N_13295);
and U14192 (N_14192,N_13195,N_13310);
and U14193 (N_14193,N_12864,N_13374);
nor U14194 (N_14194,N_12849,N_13438);
nor U14195 (N_14195,N_13018,N_13112);
nand U14196 (N_14196,N_13496,N_12814);
nor U14197 (N_14197,N_13438,N_13157);
xnor U14198 (N_14198,N_12960,N_13260);
xor U14199 (N_14199,N_12938,N_13490);
xor U14200 (N_14200,N_13156,N_13459);
nor U14201 (N_14201,N_12958,N_12950);
xor U14202 (N_14202,N_13291,N_13293);
or U14203 (N_14203,N_13344,N_12903);
nor U14204 (N_14204,N_13152,N_13281);
and U14205 (N_14205,N_12762,N_12784);
or U14206 (N_14206,N_13273,N_13347);
nor U14207 (N_14207,N_13301,N_12801);
nor U14208 (N_14208,N_13144,N_12841);
xnor U14209 (N_14209,N_13208,N_13033);
nand U14210 (N_14210,N_13011,N_13408);
or U14211 (N_14211,N_13482,N_13399);
or U14212 (N_14212,N_12965,N_13101);
xor U14213 (N_14213,N_13270,N_12902);
xor U14214 (N_14214,N_13415,N_12908);
nor U14215 (N_14215,N_13476,N_13349);
and U14216 (N_14216,N_13334,N_12890);
xor U14217 (N_14217,N_12974,N_12831);
or U14218 (N_14218,N_13066,N_13402);
nand U14219 (N_14219,N_13402,N_13131);
xnor U14220 (N_14220,N_13182,N_13394);
nand U14221 (N_14221,N_12981,N_13042);
nand U14222 (N_14222,N_13242,N_12927);
nand U14223 (N_14223,N_12985,N_12787);
nor U14224 (N_14224,N_13001,N_12775);
xor U14225 (N_14225,N_12758,N_13497);
xor U14226 (N_14226,N_13212,N_13332);
or U14227 (N_14227,N_12846,N_13335);
xor U14228 (N_14228,N_13459,N_13483);
nor U14229 (N_14229,N_12751,N_12850);
or U14230 (N_14230,N_12775,N_13156);
or U14231 (N_14231,N_13198,N_13129);
nor U14232 (N_14232,N_13367,N_12950);
or U14233 (N_14233,N_13301,N_13278);
nand U14234 (N_14234,N_13093,N_13098);
nand U14235 (N_14235,N_13342,N_12864);
nor U14236 (N_14236,N_13185,N_13416);
nor U14237 (N_14237,N_13379,N_13103);
nand U14238 (N_14238,N_13025,N_12851);
nor U14239 (N_14239,N_13472,N_13211);
and U14240 (N_14240,N_12830,N_13143);
xnor U14241 (N_14241,N_13023,N_13377);
nor U14242 (N_14242,N_13493,N_13214);
and U14243 (N_14243,N_13013,N_13367);
or U14244 (N_14244,N_13490,N_13390);
and U14245 (N_14245,N_12990,N_12801);
nor U14246 (N_14246,N_13073,N_13066);
nor U14247 (N_14247,N_13286,N_13230);
and U14248 (N_14248,N_12895,N_12971);
nand U14249 (N_14249,N_13388,N_12823);
nor U14250 (N_14250,N_13506,N_14142);
nor U14251 (N_14251,N_13630,N_14218);
and U14252 (N_14252,N_13890,N_13863);
or U14253 (N_14253,N_13978,N_14161);
or U14254 (N_14254,N_13538,N_13713);
nor U14255 (N_14255,N_14165,N_13677);
or U14256 (N_14256,N_13986,N_13741);
or U14257 (N_14257,N_13721,N_13517);
nand U14258 (N_14258,N_13844,N_14172);
and U14259 (N_14259,N_13503,N_13722);
xnor U14260 (N_14260,N_14222,N_13619);
xnor U14261 (N_14261,N_14096,N_13892);
and U14262 (N_14262,N_13738,N_14125);
or U14263 (N_14263,N_13771,N_14101);
and U14264 (N_14264,N_14006,N_13674);
xnor U14265 (N_14265,N_13940,N_13655);
nor U14266 (N_14266,N_13651,N_13899);
nand U14267 (N_14267,N_13874,N_13633);
xor U14268 (N_14268,N_13583,N_13923);
nor U14269 (N_14269,N_13531,N_13769);
or U14270 (N_14270,N_14034,N_14014);
and U14271 (N_14271,N_13696,N_14091);
and U14272 (N_14272,N_14107,N_14239);
nand U14273 (N_14273,N_14039,N_13942);
nor U14274 (N_14274,N_14221,N_13973);
xor U14275 (N_14275,N_14191,N_13746);
and U14276 (N_14276,N_14225,N_14122);
xor U14277 (N_14277,N_13909,N_13849);
nand U14278 (N_14278,N_13921,N_13620);
nand U14279 (N_14279,N_13637,N_14187);
xor U14280 (N_14280,N_13665,N_14054);
and U14281 (N_14281,N_13784,N_13649);
xnor U14282 (N_14282,N_13935,N_13879);
nand U14283 (N_14283,N_13594,N_13822);
and U14284 (N_14284,N_13829,N_13635);
xor U14285 (N_14285,N_14179,N_13616);
xor U14286 (N_14286,N_14077,N_14242);
nand U14287 (N_14287,N_14140,N_13680);
and U14288 (N_14288,N_14195,N_13774);
or U14289 (N_14289,N_13929,N_13958);
or U14290 (N_14290,N_13737,N_13964);
or U14291 (N_14291,N_13652,N_14105);
nand U14292 (N_14292,N_13623,N_13650);
nand U14293 (N_14293,N_13579,N_14231);
nand U14294 (N_14294,N_14013,N_14023);
nand U14295 (N_14295,N_14234,N_14152);
or U14296 (N_14296,N_14015,N_13584);
or U14297 (N_14297,N_13988,N_13937);
nor U14298 (N_14298,N_13563,N_13606);
and U14299 (N_14299,N_13562,N_14134);
nor U14300 (N_14300,N_13907,N_13931);
nor U14301 (N_14301,N_13814,N_14197);
xor U14302 (N_14302,N_14026,N_14228);
nand U14303 (N_14303,N_13757,N_14076);
nor U14304 (N_14304,N_13881,N_14064);
or U14305 (N_14305,N_13780,N_14022);
nor U14306 (N_14306,N_14067,N_13885);
nor U14307 (N_14307,N_13580,N_14080);
nor U14308 (N_14308,N_13704,N_13922);
or U14309 (N_14309,N_13873,N_13858);
xor U14310 (N_14310,N_13683,N_14240);
and U14311 (N_14311,N_13785,N_13758);
nand U14312 (N_14312,N_13577,N_14097);
nor U14313 (N_14313,N_13513,N_13836);
nor U14314 (N_14314,N_13880,N_14035);
nand U14315 (N_14315,N_14248,N_13735);
nor U14316 (N_14316,N_13898,N_14065);
nand U14317 (N_14317,N_13807,N_14198);
xor U14318 (N_14318,N_14209,N_14170);
xor U14319 (N_14319,N_13550,N_13537);
or U14320 (N_14320,N_14073,N_13667);
xnor U14321 (N_14321,N_13726,N_13906);
nand U14322 (N_14322,N_14144,N_13671);
nand U14323 (N_14323,N_13926,N_13859);
or U14324 (N_14324,N_13753,N_13621);
or U14325 (N_14325,N_13888,N_13972);
nor U14326 (N_14326,N_13501,N_14059);
or U14327 (N_14327,N_13558,N_14051);
nor U14328 (N_14328,N_14183,N_13653);
xor U14329 (N_14329,N_13789,N_14178);
or U14330 (N_14330,N_14009,N_13871);
nand U14331 (N_14331,N_13763,N_13661);
nand U14332 (N_14332,N_13997,N_14057);
and U14333 (N_14333,N_13614,N_14008);
and U14334 (N_14334,N_13936,N_13961);
or U14335 (N_14335,N_13541,N_13751);
or U14336 (N_14336,N_14048,N_14226);
and U14337 (N_14337,N_13967,N_13511);
xor U14338 (N_14338,N_14223,N_13542);
and U14339 (N_14339,N_13524,N_14095);
nand U14340 (N_14340,N_13723,N_14061);
or U14341 (N_14341,N_13835,N_13566);
nand U14342 (N_14342,N_13656,N_14082);
nand U14343 (N_14343,N_14004,N_13920);
and U14344 (N_14344,N_13872,N_13512);
and U14345 (N_14345,N_14189,N_13910);
or U14346 (N_14346,N_13816,N_14081);
nand U14347 (N_14347,N_13521,N_13688);
nor U14348 (N_14348,N_13854,N_13720);
and U14349 (N_14349,N_14164,N_13870);
and U14350 (N_14350,N_13518,N_13628);
nand U14351 (N_14351,N_13500,N_14216);
and U14352 (N_14352,N_14150,N_13846);
and U14353 (N_14353,N_13514,N_13897);
xor U14354 (N_14354,N_14233,N_14167);
nand U14355 (N_14355,N_13770,N_13947);
xnor U14356 (N_14356,N_13868,N_13504);
nand U14357 (N_14357,N_14078,N_13752);
nor U14358 (N_14358,N_13826,N_13794);
nor U14359 (N_14359,N_14177,N_14068);
nor U14360 (N_14360,N_13675,N_14205);
nor U14361 (N_14361,N_13841,N_14038);
xor U14362 (N_14362,N_13773,N_13918);
nor U14363 (N_14363,N_13901,N_13945);
nor U14364 (N_14364,N_13535,N_13581);
xor U14365 (N_14365,N_14135,N_13869);
nor U14366 (N_14366,N_13730,N_13719);
xor U14367 (N_14367,N_13977,N_13728);
or U14368 (N_14368,N_13520,N_13954);
nand U14369 (N_14369,N_14090,N_14083);
or U14370 (N_14370,N_14049,N_13896);
xnor U14371 (N_14371,N_14027,N_14046);
nor U14372 (N_14372,N_14235,N_13647);
nand U14373 (N_14373,N_13747,N_13793);
nor U14374 (N_14374,N_13734,N_14238);
and U14375 (N_14375,N_13618,N_14085);
and U14376 (N_14376,N_14247,N_14071);
nand U14377 (N_14377,N_13700,N_13692);
and U14378 (N_14378,N_13694,N_14237);
and U14379 (N_14379,N_13556,N_13915);
nor U14380 (N_14380,N_13928,N_13768);
nor U14381 (N_14381,N_13553,N_13695);
nand U14382 (N_14382,N_14062,N_13642);
or U14383 (N_14383,N_14110,N_13743);
nand U14384 (N_14384,N_13812,N_13919);
or U14385 (N_14385,N_13611,N_13851);
and U14386 (N_14386,N_14158,N_13956);
nor U14387 (N_14387,N_13686,N_13711);
nand U14388 (N_14388,N_13838,N_13781);
or U14389 (N_14389,N_13893,N_14184);
nor U14390 (N_14390,N_13855,N_13969);
xor U14391 (N_14391,N_14182,N_13507);
nand U14392 (N_14392,N_13914,N_13508);
xor U14393 (N_14393,N_14200,N_13895);
nor U14394 (N_14394,N_14117,N_13707);
and U14395 (N_14395,N_13522,N_14249);
nand U14396 (N_14396,N_14214,N_13548);
and U14397 (N_14397,N_13609,N_13819);
and U14398 (N_14398,N_13555,N_13660);
xor U14399 (N_14399,N_13775,N_13551);
and U14400 (N_14400,N_13975,N_14243);
or U14401 (N_14401,N_14201,N_13632);
or U14402 (N_14402,N_13733,N_13989);
xnor U14403 (N_14403,N_13999,N_13799);
nor U14404 (N_14404,N_14190,N_13803);
nand U14405 (N_14405,N_13547,N_14169);
xor U14406 (N_14406,N_14147,N_14230);
and U14407 (N_14407,N_13779,N_13693);
nand U14408 (N_14408,N_13877,N_13591);
or U14409 (N_14409,N_13845,N_14012);
nand U14410 (N_14410,N_14100,N_14166);
nand U14411 (N_14411,N_14180,N_13891);
and U14412 (N_14412,N_14132,N_13842);
and U14413 (N_14413,N_13976,N_14194);
or U14414 (N_14414,N_14120,N_13528);
nor U14415 (N_14415,N_13904,N_14136);
xor U14416 (N_14416,N_13817,N_13708);
xnor U14417 (N_14417,N_13509,N_14007);
nor U14418 (N_14418,N_13861,N_14176);
xnor U14419 (N_14419,N_13599,N_13767);
or U14420 (N_14420,N_14126,N_13903);
nand U14421 (N_14421,N_14219,N_13588);
nor U14422 (N_14422,N_13745,N_14138);
and U14423 (N_14423,N_13965,N_13949);
xor U14424 (N_14424,N_13805,N_13602);
xnor U14425 (N_14425,N_14086,N_13668);
nand U14426 (N_14426,N_13857,N_13590);
xnor U14427 (N_14427,N_13532,N_13523);
nand U14428 (N_14428,N_14050,N_14084);
nand U14429 (N_14429,N_13543,N_14186);
or U14430 (N_14430,N_13603,N_13610);
or U14431 (N_14431,N_14188,N_14056);
xor U14432 (N_14432,N_13608,N_13552);
and U14433 (N_14433,N_13529,N_13955);
xor U14434 (N_14434,N_14145,N_13716);
xor U14435 (N_14435,N_14207,N_13516);
nor U14436 (N_14436,N_13974,N_13810);
nor U14437 (N_14437,N_14011,N_13607);
or U14438 (N_14438,N_13981,N_14127);
xor U14439 (N_14439,N_13670,N_13678);
nor U14440 (N_14440,N_13724,N_14019);
nand U14441 (N_14441,N_13934,N_14149);
xor U14442 (N_14442,N_13963,N_13549);
xnor U14443 (N_14443,N_14020,N_13802);
nand U14444 (N_14444,N_13944,N_14088);
xnor U14445 (N_14445,N_13882,N_13824);
xor U14446 (N_14446,N_14215,N_14045);
and U14447 (N_14447,N_13570,N_13691);
and U14448 (N_14448,N_13941,N_13557);
nand U14449 (N_14449,N_13995,N_14024);
or U14450 (N_14450,N_13644,N_13712);
xnor U14451 (N_14451,N_14112,N_13765);
xnor U14452 (N_14452,N_13883,N_13962);
nand U14453 (N_14453,N_13762,N_14016);
nand U14454 (N_14454,N_13917,N_13801);
nor U14455 (N_14455,N_13592,N_14017);
and U14456 (N_14456,N_13828,N_13748);
and U14457 (N_14457,N_14217,N_13596);
and U14458 (N_14458,N_13864,N_13866);
nor U14459 (N_14459,N_13515,N_14063);
nor U14460 (N_14460,N_14060,N_13648);
and U14461 (N_14461,N_13772,N_13994);
nand U14462 (N_14462,N_13815,N_13848);
nor U14463 (N_14463,N_13933,N_13565);
nor U14464 (N_14464,N_14181,N_13684);
or U14465 (N_14465,N_13646,N_14104);
and U14466 (N_14466,N_13821,N_14154);
xor U14467 (N_14467,N_13818,N_13887);
or U14468 (N_14468,N_14241,N_13959);
or U14469 (N_14469,N_13715,N_13798);
and U14470 (N_14470,N_13783,N_14155);
and U14471 (N_14471,N_14093,N_13913);
xnor U14472 (N_14472,N_13834,N_14156);
and U14473 (N_14473,N_14224,N_13702);
or U14474 (N_14474,N_13672,N_13908);
nand U14475 (N_14475,N_14102,N_13571);
xnor U14476 (N_14476,N_13951,N_14058);
nand U14477 (N_14477,N_13519,N_14028);
xor U14478 (N_14478,N_13952,N_14114);
xor U14479 (N_14479,N_13982,N_13878);
or U14480 (N_14480,N_13573,N_14032);
or U14481 (N_14481,N_13681,N_14157);
or U14482 (N_14482,N_13832,N_13984);
and U14483 (N_14483,N_13604,N_13640);
or U14484 (N_14484,N_13840,N_13830);
nand U14485 (N_14485,N_13886,N_14131);
or U14486 (N_14486,N_14043,N_13791);
and U14487 (N_14487,N_13534,N_13698);
or U14488 (N_14488,N_14030,N_13643);
nand U14489 (N_14489,N_13902,N_13561);
nand U14490 (N_14490,N_13657,N_14160);
or U14491 (N_14491,N_13939,N_13809);
nor U14492 (N_14492,N_14113,N_14041);
nor U14493 (N_14493,N_13797,N_14159);
nor U14494 (N_14494,N_13597,N_13572);
and U14495 (N_14495,N_13950,N_13867);
nand U14496 (N_14496,N_13559,N_13687);
nor U14497 (N_14497,N_14137,N_13813);
xor U14498 (N_14498,N_14106,N_13862);
and U14499 (N_14499,N_13568,N_13634);
xnor U14500 (N_14500,N_13585,N_14040);
and U14501 (N_14501,N_13613,N_13759);
nand U14502 (N_14502,N_13615,N_13777);
nor U14503 (N_14503,N_14151,N_14133);
and U14504 (N_14504,N_13957,N_13740);
and U14505 (N_14505,N_13598,N_13690);
nand U14506 (N_14506,N_13676,N_14111);
or U14507 (N_14507,N_13966,N_13865);
xnor U14508 (N_14508,N_14213,N_13729);
and U14509 (N_14509,N_13662,N_13587);
or U14510 (N_14510,N_14002,N_14192);
and U14511 (N_14511,N_13586,N_14174);
nand U14512 (N_14512,N_13792,N_14236);
nand U14513 (N_14513,N_13948,N_14042);
nor U14514 (N_14514,N_13725,N_14089);
xnor U14515 (N_14515,N_14119,N_13998);
and U14516 (N_14516,N_13669,N_13847);
nand U14517 (N_14517,N_13820,N_13663);
nand U14518 (N_14518,N_13732,N_13755);
nor U14519 (N_14519,N_13742,N_13560);
or U14520 (N_14520,N_13536,N_13985);
nor U14521 (N_14521,N_13946,N_14003);
xor U14522 (N_14522,N_13564,N_14141);
and U14523 (N_14523,N_14116,N_13932);
and U14524 (N_14524,N_14148,N_14070);
and U14525 (N_14525,N_13795,N_13709);
or U14526 (N_14526,N_13979,N_14206);
nand U14527 (N_14527,N_14025,N_13626);
nand U14528 (N_14528,N_13502,N_14052);
nand U14529 (N_14529,N_13960,N_14099);
xor U14530 (N_14530,N_14108,N_13980);
xnor U14531 (N_14531,N_13790,N_13894);
and U14532 (N_14532,N_13622,N_14210);
or U14533 (N_14533,N_13900,N_13544);
or U14534 (N_14534,N_13811,N_13505);
and U14535 (N_14535,N_13673,N_14044);
nor U14536 (N_14536,N_13612,N_13576);
nor U14537 (N_14537,N_14001,N_13582);
and U14538 (N_14538,N_14204,N_13595);
xor U14539 (N_14539,N_13852,N_14199);
xnor U14540 (N_14540,N_14033,N_13526);
or U14541 (N_14541,N_14109,N_13617);
nand U14542 (N_14542,N_14053,N_14153);
or U14543 (N_14543,N_13916,N_14162);
and U14544 (N_14544,N_13530,N_14245);
or U14545 (N_14545,N_13776,N_13574);
or U14546 (N_14546,N_13736,N_14130);
or U14547 (N_14547,N_13510,N_13717);
and U14548 (N_14548,N_13843,N_13525);
xor U14549 (N_14549,N_13567,N_13823);
or U14550 (N_14550,N_14129,N_13860);
xnor U14551 (N_14551,N_13839,N_14208);
and U14552 (N_14552,N_13968,N_13600);
nor U14553 (N_14553,N_14202,N_14203);
nand U14554 (N_14554,N_14168,N_13833);
and U14555 (N_14555,N_13601,N_13546);
and U14556 (N_14556,N_13953,N_14075);
nand U14557 (N_14557,N_13699,N_14098);
nor U14558 (N_14558,N_13911,N_13912);
xnor U14559 (N_14559,N_13545,N_14246);
or U14560 (N_14560,N_13971,N_13905);
nor U14561 (N_14561,N_13706,N_13625);
xor U14562 (N_14562,N_13987,N_13788);
nand U14563 (N_14563,N_14128,N_14047);
nand U14564 (N_14564,N_13727,N_14029);
and U14565 (N_14565,N_13990,N_13991);
xnor U14566 (N_14566,N_14069,N_13714);
xor U14567 (N_14567,N_13787,N_14079);
nand U14568 (N_14568,N_13569,N_13539);
xnor U14569 (N_14569,N_13605,N_13970);
nand U14570 (N_14570,N_14010,N_13850);
and U14571 (N_14571,N_14087,N_13837);
and U14572 (N_14572,N_13527,N_13697);
or U14573 (N_14573,N_13624,N_13993);
and U14574 (N_14574,N_13631,N_13756);
xor U14575 (N_14575,N_13554,N_13856);
and U14576 (N_14576,N_14232,N_13666);
nand U14577 (N_14577,N_14092,N_14072);
nor U14578 (N_14578,N_13996,N_14121);
and U14579 (N_14579,N_14037,N_14139);
and U14580 (N_14580,N_14163,N_14227);
or U14581 (N_14581,N_13705,N_13924);
xor U14582 (N_14582,N_13876,N_14036);
nor U14583 (N_14583,N_13808,N_13578);
xor U14584 (N_14584,N_13800,N_13943);
nand U14585 (N_14585,N_14196,N_14021);
nand U14586 (N_14586,N_14212,N_13589);
and U14587 (N_14587,N_13701,N_13710);
and U14588 (N_14588,N_13927,N_14066);
nand U14589 (N_14589,N_14193,N_13760);
nor U14590 (N_14590,N_13749,N_13764);
nand U14591 (N_14591,N_13627,N_14171);
or U14592 (N_14592,N_14146,N_13641);
or U14593 (N_14593,N_13718,N_14244);
or U14594 (N_14594,N_13831,N_13639);
xor U14595 (N_14595,N_13884,N_13638);
nand U14596 (N_14596,N_13659,N_13983);
and U14597 (N_14597,N_13739,N_13782);
nor U14598 (N_14598,N_13654,N_13925);
and U14599 (N_14599,N_13685,N_14175);
and U14600 (N_14600,N_14124,N_13825);
xnor U14601 (N_14601,N_13804,N_14185);
or U14602 (N_14602,N_14005,N_13682);
nand U14603 (N_14603,N_13786,N_13766);
nand U14604 (N_14604,N_14118,N_14103);
and U14605 (N_14605,N_13629,N_14031);
or U14606 (N_14606,N_14123,N_14173);
or U14607 (N_14607,N_13636,N_14143);
or U14608 (N_14608,N_13761,N_14055);
or U14609 (N_14609,N_13664,N_13827);
nand U14610 (N_14610,N_13540,N_14094);
xor U14611 (N_14611,N_13731,N_13593);
and U14612 (N_14612,N_13992,N_13778);
xnor U14613 (N_14613,N_14220,N_13875);
nor U14614 (N_14614,N_13938,N_13750);
nand U14615 (N_14615,N_13533,N_13658);
nor U14616 (N_14616,N_13575,N_13889);
xnor U14617 (N_14617,N_14018,N_13853);
nand U14618 (N_14618,N_13796,N_14229);
nor U14619 (N_14619,N_13930,N_14211);
and U14620 (N_14620,N_13703,N_13679);
and U14621 (N_14621,N_14000,N_13689);
nand U14622 (N_14622,N_13645,N_14074);
xor U14623 (N_14623,N_13754,N_14115);
nand U14624 (N_14624,N_13806,N_13744);
nand U14625 (N_14625,N_13803,N_13513);
nand U14626 (N_14626,N_14190,N_13510);
xnor U14627 (N_14627,N_13845,N_13874);
or U14628 (N_14628,N_14026,N_13707);
nand U14629 (N_14629,N_14133,N_13910);
xor U14630 (N_14630,N_13897,N_13559);
nand U14631 (N_14631,N_14075,N_13605);
xor U14632 (N_14632,N_13658,N_14135);
or U14633 (N_14633,N_13989,N_14104);
or U14634 (N_14634,N_13805,N_13948);
or U14635 (N_14635,N_13832,N_13761);
or U14636 (N_14636,N_13670,N_13680);
or U14637 (N_14637,N_14037,N_13525);
nand U14638 (N_14638,N_13838,N_13833);
xnor U14639 (N_14639,N_13872,N_13908);
nand U14640 (N_14640,N_13680,N_13617);
nor U14641 (N_14641,N_13779,N_13977);
nand U14642 (N_14642,N_13938,N_13811);
xor U14643 (N_14643,N_13584,N_14212);
xor U14644 (N_14644,N_13921,N_14068);
or U14645 (N_14645,N_14222,N_13635);
or U14646 (N_14646,N_14054,N_14122);
and U14647 (N_14647,N_14224,N_13607);
nor U14648 (N_14648,N_13502,N_14119);
nor U14649 (N_14649,N_13883,N_13501);
nor U14650 (N_14650,N_13742,N_13806);
or U14651 (N_14651,N_14248,N_13993);
xor U14652 (N_14652,N_14199,N_13885);
or U14653 (N_14653,N_14175,N_13775);
nand U14654 (N_14654,N_14095,N_14013);
nand U14655 (N_14655,N_14018,N_14220);
nor U14656 (N_14656,N_13785,N_13529);
or U14657 (N_14657,N_13795,N_13674);
nand U14658 (N_14658,N_13828,N_14198);
nand U14659 (N_14659,N_13589,N_13692);
xor U14660 (N_14660,N_14077,N_14206);
and U14661 (N_14661,N_14046,N_13633);
and U14662 (N_14662,N_13640,N_13907);
nor U14663 (N_14663,N_13581,N_13728);
nor U14664 (N_14664,N_13901,N_13822);
and U14665 (N_14665,N_13947,N_13504);
nand U14666 (N_14666,N_13624,N_14222);
or U14667 (N_14667,N_13844,N_13746);
nor U14668 (N_14668,N_14183,N_13932);
nand U14669 (N_14669,N_13574,N_13606);
nand U14670 (N_14670,N_14065,N_13995);
and U14671 (N_14671,N_14183,N_13582);
or U14672 (N_14672,N_13985,N_13786);
and U14673 (N_14673,N_13616,N_14157);
xnor U14674 (N_14674,N_13689,N_14221);
xor U14675 (N_14675,N_14156,N_14099);
and U14676 (N_14676,N_13813,N_13612);
nor U14677 (N_14677,N_13918,N_13887);
nor U14678 (N_14678,N_13897,N_13719);
nand U14679 (N_14679,N_13668,N_13770);
xor U14680 (N_14680,N_14038,N_13602);
or U14681 (N_14681,N_14098,N_13693);
nor U14682 (N_14682,N_14247,N_13877);
and U14683 (N_14683,N_13966,N_14104);
nor U14684 (N_14684,N_13596,N_13831);
or U14685 (N_14685,N_14204,N_13921);
or U14686 (N_14686,N_13966,N_14192);
and U14687 (N_14687,N_13680,N_13838);
and U14688 (N_14688,N_14160,N_14220);
xor U14689 (N_14689,N_13688,N_13536);
and U14690 (N_14690,N_13756,N_14165);
xor U14691 (N_14691,N_13640,N_13529);
and U14692 (N_14692,N_14220,N_14143);
xnor U14693 (N_14693,N_13665,N_13835);
nand U14694 (N_14694,N_13661,N_13881);
or U14695 (N_14695,N_14152,N_13706);
nor U14696 (N_14696,N_14207,N_13761);
or U14697 (N_14697,N_14100,N_13807);
or U14698 (N_14698,N_13695,N_14169);
or U14699 (N_14699,N_14081,N_14086);
nand U14700 (N_14700,N_13932,N_13608);
nand U14701 (N_14701,N_13746,N_13828);
or U14702 (N_14702,N_13811,N_13777);
nand U14703 (N_14703,N_13534,N_13584);
xor U14704 (N_14704,N_14132,N_13793);
nor U14705 (N_14705,N_14125,N_13546);
and U14706 (N_14706,N_13583,N_13747);
or U14707 (N_14707,N_14132,N_13725);
nand U14708 (N_14708,N_13586,N_14100);
nand U14709 (N_14709,N_14136,N_13679);
and U14710 (N_14710,N_14180,N_14148);
and U14711 (N_14711,N_13645,N_14106);
nand U14712 (N_14712,N_13894,N_14079);
and U14713 (N_14713,N_13972,N_13758);
xor U14714 (N_14714,N_14166,N_13872);
and U14715 (N_14715,N_13792,N_13740);
and U14716 (N_14716,N_14013,N_13623);
nor U14717 (N_14717,N_13774,N_13577);
nand U14718 (N_14718,N_13512,N_13858);
or U14719 (N_14719,N_13938,N_14131);
or U14720 (N_14720,N_14183,N_13566);
xor U14721 (N_14721,N_13849,N_13870);
nor U14722 (N_14722,N_14008,N_14144);
or U14723 (N_14723,N_14074,N_13849);
or U14724 (N_14724,N_14073,N_13682);
nand U14725 (N_14725,N_13909,N_13735);
xnor U14726 (N_14726,N_13642,N_13584);
or U14727 (N_14727,N_13857,N_13788);
nand U14728 (N_14728,N_14075,N_13859);
nor U14729 (N_14729,N_13508,N_13681);
nor U14730 (N_14730,N_13906,N_14053);
and U14731 (N_14731,N_14057,N_13799);
xor U14732 (N_14732,N_13655,N_14177);
xnor U14733 (N_14733,N_13501,N_13992);
xnor U14734 (N_14734,N_13531,N_13842);
or U14735 (N_14735,N_13790,N_13911);
or U14736 (N_14736,N_13910,N_13590);
and U14737 (N_14737,N_13526,N_13604);
nor U14738 (N_14738,N_13844,N_13569);
nor U14739 (N_14739,N_14016,N_13889);
nand U14740 (N_14740,N_14164,N_13638);
nor U14741 (N_14741,N_14122,N_13713);
and U14742 (N_14742,N_14228,N_14211);
nor U14743 (N_14743,N_13532,N_14000);
and U14744 (N_14744,N_14100,N_13666);
nand U14745 (N_14745,N_13561,N_13959);
nor U14746 (N_14746,N_14106,N_13880);
and U14747 (N_14747,N_13519,N_14223);
nand U14748 (N_14748,N_13615,N_13535);
and U14749 (N_14749,N_13885,N_13724);
nand U14750 (N_14750,N_13598,N_13572);
xnor U14751 (N_14751,N_14048,N_13731);
and U14752 (N_14752,N_13643,N_14180);
and U14753 (N_14753,N_13680,N_14138);
or U14754 (N_14754,N_13786,N_14081);
nand U14755 (N_14755,N_14190,N_13794);
xor U14756 (N_14756,N_13709,N_13516);
nand U14757 (N_14757,N_13717,N_13626);
or U14758 (N_14758,N_14125,N_13653);
xor U14759 (N_14759,N_13798,N_13870);
or U14760 (N_14760,N_13983,N_13753);
nor U14761 (N_14761,N_13602,N_13624);
xnor U14762 (N_14762,N_13783,N_13954);
nand U14763 (N_14763,N_13709,N_13654);
nand U14764 (N_14764,N_13986,N_14156);
nand U14765 (N_14765,N_13711,N_14180);
nor U14766 (N_14766,N_13847,N_14003);
xnor U14767 (N_14767,N_13716,N_13945);
or U14768 (N_14768,N_13599,N_13597);
and U14769 (N_14769,N_13759,N_14049);
and U14770 (N_14770,N_13668,N_14183);
nor U14771 (N_14771,N_14136,N_13920);
or U14772 (N_14772,N_14090,N_14056);
xnor U14773 (N_14773,N_13942,N_14085);
nor U14774 (N_14774,N_13688,N_13560);
and U14775 (N_14775,N_13846,N_13837);
or U14776 (N_14776,N_13644,N_13635);
xnor U14777 (N_14777,N_14143,N_13997);
or U14778 (N_14778,N_14035,N_14041);
and U14779 (N_14779,N_13662,N_13942);
xnor U14780 (N_14780,N_13649,N_13639);
and U14781 (N_14781,N_13704,N_14042);
nor U14782 (N_14782,N_13554,N_13928);
and U14783 (N_14783,N_14113,N_13963);
and U14784 (N_14784,N_13774,N_13971);
nor U14785 (N_14785,N_13881,N_13855);
or U14786 (N_14786,N_13879,N_13930);
xor U14787 (N_14787,N_14168,N_13896);
nor U14788 (N_14788,N_14081,N_13747);
nor U14789 (N_14789,N_14214,N_13998);
nor U14790 (N_14790,N_14075,N_13855);
nor U14791 (N_14791,N_13858,N_13914);
nor U14792 (N_14792,N_13898,N_13674);
nor U14793 (N_14793,N_13844,N_13709);
and U14794 (N_14794,N_13650,N_13651);
nor U14795 (N_14795,N_14108,N_13900);
and U14796 (N_14796,N_13531,N_13863);
xnor U14797 (N_14797,N_13966,N_13752);
and U14798 (N_14798,N_14178,N_14062);
nand U14799 (N_14799,N_13857,N_14210);
nand U14800 (N_14800,N_13820,N_14118);
or U14801 (N_14801,N_13855,N_13545);
xnor U14802 (N_14802,N_13847,N_13607);
or U14803 (N_14803,N_14134,N_14224);
nor U14804 (N_14804,N_14006,N_13595);
nand U14805 (N_14805,N_13790,N_13733);
and U14806 (N_14806,N_14055,N_13825);
or U14807 (N_14807,N_13538,N_13502);
and U14808 (N_14808,N_13946,N_13612);
xor U14809 (N_14809,N_13713,N_14161);
and U14810 (N_14810,N_13771,N_14234);
xor U14811 (N_14811,N_13923,N_14052);
or U14812 (N_14812,N_13747,N_13978);
nor U14813 (N_14813,N_13762,N_13927);
nand U14814 (N_14814,N_14167,N_14172);
xnor U14815 (N_14815,N_14033,N_13651);
and U14816 (N_14816,N_13959,N_14007);
or U14817 (N_14817,N_13620,N_13591);
nand U14818 (N_14818,N_13534,N_14163);
xnor U14819 (N_14819,N_13602,N_13628);
nand U14820 (N_14820,N_13869,N_13937);
nor U14821 (N_14821,N_14092,N_13870);
nand U14822 (N_14822,N_14211,N_14028);
nor U14823 (N_14823,N_13866,N_13894);
nor U14824 (N_14824,N_13953,N_13962);
and U14825 (N_14825,N_13719,N_13890);
nor U14826 (N_14826,N_14179,N_13555);
xnor U14827 (N_14827,N_13517,N_13689);
xnor U14828 (N_14828,N_13993,N_14107);
or U14829 (N_14829,N_14230,N_13739);
xor U14830 (N_14830,N_13765,N_13706);
or U14831 (N_14831,N_13661,N_13640);
nor U14832 (N_14832,N_13623,N_13840);
or U14833 (N_14833,N_13899,N_13685);
and U14834 (N_14834,N_13992,N_13866);
nor U14835 (N_14835,N_14217,N_14226);
nand U14836 (N_14836,N_13694,N_13861);
nor U14837 (N_14837,N_14014,N_13818);
nor U14838 (N_14838,N_13658,N_13573);
and U14839 (N_14839,N_13746,N_13568);
or U14840 (N_14840,N_13502,N_14032);
xnor U14841 (N_14841,N_13638,N_13589);
or U14842 (N_14842,N_13900,N_14077);
nand U14843 (N_14843,N_14007,N_13698);
nor U14844 (N_14844,N_13599,N_13669);
xnor U14845 (N_14845,N_13926,N_13741);
xor U14846 (N_14846,N_13820,N_13551);
and U14847 (N_14847,N_13761,N_13836);
xor U14848 (N_14848,N_13669,N_13805);
xor U14849 (N_14849,N_13674,N_13630);
nor U14850 (N_14850,N_13544,N_13630);
nor U14851 (N_14851,N_14114,N_13715);
nand U14852 (N_14852,N_13802,N_13747);
and U14853 (N_14853,N_13736,N_14004);
or U14854 (N_14854,N_14191,N_13814);
nand U14855 (N_14855,N_13513,N_13880);
nand U14856 (N_14856,N_13879,N_13527);
nor U14857 (N_14857,N_13979,N_14168);
xnor U14858 (N_14858,N_13913,N_13796);
and U14859 (N_14859,N_14157,N_14206);
xnor U14860 (N_14860,N_13589,N_14162);
xor U14861 (N_14861,N_13509,N_13787);
xor U14862 (N_14862,N_13988,N_13651);
and U14863 (N_14863,N_13625,N_14039);
nand U14864 (N_14864,N_13768,N_14039);
and U14865 (N_14865,N_13632,N_13598);
and U14866 (N_14866,N_13752,N_13822);
and U14867 (N_14867,N_14244,N_14041);
or U14868 (N_14868,N_13743,N_14151);
and U14869 (N_14869,N_14100,N_13580);
xor U14870 (N_14870,N_13971,N_13546);
nand U14871 (N_14871,N_13949,N_13920);
or U14872 (N_14872,N_13977,N_13846);
nand U14873 (N_14873,N_13973,N_14188);
and U14874 (N_14874,N_13826,N_13563);
or U14875 (N_14875,N_13769,N_14021);
xnor U14876 (N_14876,N_13559,N_13679);
nor U14877 (N_14877,N_13648,N_13525);
nor U14878 (N_14878,N_13749,N_14015);
nor U14879 (N_14879,N_13870,N_14176);
and U14880 (N_14880,N_13916,N_13719);
xnor U14881 (N_14881,N_14087,N_13895);
and U14882 (N_14882,N_13688,N_13607);
nand U14883 (N_14883,N_13617,N_13837);
or U14884 (N_14884,N_13707,N_14120);
or U14885 (N_14885,N_13860,N_14069);
or U14886 (N_14886,N_13821,N_13758);
or U14887 (N_14887,N_14100,N_14216);
and U14888 (N_14888,N_13999,N_13960);
nand U14889 (N_14889,N_13862,N_13525);
nand U14890 (N_14890,N_14113,N_13609);
nor U14891 (N_14891,N_13769,N_13909);
and U14892 (N_14892,N_13904,N_13541);
xor U14893 (N_14893,N_14079,N_13556);
xor U14894 (N_14894,N_14233,N_13907);
nor U14895 (N_14895,N_13589,N_13636);
or U14896 (N_14896,N_13819,N_14075);
xnor U14897 (N_14897,N_14192,N_13815);
and U14898 (N_14898,N_13536,N_13955);
or U14899 (N_14899,N_13725,N_14075);
nor U14900 (N_14900,N_14110,N_13691);
nor U14901 (N_14901,N_13924,N_13784);
xnor U14902 (N_14902,N_14199,N_13605);
or U14903 (N_14903,N_13719,N_14091);
or U14904 (N_14904,N_14235,N_13768);
nand U14905 (N_14905,N_14227,N_13925);
and U14906 (N_14906,N_13635,N_13773);
and U14907 (N_14907,N_13909,N_13712);
xor U14908 (N_14908,N_14146,N_14135);
nand U14909 (N_14909,N_13510,N_13764);
xor U14910 (N_14910,N_13859,N_13691);
nor U14911 (N_14911,N_13711,N_13543);
nand U14912 (N_14912,N_13886,N_14214);
and U14913 (N_14913,N_13720,N_13953);
or U14914 (N_14914,N_14248,N_13681);
xnor U14915 (N_14915,N_13508,N_14038);
and U14916 (N_14916,N_13635,N_14224);
nand U14917 (N_14917,N_14141,N_14246);
or U14918 (N_14918,N_14006,N_13621);
nor U14919 (N_14919,N_14197,N_14185);
and U14920 (N_14920,N_14232,N_14004);
xor U14921 (N_14921,N_13563,N_13823);
and U14922 (N_14922,N_13888,N_13770);
nand U14923 (N_14923,N_14238,N_13954);
or U14924 (N_14924,N_14045,N_14017);
xnor U14925 (N_14925,N_14153,N_13925);
and U14926 (N_14926,N_13673,N_14017);
nand U14927 (N_14927,N_13977,N_13612);
nor U14928 (N_14928,N_14091,N_14236);
and U14929 (N_14929,N_13985,N_13980);
nand U14930 (N_14930,N_13606,N_14123);
or U14931 (N_14931,N_14226,N_14183);
or U14932 (N_14932,N_13956,N_13586);
nor U14933 (N_14933,N_14085,N_13796);
xnor U14934 (N_14934,N_13662,N_13769);
and U14935 (N_14935,N_14077,N_13959);
nand U14936 (N_14936,N_14041,N_13888);
xor U14937 (N_14937,N_14084,N_13708);
nor U14938 (N_14938,N_13809,N_14068);
xnor U14939 (N_14939,N_13699,N_14139);
xnor U14940 (N_14940,N_13810,N_14168);
nor U14941 (N_14941,N_13686,N_13535);
and U14942 (N_14942,N_13724,N_13887);
or U14943 (N_14943,N_14129,N_13903);
and U14944 (N_14944,N_13996,N_13584);
nand U14945 (N_14945,N_13571,N_13774);
or U14946 (N_14946,N_14244,N_14158);
or U14947 (N_14947,N_13505,N_13787);
nor U14948 (N_14948,N_13876,N_14025);
or U14949 (N_14949,N_14185,N_14142);
and U14950 (N_14950,N_13514,N_13802);
xor U14951 (N_14951,N_13694,N_14147);
or U14952 (N_14952,N_14003,N_14033);
nand U14953 (N_14953,N_13626,N_13579);
nand U14954 (N_14954,N_13943,N_13915);
xor U14955 (N_14955,N_14207,N_13751);
xnor U14956 (N_14956,N_14111,N_13560);
xor U14957 (N_14957,N_13561,N_13567);
nor U14958 (N_14958,N_14247,N_13910);
nor U14959 (N_14959,N_13822,N_13504);
xor U14960 (N_14960,N_14087,N_13988);
and U14961 (N_14961,N_13922,N_14181);
nor U14962 (N_14962,N_13861,N_14000);
or U14963 (N_14963,N_14191,N_13787);
and U14964 (N_14964,N_13671,N_13728);
nor U14965 (N_14965,N_13967,N_13939);
nor U14966 (N_14966,N_13643,N_13815);
nand U14967 (N_14967,N_14089,N_13552);
and U14968 (N_14968,N_14171,N_13732);
or U14969 (N_14969,N_14168,N_13582);
xnor U14970 (N_14970,N_14106,N_13737);
xnor U14971 (N_14971,N_13777,N_13755);
xor U14972 (N_14972,N_13518,N_13543);
and U14973 (N_14973,N_13724,N_14027);
nand U14974 (N_14974,N_14129,N_13999);
and U14975 (N_14975,N_14159,N_13777);
and U14976 (N_14976,N_13577,N_13910);
xor U14977 (N_14977,N_13921,N_14203);
nand U14978 (N_14978,N_13949,N_14076);
or U14979 (N_14979,N_14112,N_14144);
or U14980 (N_14980,N_14186,N_13628);
and U14981 (N_14981,N_13973,N_13847);
xor U14982 (N_14982,N_13757,N_13515);
and U14983 (N_14983,N_13822,N_13965);
nor U14984 (N_14984,N_13904,N_14176);
nand U14985 (N_14985,N_14211,N_13650);
xnor U14986 (N_14986,N_13563,N_13560);
nor U14987 (N_14987,N_14053,N_13564);
nor U14988 (N_14988,N_13829,N_13890);
and U14989 (N_14989,N_13591,N_13978);
and U14990 (N_14990,N_14020,N_14222);
or U14991 (N_14991,N_14185,N_13867);
nand U14992 (N_14992,N_13852,N_13718);
or U14993 (N_14993,N_13822,N_13665);
nand U14994 (N_14994,N_13793,N_13720);
and U14995 (N_14995,N_13953,N_14121);
and U14996 (N_14996,N_14161,N_14135);
or U14997 (N_14997,N_13857,N_13612);
nor U14998 (N_14998,N_14120,N_13902);
and U14999 (N_14999,N_13635,N_13726);
xnor UO_0 (O_0,N_14978,N_14789);
and UO_1 (O_1,N_14563,N_14540);
nor UO_2 (O_2,N_14701,N_14345);
or UO_3 (O_3,N_14323,N_14778);
nor UO_4 (O_4,N_14430,N_14426);
or UO_5 (O_5,N_14849,N_14530);
nor UO_6 (O_6,N_14310,N_14749);
xor UO_7 (O_7,N_14950,N_14918);
and UO_8 (O_8,N_14954,N_14851);
xor UO_9 (O_9,N_14254,N_14301);
xor UO_10 (O_10,N_14696,N_14419);
and UO_11 (O_11,N_14815,N_14311);
xor UO_12 (O_12,N_14413,N_14390);
xor UO_13 (O_13,N_14606,N_14469);
nor UO_14 (O_14,N_14486,N_14770);
or UO_15 (O_15,N_14689,N_14598);
xnor UO_16 (O_16,N_14882,N_14391);
nor UO_17 (O_17,N_14425,N_14512);
xnor UO_18 (O_18,N_14304,N_14927);
or UO_19 (O_19,N_14875,N_14546);
xnor UO_20 (O_20,N_14854,N_14731);
nand UO_21 (O_21,N_14772,N_14891);
xor UO_22 (O_22,N_14946,N_14832);
xnor UO_23 (O_23,N_14578,N_14841);
nand UO_24 (O_24,N_14559,N_14520);
nand UO_25 (O_25,N_14613,N_14935);
or UO_26 (O_26,N_14788,N_14605);
nand UO_27 (O_27,N_14475,N_14829);
xnor UO_28 (O_28,N_14526,N_14402);
or UO_29 (O_29,N_14279,N_14300);
nor UO_30 (O_30,N_14353,N_14900);
xnor UO_31 (O_31,N_14330,N_14289);
or UO_32 (O_32,N_14556,N_14705);
nand UO_33 (O_33,N_14564,N_14790);
and UO_34 (O_34,N_14907,N_14420);
nand UO_35 (O_35,N_14607,N_14913);
xnor UO_36 (O_36,N_14270,N_14378);
nor UO_37 (O_37,N_14591,N_14926);
xnor UO_38 (O_38,N_14836,N_14478);
nor UO_39 (O_39,N_14305,N_14883);
xor UO_40 (O_40,N_14320,N_14461);
nor UO_41 (O_41,N_14684,N_14779);
nor UO_42 (O_42,N_14912,N_14516);
or UO_43 (O_43,N_14892,N_14862);
nor UO_44 (O_44,N_14975,N_14853);
nor UO_45 (O_45,N_14754,N_14716);
or UO_46 (O_46,N_14359,N_14893);
or UO_47 (O_47,N_14594,N_14711);
nor UO_48 (O_48,N_14357,N_14870);
or UO_49 (O_49,N_14455,N_14423);
nor UO_50 (O_50,N_14427,N_14643);
or UO_51 (O_51,N_14660,N_14804);
and UO_52 (O_52,N_14690,N_14915);
nor UO_53 (O_53,N_14321,N_14707);
xnor UO_54 (O_54,N_14636,N_14457);
nand UO_55 (O_55,N_14999,N_14681);
and UO_56 (O_56,N_14931,N_14414);
or UO_57 (O_57,N_14970,N_14566);
nand UO_58 (O_58,N_14452,N_14617);
xor UO_59 (O_59,N_14485,N_14542);
nand UO_60 (O_60,N_14316,N_14615);
nor UO_61 (O_61,N_14953,N_14980);
or UO_62 (O_62,N_14940,N_14773);
and UO_63 (O_63,N_14302,N_14651);
xnor UO_64 (O_64,N_14751,N_14326);
or UO_65 (O_65,N_14582,N_14968);
and UO_66 (O_66,N_14969,N_14264);
or UO_67 (O_67,N_14547,N_14428);
and UO_68 (O_68,N_14818,N_14332);
nor UO_69 (O_69,N_14290,N_14502);
xnor UO_70 (O_70,N_14794,N_14745);
nor UO_71 (O_71,N_14858,N_14928);
or UO_72 (O_72,N_14528,N_14462);
and UO_73 (O_73,N_14676,N_14960);
nand UO_74 (O_74,N_14618,N_14753);
nand UO_75 (O_75,N_14394,N_14449);
and UO_76 (O_76,N_14331,N_14645);
xnor UO_77 (O_77,N_14816,N_14787);
nor UO_78 (O_78,N_14780,N_14421);
or UO_79 (O_79,N_14863,N_14833);
xor UO_80 (O_80,N_14842,N_14755);
nand UO_81 (O_81,N_14679,N_14336);
nor UO_82 (O_82,N_14922,N_14495);
nor UO_83 (O_83,N_14990,N_14810);
nor UO_84 (O_84,N_14532,N_14997);
nor UO_85 (O_85,N_14799,N_14719);
xor UO_86 (O_86,N_14687,N_14860);
nand UO_87 (O_87,N_14667,N_14781);
nor UO_88 (O_88,N_14588,N_14592);
or UO_89 (O_89,N_14878,N_14898);
and UO_90 (O_90,N_14683,N_14675);
nand UO_91 (O_91,N_14261,N_14333);
or UO_92 (O_92,N_14470,N_14776);
xor UO_93 (O_93,N_14351,N_14347);
nand UO_94 (O_94,N_14920,N_14864);
and UO_95 (O_95,N_14814,N_14429);
nand UO_96 (O_96,N_14252,N_14974);
or UO_97 (O_97,N_14471,N_14367);
nor UO_98 (O_98,N_14368,N_14611);
or UO_99 (O_99,N_14263,N_14318);
nand UO_100 (O_100,N_14957,N_14435);
xor UO_101 (O_101,N_14541,N_14843);
nor UO_102 (O_102,N_14399,N_14568);
nor UO_103 (O_103,N_14880,N_14576);
nand UO_104 (O_104,N_14637,N_14694);
nand UO_105 (O_105,N_14406,N_14871);
and UO_106 (O_106,N_14847,N_14947);
or UO_107 (O_107,N_14856,N_14702);
xnor UO_108 (O_108,N_14884,N_14819);
or UO_109 (O_109,N_14734,N_14567);
xor UO_110 (O_110,N_14560,N_14937);
and UO_111 (O_111,N_14805,N_14389);
nor UO_112 (O_112,N_14396,N_14817);
nor UO_113 (O_113,N_14522,N_14793);
nor UO_114 (O_114,N_14986,N_14303);
xnor UO_115 (O_115,N_14839,N_14756);
xnor UO_116 (O_116,N_14655,N_14285);
or UO_117 (O_117,N_14855,N_14941);
xnor UO_118 (O_118,N_14708,N_14837);
xor UO_119 (O_119,N_14629,N_14872);
and UO_120 (O_120,N_14733,N_14993);
nand UO_121 (O_121,N_14742,N_14801);
xnor UO_122 (O_122,N_14967,N_14657);
nand UO_123 (O_123,N_14595,N_14561);
nand UO_124 (O_124,N_14360,N_14584);
nand UO_125 (O_125,N_14570,N_14439);
nor UO_126 (O_126,N_14544,N_14812);
xnor UO_127 (O_127,N_14649,N_14890);
xnor UO_128 (O_128,N_14991,N_14340);
nand UO_129 (O_129,N_14677,N_14253);
nand UO_130 (O_130,N_14639,N_14809);
nor UO_131 (O_131,N_14740,N_14981);
and UO_132 (O_132,N_14943,N_14944);
xor UO_133 (O_133,N_14736,N_14700);
nand UO_134 (O_134,N_14472,N_14766);
and UO_135 (O_135,N_14897,N_14998);
xor UO_136 (O_136,N_14866,N_14460);
and UO_137 (O_137,N_14515,N_14807);
xor UO_138 (O_138,N_14258,N_14724);
or UO_139 (O_139,N_14747,N_14325);
xnor UO_140 (O_140,N_14930,N_14436);
nand UO_141 (O_141,N_14835,N_14976);
or UO_142 (O_142,N_14418,N_14401);
nor UO_143 (O_143,N_14796,N_14664);
nand UO_144 (O_144,N_14294,N_14373);
or UO_145 (O_145,N_14374,N_14334);
xnor UO_146 (O_146,N_14939,N_14830);
xor UO_147 (O_147,N_14342,N_14350);
or UO_148 (O_148,N_14480,N_14840);
nor UO_149 (O_149,N_14506,N_14762);
xor UO_150 (O_150,N_14824,N_14671);
and UO_151 (O_151,N_14370,N_14888);
nor UO_152 (O_152,N_14669,N_14621);
or UO_153 (O_153,N_14717,N_14309);
xor UO_154 (O_154,N_14795,N_14752);
xnor UO_155 (O_155,N_14723,N_14324);
or UO_156 (O_156,N_14417,N_14441);
nand UO_157 (O_157,N_14732,N_14955);
or UO_158 (O_158,N_14298,N_14276);
nor UO_159 (O_159,N_14473,N_14813);
and UO_160 (O_160,N_14963,N_14977);
and UO_161 (O_161,N_14599,N_14328);
or UO_162 (O_162,N_14277,N_14295);
xor UO_163 (O_163,N_14317,N_14499);
nor UO_164 (O_164,N_14834,N_14273);
or UO_165 (O_165,N_14562,N_14500);
or UO_166 (O_166,N_14785,N_14392);
and UO_167 (O_167,N_14909,N_14821);
or UO_168 (O_168,N_14476,N_14886);
nand UO_169 (O_169,N_14524,N_14791);
nor UO_170 (O_170,N_14251,N_14760);
xor UO_171 (O_171,N_14250,N_14782);
nand UO_172 (O_172,N_14597,N_14474);
or UO_173 (O_173,N_14774,N_14466);
xnor UO_174 (O_174,N_14456,N_14343);
nor UO_175 (O_175,N_14635,N_14658);
or UO_176 (O_176,N_14691,N_14800);
and UO_177 (O_177,N_14400,N_14982);
and UO_178 (O_178,N_14715,N_14539);
and UO_179 (O_179,N_14765,N_14558);
nand UO_180 (O_180,N_14728,N_14518);
and UO_181 (O_181,N_14641,N_14627);
and UO_182 (O_182,N_14306,N_14577);
nand UO_183 (O_183,N_14281,N_14513);
and UO_184 (O_184,N_14623,N_14291);
and UO_185 (O_185,N_14678,N_14356);
nand UO_186 (O_186,N_14438,N_14407);
xnor UO_187 (O_187,N_14983,N_14448);
xnor UO_188 (O_188,N_14299,N_14758);
nand UO_189 (O_189,N_14868,N_14811);
or UO_190 (O_190,N_14265,N_14372);
and UO_191 (O_191,N_14464,N_14602);
xnor UO_192 (O_192,N_14625,N_14958);
and UO_193 (O_193,N_14395,N_14867);
and UO_194 (O_194,N_14579,N_14424);
nand UO_195 (O_195,N_14646,N_14271);
nand UO_196 (O_196,N_14786,N_14881);
nor UO_197 (O_197,N_14846,N_14668);
or UO_198 (O_198,N_14550,N_14349);
and UO_199 (O_199,N_14533,N_14269);
and UO_200 (O_200,N_14896,N_14257);
xnor UO_201 (O_201,N_14501,N_14477);
nor UO_202 (O_202,N_14962,N_14553);
nand UO_203 (O_203,N_14445,N_14344);
and UO_204 (O_204,N_14852,N_14315);
and UO_205 (O_205,N_14590,N_14925);
xnor UO_206 (O_206,N_14797,N_14322);
nor UO_207 (O_207,N_14911,N_14514);
nand UO_208 (O_208,N_14844,N_14670);
xnor UO_209 (O_209,N_14859,N_14916);
and UO_210 (O_210,N_14828,N_14600);
nand UO_211 (O_211,N_14517,N_14624);
nor UO_212 (O_212,N_14965,N_14296);
and UO_213 (O_213,N_14726,N_14415);
nor UO_214 (O_214,N_14693,N_14848);
nor UO_215 (O_215,N_14468,N_14654);
and UO_216 (O_216,N_14910,N_14293);
or UO_217 (O_217,N_14572,N_14437);
nor UO_218 (O_218,N_14640,N_14255);
xnor UO_219 (O_219,N_14934,N_14822);
or UO_220 (O_220,N_14527,N_14434);
nand UO_221 (O_221,N_14308,N_14709);
xor UO_222 (O_222,N_14885,N_14995);
xnor UO_223 (O_223,N_14631,N_14284);
xor UO_224 (O_224,N_14535,N_14899);
and UO_225 (O_225,N_14362,N_14771);
or UO_226 (O_226,N_14901,N_14735);
and UO_227 (O_227,N_14652,N_14352);
nor UO_228 (O_228,N_14404,N_14511);
or UO_229 (O_229,N_14361,N_14387);
and UO_230 (O_230,N_14966,N_14497);
or UO_231 (O_231,N_14659,N_14783);
xor UO_232 (O_232,N_14992,N_14551);
nand UO_233 (O_233,N_14385,N_14329);
and UO_234 (O_234,N_14902,N_14686);
and UO_235 (O_235,N_14924,N_14650);
and UO_236 (O_236,N_14921,N_14680);
xor UO_237 (O_237,N_14951,N_14431);
or UO_238 (O_238,N_14877,N_14750);
or UO_239 (O_239,N_14382,N_14432);
nor UO_240 (O_240,N_14288,N_14917);
xor UO_241 (O_241,N_14763,N_14297);
or UO_242 (O_242,N_14938,N_14908);
nand UO_243 (O_243,N_14491,N_14587);
or UO_244 (O_244,N_14622,N_14620);
or UO_245 (O_245,N_14876,N_14710);
and UO_246 (O_246,N_14952,N_14626);
and UO_247 (O_247,N_14525,N_14757);
nor UO_248 (O_248,N_14831,N_14739);
nor UO_249 (O_249,N_14256,N_14339);
nor UO_250 (O_250,N_14555,N_14447);
nand UO_251 (O_251,N_14531,N_14337);
and UO_252 (O_252,N_14534,N_14274);
xnor UO_253 (O_253,N_14879,N_14388);
xor UO_254 (O_254,N_14610,N_14905);
nor UO_255 (O_255,N_14292,N_14985);
or UO_256 (O_256,N_14384,N_14722);
xor UO_257 (O_257,N_14416,N_14412);
nand UO_258 (O_258,N_14453,N_14503);
and UO_259 (O_259,N_14695,N_14487);
and UO_260 (O_260,N_14383,N_14873);
and UO_261 (O_261,N_14727,N_14792);
nand UO_262 (O_262,N_14267,N_14820);
nand UO_263 (O_263,N_14479,N_14523);
and UO_264 (O_264,N_14529,N_14612);
nor UO_265 (O_265,N_14633,N_14699);
or UO_266 (O_266,N_14496,N_14730);
or UO_267 (O_267,N_14319,N_14914);
nand UO_268 (O_268,N_14825,N_14327);
nand UO_269 (O_269,N_14386,N_14397);
or UO_270 (O_270,N_14259,N_14364);
or UO_271 (O_271,N_14569,N_14580);
xnor UO_272 (O_272,N_14433,N_14614);
xnor UO_273 (O_273,N_14704,N_14307);
or UO_274 (O_274,N_14379,N_14565);
xnor UO_275 (O_275,N_14554,N_14672);
nor UO_276 (O_276,N_14278,N_14906);
xnor UO_277 (O_277,N_14663,N_14573);
nand UO_278 (O_278,N_14647,N_14823);
or UO_279 (O_279,N_14984,N_14838);
xor UO_280 (O_280,N_14536,N_14411);
nand UO_281 (O_281,N_14262,N_14987);
xnor UO_282 (O_282,N_14948,N_14405);
and UO_283 (O_283,N_14688,N_14904);
nor UO_284 (O_284,N_14761,N_14994);
xnor UO_285 (O_285,N_14371,N_14521);
xnor UO_286 (O_286,N_14537,N_14355);
nand UO_287 (O_287,N_14363,N_14630);
xor UO_288 (O_288,N_14609,N_14408);
nor UO_289 (O_289,N_14467,N_14409);
nand UO_290 (O_290,N_14768,N_14377);
nand UO_291 (O_291,N_14619,N_14354);
or UO_292 (O_292,N_14489,N_14973);
or UO_293 (O_293,N_14826,N_14936);
and UO_294 (O_294,N_14313,N_14545);
and UO_295 (O_295,N_14272,N_14996);
nor UO_296 (O_296,N_14803,N_14510);
xor UO_297 (O_297,N_14737,N_14596);
nand UO_298 (O_298,N_14450,N_14483);
or UO_299 (O_299,N_14692,N_14451);
nand UO_300 (O_300,N_14956,N_14703);
and UO_301 (O_301,N_14575,N_14632);
nor UO_302 (O_302,N_14463,N_14446);
and UO_303 (O_303,N_14923,N_14410);
nand UO_304 (O_304,N_14519,N_14748);
xnor UO_305 (O_305,N_14581,N_14538);
or UO_306 (O_306,N_14484,N_14380);
nor UO_307 (O_307,N_14286,N_14718);
and UO_308 (O_308,N_14932,N_14698);
nor UO_309 (O_309,N_14806,N_14959);
nor UO_310 (O_310,N_14422,N_14656);
and UO_311 (O_311,N_14850,N_14571);
or UO_312 (O_312,N_14759,N_14509);
or UO_313 (O_313,N_14802,N_14662);
xnor UO_314 (O_314,N_14552,N_14498);
and UO_315 (O_315,N_14348,N_14585);
and UO_316 (O_316,N_14505,N_14653);
xnor UO_317 (O_317,N_14775,N_14769);
nor UO_318 (O_318,N_14583,N_14381);
nand UO_319 (O_319,N_14601,N_14403);
or UO_320 (O_320,N_14644,N_14971);
or UO_321 (O_321,N_14282,N_14507);
nand UO_322 (O_322,N_14725,N_14933);
xor UO_323 (O_323,N_14266,N_14665);
nor UO_324 (O_324,N_14398,N_14714);
nor UO_325 (O_325,N_14894,N_14845);
xnor UO_326 (O_326,N_14697,N_14260);
nor UO_327 (O_327,N_14440,N_14685);
and UO_328 (O_328,N_14312,N_14949);
nand UO_329 (O_329,N_14508,N_14493);
and UO_330 (O_330,N_14442,N_14548);
nor UO_331 (O_331,N_14488,N_14903);
nor UO_332 (O_332,N_14746,N_14706);
nor UO_333 (O_333,N_14604,N_14335);
and UO_334 (O_334,N_14492,N_14638);
or UO_335 (O_335,N_14713,N_14574);
and UO_336 (O_336,N_14857,N_14942);
and UO_337 (O_337,N_14895,N_14314);
or UO_338 (O_338,N_14764,N_14972);
xor UO_339 (O_339,N_14366,N_14459);
nand UO_340 (O_340,N_14738,N_14586);
or UO_341 (O_341,N_14865,N_14504);
nand UO_342 (O_342,N_14543,N_14808);
or UO_343 (O_343,N_14275,N_14481);
nand UO_344 (O_344,N_14784,N_14767);
xnor UO_345 (O_345,N_14557,N_14798);
xor UO_346 (O_346,N_14376,N_14929);
or UO_347 (O_347,N_14375,N_14827);
and UO_348 (O_348,N_14280,N_14444);
nor UO_349 (O_349,N_14589,N_14741);
or UO_350 (O_350,N_14989,N_14961);
or UO_351 (O_351,N_14268,N_14721);
nor UO_352 (O_352,N_14341,N_14454);
nor UO_353 (O_353,N_14358,N_14712);
or UO_354 (O_354,N_14964,N_14346);
xor UO_355 (O_355,N_14869,N_14369);
nand UO_356 (O_356,N_14874,N_14628);
or UO_357 (O_357,N_14593,N_14634);
or UO_358 (O_358,N_14490,N_14861);
nor UO_359 (O_359,N_14482,N_14720);
and UO_360 (O_360,N_14494,N_14729);
and UO_361 (O_361,N_14603,N_14682);
nor UO_362 (O_362,N_14287,N_14744);
xor UO_363 (O_363,N_14666,N_14648);
nor UO_364 (O_364,N_14889,N_14616);
and UO_365 (O_365,N_14661,N_14283);
and UO_366 (O_366,N_14393,N_14673);
or UO_367 (O_367,N_14743,N_14365);
or UO_368 (O_368,N_14465,N_14642);
or UO_369 (O_369,N_14443,N_14338);
nand UO_370 (O_370,N_14979,N_14608);
or UO_371 (O_371,N_14674,N_14777);
nand UO_372 (O_372,N_14549,N_14919);
nand UO_373 (O_373,N_14988,N_14887);
or UO_374 (O_374,N_14458,N_14945);
xnor UO_375 (O_375,N_14279,N_14456);
nor UO_376 (O_376,N_14389,N_14408);
nor UO_377 (O_377,N_14438,N_14296);
or UO_378 (O_378,N_14780,N_14839);
and UO_379 (O_379,N_14800,N_14408);
nor UO_380 (O_380,N_14536,N_14954);
or UO_381 (O_381,N_14569,N_14398);
xor UO_382 (O_382,N_14625,N_14662);
nand UO_383 (O_383,N_14313,N_14767);
nor UO_384 (O_384,N_14482,N_14255);
and UO_385 (O_385,N_14975,N_14288);
nand UO_386 (O_386,N_14493,N_14769);
nor UO_387 (O_387,N_14974,N_14976);
or UO_388 (O_388,N_14477,N_14757);
nand UO_389 (O_389,N_14453,N_14756);
and UO_390 (O_390,N_14461,N_14785);
or UO_391 (O_391,N_14646,N_14945);
nor UO_392 (O_392,N_14624,N_14806);
or UO_393 (O_393,N_14808,N_14966);
xnor UO_394 (O_394,N_14982,N_14643);
xor UO_395 (O_395,N_14584,N_14660);
xnor UO_396 (O_396,N_14992,N_14614);
nand UO_397 (O_397,N_14396,N_14921);
or UO_398 (O_398,N_14652,N_14372);
nand UO_399 (O_399,N_14941,N_14384);
xor UO_400 (O_400,N_14478,N_14389);
nor UO_401 (O_401,N_14728,N_14511);
xnor UO_402 (O_402,N_14565,N_14908);
nor UO_403 (O_403,N_14506,N_14485);
or UO_404 (O_404,N_14943,N_14604);
and UO_405 (O_405,N_14565,N_14981);
and UO_406 (O_406,N_14357,N_14833);
or UO_407 (O_407,N_14764,N_14496);
nand UO_408 (O_408,N_14931,N_14809);
xor UO_409 (O_409,N_14882,N_14480);
xnor UO_410 (O_410,N_14739,N_14969);
nor UO_411 (O_411,N_14612,N_14803);
xor UO_412 (O_412,N_14687,N_14634);
nand UO_413 (O_413,N_14671,N_14629);
or UO_414 (O_414,N_14848,N_14586);
nor UO_415 (O_415,N_14792,N_14881);
nand UO_416 (O_416,N_14790,N_14915);
and UO_417 (O_417,N_14294,N_14562);
and UO_418 (O_418,N_14891,N_14879);
or UO_419 (O_419,N_14760,N_14947);
nor UO_420 (O_420,N_14985,N_14905);
xnor UO_421 (O_421,N_14403,N_14295);
nor UO_422 (O_422,N_14845,N_14745);
and UO_423 (O_423,N_14563,N_14286);
or UO_424 (O_424,N_14843,N_14302);
or UO_425 (O_425,N_14733,N_14954);
or UO_426 (O_426,N_14988,N_14886);
or UO_427 (O_427,N_14921,N_14730);
and UO_428 (O_428,N_14585,N_14367);
and UO_429 (O_429,N_14618,N_14400);
nand UO_430 (O_430,N_14700,N_14952);
xnor UO_431 (O_431,N_14556,N_14806);
xor UO_432 (O_432,N_14811,N_14711);
xor UO_433 (O_433,N_14325,N_14448);
or UO_434 (O_434,N_14957,N_14443);
nand UO_435 (O_435,N_14533,N_14647);
and UO_436 (O_436,N_14930,N_14544);
nand UO_437 (O_437,N_14677,N_14797);
or UO_438 (O_438,N_14695,N_14328);
xnor UO_439 (O_439,N_14524,N_14334);
nor UO_440 (O_440,N_14568,N_14646);
or UO_441 (O_441,N_14466,N_14648);
nand UO_442 (O_442,N_14280,N_14985);
or UO_443 (O_443,N_14836,N_14590);
xnor UO_444 (O_444,N_14388,N_14717);
nand UO_445 (O_445,N_14602,N_14767);
nor UO_446 (O_446,N_14739,N_14329);
xor UO_447 (O_447,N_14542,N_14338);
nor UO_448 (O_448,N_14288,N_14896);
nor UO_449 (O_449,N_14620,N_14298);
xor UO_450 (O_450,N_14907,N_14954);
and UO_451 (O_451,N_14770,N_14442);
and UO_452 (O_452,N_14854,N_14638);
and UO_453 (O_453,N_14344,N_14313);
xor UO_454 (O_454,N_14694,N_14741);
nor UO_455 (O_455,N_14266,N_14518);
nand UO_456 (O_456,N_14987,N_14934);
or UO_457 (O_457,N_14851,N_14848);
nor UO_458 (O_458,N_14521,N_14827);
xnor UO_459 (O_459,N_14420,N_14368);
nand UO_460 (O_460,N_14271,N_14678);
nor UO_461 (O_461,N_14607,N_14554);
or UO_462 (O_462,N_14532,N_14685);
nor UO_463 (O_463,N_14965,N_14396);
nand UO_464 (O_464,N_14806,N_14918);
xor UO_465 (O_465,N_14708,N_14754);
nand UO_466 (O_466,N_14364,N_14543);
nand UO_467 (O_467,N_14898,N_14563);
nand UO_468 (O_468,N_14980,N_14922);
nor UO_469 (O_469,N_14359,N_14338);
xor UO_470 (O_470,N_14677,N_14880);
nand UO_471 (O_471,N_14539,N_14308);
nand UO_472 (O_472,N_14499,N_14505);
xor UO_473 (O_473,N_14386,N_14389);
and UO_474 (O_474,N_14526,N_14737);
nand UO_475 (O_475,N_14746,N_14819);
or UO_476 (O_476,N_14915,N_14800);
nand UO_477 (O_477,N_14686,N_14407);
nor UO_478 (O_478,N_14308,N_14704);
or UO_479 (O_479,N_14655,N_14918);
or UO_480 (O_480,N_14819,N_14260);
nand UO_481 (O_481,N_14687,N_14371);
or UO_482 (O_482,N_14401,N_14953);
nor UO_483 (O_483,N_14880,N_14466);
and UO_484 (O_484,N_14681,N_14426);
nand UO_485 (O_485,N_14655,N_14385);
xnor UO_486 (O_486,N_14276,N_14471);
nor UO_487 (O_487,N_14839,N_14361);
xnor UO_488 (O_488,N_14252,N_14868);
xnor UO_489 (O_489,N_14897,N_14670);
or UO_490 (O_490,N_14885,N_14323);
nand UO_491 (O_491,N_14991,N_14354);
and UO_492 (O_492,N_14789,N_14717);
xor UO_493 (O_493,N_14922,N_14281);
nor UO_494 (O_494,N_14432,N_14609);
or UO_495 (O_495,N_14286,N_14295);
nor UO_496 (O_496,N_14338,N_14394);
nand UO_497 (O_497,N_14749,N_14443);
or UO_498 (O_498,N_14591,N_14837);
nor UO_499 (O_499,N_14539,N_14278);
nand UO_500 (O_500,N_14425,N_14696);
xor UO_501 (O_501,N_14649,N_14997);
and UO_502 (O_502,N_14454,N_14843);
nand UO_503 (O_503,N_14323,N_14692);
or UO_504 (O_504,N_14301,N_14882);
nand UO_505 (O_505,N_14604,N_14287);
and UO_506 (O_506,N_14708,N_14795);
and UO_507 (O_507,N_14503,N_14795);
nand UO_508 (O_508,N_14597,N_14900);
nand UO_509 (O_509,N_14294,N_14577);
xor UO_510 (O_510,N_14592,N_14985);
and UO_511 (O_511,N_14521,N_14909);
xnor UO_512 (O_512,N_14472,N_14338);
and UO_513 (O_513,N_14470,N_14558);
or UO_514 (O_514,N_14262,N_14524);
nand UO_515 (O_515,N_14590,N_14260);
or UO_516 (O_516,N_14780,N_14582);
or UO_517 (O_517,N_14505,N_14691);
and UO_518 (O_518,N_14900,N_14586);
nor UO_519 (O_519,N_14415,N_14957);
and UO_520 (O_520,N_14404,N_14846);
nand UO_521 (O_521,N_14531,N_14723);
nor UO_522 (O_522,N_14581,N_14713);
xor UO_523 (O_523,N_14978,N_14908);
xor UO_524 (O_524,N_14726,N_14770);
and UO_525 (O_525,N_14995,N_14946);
nand UO_526 (O_526,N_14795,N_14920);
nor UO_527 (O_527,N_14563,N_14702);
nand UO_528 (O_528,N_14604,N_14503);
and UO_529 (O_529,N_14594,N_14901);
or UO_530 (O_530,N_14303,N_14764);
xor UO_531 (O_531,N_14317,N_14359);
nor UO_532 (O_532,N_14752,N_14948);
xnor UO_533 (O_533,N_14795,N_14970);
nand UO_534 (O_534,N_14585,N_14586);
xnor UO_535 (O_535,N_14322,N_14378);
nor UO_536 (O_536,N_14981,N_14281);
xor UO_537 (O_537,N_14250,N_14786);
nand UO_538 (O_538,N_14953,N_14796);
or UO_539 (O_539,N_14893,N_14372);
and UO_540 (O_540,N_14953,N_14685);
and UO_541 (O_541,N_14631,N_14407);
nor UO_542 (O_542,N_14411,N_14714);
xnor UO_543 (O_543,N_14374,N_14961);
or UO_544 (O_544,N_14865,N_14720);
or UO_545 (O_545,N_14585,N_14890);
xnor UO_546 (O_546,N_14736,N_14929);
or UO_547 (O_547,N_14505,N_14408);
or UO_548 (O_548,N_14497,N_14631);
or UO_549 (O_549,N_14720,N_14650);
xor UO_550 (O_550,N_14550,N_14538);
xor UO_551 (O_551,N_14874,N_14530);
nand UO_552 (O_552,N_14819,N_14288);
nand UO_553 (O_553,N_14295,N_14632);
and UO_554 (O_554,N_14421,N_14784);
nor UO_555 (O_555,N_14770,N_14836);
xor UO_556 (O_556,N_14605,N_14743);
nor UO_557 (O_557,N_14690,N_14253);
nand UO_558 (O_558,N_14289,N_14311);
and UO_559 (O_559,N_14912,N_14660);
nor UO_560 (O_560,N_14747,N_14756);
or UO_561 (O_561,N_14543,N_14653);
xor UO_562 (O_562,N_14432,N_14936);
and UO_563 (O_563,N_14401,N_14638);
nand UO_564 (O_564,N_14869,N_14809);
nor UO_565 (O_565,N_14566,N_14586);
nor UO_566 (O_566,N_14662,N_14744);
nor UO_567 (O_567,N_14938,N_14394);
xor UO_568 (O_568,N_14889,N_14463);
and UO_569 (O_569,N_14726,N_14894);
nor UO_570 (O_570,N_14609,N_14662);
or UO_571 (O_571,N_14454,N_14271);
nor UO_572 (O_572,N_14614,N_14758);
and UO_573 (O_573,N_14748,N_14580);
xor UO_574 (O_574,N_14867,N_14487);
xor UO_575 (O_575,N_14370,N_14377);
nor UO_576 (O_576,N_14573,N_14639);
nand UO_577 (O_577,N_14805,N_14776);
or UO_578 (O_578,N_14754,N_14527);
or UO_579 (O_579,N_14942,N_14617);
xnor UO_580 (O_580,N_14756,N_14492);
xnor UO_581 (O_581,N_14684,N_14726);
nor UO_582 (O_582,N_14353,N_14865);
or UO_583 (O_583,N_14268,N_14740);
or UO_584 (O_584,N_14415,N_14366);
and UO_585 (O_585,N_14676,N_14429);
nor UO_586 (O_586,N_14939,N_14387);
or UO_587 (O_587,N_14679,N_14439);
xnor UO_588 (O_588,N_14678,N_14944);
xor UO_589 (O_589,N_14283,N_14616);
nand UO_590 (O_590,N_14761,N_14913);
and UO_591 (O_591,N_14980,N_14710);
and UO_592 (O_592,N_14410,N_14508);
nand UO_593 (O_593,N_14737,N_14521);
nand UO_594 (O_594,N_14621,N_14930);
nor UO_595 (O_595,N_14678,N_14634);
nand UO_596 (O_596,N_14980,N_14884);
xnor UO_597 (O_597,N_14323,N_14730);
xor UO_598 (O_598,N_14731,N_14573);
nor UO_599 (O_599,N_14879,N_14632);
nor UO_600 (O_600,N_14512,N_14838);
nand UO_601 (O_601,N_14849,N_14902);
nor UO_602 (O_602,N_14892,N_14811);
nor UO_603 (O_603,N_14372,N_14739);
and UO_604 (O_604,N_14393,N_14809);
and UO_605 (O_605,N_14525,N_14747);
xnor UO_606 (O_606,N_14879,N_14704);
xnor UO_607 (O_607,N_14613,N_14297);
nand UO_608 (O_608,N_14796,N_14891);
nand UO_609 (O_609,N_14361,N_14733);
nand UO_610 (O_610,N_14408,N_14307);
or UO_611 (O_611,N_14466,N_14424);
nor UO_612 (O_612,N_14851,N_14286);
xor UO_613 (O_613,N_14283,N_14818);
and UO_614 (O_614,N_14403,N_14923);
or UO_615 (O_615,N_14683,N_14264);
and UO_616 (O_616,N_14281,N_14316);
xnor UO_617 (O_617,N_14739,N_14816);
or UO_618 (O_618,N_14564,N_14897);
or UO_619 (O_619,N_14436,N_14399);
nand UO_620 (O_620,N_14995,N_14268);
nand UO_621 (O_621,N_14969,N_14618);
xor UO_622 (O_622,N_14833,N_14695);
or UO_623 (O_623,N_14562,N_14341);
xor UO_624 (O_624,N_14280,N_14483);
nor UO_625 (O_625,N_14758,N_14700);
nor UO_626 (O_626,N_14580,N_14440);
and UO_627 (O_627,N_14708,N_14385);
and UO_628 (O_628,N_14445,N_14915);
or UO_629 (O_629,N_14871,N_14783);
xnor UO_630 (O_630,N_14841,N_14686);
nand UO_631 (O_631,N_14903,N_14521);
or UO_632 (O_632,N_14984,N_14732);
or UO_633 (O_633,N_14950,N_14840);
nor UO_634 (O_634,N_14742,N_14802);
nand UO_635 (O_635,N_14583,N_14790);
or UO_636 (O_636,N_14658,N_14323);
xnor UO_637 (O_637,N_14964,N_14453);
nand UO_638 (O_638,N_14574,N_14648);
nand UO_639 (O_639,N_14971,N_14560);
or UO_640 (O_640,N_14357,N_14822);
xor UO_641 (O_641,N_14995,N_14652);
nor UO_642 (O_642,N_14361,N_14523);
xor UO_643 (O_643,N_14272,N_14463);
xnor UO_644 (O_644,N_14414,N_14516);
or UO_645 (O_645,N_14373,N_14817);
nor UO_646 (O_646,N_14729,N_14866);
xnor UO_647 (O_647,N_14947,N_14554);
nand UO_648 (O_648,N_14903,N_14359);
xor UO_649 (O_649,N_14926,N_14268);
nand UO_650 (O_650,N_14909,N_14293);
and UO_651 (O_651,N_14920,N_14995);
xor UO_652 (O_652,N_14321,N_14716);
and UO_653 (O_653,N_14479,N_14662);
and UO_654 (O_654,N_14644,N_14258);
and UO_655 (O_655,N_14855,N_14679);
nand UO_656 (O_656,N_14901,N_14495);
or UO_657 (O_657,N_14721,N_14452);
nor UO_658 (O_658,N_14688,N_14327);
and UO_659 (O_659,N_14584,N_14753);
and UO_660 (O_660,N_14324,N_14957);
nand UO_661 (O_661,N_14796,N_14983);
or UO_662 (O_662,N_14950,N_14855);
nor UO_663 (O_663,N_14676,N_14898);
and UO_664 (O_664,N_14994,N_14402);
and UO_665 (O_665,N_14605,N_14319);
or UO_666 (O_666,N_14824,N_14600);
nand UO_667 (O_667,N_14633,N_14362);
nor UO_668 (O_668,N_14555,N_14265);
xor UO_669 (O_669,N_14884,N_14410);
and UO_670 (O_670,N_14517,N_14255);
nand UO_671 (O_671,N_14421,N_14556);
or UO_672 (O_672,N_14499,N_14840);
or UO_673 (O_673,N_14890,N_14310);
and UO_674 (O_674,N_14846,N_14769);
and UO_675 (O_675,N_14665,N_14467);
and UO_676 (O_676,N_14508,N_14821);
xor UO_677 (O_677,N_14746,N_14957);
xnor UO_678 (O_678,N_14499,N_14990);
and UO_679 (O_679,N_14958,N_14874);
nor UO_680 (O_680,N_14347,N_14436);
nand UO_681 (O_681,N_14258,N_14745);
and UO_682 (O_682,N_14521,N_14984);
and UO_683 (O_683,N_14806,N_14935);
nor UO_684 (O_684,N_14251,N_14590);
nor UO_685 (O_685,N_14796,N_14637);
nand UO_686 (O_686,N_14633,N_14385);
and UO_687 (O_687,N_14377,N_14701);
or UO_688 (O_688,N_14708,N_14880);
nor UO_689 (O_689,N_14991,N_14441);
xnor UO_690 (O_690,N_14333,N_14552);
xnor UO_691 (O_691,N_14616,N_14335);
and UO_692 (O_692,N_14335,N_14421);
nor UO_693 (O_693,N_14690,N_14272);
or UO_694 (O_694,N_14620,N_14522);
nor UO_695 (O_695,N_14622,N_14916);
and UO_696 (O_696,N_14827,N_14769);
nand UO_697 (O_697,N_14707,N_14290);
and UO_698 (O_698,N_14717,N_14926);
or UO_699 (O_699,N_14252,N_14831);
or UO_700 (O_700,N_14663,N_14694);
nand UO_701 (O_701,N_14296,N_14343);
nand UO_702 (O_702,N_14765,N_14387);
xor UO_703 (O_703,N_14796,N_14291);
and UO_704 (O_704,N_14779,N_14622);
nor UO_705 (O_705,N_14527,N_14858);
or UO_706 (O_706,N_14321,N_14875);
or UO_707 (O_707,N_14454,N_14575);
nand UO_708 (O_708,N_14750,N_14415);
or UO_709 (O_709,N_14730,N_14494);
nand UO_710 (O_710,N_14855,N_14927);
or UO_711 (O_711,N_14347,N_14272);
or UO_712 (O_712,N_14802,N_14583);
xor UO_713 (O_713,N_14827,N_14442);
nand UO_714 (O_714,N_14381,N_14613);
or UO_715 (O_715,N_14819,N_14829);
or UO_716 (O_716,N_14328,N_14754);
nor UO_717 (O_717,N_14404,N_14543);
and UO_718 (O_718,N_14807,N_14602);
and UO_719 (O_719,N_14293,N_14859);
or UO_720 (O_720,N_14677,N_14517);
xnor UO_721 (O_721,N_14721,N_14979);
nand UO_722 (O_722,N_14293,N_14341);
nand UO_723 (O_723,N_14827,N_14572);
or UO_724 (O_724,N_14519,N_14723);
and UO_725 (O_725,N_14347,N_14988);
xnor UO_726 (O_726,N_14810,N_14888);
and UO_727 (O_727,N_14763,N_14352);
or UO_728 (O_728,N_14745,N_14402);
and UO_729 (O_729,N_14866,N_14675);
nor UO_730 (O_730,N_14902,N_14937);
and UO_731 (O_731,N_14280,N_14473);
nand UO_732 (O_732,N_14260,N_14621);
and UO_733 (O_733,N_14817,N_14381);
or UO_734 (O_734,N_14520,N_14272);
or UO_735 (O_735,N_14683,N_14508);
or UO_736 (O_736,N_14900,N_14400);
nor UO_737 (O_737,N_14542,N_14987);
nor UO_738 (O_738,N_14812,N_14833);
nand UO_739 (O_739,N_14718,N_14270);
xor UO_740 (O_740,N_14450,N_14821);
and UO_741 (O_741,N_14766,N_14795);
or UO_742 (O_742,N_14893,N_14408);
and UO_743 (O_743,N_14507,N_14590);
or UO_744 (O_744,N_14316,N_14687);
or UO_745 (O_745,N_14542,N_14696);
nor UO_746 (O_746,N_14714,N_14421);
nor UO_747 (O_747,N_14474,N_14643);
nand UO_748 (O_748,N_14583,N_14382);
and UO_749 (O_749,N_14257,N_14635);
nor UO_750 (O_750,N_14437,N_14588);
and UO_751 (O_751,N_14631,N_14703);
and UO_752 (O_752,N_14310,N_14297);
xnor UO_753 (O_753,N_14354,N_14348);
nand UO_754 (O_754,N_14273,N_14568);
or UO_755 (O_755,N_14754,N_14587);
nor UO_756 (O_756,N_14852,N_14741);
nand UO_757 (O_757,N_14481,N_14944);
or UO_758 (O_758,N_14922,N_14517);
or UO_759 (O_759,N_14738,N_14972);
nor UO_760 (O_760,N_14676,N_14637);
xnor UO_761 (O_761,N_14622,N_14495);
nor UO_762 (O_762,N_14934,N_14291);
xor UO_763 (O_763,N_14918,N_14844);
nor UO_764 (O_764,N_14911,N_14971);
nand UO_765 (O_765,N_14368,N_14735);
and UO_766 (O_766,N_14825,N_14754);
and UO_767 (O_767,N_14432,N_14822);
and UO_768 (O_768,N_14847,N_14621);
or UO_769 (O_769,N_14638,N_14440);
or UO_770 (O_770,N_14693,N_14984);
or UO_771 (O_771,N_14820,N_14736);
xor UO_772 (O_772,N_14517,N_14330);
and UO_773 (O_773,N_14347,N_14910);
and UO_774 (O_774,N_14513,N_14368);
xnor UO_775 (O_775,N_14598,N_14738);
nand UO_776 (O_776,N_14760,N_14517);
xnor UO_777 (O_777,N_14327,N_14635);
or UO_778 (O_778,N_14388,N_14623);
nand UO_779 (O_779,N_14286,N_14712);
or UO_780 (O_780,N_14668,N_14978);
or UO_781 (O_781,N_14887,N_14590);
and UO_782 (O_782,N_14716,N_14929);
or UO_783 (O_783,N_14356,N_14531);
xnor UO_784 (O_784,N_14718,N_14675);
or UO_785 (O_785,N_14484,N_14653);
xor UO_786 (O_786,N_14664,N_14843);
nand UO_787 (O_787,N_14392,N_14758);
nand UO_788 (O_788,N_14256,N_14653);
xnor UO_789 (O_789,N_14710,N_14347);
xnor UO_790 (O_790,N_14507,N_14530);
nand UO_791 (O_791,N_14341,N_14423);
and UO_792 (O_792,N_14907,N_14857);
and UO_793 (O_793,N_14557,N_14833);
and UO_794 (O_794,N_14678,N_14375);
nor UO_795 (O_795,N_14656,N_14526);
nand UO_796 (O_796,N_14366,N_14411);
and UO_797 (O_797,N_14983,N_14887);
xnor UO_798 (O_798,N_14541,N_14926);
nor UO_799 (O_799,N_14837,N_14484);
nor UO_800 (O_800,N_14702,N_14425);
nor UO_801 (O_801,N_14717,N_14570);
nor UO_802 (O_802,N_14282,N_14498);
or UO_803 (O_803,N_14971,N_14923);
or UO_804 (O_804,N_14929,N_14422);
nand UO_805 (O_805,N_14620,N_14986);
xnor UO_806 (O_806,N_14664,N_14693);
or UO_807 (O_807,N_14558,N_14889);
xor UO_808 (O_808,N_14928,N_14261);
nand UO_809 (O_809,N_14693,N_14685);
and UO_810 (O_810,N_14553,N_14850);
nand UO_811 (O_811,N_14987,N_14919);
and UO_812 (O_812,N_14611,N_14309);
and UO_813 (O_813,N_14681,N_14488);
and UO_814 (O_814,N_14569,N_14579);
and UO_815 (O_815,N_14558,N_14543);
nor UO_816 (O_816,N_14488,N_14852);
nand UO_817 (O_817,N_14414,N_14342);
nor UO_818 (O_818,N_14708,N_14943);
xnor UO_819 (O_819,N_14375,N_14731);
nor UO_820 (O_820,N_14561,N_14378);
nand UO_821 (O_821,N_14393,N_14845);
and UO_822 (O_822,N_14927,N_14774);
nor UO_823 (O_823,N_14856,N_14524);
or UO_824 (O_824,N_14662,N_14677);
xnor UO_825 (O_825,N_14404,N_14922);
or UO_826 (O_826,N_14736,N_14726);
nand UO_827 (O_827,N_14908,N_14372);
nand UO_828 (O_828,N_14343,N_14499);
xor UO_829 (O_829,N_14790,N_14935);
xnor UO_830 (O_830,N_14463,N_14931);
or UO_831 (O_831,N_14320,N_14482);
xor UO_832 (O_832,N_14814,N_14974);
xnor UO_833 (O_833,N_14694,N_14429);
nor UO_834 (O_834,N_14478,N_14599);
nand UO_835 (O_835,N_14675,N_14836);
xnor UO_836 (O_836,N_14858,N_14709);
nand UO_837 (O_837,N_14804,N_14558);
and UO_838 (O_838,N_14461,N_14968);
xnor UO_839 (O_839,N_14460,N_14434);
and UO_840 (O_840,N_14940,N_14619);
xor UO_841 (O_841,N_14594,N_14676);
nor UO_842 (O_842,N_14603,N_14847);
nor UO_843 (O_843,N_14485,N_14660);
or UO_844 (O_844,N_14808,N_14812);
or UO_845 (O_845,N_14402,N_14878);
xnor UO_846 (O_846,N_14668,N_14865);
xnor UO_847 (O_847,N_14487,N_14261);
xnor UO_848 (O_848,N_14471,N_14622);
or UO_849 (O_849,N_14281,N_14526);
and UO_850 (O_850,N_14632,N_14813);
nand UO_851 (O_851,N_14254,N_14620);
nor UO_852 (O_852,N_14839,N_14480);
xnor UO_853 (O_853,N_14423,N_14535);
xor UO_854 (O_854,N_14627,N_14501);
or UO_855 (O_855,N_14368,N_14631);
nor UO_856 (O_856,N_14991,N_14848);
and UO_857 (O_857,N_14335,N_14533);
or UO_858 (O_858,N_14901,N_14837);
nor UO_859 (O_859,N_14653,N_14548);
and UO_860 (O_860,N_14642,N_14412);
and UO_861 (O_861,N_14898,N_14707);
and UO_862 (O_862,N_14988,N_14596);
and UO_863 (O_863,N_14477,N_14892);
nand UO_864 (O_864,N_14923,N_14456);
and UO_865 (O_865,N_14255,N_14461);
nand UO_866 (O_866,N_14378,N_14318);
and UO_867 (O_867,N_14747,N_14768);
nor UO_868 (O_868,N_14616,N_14876);
or UO_869 (O_869,N_14618,N_14906);
xor UO_870 (O_870,N_14979,N_14410);
or UO_871 (O_871,N_14251,N_14914);
or UO_872 (O_872,N_14458,N_14826);
or UO_873 (O_873,N_14778,N_14429);
or UO_874 (O_874,N_14928,N_14424);
or UO_875 (O_875,N_14516,N_14281);
and UO_876 (O_876,N_14756,N_14379);
nand UO_877 (O_877,N_14501,N_14619);
nor UO_878 (O_878,N_14504,N_14413);
or UO_879 (O_879,N_14545,N_14827);
and UO_880 (O_880,N_14376,N_14745);
nand UO_881 (O_881,N_14783,N_14960);
or UO_882 (O_882,N_14498,N_14365);
nor UO_883 (O_883,N_14644,N_14578);
nor UO_884 (O_884,N_14887,N_14872);
nand UO_885 (O_885,N_14645,N_14998);
nor UO_886 (O_886,N_14392,N_14432);
nor UO_887 (O_887,N_14551,N_14921);
nand UO_888 (O_888,N_14612,N_14561);
or UO_889 (O_889,N_14835,N_14766);
or UO_890 (O_890,N_14992,N_14482);
and UO_891 (O_891,N_14582,N_14321);
xnor UO_892 (O_892,N_14432,N_14348);
or UO_893 (O_893,N_14869,N_14332);
nor UO_894 (O_894,N_14681,N_14929);
nand UO_895 (O_895,N_14630,N_14383);
or UO_896 (O_896,N_14638,N_14990);
nor UO_897 (O_897,N_14343,N_14563);
xnor UO_898 (O_898,N_14402,N_14903);
and UO_899 (O_899,N_14721,N_14758);
or UO_900 (O_900,N_14647,N_14897);
and UO_901 (O_901,N_14298,N_14845);
xnor UO_902 (O_902,N_14909,N_14585);
or UO_903 (O_903,N_14277,N_14795);
and UO_904 (O_904,N_14720,N_14732);
xor UO_905 (O_905,N_14591,N_14604);
and UO_906 (O_906,N_14352,N_14935);
xnor UO_907 (O_907,N_14767,N_14350);
nand UO_908 (O_908,N_14453,N_14884);
xor UO_909 (O_909,N_14957,N_14400);
or UO_910 (O_910,N_14480,N_14917);
nor UO_911 (O_911,N_14554,N_14557);
nor UO_912 (O_912,N_14501,N_14636);
and UO_913 (O_913,N_14386,N_14464);
nand UO_914 (O_914,N_14360,N_14876);
nand UO_915 (O_915,N_14935,N_14976);
and UO_916 (O_916,N_14921,N_14928);
xor UO_917 (O_917,N_14953,N_14791);
nor UO_918 (O_918,N_14593,N_14444);
nand UO_919 (O_919,N_14596,N_14704);
nor UO_920 (O_920,N_14564,N_14352);
nand UO_921 (O_921,N_14865,N_14442);
nor UO_922 (O_922,N_14272,N_14339);
nand UO_923 (O_923,N_14712,N_14860);
xor UO_924 (O_924,N_14731,N_14813);
or UO_925 (O_925,N_14898,N_14965);
xor UO_926 (O_926,N_14994,N_14474);
nand UO_927 (O_927,N_14487,N_14579);
and UO_928 (O_928,N_14772,N_14533);
nand UO_929 (O_929,N_14744,N_14438);
nand UO_930 (O_930,N_14941,N_14412);
nand UO_931 (O_931,N_14301,N_14540);
nor UO_932 (O_932,N_14728,N_14474);
nand UO_933 (O_933,N_14938,N_14520);
and UO_934 (O_934,N_14729,N_14452);
nor UO_935 (O_935,N_14913,N_14522);
or UO_936 (O_936,N_14933,N_14731);
or UO_937 (O_937,N_14460,N_14523);
nand UO_938 (O_938,N_14487,N_14599);
and UO_939 (O_939,N_14611,N_14434);
or UO_940 (O_940,N_14833,N_14785);
xor UO_941 (O_941,N_14562,N_14968);
or UO_942 (O_942,N_14457,N_14789);
nor UO_943 (O_943,N_14474,N_14325);
nand UO_944 (O_944,N_14530,N_14534);
nand UO_945 (O_945,N_14941,N_14776);
xnor UO_946 (O_946,N_14312,N_14989);
xor UO_947 (O_947,N_14544,N_14659);
nor UO_948 (O_948,N_14994,N_14473);
nand UO_949 (O_949,N_14575,N_14393);
or UO_950 (O_950,N_14590,N_14570);
xnor UO_951 (O_951,N_14455,N_14983);
xnor UO_952 (O_952,N_14932,N_14887);
nor UO_953 (O_953,N_14786,N_14747);
nand UO_954 (O_954,N_14544,N_14351);
nor UO_955 (O_955,N_14553,N_14281);
nor UO_956 (O_956,N_14952,N_14425);
nor UO_957 (O_957,N_14680,N_14260);
xor UO_958 (O_958,N_14623,N_14958);
xnor UO_959 (O_959,N_14993,N_14876);
or UO_960 (O_960,N_14925,N_14992);
xor UO_961 (O_961,N_14368,N_14737);
nand UO_962 (O_962,N_14883,N_14916);
nor UO_963 (O_963,N_14832,N_14346);
xor UO_964 (O_964,N_14795,N_14800);
and UO_965 (O_965,N_14323,N_14273);
nor UO_966 (O_966,N_14620,N_14788);
nand UO_967 (O_967,N_14567,N_14623);
or UO_968 (O_968,N_14700,N_14663);
xnor UO_969 (O_969,N_14886,N_14906);
nor UO_970 (O_970,N_14884,N_14256);
xor UO_971 (O_971,N_14677,N_14967);
xnor UO_972 (O_972,N_14575,N_14854);
and UO_973 (O_973,N_14806,N_14745);
nand UO_974 (O_974,N_14511,N_14919);
and UO_975 (O_975,N_14361,N_14765);
xnor UO_976 (O_976,N_14428,N_14727);
or UO_977 (O_977,N_14311,N_14443);
and UO_978 (O_978,N_14694,N_14919);
xnor UO_979 (O_979,N_14721,N_14458);
or UO_980 (O_980,N_14665,N_14417);
xnor UO_981 (O_981,N_14751,N_14367);
nor UO_982 (O_982,N_14522,N_14419);
and UO_983 (O_983,N_14250,N_14773);
xor UO_984 (O_984,N_14581,N_14510);
or UO_985 (O_985,N_14476,N_14537);
and UO_986 (O_986,N_14575,N_14683);
or UO_987 (O_987,N_14398,N_14937);
nor UO_988 (O_988,N_14641,N_14753);
nand UO_989 (O_989,N_14435,N_14301);
xor UO_990 (O_990,N_14444,N_14551);
or UO_991 (O_991,N_14993,N_14656);
nor UO_992 (O_992,N_14684,N_14743);
xnor UO_993 (O_993,N_14468,N_14287);
nor UO_994 (O_994,N_14665,N_14452);
nor UO_995 (O_995,N_14826,N_14280);
and UO_996 (O_996,N_14725,N_14374);
nand UO_997 (O_997,N_14404,N_14296);
or UO_998 (O_998,N_14688,N_14644);
xor UO_999 (O_999,N_14708,N_14781);
xnor UO_1000 (O_1000,N_14469,N_14844);
nand UO_1001 (O_1001,N_14810,N_14989);
or UO_1002 (O_1002,N_14978,N_14781);
nand UO_1003 (O_1003,N_14552,N_14399);
nor UO_1004 (O_1004,N_14560,N_14304);
xnor UO_1005 (O_1005,N_14539,N_14425);
nor UO_1006 (O_1006,N_14862,N_14307);
xor UO_1007 (O_1007,N_14326,N_14830);
xnor UO_1008 (O_1008,N_14784,N_14781);
xor UO_1009 (O_1009,N_14746,N_14446);
or UO_1010 (O_1010,N_14731,N_14820);
and UO_1011 (O_1011,N_14619,N_14460);
and UO_1012 (O_1012,N_14656,N_14490);
nor UO_1013 (O_1013,N_14394,N_14999);
xor UO_1014 (O_1014,N_14561,N_14349);
and UO_1015 (O_1015,N_14293,N_14422);
and UO_1016 (O_1016,N_14559,N_14919);
nand UO_1017 (O_1017,N_14937,N_14559);
and UO_1018 (O_1018,N_14585,N_14955);
and UO_1019 (O_1019,N_14816,N_14610);
nand UO_1020 (O_1020,N_14324,N_14848);
nor UO_1021 (O_1021,N_14763,N_14277);
nand UO_1022 (O_1022,N_14430,N_14296);
and UO_1023 (O_1023,N_14528,N_14789);
or UO_1024 (O_1024,N_14296,N_14250);
or UO_1025 (O_1025,N_14903,N_14552);
nor UO_1026 (O_1026,N_14254,N_14401);
and UO_1027 (O_1027,N_14272,N_14670);
nand UO_1028 (O_1028,N_14569,N_14269);
and UO_1029 (O_1029,N_14685,N_14470);
xor UO_1030 (O_1030,N_14842,N_14827);
nand UO_1031 (O_1031,N_14921,N_14344);
nand UO_1032 (O_1032,N_14912,N_14717);
and UO_1033 (O_1033,N_14525,N_14765);
nand UO_1034 (O_1034,N_14406,N_14748);
and UO_1035 (O_1035,N_14729,N_14777);
nand UO_1036 (O_1036,N_14731,N_14333);
and UO_1037 (O_1037,N_14976,N_14945);
nor UO_1038 (O_1038,N_14714,N_14522);
nand UO_1039 (O_1039,N_14701,N_14442);
nand UO_1040 (O_1040,N_14921,N_14492);
and UO_1041 (O_1041,N_14625,N_14754);
nor UO_1042 (O_1042,N_14716,N_14750);
or UO_1043 (O_1043,N_14896,N_14635);
nand UO_1044 (O_1044,N_14277,N_14451);
xnor UO_1045 (O_1045,N_14652,N_14700);
nand UO_1046 (O_1046,N_14969,N_14885);
xor UO_1047 (O_1047,N_14436,N_14643);
nand UO_1048 (O_1048,N_14376,N_14887);
xor UO_1049 (O_1049,N_14388,N_14729);
and UO_1050 (O_1050,N_14860,N_14353);
or UO_1051 (O_1051,N_14279,N_14900);
or UO_1052 (O_1052,N_14753,N_14704);
or UO_1053 (O_1053,N_14392,N_14943);
and UO_1054 (O_1054,N_14929,N_14690);
nand UO_1055 (O_1055,N_14577,N_14673);
or UO_1056 (O_1056,N_14792,N_14842);
xnor UO_1057 (O_1057,N_14990,N_14880);
nor UO_1058 (O_1058,N_14321,N_14754);
and UO_1059 (O_1059,N_14266,N_14320);
xor UO_1060 (O_1060,N_14507,N_14452);
xor UO_1061 (O_1061,N_14932,N_14745);
or UO_1062 (O_1062,N_14264,N_14847);
nor UO_1063 (O_1063,N_14399,N_14573);
and UO_1064 (O_1064,N_14510,N_14522);
nand UO_1065 (O_1065,N_14940,N_14335);
xnor UO_1066 (O_1066,N_14885,N_14664);
nor UO_1067 (O_1067,N_14446,N_14760);
xnor UO_1068 (O_1068,N_14532,N_14934);
and UO_1069 (O_1069,N_14772,N_14513);
nor UO_1070 (O_1070,N_14400,N_14959);
xnor UO_1071 (O_1071,N_14920,N_14504);
xor UO_1072 (O_1072,N_14960,N_14603);
xor UO_1073 (O_1073,N_14553,N_14708);
nand UO_1074 (O_1074,N_14276,N_14499);
and UO_1075 (O_1075,N_14431,N_14286);
nor UO_1076 (O_1076,N_14528,N_14389);
nand UO_1077 (O_1077,N_14740,N_14886);
and UO_1078 (O_1078,N_14697,N_14302);
and UO_1079 (O_1079,N_14562,N_14773);
xnor UO_1080 (O_1080,N_14724,N_14390);
xor UO_1081 (O_1081,N_14336,N_14380);
nand UO_1082 (O_1082,N_14312,N_14813);
xor UO_1083 (O_1083,N_14602,N_14569);
nand UO_1084 (O_1084,N_14323,N_14397);
nor UO_1085 (O_1085,N_14945,N_14754);
nor UO_1086 (O_1086,N_14265,N_14626);
xor UO_1087 (O_1087,N_14635,N_14571);
nor UO_1088 (O_1088,N_14395,N_14491);
xor UO_1089 (O_1089,N_14928,N_14382);
xnor UO_1090 (O_1090,N_14987,N_14317);
nor UO_1091 (O_1091,N_14402,N_14408);
xor UO_1092 (O_1092,N_14466,N_14401);
xnor UO_1093 (O_1093,N_14439,N_14682);
nor UO_1094 (O_1094,N_14711,N_14966);
xnor UO_1095 (O_1095,N_14373,N_14447);
xor UO_1096 (O_1096,N_14766,N_14726);
and UO_1097 (O_1097,N_14669,N_14325);
and UO_1098 (O_1098,N_14946,N_14410);
xnor UO_1099 (O_1099,N_14687,N_14422);
and UO_1100 (O_1100,N_14942,N_14843);
and UO_1101 (O_1101,N_14543,N_14585);
or UO_1102 (O_1102,N_14638,N_14828);
xor UO_1103 (O_1103,N_14812,N_14876);
nor UO_1104 (O_1104,N_14384,N_14829);
or UO_1105 (O_1105,N_14734,N_14721);
nand UO_1106 (O_1106,N_14601,N_14753);
and UO_1107 (O_1107,N_14570,N_14913);
or UO_1108 (O_1108,N_14769,N_14790);
nor UO_1109 (O_1109,N_14904,N_14368);
nor UO_1110 (O_1110,N_14605,N_14913);
and UO_1111 (O_1111,N_14590,N_14859);
nor UO_1112 (O_1112,N_14389,N_14924);
nor UO_1113 (O_1113,N_14407,N_14832);
nand UO_1114 (O_1114,N_14458,N_14892);
xnor UO_1115 (O_1115,N_14492,N_14597);
or UO_1116 (O_1116,N_14748,N_14995);
nor UO_1117 (O_1117,N_14414,N_14552);
xnor UO_1118 (O_1118,N_14833,N_14842);
nand UO_1119 (O_1119,N_14693,N_14701);
xnor UO_1120 (O_1120,N_14591,N_14858);
xor UO_1121 (O_1121,N_14714,N_14518);
and UO_1122 (O_1122,N_14924,N_14876);
and UO_1123 (O_1123,N_14685,N_14359);
and UO_1124 (O_1124,N_14387,N_14261);
and UO_1125 (O_1125,N_14303,N_14429);
nor UO_1126 (O_1126,N_14617,N_14500);
nand UO_1127 (O_1127,N_14866,N_14279);
nor UO_1128 (O_1128,N_14408,N_14820);
xor UO_1129 (O_1129,N_14360,N_14952);
or UO_1130 (O_1130,N_14707,N_14379);
or UO_1131 (O_1131,N_14707,N_14317);
xor UO_1132 (O_1132,N_14770,N_14580);
xnor UO_1133 (O_1133,N_14931,N_14402);
xor UO_1134 (O_1134,N_14286,N_14359);
or UO_1135 (O_1135,N_14287,N_14876);
nor UO_1136 (O_1136,N_14636,N_14353);
nand UO_1137 (O_1137,N_14474,N_14500);
or UO_1138 (O_1138,N_14844,N_14910);
nor UO_1139 (O_1139,N_14523,N_14543);
or UO_1140 (O_1140,N_14823,N_14622);
nor UO_1141 (O_1141,N_14757,N_14428);
or UO_1142 (O_1142,N_14711,N_14655);
and UO_1143 (O_1143,N_14258,N_14882);
xnor UO_1144 (O_1144,N_14686,N_14972);
xor UO_1145 (O_1145,N_14760,N_14614);
xnor UO_1146 (O_1146,N_14598,N_14259);
or UO_1147 (O_1147,N_14765,N_14986);
and UO_1148 (O_1148,N_14874,N_14749);
xnor UO_1149 (O_1149,N_14518,N_14333);
and UO_1150 (O_1150,N_14347,N_14523);
nand UO_1151 (O_1151,N_14419,N_14545);
nand UO_1152 (O_1152,N_14568,N_14616);
and UO_1153 (O_1153,N_14764,N_14306);
and UO_1154 (O_1154,N_14530,N_14935);
and UO_1155 (O_1155,N_14901,N_14341);
nand UO_1156 (O_1156,N_14665,N_14325);
or UO_1157 (O_1157,N_14319,N_14262);
or UO_1158 (O_1158,N_14380,N_14866);
nand UO_1159 (O_1159,N_14281,N_14610);
nor UO_1160 (O_1160,N_14817,N_14617);
xnor UO_1161 (O_1161,N_14299,N_14908);
xor UO_1162 (O_1162,N_14314,N_14719);
xnor UO_1163 (O_1163,N_14760,N_14487);
and UO_1164 (O_1164,N_14916,N_14430);
xnor UO_1165 (O_1165,N_14360,N_14555);
nor UO_1166 (O_1166,N_14824,N_14407);
nor UO_1167 (O_1167,N_14397,N_14307);
xor UO_1168 (O_1168,N_14892,N_14558);
nor UO_1169 (O_1169,N_14712,N_14641);
xor UO_1170 (O_1170,N_14836,N_14349);
xnor UO_1171 (O_1171,N_14528,N_14315);
and UO_1172 (O_1172,N_14381,N_14256);
or UO_1173 (O_1173,N_14977,N_14857);
and UO_1174 (O_1174,N_14908,N_14556);
nand UO_1175 (O_1175,N_14955,N_14597);
nand UO_1176 (O_1176,N_14574,N_14422);
or UO_1177 (O_1177,N_14598,N_14784);
xnor UO_1178 (O_1178,N_14505,N_14581);
nor UO_1179 (O_1179,N_14720,N_14468);
nor UO_1180 (O_1180,N_14879,N_14590);
xor UO_1181 (O_1181,N_14342,N_14799);
or UO_1182 (O_1182,N_14777,N_14995);
and UO_1183 (O_1183,N_14991,N_14590);
and UO_1184 (O_1184,N_14328,N_14968);
nand UO_1185 (O_1185,N_14515,N_14605);
and UO_1186 (O_1186,N_14535,N_14294);
and UO_1187 (O_1187,N_14534,N_14346);
or UO_1188 (O_1188,N_14976,N_14895);
xor UO_1189 (O_1189,N_14657,N_14842);
or UO_1190 (O_1190,N_14532,N_14754);
nor UO_1191 (O_1191,N_14916,N_14565);
or UO_1192 (O_1192,N_14899,N_14497);
or UO_1193 (O_1193,N_14381,N_14853);
and UO_1194 (O_1194,N_14844,N_14882);
and UO_1195 (O_1195,N_14639,N_14846);
nand UO_1196 (O_1196,N_14507,N_14589);
nand UO_1197 (O_1197,N_14643,N_14660);
nor UO_1198 (O_1198,N_14646,N_14427);
xor UO_1199 (O_1199,N_14604,N_14690);
nand UO_1200 (O_1200,N_14272,N_14535);
nand UO_1201 (O_1201,N_14309,N_14407);
nand UO_1202 (O_1202,N_14314,N_14893);
xor UO_1203 (O_1203,N_14932,N_14290);
nor UO_1204 (O_1204,N_14647,N_14785);
xor UO_1205 (O_1205,N_14780,N_14401);
and UO_1206 (O_1206,N_14768,N_14532);
xor UO_1207 (O_1207,N_14266,N_14527);
xnor UO_1208 (O_1208,N_14696,N_14459);
and UO_1209 (O_1209,N_14291,N_14984);
or UO_1210 (O_1210,N_14757,N_14770);
and UO_1211 (O_1211,N_14708,N_14616);
xor UO_1212 (O_1212,N_14793,N_14878);
and UO_1213 (O_1213,N_14758,N_14646);
nor UO_1214 (O_1214,N_14958,N_14908);
nor UO_1215 (O_1215,N_14579,N_14927);
or UO_1216 (O_1216,N_14884,N_14273);
xor UO_1217 (O_1217,N_14934,N_14303);
nor UO_1218 (O_1218,N_14831,N_14622);
and UO_1219 (O_1219,N_14925,N_14427);
or UO_1220 (O_1220,N_14658,N_14287);
or UO_1221 (O_1221,N_14721,N_14711);
nand UO_1222 (O_1222,N_14845,N_14852);
xnor UO_1223 (O_1223,N_14914,N_14607);
xnor UO_1224 (O_1224,N_14407,N_14587);
and UO_1225 (O_1225,N_14319,N_14624);
nand UO_1226 (O_1226,N_14545,N_14440);
nand UO_1227 (O_1227,N_14513,N_14267);
nand UO_1228 (O_1228,N_14660,N_14790);
and UO_1229 (O_1229,N_14311,N_14363);
and UO_1230 (O_1230,N_14850,N_14439);
and UO_1231 (O_1231,N_14551,N_14742);
and UO_1232 (O_1232,N_14305,N_14439);
or UO_1233 (O_1233,N_14987,N_14822);
xnor UO_1234 (O_1234,N_14304,N_14317);
nor UO_1235 (O_1235,N_14805,N_14454);
or UO_1236 (O_1236,N_14675,N_14952);
or UO_1237 (O_1237,N_14683,N_14512);
or UO_1238 (O_1238,N_14469,N_14506);
xnor UO_1239 (O_1239,N_14270,N_14322);
and UO_1240 (O_1240,N_14523,N_14976);
xor UO_1241 (O_1241,N_14573,N_14525);
nor UO_1242 (O_1242,N_14582,N_14611);
or UO_1243 (O_1243,N_14426,N_14640);
or UO_1244 (O_1244,N_14887,N_14583);
nand UO_1245 (O_1245,N_14325,N_14353);
xnor UO_1246 (O_1246,N_14545,N_14526);
xnor UO_1247 (O_1247,N_14867,N_14977);
and UO_1248 (O_1248,N_14398,N_14819);
xnor UO_1249 (O_1249,N_14412,N_14568);
nor UO_1250 (O_1250,N_14787,N_14735);
or UO_1251 (O_1251,N_14647,N_14983);
and UO_1252 (O_1252,N_14402,N_14872);
nand UO_1253 (O_1253,N_14325,N_14804);
nor UO_1254 (O_1254,N_14862,N_14503);
and UO_1255 (O_1255,N_14728,N_14842);
nor UO_1256 (O_1256,N_14481,N_14569);
or UO_1257 (O_1257,N_14283,N_14810);
or UO_1258 (O_1258,N_14799,N_14730);
and UO_1259 (O_1259,N_14992,N_14587);
xor UO_1260 (O_1260,N_14475,N_14371);
nand UO_1261 (O_1261,N_14676,N_14699);
and UO_1262 (O_1262,N_14308,N_14897);
nor UO_1263 (O_1263,N_14843,N_14622);
and UO_1264 (O_1264,N_14808,N_14835);
and UO_1265 (O_1265,N_14711,N_14479);
or UO_1266 (O_1266,N_14623,N_14736);
nor UO_1267 (O_1267,N_14769,N_14382);
nor UO_1268 (O_1268,N_14761,N_14436);
or UO_1269 (O_1269,N_14361,N_14767);
and UO_1270 (O_1270,N_14646,N_14287);
xnor UO_1271 (O_1271,N_14501,N_14350);
and UO_1272 (O_1272,N_14518,N_14439);
and UO_1273 (O_1273,N_14884,N_14528);
xnor UO_1274 (O_1274,N_14924,N_14695);
nor UO_1275 (O_1275,N_14532,N_14508);
and UO_1276 (O_1276,N_14665,N_14352);
xnor UO_1277 (O_1277,N_14384,N_14438);
and UO_1278 (O_1278,N_14474,N_14501);
nand UO_1279 (O_1279,N_14576,N_14382);
and UO_1280 (O_1280,N_14533,N_14894);
and UO_1281 (O_1281,N_14508,N_14709);
nor UO_1282 (O_1282,N_14871,N_14841);
xnor UO_1283 (O_1283,N_14927,N_14833);
xor UO_1284 (O_1284,N_14646,N_14800);
or UO_1285 (O_1285,N_14304,N_14861);
and UO_1286 (O_1286,N_14941,N_14475);
and UO_1287 (O_1287,N_14643,N_14586);
or UO_1288 (O_1288,N_14404,N_14703);
nor UO_1289 (O_1289,N_14451,N_14476);
and UO_1290 (O_1290,N_14928,N_14287);
or UO_1291 (O_1291,N_14883,N_14809);
nand UO_1292 (O_1292,N_14920,N_14339);
and UO_1293 (O_1293,N_14259,N_14410);
nor UO_1294 (O_1294,N_14803,N_14369);
and UO_1295 (O_1295,N_14858,N_14722);
and UO_1296 (O_1296,N_14626,N_14510);
xnor UO_1297 (O_1297,N_14502,N_14575);
xor UO_1298 (O_1298,N_14952,N_14305);
and UO_1299 (O_1299,N_14997,N_14644);
and UO_1300 (O_1300,N_14698,N_14617);
nand UO_1301 (O_1301,N_14811,N_14440);
nor UO_1302 (O_1302,N_14784,N_14835);
and UO_1303 (O_1303,N_14467,N_14860);
nand UO_1304 (O_1304,N_14439,N_14839);
xor UO_1305 (O_1305,N_14261,N_14650);
or UO_1306 (O_1306,N_14590,N_14749);
xor UO_1307 (O_1307,N_14305,N_14802);
nor UO_1308 (O_1308,N_14372,N_14673);
and UO_1309 (O_1309,N_14774,N_14808);
and UO_1310 (O_1310,N_14510,N_14273);
xor UO_1311 (O_1311,N_14579,N_14605);
nor UO_1312 (O_1312,N_14699,N_14358);
nand UO_1313 (O_1313,N_14965,N_14903);
nand UO_1314 (O_1314,N_14816,N_14676);
nor UO_1315 (O_1315,N_14581,N_14312);
nand UO_1316 (O_1316,N_14328,N_14384);
or UO_1317 (O_1317,N_14761,N_14940);
xor UO_1318 (O_1318,N_14781,N_14272);
nand UO_1319 (O_1319,N_14685,N_14783);
nand UO_1320 (O_1320,N_14691,N_14435);
nand UO_1321 (O_1321,N_14775,N_14358);
nand UO_1322 (O_1322,N_14317,N_14392);
xor UO_1323 (O_1323,N_14645,N_14886);
nor UO_1324 (O_1324,N_14518,N_14657);
xnor UO_1325 (O_1325,N_14973,N_14704);
nor UO_1326 (O_1326,N_14364,N_14938);
and UO_1327 (O_1327,N_14817,N_14988);
and UO_1328 (O_1328,N_14924,N_14500);
and UO_1329 (O_1329,N_14644,N_14338);
or UO_1330 (O_1330,N_14371,N_14977);
nand UO_1331 (O_1331,N_14251,N_14837);
nand UO_1332 (O_1332,N_14605,N_14694);
or UO_1333 (O_1333,N_14697,N_14981);
and UO_1334 (O_1334,N_14648,N_14520);
nor UO_1335 (O_1335,N_14848,N_14337);
or UO_1336 (O_1336,N_14826,N_14639);
nand UO_1337 (O_1337,N_14503,N_14647);
and UO_1338 (O_1338,N_14585,N_14728);
nor UO_1339 (O_1339,N_14885,N_14962);
xor UO_1340 (O_1340,N_14832,N_14591);
or UO_1341 (O_1341,N_14529,N_14729);
xnor UO_1342 (O_1342,N_14509,N_14720);
and UO_1343 (O_1343,N_14816,N_14329);
and UO_1344 (O_1344,N_14990,N_14966);
and UO_1345 (O_1345,N_14264,N_14654);
or UO_1346 (O_1346,N_14587,N_14374);
nand UO_1347 (O_1347,N_14467,N_14688);
nand UO_1348 (O_1348,N_14542,N_14645);
and UO_1349 (O_1349,N_14312,N_14567);
nor UO_1350 (O_1350,N_14997,N_14403);
and UO_1351 (O_1351,N_14997,N_14629);
xnor UO_1352 (O_1352,N_14325,N_14594);
nand UO_1353 (O_1353,N_14658,N_14354);
nor UO_1354 (O_1354,N_14450,N_14636);
nand UO_1355 (O_1355,N_14444,N_14584);
nand UO_1356 (O_1356,N_14551,N_14689);
or UO_1357 (O_1357,N_14416,N_14307);
xnor UO_1358 (O_1358,N_14851,N_14867);
and UO_1359 (O_1359,N_14397,N_14955);
xnor UO_1360 (O_1360,N_14484,N_14920);
nand UO_1361 (O_1361,N_14786,N_14300);
or UO_1362 (O_1362,N_14397,N_14872);
xnor UO_1363 (O_1363,N_14600,N_14521);
nand UO_1364 (O_1364,N_14657,N_14887);
xnor UO_1365 (O_1365,N_14600,N_14456);
or UO_1366 (O_1366,N_14615,N_14290);
and UO_1367 (O_1367,N_14770,N_14325);
xnor UO_1368 (O_1368,N_14352,N_14514);
and UO_1369 (O_1369,N_14369,N_14468);
nand UO_1370 (O_1370,N_14556,N_14657);
xor UO_1371 (O_1371,N_14931,N_14509);
or UO_1372 (O_1372,N_14648,N_14845);
or UO_1373 (O_1373,N_14755,N_14865);
nand UO_1374 (O_1374,N_14351,N_14799);
xor UO_1375 (O_1375,N_14352,N_14889);
nor UO_1376 (O_1376,N_14279,N_14414);
nor UO_1377 (O_1377,N_14607,N_14399);
nand UO_1378 (O_1378,N_14933,N_14648);
or UO_1379 (O_1379,N_14872,N_14483);
nand UO_1380 (O_1380,N_14403,N_14603);
xnor UO_1381 (O_1381,N_14892,N_14725);
or UO_1382 (O_1382,N_14307,N_14879);
xnor UO_1383 (O_1383,N_14701,N_14444);
and UO_1384 (O_1384,N_14859,N_14756);
nand UO_1385 (O_1385,N_14697,N_14794);
nor UO_1386 (O_1386,N_14717,N_14341);
or UO_1387 (O_1387,N_14772,N_14754);
and UO_1388 (O_1388,N_14359,N_14927);
nor UO_1389 (O_1389,N_14563,N_14356);
or UO_1390 (O_1390,N_14426,N_14274);
or UO_1391 (O_1391,N_14657,N_14336);
nor UO_1392 (O_1392,N_14664,N_14396);
or UO_1393 (O_1393,N_14279,N_14371);
or UO_1394 (O_1394,N_14298,N_14478);
xor UO_1395 (O_1395,N_14971,N_14364);
xnor UO_1396 (O_1396,N_14542,N_14820);
xor UO_1397 (O_1397,N_14625,N_14803);
xor UO_1398 (O_1398,N_14343,N_14916);
nor UO_1399 (O_1399,N_14976,N_14380);
xnor UO_1400 (O_1400,N_14725,N_14649);
nand UO_1401 (O_1401,N_14661,N_14407);
or UO_1402 (O_1402,N_14923,N_14938);
nand UO_1403 (O_1403,N_14481,N_14381);
xnor UO_1404 (O_1404,N_14408,N_14608);
or UO_1405 (O_1405,N_14503,N_14307);
nand UO_1406 (O_1406,N_14600,N_14791);
xor UO_1407 (O_1407,N_14967,N_14476);
and UO_1408 (O_1408,N_14964,N_14938);
xor UO_1409 (O_1409,N_14412,N_14921);
and UO_1410 (O_1410,N_14701,N_14300);
nand UO_1411 (O_1411,N_14547,N_14808);
nand UO_1412 (O_1412,N_14689,N_14515);
xor UO_1413 (O_1413,N_14980,N_14658);
and UO_1414 (O_1414,N_14277,N_14857);
and UO_1415 (O_1415,N_14401,N_14864);
or UO_1416 (O_1416,N_14609,N_14264);
nand UO_1417 (O_1417,N_14529,N_14325);
or UO_1418 (O_1418,N_14544,N_14426);
or UO_1419 (O_1419,N_14768,N_14870);
nand UO_1420 (O_1420,N_14592,N_14732);
nor UO_1421 (O_1421,N_14681,N_14376);
nor UO_1422 (O_1422,N_14969,N_14797);
nor UO_1423 (O_1423,N_14816,N_14348);
xor UO_1424 (O_1424,N_14786,N_14936);
xor UO_1425 (O_1425,N_14900,N_14280);
and UO_1426 (O_1426,N_14723,N_14656);
nand UO_1427 (O_1427,N_14987,N_14350);
or UO_1428 (O_1428,N_14976,N_14312);
and UO_1429 (O_1429,N_14965,N_14978);
xnor UO_1430 (O_1430,N_14703,N_14981);
and UO_1431 (O_1431,N_14407,N_14916);
nor UO_1432 (O_1432,N_14776,N_14381);
or UO_1433 (O_1433,N_14288,N_14298);
and UO_1434 (O_1434,N_14776,N_14497);
nand UO_1435 (O_1435,N_14385,N_14612);
and UO_1436 (O_1436,N_14808,N_14363);
or UO_1437 (O_1437,N_14265,N_14410);
and UO_1438 (O_1438,N_14634,N_14359);
nand UO_1439 (O_1439,N_14700,N_14556);
or UO_1440 (O_1440,N_14494,N_14575);
xnor UO_1441 (O_1441,N_14742,N_14751);
nand UO_1442 (O_1442,N_14298,N_14986);
nand UO_1443 (O_1443,N_14442,N_14610);
or UO_1444 (O_1444,N_14908,N_14307);
nor UO_1445 (O_1445,N_14807,N_14726);
nand UO_1446 (O_1446,N_14881,N_14824);
nor UO_1447 (O_1447,N_14873,N_14658);
xnor UO_1448 (O_1448,N_14379,N_14484);
nand UO_1449 (O_1449,N_14477,N_14420);
and UO_1450 (O_1450,N_14376,N_14509);
nand UO_1451 (O_1451,N_14784,N_14353);
xnor UO_1452 (O_1452,N_14759,N_14385);
nor UO_1453 (O_1453,N_14318,N_14461);
and UO_1454 (O_1454,N_14561,N_14924);
nor UO_1455 (O_1455,N_14431,N_14329);
nor UO_1456 (O_1456,N_14815,N_14813);
nand UO_1457 (O_1457,N_14597,N_14796);
and UO_1458 (O_1458,N_14914,N_14977);
or UO_1459 (O_1459,N_14279,N_14609);
nand UO_1460 (O_1460,N_14253,N_14683);
and UO_1461 (O_1461,N_14915,N_14911);
or UO_1462 (O_1462,N_14336,N_14260);
nand UO_1463 (O_1463,N_14409,N_14667);
xnor UO_1464 (O_1464,N_14743,N_14814);
nor UO_1465 (O_1465,N_14958,N_14406);
nand UO_1466 (O_1466,N_14708,N_14490);
xor UO_1467 (O_1467,N_14887,N_14981);
and UO_1468 (O_1468,N_14923,N_14972);
nor UO_1469 (O_1469,N_14781,N_14612);
nand UO_1470 (O_1470,N_14715,N_14288);
and UO_1471 (O_1471,N_14996,N_14259);
nor UO_1472 (O_1472,N_14645,N_14685);
or UO_1473 (O_1473,N_14317,N_14803);
xor UO_1474 (O_1474,N_14677,N_14454);
nand UO_1475 (O_1475,N_14852,N_14269);
or UO_1476 (O_1476,N_14799,N_14538);
nand UO_1477 (O_1477,N_14552,N_14975);
xor UO_1478 (O_1478,N_14410,N_14656);
nor UO_1479 (O_1479,N_14881,N_14674);
nor UO_1480 (O_1480,N_14582,N_14837);
nor UO_1481 (O_1481,N_14556,N_14706);
nand UO_1482 (O_1482,N_14674,N_14305);
or UO_1483 (O_1483,N_14759,N_14396);
xor UO_1484 (O_1484,N_14301,N_14481);
nand UO_1485 (O_1485,N_14739,N_14765);
xnor UO_1486 (O_1486,N_14748,N_14262);
and UO_1487 (O_1487,N_14591,N_14393);
nand UO_1488 (O_1488,N_14420,N_14383);
or UO_1489 (O_1489,N_14277,N_14952);
nor UO_1490 (O_1490,N_14615,N_14744);
and UO_1491 (O_1491,N_14468,N_14563);
xnor UO_1492 (O_1492,N_14793,N_14461);
nor UO_1493 (O_1493,N_14342,N_14513);
nand UO_1494 (O_1494,N_14651,N_14778);
or UO_1495 (O_1495,N_14677,N_14425);
xnor UO_1496 (O_1496,N_14311,N_14743);
nand UO_1497 (O_1497,N_14880,N_14253);
or UO_1498 (O_1498,N_14557,N_14955);
nand UO_1499 (O_1499,N_14713,N_14778);
xnor UO_1500 (O_1500,N_14402,N_14279);
and UO_1501 (O_1501,N_14747,N_14664);
nand UO_1502 (O_1502,N_14486,N_14306);
and UO_1503 (O_1503,N_14827,N_14532);
xnor UO_1504 (O_1504,N_14888,N_14751);
nand UO_1505 (O_1505,N_14697,N_14783);
and UO_1506 (O_1506,N_14316,N_14818);
xor UO_1507 (O_1507,N_14764,N_14553);
nor UO_1508 (O_1508,N_14451,N_14259);
and UO_1509 (O_1509,N_14925,N_14659);
nor UO_1510 (O_1510,N_14779,N_14429);
and UO_1511 (O_1511,N_14816,N_14834);
xor UO_1512 (O_1512,N_14768,N_14853);
nor UO_1513 (O_1513,N_14623,N_14894);
nor UO_1514 (O_1514,N_14586,N_14339);
nand UO_1515 (O_1515,N_14778,N_14715);
and UO_1516 (O_1516,N_14818,N_14740);
nor UO_1517 (O_1517,N_14500,N_14798);
or UO_1518 (O_1518,N_14871,N_14359);
xor UO_1519 (O_1519,N_14662,N_14304);
nor UO_1520 (O_1520,N_14744,N_14709);
nor UO_1521 (O_1521,N_14837,N_14662);
and UO_1522 (O_1522,N_14611,N_14739);
or UO_1523 (O_1523,N_14457,N_14292);
nand UO_1524 (O_1524,N_14413,N_14940);
nor UO_1525 (O_1525,N_14846,N_14383);
or UO_1526 (O_1526,N_14368,N_14419);
nand UO_1527 (O_1527,N_14451,N_14440);
and UO_1528 (O_1528,N_14732,N_14467);
and UO_1529 (O_1529,N_14414,N_14575);
nor UO_1530 (O_1530,N_14692,N_14690);
nor UO_1531 (O_1531,N_14558,N_14999);
and UO_1532 (O_1532,N_14834,N_14546);
nand UO_1533 (O_1533,N_14467,N_14364);
nor UO_1534 (O_1534,N_14625,N_14752);
nor UO_1535 (O_1535,N_14597,N_14289);
nor UO_1536 (O_1536,N_14951,N_14404);
or UO_1537 (O_1537,N_14773,N_14342);
nor UO_1538 (O_1538,N_14704,N_14931);
nand UO_1539 (O_1539,N_14698,N_14815);
nor UO_1540 (O_1540,N_14921,N_14487);
or UO_1541 (O_1541,N_14352,N_14910);
xor UO_1542 (O_1542,N_14385,N_14687);
nor UO_1543 (O_1543,N_14394,N_14738);
xnor UO_1544 (O_1544,N_14781,N_14852);
or UO_1545 (O_1545,N_14338,N_14437);
xor UO_1546 (O_1546,N_14610,N_14608);
xnor UO_1547 (O_1547,N_14704,N_14366);
nor UO_1548 (O_1548,N_14989,N_14951);
or UO_1549 (O_1549,N_14949,N_14275);
nor UO_1550 (O_1550,N_14775,N_14744);
and UO_1551 (O_1551,N_14408,N_14709);
and UO_1552 (O_1552,N_14979,N_14783);
nor UO_1553 (O_1553,N_14869,N_14745);
and UO_1554 (O_1554,N_14253,N_14357);
xor UO_1555 (O_1555,N_14701,N_14591);
and UO_1556 (O_1556,N_14542,N_14662);
and UO_1557 (O_1557,N_14615,N_14350);
or UO_1558 (O_1558,N_14440,N_14912);
nand UO_1559 (O_1559,N_14671,N_14659);
xor UO_1560 (O_1560,N_14724,N_14791);
xor UO_1561 (O_1561,N_14611,N_14314);
and UO_1562 (O_1562,N_14636,N_14936);
or UO_1563 (O_1563,N_14560,N_14321);
nand UO_1564 (O_1564,N_14326,N_14512);
and UO_1565 (O_1565,N_14951,N_14469);
nand UO_1566 (O_1566,N_14911,N_14407);
and UO_1567 (O_1567,N_14774,N_14722);
xnor UO_1568 (O_1568,N_14627,N_14736);
nor UO_1569 (O_1569,N_14791,N_14902);
nand UO_1570 (O_1570,N_14327,N_14746);
xnor UO_1571 (O_1571,N_14510,N_14909);
or UO_1572 (O_1572,N_14569,N_14819);
and UO_1573 (O_1573,N_14396,N_14352);
nor UO_1574 (O_1574,N_14772,N_14710);
xor UO_1575 (O_1575,N_14539,N_14395);
nand UO_1576 (O_1576,N_14805,N_14925);
nor UO_1577 (O_1577,N_14700,N_14593);
xor UO_1578 (O_1578,N_14978,N_14882);
or UO_1579 (O_1579,N_14344,N_14361);
nor UO_1580 (O_1580,N_14270,N_14474);
or UO_1581 (O_1581,N_14870,N_14944);
xnor UO_1582 (O_1582,N_14448,N_14939);
nor UO_1583 (O_1583,N_14493,N_14434);
nand UO_1584 (O_1584,N_14890,N_14552);
nand UO_1585 (O_1585,N_14710,N_14883);
or UO_1586 (O_1586,N_14475,N_14979);
nand UO_1587 (O_1587,N_14601,N_14475);
xor UO_1588 (O_1588,N_14463,N_14837);
xor UO_1589 (O_1589,N_14458,N_14568);
nor UO_1590 (O_1590,N_14818,N_14909);
nand UO_1591 (O_1591,N_14424,N_14257);
and UO_1592 (O_1592,N_14863,N_14871);
and UO_1593 (O_1593,N_14618,N_14673);
and UO_1594 (O_1594,N_14993,N_14577);
nor UO_1595 (O_1595,N_14647,N_14889);
nor UO_1596 (O_1596,N_14755,N_14634);
nor UO_1597 (O_1597,N_14969,N_14751);
nand UO_1598 (O_1598,N_14457,N_14617);
nor UO_1599 (O_1599,N_14557,N_14665);
or UO_1600 (O_1600,N_14405,N_14962);
xnor UO_1601 (O_1601,N_14956,N_14521);
nor UO_1602 (O_1602,N_14952,N_14339);
or UO_1603 (O_1603,N_14567,N_14628);
nor UO_1604 (O_1604,N_14818,N_14703);
xnor UO_1605 (O_1605,N_14794,N_14889);
xor UO_1606 (O_1606,N_14506,N_14319);
xor UO_1607 (O_1607,N_14559,N_14851);
and UO_1608 (O_1608,N_14735,N_14510);
xor UO_1609 (O_1609,N_14281,N_14381);
nor UO_1610 (O_1610,N_14850,N_14276);
or UO_1611 (O_1611,N_14686,N_14372);
xor UO_1612 (O_1612,N_14610,N_14822);
nor UO_1613 (O_1613,N_14555,N_14936);
xnor UO_1614 (O_1614,N_14780,N_14723);
and UO_1615 (O_1615,N_14653,N_14783);
nor UO_1616 (O_1616,N_14995,N_14649);
nor UO_1617 (O_1617,N_14580,N_14394);
nand UO_1618 (O_1618,N_14334,N_14859);
xor UO_1619 (O_1619,N_14429,N_14292);
or UO_1620 (O_1620,N_14943,N_14548);
or UO_1621 (O_1621,N_14766,N_14258);
nor UO_1622 (O_1622,N_14568,N_14949);
or UO_1623 (O_1623,N_14698,N_14725);
or UO_1624 (O_1624,N_14676,N_14379);
and UO_1625 (O_1625,N_14848,N_14765);
nand UO_1626 (O_1626,N_14767,N_14327);
nor UO_1627 (O_1627,N_14819,N_14276);
nand UO_1628 (O_1628,N_14415,N_14563);
or UO_1629 (O_1629,N_14689,N_14539);
nor UO_1630 (O_1630,N_14791,N_14673);
nor UO_1631 (O_1631,N_14286,N_14946);
xnor UO_1632 (O_1632,N_14668,N_14566);
or UO_1633 (O_1633,N_14739,N_14598);
nor UO_1634 (O_1634,N_14469,N_14533);
and UO_1635 (O_1635,N_14442,N_14340);
nor UO_1636 (O_1636,N_14861,N_14754);
and UO_1637 (O_1637,N_14913,N_14897);
nand UO_1638 (O_1638,N_14814,N_14641);
nor UO_1639 (O_1639,N_14870,N_14915);
and UO_1640 (O_1640,N_14260,N_14917);
nand UO_1641 (O_1641,N_14563,N_14807);
or UO_1642 (O_1642,N_14481,N_14693);
nor UO_1643 (O_1643,N_14512,N_14353);
nand UO_1644 (O_1644,N_14828,N_14544);
nand UO_1645 (O_1645,N_14779,N_14352);
xnor UO_1646 (O_1646,N_14453,N_14542);
or UO_1647 (O_1647,N_14864,N_14721);
or UO_1648 (O_1648,N_14500,N_14729);
xor UO_1649 (O_1649,N_14540,N_14980);
xnor UO_1650 (O_1650,N_14776,N_14600);
xor UO_1651 (O_1651,N_14432,N_14799);
nor UO_1652 (O_1652,N_14836,N_14476);
or UO_1653 (O_1653,N_14362,N_14492);
and UO_1654 (O_1654,N_14386,N_14465);
or UO_1655 (O_1655,N_14644,N_14275);
or UO_1656 (O_1656,N_14370,N_14673);
and UO_1657 (O_1657,N_14881,N_14484);
or UO_1658 (O_1658,N_14736,N_14404);
nor UO_1659 (O_1659,N_14753,N_14561);
xnor UO_1660 (O_1660,N_14750,N_14906);
nor UO_1661 (O_1661,N_14892,N_14293);
nand UO_1662 (O_1662,N_14573,N_14857);
nand UO_1663 (O_1663,N_14712,N_14934);
nor UO_1664 (O_1664,N_14551,N_14691);
nor UO_1665 (O_1665,N_14877,N_14633);
or UO_1666 (O_1666,N_14498,N_14612);
nor UO_1667 (O_1667,N_14919,N_14597);
or UO_1668 (O_1668,N_14984,N_14439);
nand UO_1669 (O_1669,N_14817,N_14419);
and UO_1670 (O_1670,N_14716,N_14259);
nor UO_1671 (O_1671,N_14697,N_14396);
and UO_1672 (O_1672,N_14985,N_14304);
or UO_1673 (O_1673,N_14919,N_14471);
or UO_1674 (O_1674,N_14994,N_14400);
or UO_1675 (O_1675,N_14989,N_14252);
xor UO_1676 (O_1676,N_14987,N_14922);
nand UO_1677 (O_1677,N_14657,N_14975);
or UO_1678 (O_1678,N_14546,N_14654);
or UO_1679 (O_1679,N_14891,N_14864);
nor UO_1680 (O_1680,N_14591,N_14437);
or UO_1681 (O_1681,N_14554,N_14788);
nor UO_1682 (O_1682,N_14363,N_14742);
nor UO_1683 (O_1683,N_14532,N_14531);
xnor UO_1684 (O_1684,N_14621,N_14888);
or UO_1685 (O_1685,N_14886,N_14395);
or UO_1686 (O_1686,N_14960,N_14626);
or UO_1687 (O_1687,N_14431,N_14629);
and UO_1688 (O_1688,N_14899,N_14946);
nand UO_1689 (O_1689,N_14799,N_14402);
nor UO_1690 (O_1690,N_14903,N_14941);
and UO_1691 (O_1691,N_14366,N_14777);
xnor UO_1692 (O_1692,N_14289,N_14637);
xor UO_1693 (O_1693,N_14277,N_14741);
nand UO_1694 (O_1694,N_14385,N_14697);
nor UO_1695 (O_1695,N_14717,N_14428);
or UO_1696 (O_1696,N_14418,N_14451);
nor UO_1697 (O_1697,N_14651,N_14264);
xor UO_1698 (O_1698,N_14739,N_14769);
xor UO_1699 (O_1699,N_14291,N_14584);
and UO_1700 (O_1700,N_14446,N_14460);
and UO_1701 (O_1701,N_14535,N_14622);
and UO_1702 (O_1702,N_14674,N_14344);
or UO_1703 (O_1703,N_14945,N_14848);
or UO_1704 (O_1704,N_14801,N_14559);
nor UO_1705 (O_1705,N_14268,N_14464);
nor UO_1706 (O_1706,N_14492,N_14704);
xor UO_1707 (O_1707,N_14393,N_14808);
or UO_1708 (O_1708,N_14480,N_14888);
xor UO_1709 (O_1709,N_14732,N_14902);
xor UO_1710 (O_1710,N_14994,N_14624);
nand UO_1711 (O_1711,N_14777,N_14330);
nand UO_1712 (O_1712,N_14856,N_14924);
nand UO_1713 (O_1713,N_14783,N_14834);
and UO_1714 (O_1714,N_14789,N_14292);
and UO_1715 (O_1715,N_14460,N_14318);
and UO_1716 (O_1716,N_14606,N_14421);
nor UO_1717 (O_1717,N_14616,N_14685);
xor UO_1718 (O_1718,N_14541,N_14635);
xnor UO_1719 (O_1719,N_14779,N_14523);
nand UO_1720 (O_1720,N_14600,N_14351);
nor UO_1721 (O_1721,N_14642,N_14924);
xnor UO_1722 (O_1722,N_14494,N_14511);
and UO_1723 (O_1723,N_14954,N_14272);
nand UO_1724 (O_1724,N_14511,N_14436);
xnor UO_1725 (O_1725,N_14581,N_14361);
nand UO_1726 (O_1726,N_14821,N_14999);
xor UO_1727 (O_1727,N_14785,N_14390);
nand UO_1728 (O_1728,N_14835,N_14771);
nand UO_1729 (O_1729,N_14798,N_14523);
and UO_1730 (O_1730,N_14419,N_14664);
nand UO_1731 (O_1731,N_14654,N_14914);
xnor UO_1732 (O_1732,N_14762,N_14511);
and UO_1733 (O_1733,N_14728,N_14524);
or UO_1734 (O_1734,N_14996,N_14685);
and UO_1735 (O_1735,N_14886,N_14904);
nand UO_1736 (O_1736,N_14901,N_14742);
nor UO_1737 (O_1737,N_14961,N_14259);
xnor UO_1738 (O_1738,N_14509,N_14914);
nand UO_1739 (O_1739,N_14931,N_14677);
or UO_1740 (O_1740,N_14465,N_14546);
xor UO_1741 (O_1741,N_14507,N_14581);
and UO_1742 (O_1742,N_14960,N_14721);
nand UO_1743 (O_1743,N_14628,N_14580);
xnor UO_1744 (O_1744,N_14352,N_14727);
nor UO_1745 (O_1745,N_14373,N_14446);
xor UO_1746 (O_1746,N_14862,N_14891);
nor UO_1747 (O_1747,N_14669,N_14482);
and UO_1748 (O_1748,N_14699,N_14559);
nor UO_1749 (O_1749,N_14390,N_14370);
xnor UO_1750 (O_1750,N_14268,N_14707);
or UO_1751 (O_1751,N_14371,N_14400);
nor UO_1752 (O_1752,N_14754,N_14389);
nor UO_1753 (O_1753,N_14514,N_14509);
nor UO_1754 (O_1754,N_14855,N_14639);
nor UO_1755 (O_1755,N_14776,N_14815);
and UO_1756 (O_1756,N_14641,N_14710);
xor UO_1757 (O_1757,N_14662,N_14804);
nor UO_1758 (O_1758,N_14520,N_14974);
nand UO_1759 (O_1759,N_14547,N_14762);
xor UO_1760 (O_1760,N_14291,N_14403);
nand UO_1761 (O_1761,N_14962,N_14649);
nand UO_1762 (O_1762,N_14528,N_14318);
or UO_1763 (O_1763,N_14546,N_14758);
and UO_1764 (O_1764,N_14646,N_14588);
nor UO_1765 (O_1765,N_14788,N_14327);
nor UO_1766 (O_1766,N_14529,N_14911);
and UO_1767 (O_1767,N_14864,N_14329);
or UO_1768 (O_1768,N_14608,N_14950);
xor UO_1769 (O_1769,N_14813,N_14288);
and UO_1770 (O_1770,N_14487,N_14794);
and UO_1771 (O_1771,N_14265,N_14772);
nand UO_1772 (O_1772,N_14409,N_14602);
nor UO_1773 (O_1773,N_14759,N_14572);
nor UO_1774 (O_1774,N_14976,N_14782);
nor UO_1775 (O_1775,N_14290,N_14377);
or UO_1776 (O_1776,N_14358,N_14597);
xnor UO_1777 (O_1777,N_14418,N_14354);
xnor UO_1778 (O_1778,N_14539,N_14510);
nand UO_1779 (O_1779,N_14627,N_14760);
and UO_1780 (O_1780,N_14397,N_14268);
and UO_1781 (O_1781,N_14634,N_14569);
xnor UO_1782 (O_1782,N_14894,N_14309);
nand UO_1783 (O_1783,N_14690,N_14751);
and UO_1784 (O_1784,N_14903,N_14758);
nand UO_1785 (O_1785,N_14840,N_14374);
nor UO_1786 (O_1786,N_14434,N_14267);
or UO_1787 (O_1787,N_14997,N_14708);
xnor UO_1788 (O_1788,N_14816,N_14917);
nand UO_1789 (O_1789,N_14638,N_14430);
xor UO_1790 (O_1790,N_14534,N_14965);
or UO_1791 (O_1791,N_14512,N_14337);
xnor UO_1792 (O_1792,N_14535,N_14608);
nand UO_1793 (O_1793,N_14933,N_14854);
and UO_1794 (O_1794,N_14371,N_14287);
nand UO_1795 (O_1795,N_14591,N_14995);
xnor UO_1796 (O_1796,N_14388,N_14494);
or UO_1797 (O_1797,N_14597,N_14809);
and UO_1798 (O_1798,N_14733,N_14991);
and UO_1799 (O_1799,N_14981,N_14363);
nor UO_1800 (O_1800,N_14837,N_14278);
nand UO_1801 (O_1801,N_14486,N_14858);
nand UO_1802 (O_1802,N_14862,N_14521);
nand UO_1803 (O_1803,N_14849,N_14762);
xor UO_1804 (O_1804,N_14952,N_14458);
and UO_1805 (O_1805,N_14778,N_14901);
or UO_1806 (O_1806,N_14802,N_14513);
or UO_1807 (O_1807,N_14457,N_14304);
nand UO_1808 (O_1808,N_14751,N_14397);
nor UO_1809 (O_1809,N_14617,N_14957);
xor UO_1810 (O_1810,N_14959,N_14310);
and UO_1811 (O_1811,N_14584,N_14836);
xor UO_1812 (O_1812,N_14695,N_14610);
xnor UO_1813 (O_1813,N_14387,N_14959);
and UO_1814 (O_1814,N_14675,N_14483);
or UO_1815 (O_1815,N_14856,N_14293);
xnor UO_1816 (O_1816,N_14436,N_14742);
and UO_1817 (O_1817,N_14397,N_14502);
and UO_1818 (O_1818,N_14552,N_14743);
or UO_1819 (O_1819,N_14725,N_14520);
nor UO_1820 (O_1820,N_14470,N_14843);
and UO_1821 (O_1821,N_14840,N_14790);
and UO_1822 (O_1822,N_14646,N_14467);
or UO_1823 (O_1823,N_14264,N_14724);
or UO_1824 (O_1824,N_14525,N_14744);
and UO_1825 (O_1825,N_14817,N_14603);
nand UO_1826 (O_1826,N_14717,N_14646);
and UO_1827 (O_1827,N_14411,N_14703);
xor UO_1828 (O_1828,N_14774,N_14356);
nor UO_1829 (O_1829,N_14269,N_14345);
xor UO_1830 (O_1830,N_14551,N_14683);
or UO_1831 (O_1831,N_14359,N_14813);
or UO_1832 (O_1832,N_14506,N_14622);
or UO_1833 (O_1833,N_14941,N_14926);
xor UO_1834 (O_1834,N_14631,N_14591);
nor UO_1835 (O_1835,N_14527,N_14812);
nand UO_1836 (O_1836,N_14461,N_14703);
nor UO_1837 (O_1837,N_14800,N_14686);
or UO_1838 (O_1838,N_14277,N_14739);
xor UO_1839 (O_1839,N_14524,N_14982);
nand UO_1840 (O_1840,N_14451,N_14286);
and UO_1841 (O_1841,N_14472,N_14925);
or UO_1842 (O_1842,N_14890,N_14299);
or UO_1843 (O_1843,N_14383,N_14771);
xnor UO_1844 (O_1844,N_14523,N_14428);
and UO_1845 (O_1845,N_14476,N_14444);
and UO_1846 (O_1846,N_14679,N_14746);
or UO_1847 (O_1847,N_14921,N_14609);
nor UO_1848 (O_1848,N_14403,N_14579);
xor UO_1849 (O_1849,N_14639,N_14401);
nor UO_1850 (O_1850,N_14728,N_14399);
and UO_1851 (O_1851,N_14564,N_14557);
or UO_1852 (O_1852,N_14845,N_14530);
or UO_1853 (O_1853,N_14828,N_14884);
xor UO_1854 (O_1854,N_14282,N_14789);
xor UO_1855 (O_1855,N_14930,N_14252);
or UO_1856 (O_1856,N_14661,N_14309);
or UO_1857 (O_1857,N_14622,N_14318);
or UO_1858 (O_1858,N_14839,N_14909);
or UO_1859 (O_1859,N_14340,N_14373);
or UO_1860 (O_1860,N_14355,N_14782);
and UO_1861 (O_1861,N_14891,N_14585);
nor UO_1862 (O_1862,N_14321,N_14616);
xnor UO_1863 (O_1863,N_14732,N_14660);
nor UO_1864 (O_1864,N_14998,N_14420);
nor UO_1865 (O_1865,N_14835,N_14915);
xnor UO_1866 (O_1866,N_14526,N_14340);
and UO_1867 (O_1867,N_14560,N_14550);
or UO_1868 (O_1868,N_14458,N_14853);
nand UO_1869 (O_1869,N_14889,N_14727);
xor UO_1870 (O_1870,N_14648,N_14265);
nor UO_1871 (O_1871,N_14564,N_14628);
nor UO_1872 (O_1872,N_14930,N_14645);
and UO_1873 (O_1873,N_14288,N_14388);
nor UO_1874 (O_1874,N_14630,N_14655);
xor UO_1875 (O_1875,N_14462,N_14788);
nand UO_1876 (O_1876,N_14780,N_14897);
and UO_1877 (O_1877,N_14729,N_14914);
nor UO_1878 (O_1878,N_14828,N_14456);
or UO_1879 (O_1879,N_14691,N_14629);
nand UO_1880 (O_1880,N_14976,N_14361);
or UO_1881 (O_1881,N_14388,N_14939);
nand UO_1882 (O_1882,N_14866,N_14473);
xor UO_1883 (O_1883,N_14988,N_14278);
nor UO_1884 (O_1884,N_14759,N_14282);
or UO_1885 (O_1885,N_14705,N_14638);
xnor UO_1886 (O_1886,N_14646,N_14929);
and UO_1887 (O_1887,N_14665,N_14705);
xor UO_1888 (O_1888,N_14822,N_14281);
xor UO_1889 (O_1889,N_14572,N_14501);
xnor UO_1890 (O_1890,N_14873,N_14268);
nand UO_1891 (O_1891,N_14835,N_14885);
or UO_1892 (O_1892,N_14512,N_14854);
nor UO_1893 (O_1893,N_14478,N_14466);
nor UO_1894 (O_1894,N_14660,N_14798);
and UO_1895 (O_1895,N_14399,N_14948);
and UO_1896 (O_1896,N_14984,N_14487);
or UO_1897 (O_1897,N_14933,N_14348);
or UO_1898 (O_1898,N_14475,N_14659);
nor UO_1899 (O_1899,N_14431,N_14697);
nor UO_1900 (O_1900,N_14640,N_14474);
nand UO_1901 (O_1901,N_14303,N_14481);
or UO_1902 (O_1902,N_14835,N_14783);
xor UO_1903 (O_1903,N_14931,N_14710);
and UO_1904 (O_1904,N_14796,N_14895);
nor UO_1905 (O_1905,N_14778,N_14341);
nand UO_1906 (O_1906,N_14341,N_14518);
nand UO_1907 (O_1907,N_14477,N_14901);
and UO_1908 (O_1908,N_14864,N_14456);
xnor UO_1909 (O_1909,N_14816,N_14697);
or UO_1910 (O_1910,N_14651,N_14935);
nand UO_1911 (O_1911,N_14515,N_14290);
nor UO_1912 (O_1912,N_14870,N_14880);
and UO_1913 (O_1913,N_14455,N_14914);
or UO_1914 (O_1914,N_14937,N_14508);
and UO_1915 (O_1915,N_14861,N_14757);
nor UO_1916 (O_1916,N_14894,N_14924);
nand UO_1917 (O_1917,N_14496,N_14428);
xor UO_1918 (O_1918,N_14725,N_14938);
nand UO_1919 (O_1919,N_14871,N_14980);
xnor UO_1920 (O_1920,N_14280,N_14559);
and UO_1921 (O_1921,N_14676,N_14608);
xnor UO_1922 (O_1922,N_14825,N_14910);
or UO_1923 (O_1923,N_14669,N_14899);
or UO_1924 (O_1924,N_14617,N_14505);
nor UO_1925 (O_1925,N_14764,N_14610);
nor UO_1926 (O_1926,N_14278,N_14644);
nor UO_1927 (O_1927,N_14911,N_14603);
and UO_1928 (O_1928,N_14395,N_14554);
nor UO_1929 (O_1929,N_14768,N_14484);
xnor UO_1930 (O_1930,N_14645,N_14480);
and UO_1931 (O_1931,N_14597,N_14761);
and UO_1932 (O_1932,N_14504,N_14831);
and UO_1933 (O_1933,N_14912,N_14348);
nand UO_1934 (O_1934,N_14420,N_14900);
xor UO_1935 (O_1935,N_14761,N_14530);
or UO_1936 (O_1936,N_14392,N_14315);
or UO_1937 (O_1937,N_14263,N_14305);
xor UO_1938 (O_1938,N_14984,N_14848);
nand UO_1939 (O_1939,N_14903,N_14679);
nand UO_1940 (O_1940,N_14786,N_14483);
xnor UO_1941 (O_1941,N_14516,N_14517);
and UO_1942 (O_1942,N_14438,N_14499);
xnor UO_1943 (O_1943,N_14774,N_14433);
nand UO_1944 (O_1944,N_14502,N_14481);
xor UO_1945 (O_1945,N_14804,N_14485);
and UO_1946 (O_1946,N_14852,N_14417);
or UO_1947 (O_1947,N_14909,N_14753);
nor UO_1948 (O_1948,N_14867,N_14614);
or UO_1949 (O_1949,N_14925,N_14361);
xnor UO_1950 (O_1950,N_14498,N_14990);
or UO_1951 (O_1951,N_14720,N_14960);
nor UO_1952 (O_1952,N_14896,N_14535);
and UO_1953 (O_1953,N_14936,N_14906);
and UO_1954 (O_1954,N_14539,N_14978);
nor UO_1955 (O_1955,N_14456,N_14265);
nand UO_1956 (O_1956,N_14581,N_14575);
nor UO_1957 (O_1957,N_14497,N_14917);
and UO_1958 (O_1958,N_14353,N_14692);
nor UO_1959 (O_1959,N_14433,N_14642);
xnor UO_1960 (O_1960,N_14802,N_14514);
nand UO_1961 (O_1961,N_14748,N_14872);
nand UO_1962 (O_1962,N_14834,N_14952);
and UO_1963 (O_1963,N_14459,N_14537);
or UO_1964 (O_1964,N_14629,N_14377);
xor UO_1965 (O_1965,N_14927,N_14737);
nor UO_1966 (O_1966,N_14843,N_14500);
xor UO_1967 (O_1967,N_14253,N_14760);
nand UO_1968 (O_1968,N_14311,N_14691);
or UO_1969 (O_1969,N_14835,N_14268);
nor UO_1970 (O_1970,N_14844,N_14561);
nor UO_1971 (O_1971,N_14686,N_14758);
nand UO_1972 (O_1972,N_14383,N_14892);
xnor UO_1973 (O_1973,N_14275,N_14476);
or UO_1974 (O_1974,N_14823,N_14728);
nor UO_1975 (O_1975,N_14391,N_14359);
nand UO_1976 (O_1976,N_14460,N_14595);
or UO_1977 (O_1977,N_14898,N_14945);
or UO_1978 (O_1978,N_14573,N_14628);
or UO_1979 (O_1979,N_14788,N_14350);
nand UO_1980 (O_1980,N_14317,N_14372);
nand UO_1981 (O_1981,N_14916,N_14813);
xor UO_1982 (O_1982,N_14886,N_14491);
nand UO_1983 (O_1983,N_14729,N_14582);
and UO_1984 (O_1984,N_14304,N_14276);
nand UO_1985 (O_1985,N_14533,N_14342);
xnor UO_1986 (O_1986,N_14748,N_14414);
nand UO_1987 (O_1987,N_14758,N_14956);
or UO_1988 (O_1988,N_14752,N_14289);
nand UO_1989 (O_1989,N_14865,N_14678);
nand UO_1990 (O_1990,N_14525,N_14978);
and UO_1991 (O_1991,N_14512,N_14450);
or UO_1992 (O_1992,N_14894,N_14254);
nand UO_1993 (O_1993,N_14548,N_14315);
nand UO_1994 (O_1994,N_14541,N_14880);
xor UO_1995 (O_1995,N_14642,N_14746);
nor UO_1996 (O_1996,N_14361,N_14469);
and UO_1997 (O_1997,N_14583,N_14522);
or UO_1998 (O_1998,N_14274,N_14811);
nand UO_1999 (O_1999,N_14548,N_14872);
endmodule