module basic_1000_10000_1500_20_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_205,In_495);
nor U1 (N_1,In_441,In_869);
nand U2 (N_2,In_927,In_85);
and U3 (N_3,In_176,In_337);
and U4 (N_4,In_803,In_500);
or U5 (N_5,In_108,In_276);
or U6 (N_6,In_533,In_664);
or U7 (N_7,In_261,In_364);
nand U8 (N_8,In_314,In_751);
nor U9 (N_9,In_582,In_581);
and U10 (N_10,In_335,In_850);
nand U11 (N_11,In_826,In_901);
xor U12 (N_12,In_838,In_550);
and U13 (N_13,In_687,In_657);
xnor U14 (N_14,In_759,In_374);
and U15 (N_15,In_969,In_580);
nor U16 (N_16,In_267,In_216);
nor U17 (N_17,In_942,In_941);
nand U18 (N_18,In_928,In_917);
nand U19 (N_19,In_483,In_493);
or U20 (N_20,In_697,In_924);
nand U21 (N_21,In_312,In_332);
or U22 (N_22,In_933,In_719);
xnor U23 (N_23,In_457,In_251);
xor U24 (N_24,In_490,In_561);
nor U25 (N_25,In_865,In_682);
or U26 (N_26,In_883,In_227);
or U27 (N_27,In_867,In_782);
nor U28 (N_28,In_275,In_674);
and U29 (N_29,In_943,In_834);
and U30 (N_30,In_553,In_793);
or U31 (N_31,In_497,In_667);
nor U32 (N_32,In_963,In_385);
nor U33 (N_33,In_857,In_406);
nor U34 (N_34,In_158,In_926);
and U35 (N_35,In_136,In_295);
xor U36 (N_36,In_821,In_117);
or U37 (N_37,In_703,In_583);
and U38 (N_38,In_436,In_240);
xnor U39 (N_39,In_134,In_1);
nor U40 (N_40,In_822,In_661);
nand U41 (N_41,In_115,In_98);
xnor U42 (N_42,In_617,In_895);
or U43 (N_43,In_445,In_338);
nand U44 (N_44,In_146,In_74);
or U45 (N_45,In_952,In_496);
or U46 (N_46,In_831,In_579);
or U47 (N_47,In_846,In_481);
or U48 (N_48,In_325,In_945);
nor U49 (N_49,In_989,In_570);
or U50 (N_50,In_363,In_26);
xnor U51 (N_51,In_587,In_959);
or U52 (N_52,In_451,In_344);
nor U53 (N_53,In_265,In_705);
nor U54 (N_54,In_139,In_182);
nand U55 (N_55,In_534,In_415);
xor U56 (N_56,In_77,In_257);
nor U57 (N_57,In_112,In_619);
and U58 (N_58,In_828,In_426);
xor U59 (N_59,In_516,In_286);
nor U60 (N_60,In_489,In_913);
nand U61 (N_61,In_998,In_418);
and U62 (N_62,In_485,In_27);
or U63 (N_63,In_966,In_238);
or U64 (N_64,In_129,In_671);
nand U65 (N_65,In_137,In_646);
or U66 (N_66,In_212,In_175);
and U67 (N_67,In_37,In_863);
nor U68 (N_68,In_815,In_892);
xor U69 (N_69,In_551,In_890);
nand U70 (N_70,In_605,In_44);
xnor U71 (N_71,In_925,In_342);
xor U72 (N_72,In_488,In_28);
and U73 (N_73,In_362,In_764);
xnor U74 (N_74,In_233,In_844);
xor U75 (N_75,In_35,In_403);
nand U76 (N_76,In_186,In_565);
xnor U77 (N_77,In_856,In_676);
xnor U78 (N_78,In_101,In_306);
xnor U79 (N_79,In_210,In_401);
or U80 (N_80,In_15,In_552);
and U81 (N_81,In_820,In_904);
xnor U82 (N_82,In_128,In_615);
nor U83 (N_83,In_673,In_556);
nand U84 (N_84,In_243,In_593);
and U85 (N_85,In_547,In_596);
xnor U86 (N_86,In_150,In_590);
and U87 (N_87,In_313,In_263);
and U88 (N_88,In_383,In_49);
or U89 (N_89,In_694,In_521);
nor U90 (N_90,In_100,In_684);
and U91 (N_91,In_473,In_635);
nor U92 (N_92,In_690,In_519);
and U93 (N_93,In_854,In_459);
xnor U94 (N_94,In_626,In_909);
and U95 (N_95,In_991,In_310);
nor U96 (N_96,In_650,In_638);
or U97 (N_97,In_272,In_382);
and U98 (N_98,In_894,In_125);
nand U99 (N_99,In_994,In_370);
nor U100 (N_100,In_499,In_555);
nand U101 (N_101,In_754,In_36);
or U102 (N_102,In_598,In_858);
or U103 (N_103,In_118,In_178);
nor U104 (N_104,In_948,In_223);
xnor U105 (N_105,In_911,In_824);
and U106 (N_106,In_962,In_506);
xor U107 (N_107,In_217,In_806);
nand U108 (N_108,In_123,In_404);
nor U109 (N_109,In_111,In_900);
and U110 (N_110,In_498,In_620);
nand U111 (N_111,In_207,In_92);
nand U112 (N_112,In_64,In_466);
xor U113 (N_113,In_277,In_899);
nor U114 (N_114,In_405,In_59);
and U115 (N_115,In_375,In_818);
xor U116 (N_116,In_870,In_264);
and U117 (N_117,In_234,In_780);
nand U118 (N_118,In_573,In_938);
nor U119 (N_119,In_634,In_842);
or U120 (N_120,In_975,In_0);
or U121 (N_121,In_808,In_778);
nor U122 (N_122,In_503,In_199);
or U123 (N_123,In_138,In_285);
and U124 (N_124,In_987,In_774);
nor U125 (N_125,In_679,In_878);
and U126 (N_126,In_66,In_731);
xnor U127 (N_127,In_392,In_612);
or U128 (N_128,In_181,In_226);
and U129 (N_129,In_305,In_96);
nand U130 (N_130,In_607,In_680);
nor U131 (N_131,In_662,In_931);
xor U132 (N_132,In_361,In_843);
xor U133 (N_133,In_688,In_34);
nor U134 (N_134,In_651,In_877);
nor U135 (N_135,In_318,In_311);
or U136 (N_136,In_777,In_514);
or U137 (N_137,In_916,In_20);
or U138 (N_138,In_773,In_696);
nand U139 (N_139,In_980,In_906);
or U140 (N_140,In_287,In_429);
nor U141 (N_141,In_558,In_54);
xor U142 (N_142,In_756,In_781);
xor U143 (N_143,In_745,In_654);
nand U144 (N_144,In_208,In_341);
nor U145 (N_145,In_542,In_154);
nand U146 (N_146,In_474,In_354);
nor U147 (N_147,In_185,In_527);
and U148 (N_148,In_475,In_653);
xor U149 (N_149,In_188,In_470);
nor U150 (N_150,In_455,In_25);
nand U151 (N_151,In_611,In_725);
and U152 (N_152,In_730,In_113);
or U153 (N_153,In_12,In_203);
nor U154 (N_154,In_359,In_577);
and U155 (N_155,In_187,In_666);
nor U156 (N_156,In_701,In_672);
nor U157 (N_157,In_446,In_790);
xor U158 (N_158,In_538,In_127);
nand U159 (N_159,In_640,In_560);
nor U160 (N_160,In_559,In_507);
nand U161 (N_161,In_576,In_548);
or U162 (N_162,In_65,In_645);
xor U163 (N_163,In_410,In_698);
nand U164 (N_164,In_961,In_55);
xor U165 (N_165,In_174,In_215);
and U166 (N_166,In_126,In_367);
nor U167 (N_167,In_431,In_592);
or U168 (N_168,In_61,In_949);
xnor U169 (N_169,In_353,In_135);
nor U170 (N_170,In_740,In_494);
nand U171 (N_171,In_202,In_152);
nor U172 (N_172,In_695,In_861);
nand U173 (N_173,In_245,In_308);
nand U174 (N_174,In_144,In_586);
xor U175 (N_175,In_523,In_183);
nand U176 (N_176,In_141,In_380);
or U177 (N_177,In_201,In_124);
xor U178 (N_178,In_32,In_486);
nor U179 (N_179,In_702,In_440);
xor U180 (N_180,In_38,In_737);
and U181 (N_181,In_990,In_813);
xnor U182 (N_182,In_315,In_706);
or U183 (N_183,In_224,In_785);
or U184 (N_184,In_588,In_81);
nor U185 (N_185,In_394,In_866);
and U186 (N_186,In_231,In_369);
and U187 (N_187,In_452,In_11);
nor U188 (N_188,In_422,In_454);
nor U189 (N_189,In_816,In_602);
nand U190 (N_190,In_63,In_148);
or U191 (N_191,In_478,In_316);
xor U192 (N_192,In_840,In_841);
or U193 (N_193,In_169,In_402);
nand U194 (N_194,In_232,In_629);
xor U195 (N_195,In_322,In_438);
xor U196 (N_196,In_919,In_220);
or U197 (N_197,In_562,In_746);
nor U198 (N_198,In_734,In_755);
xor U199 (N_199,In_214,In_256);
nor U200 (N_200,In_235,In_735);
xor U201 (N_201,In_196,In_145);
nand U202 (N_202,In_563,In_116);
and U203 (N_203,In_419,In_366);
nand U204 (N_204,In_625,In_918);
xnor U205 (N_205,In_253,In_509);
or U206 (N_206,In_979,In_472);
nor U207 (N_207,In_512,In_347);
nor U208 (N_208,In_397,In_198);
xnor U209 (N_209,In_896,In_633);
xnor U210 (N_210,In_923,In_847);
or U211 (N_211,In_434,In_86);
nand U212 (N_212,In_43,In_655);
nor U213 (N_213,In_167,In_53);
and U214 (N_214,In_423,In_761);
or U215 (N_215,In_520,In_995);
nor U216 (N_216,In_304,In_326);
nor U217 (N_217,In_665,In_627);
nor U218 (N_218,In_594,In_432);
and U219 (N_219,In_31,In_798);
nor U220 (N_220,In_950,In_302);
nand U221 (N_221,In_330,In_750);
nor U222 (N_222,In_689,In_329);
xor U223 (N_223,In_898,In_51);
nor U224 (N_224,In_502,In_853);
or U225 (N_225,In_744,In_881);
and U226 (N_226,In_225,In_518);
and U227 (N_227,In_46,In_190);
nor U228 (N_228,In_545,In_307);
and U229 (N_229,In_606,In_106);
and U230 (N_230,In_464,In_334);
nand U231 (N_231,In_531,In_864);
nand U232 (N_232,In_835,In_168);
or U233 (N_233,In_642,In_915);
xnor U234 (N_234,In_340,In_951);
and U235 (N_235,In_639,In_376);
nand U236 (N_236,In_525,In_78);
nor U237 (N_237,In_298,In_427);
or U238 (N_238,In_571,In_250);
nand U239 (N_239,In_75,In_24);
nor U240 (N_240,In_537,In_271);
nand U241 (N_241,In_317,In_350);
xor U242 (N_242,In_663,In_789);
or U243 (N_243,In_155,In_609);
or U244 (N_244,In_707,In_549);
xor U245 (N_245,In_411,In_783);
or U246 (N_246,In_536,In_184);
and U247 (N_247,In_300,In_603);
nor U248 (N_248,In_160,In_328);
xnor U249 (N_249,In_76,In_814);
xor U250 (N_250,In_297,In_442);
nand U251 (N_251,In_544,In_630);
xor U252 (N_252,In_324,In_871);
xor U253 (N_253,In_652,In_218);
nand U254 (N_254,In_41,In_56);
nand U255 (N_255,In_487,In_618);
or U256 (N_256,In_616,In_830);
or U257 (N_257,In_902,In_433);
nor U258 (N_258,In_22,In_880);
or U259 (N_259,In_749,In_14);
and U260 (N_260,In_191,In_400);
xnor U261 (N_261,In_58,In_600);
and U262 (N_262,In_491,In_412);
xnor U263 (N_263,In_424,In_296);
nor U264 (N_264,In_739,In_303);
nand U265 (N_265,In_517,In_274);
xnor U266 (N_266,In_159,In_767);
or U267 (N_267,In_805,In_289);
nand U268 (N_268,In_40,In_102);
or U269 (N_269,In_732,In_794);
xnor U270 (N_270,In_244,In_281);
and U271 (N_271,In_5,In_956);
nor U272 (N_272,In_832,In_396);
nand U273 (N_273,In_399,In_930);
nor U274 (N_274,In_430,In_988);
nand U275 (N_275,In_492,In_60);
or U276 (N_276,In_566,In_458);
or U277 (N_277,In_122,In_823);
nand U278 (N_278,In_910,In_29);
nor U279 (N_279,In_775,In_110);
or U280 (N_280,In_278,In_88);
or U281 (N_281,In_413,In_685);
or U282 (N_282,In_985,In_83);
xor U283 (N_283,In_786,In_885);
nor U284 (N_284,In_48,In_389);
and U285 (N_285,In_797,In_284);
nor U286 (N_286,In_16,In_428);
or U287 (N_287,In_784,In_368);
and U288 (N_288,In_944,In_252);
xnor U289 (N_289,In_254,In_482);
and U290 (N_290,In_839,In_709);
nand U291 (N_291,In_408,In_192);
xnor U292 (N_292,In_393,In_779);
xor U293 (N_293,In_355,In_120);
and U294 (N_294,In_437,In_365);
xor U295 (N_295,In_69,In_868);
xor U296 (N_296,In_165,In_180);
nand U297 (N_297,In_505,In_572);
nand U298 (N_298,In_804,In_921);
nand U299 (N_299,In_940,In_425);
or U300 (N_300,In_84,In_997);
nand U301 (N_301,In_628,In_741);
xnor U302 (N_302,In_678,In_977);
nand U303 (N_303,In_456,In_301);
and U304 (N_304,In_541,In_331);
xnor U305 (N_305,In_768,In_345);
nor U306 (N_306,In_965,In_280);
nand U307 (N_307,In_132,In_70);
nor U308 (N_308,In_597,In_578);
nor U309 (N_309,In_692,In_170);
nor U310 (N_310,In_273,In_39);
and U311 (N_311,In_920,In_554);
and U312 (N_312,In_677,In_260);
nand U313 (N_313,In_333,In_753);
xor U314 (N_314,In_613,In_656);
nor U315 (N_315,In_193,In_282);
or U316 (N_316,In_197,In_460);
xnor U317 (N_317,In_151,In_972);
nand U318 (N_318,In_670,In_23);
xnor U319 (N_319,In_971,In_763);
nor U320 (N_320,In_812,In_801);
or U321 (N_321,In_131,In_601);
nand U322 (N_322,In_97,In_89);
and U323 (N_323,In_584,In_978);
nand U324 (N_324,In_153,In_686);
or U325 (N_325,In_851,In_540);
xor U326 (N_326,In_339,In_748);
nor U327 (N_327,In_147,In_172);
or U328 (N_328,In_937,In_10);
xnor U329 (N_329,In_323,In_907);
nor U330 (N_330,In_872,In_947);
or U331 (N_331,In_968,In_957);
nand U332 (N_332,In_3,In_758);
and U333 (N_333,In_348,In_378);
or U334 (N_334,In_173,In_209);
nand U335 (N_335,In_564,In_683);
and U336 (N_336,In_62,In_42);
nand U337 (N_337,In_388,In_811);
nand U338 (N_338,In_999,In_912);
or U339 (N_339,In_752,In_4);
or U340 (N_340,In_621,In_727);
or U341 (N_341,In_246,In_258);
nand U342 (N_342,In_321,In_237);
nor U343 (N_343,In_177,In_336);
nand U344 (N_344,In_421,In_2);
nor U345 (N_345,In_343,In_9);
nor U346 (N_346,In_879,In_776);
xnor U347 (N_347,In_772,In_644);
and U348 (N_348,In_142,In_713);
xor U349 (N_349,In_882,In_932);
xor U350 (N_350,In_13,In_704);
nand U351 (N_351,In_827,In_953);
nand U352 (N_352,In_130,In_888);
or U353 (N_353,In_259,In_194);
xor U354 (N_354,In_30,In_595);
nand U355 (N_355,In_795,In_221);
nand U356 (N_356,In_973,In_860);
and U357 (N_357,In_515,In_381);
xnor U358 (N_358,In_710,In_939);
xor U359 (N_359,In_668,In_420);
and U360 (N_360,In_269,In_760);
and U361 (N_361,In_510,In_79);
xnor U362 (N_362,In_463,In_200);
or U363 (N_363,In_395,In_819);
nor U364 (N_364,In_967,In_164);
xnor U365 (N_365,In_765,In_99);
and U366 (N_366,In_249,In_862);
or U367 (N_367,In_810,In_787);
xnor U368 (N_368,In_743,In_290);
xor U369 (N_369,In_723,In_501);
nor U370 (N_370,In_50,In_247);
and U371 (N_371,In_960,In_7);
and U372 (N_372,In_319,In_792);
and U373 (N_373,In_357,In_873);
xnor U374 (N_374,In_714,In_80);
nor U375 (N_375,In_157,In_104);
nand U376 (N_376,In_239,In_72);
and U377 (N_377,In_637,In_649);
and U378 (N_378,In_929,In_799);
or U379 (N_379,In_255,In_121);
xor U380 (N_380,In_480,In_386);
xnor U381 (N_381,In_817,In_539);
xor U382 (N_382,In_372,In_283);
or U383 (N_383,In_309,In_114);
and U384 (N_384,In_299,In_675);
or U385 (N_385,In_384,In_461);
nor U386 (N_386,In_802,In_522);
xor U387 (N_387,In_407,In_471);
nand U388 (N_388,In_398,In_631);
or U389 (N_389,In_721,In_736);
or U390 (N_390,In_379,In_807);
and U391 (N_391,In_585,In_693);
nand U392 (N_392,In_149,In_935);
nor U393 (N_393,In_632,In_508);
nor U394 (N_394,In_992,In_358);
nand U395 (N_395,In_204,In_195);
and U396 (N_396,In_156,In_477);
and U397 (N_397,In_884,In_19);
xor U398 (N_398,In_268,In_771);
nor U399 (N_399,In_546,In_45);
xor U400 (N_400,In_848,In_722);
nor U401 (N_401,In_465,In_691);
xor U402 (N_402,In_416,In_453);
xor U403 (N_403,In_73,In_213);
nor U404 (N_404,In_107,In_574);
nor U405 (N_405,In_293,In_94);
and U406 (N_406,In_762,In_161);
or U407 (N_407,In_874,In_417);
nand U408 (N_408,In_179,In_903);
and U409 (N_409,In_886,In_17);
xnor U410 (N_410,In_8,In_377);
or U411 (N_411,In_922,In_766);
xor U412 (N_412,In_229,In_288);
xnor U413 (N_413,In_33,In_449);
and U414 (N_414,In_993,In_716);
and U415 (N_415,In_57,In_140);
nor U416 (N_416,In_206,In_95);
nand U417 (N_417,In_717,In_467);
nor U418 (N_418,In_532,In_720);
xnor U419 (N_419,In_981,In_958);
or U420 (N_420,In_356,In_614);
nor U421 (N_421,In_849,In_568);
nand U422 (N_422,In_189,In_528);
nand U423 (N_423,In_511,In_728);
nand U424 (N_424,In_349,In_769);
nor U425 (N_425,In_591,In_791);
nand U426 (N_426,In_976,In_530);
xnor U427 (N_427,In_715,In_875);
and U428 (N_428,In_543,In_435);
nor U429 (N_429,In_575,In_242);
xor U430 (N_430,In_796,In_462);
xor U431 (N_431,In_891,In_636);
xnor U432 (N_432,In_733,In_236);
and U433 (N_433,In_954,In_119);
or U434 (N_434,In_712,In_946);
or U435 (N_435,In_162,In_166);
nand U436 (N_436,In_373,In_230);
xnor U437 (N_437,In_529,In_788);
or U438 (N_438,In_82,In_908);
xnor U439 (N_439,In_660,In_569);
xor U440 (N_440,In_171,In_825);
or U441 (N_441,In_833,In_143);
and U442 (N_442,In_18,In_726);
and U443 (N_443,In_444,In_647);
nor U444 (N_444,In_729,In_852);
or U445 (N_445,In_67,In_387);
nand U446 (N_446,In_718,In_699);
xor U447 (N_447,In_450,In_262);
or U448 (N_448,In_266,In_608);
nand U449 (N_449,In_700,In_836);
nand U450 (N_450,In_648,In_681);
nor U451 (N_451,In_294,In_504);
nand U452 (N_452,In_469,In_447);
or U453 (N_453,In_983,In_90);
nand U454 (N_454,In_934,In_996);
or U455 (N_455,In_241,In_974);
or U456 (N_456,In_448,In_986);
xor U457 (N_457,In_711,In_622);
and U458 (N_458,In_513,In_982);
nand U459 (N_459,In_439,In_6);
nand U460 (N_460,In_800,In_708);
xor U461 (N_461,In_970,In_624);
nor U462 (N_462,In_360,In_222);
xnor U463 (N_463,In_557,In_109);
xnor U464 (N_464,In_936,In_484);
or U465 (N_465,In_747,In_279);
nor U466 (N_466,In_589,In_914);
and U467 (N_467,In_897,In_889);
xnor U468 (N_468,In_610,In_659);
and U469 (N_469,In_52,In_837);
or U470 (N_470,In_658,In_567);
xor U471 (N_471,In_443,In_219);
nand U472 (N_472,In_845,In_248);
xor U473 (N_473,In_905,In_829);
and U474 (N_474,In_526,In_391);
or U475 (N_475,In_351,In_346);
nand U476 (N_476,In_103,In_599);
nand U477 (N_477,In_211,In_163);
nand U478 (N_478,In_91,In_320);
and U479 (N_479,In_292,In_105);
and U480 (N_480,In_893,In_93);
xor U481 (N_481,In_955,In_414);
nand U482 (N_482,In_327,In_641);
and U483 (N_483,In_291,In_71);
nand U484 (N_484,In_887,In_724);
and U485 (N_485,In_524,In_535);
xnor U486 (N_486,In_738,In_371);
or U487 (N_487,In_409,In_479);
and U488 (N_488,In_859,In_476);
and U489 (N_489,In_21,In_964);
nand U490 (N_490,In_390,In_87);
or U491 (N_491,In_770,In_47);
xor U492 (N_492,In_468,In_855);
xnor U493 (N_493,In_984,In_757);
nand U494 (N_494,In_133,In_669);
or U495 (N_495,In_809,In_623);
nor U496 (N_496,In_643,In_604);
nor U497 (N_497,In_876,In_228);
nor U498 (N_498,In_742,In_352);
xnor U499 (N_499,In_270,In_68);
or U500 (N_500,N_245,N_66);
xor U501 (N_501,N_251,N_133);
nand U502 (N_502,N_486,N_303);
xor U503 (N_503,N_54,N_269);
nand U504 (N_504,N_74,N_171);
or U505 (N_505,N_292,N_489);
nand U506 (N_506,N_44,N_99);
or U507 (N_507,N_126,N_69);
xor U508 (N_508,N_5,N_268);
xnor U509 (N_509,N_234,N_252);
nor U510 (N_510,N_409,N_202);
or U511 (N_511,N_160,N_471);
nand U512 (N_512,N_33,N_186);
and U513 (N_513,N_161,N_85);
and U514 (N_514,N_187,N_240);
nor U515 (N_515,N_106,N_24);
xor U516 (N_516,N_265,N_395);
nor U517 (N_517,N_495,N_207);
nand U518 (N_518,N_346,N_79);
nand U519 (N_519,N_182,N_375);
or U520 (N_520,N_144,N_151);
xnor U521 (N_521,N_104,N_12);
and U522 (N_522,N_464,N_345);
and U523 (N_523,N_243,N_478);
xnor U524 (N_524,N_181,N_390);
and U525 (N_525,N_82,N_192);
and U526 (N_526,N_100,N_23);
and U527 (N_527,N_429,N_97);
and U528 (N_528,N_93,N_333);
xor U529 (N_529,N_98,N_154);
or U530 (N_530,N_75,N_122);
or U531 (N_531,N_418,N_255);
and U532 (N_532,N_212,N_287);
and U533 (N_533,N_308,N_6);
nor U534 (N_534,N_419,N_490);
and U535 (N_535,N_31,N_311);
nor U536 (N_536,N_452,N_455);
nor U537 (N_537,N_153,N_258);
or U538 (N_538,N_432,N_280);
nor U539 (N_539,N_189,N_147);
nor U540 (N_540,N_408,N_394);
xnor U541 (N_541,N_124,N_468);
nand U542 (N_542,N_421,N_237);
or U543 (N_543,N_244,N_101);
nand U544 (N_544,N_89,N_474);
and U545 (N_545,N_112,N_371);
and U546 (N_546,N_137,N_127);
xnor U547 (N_547,N_325,N_461);
or U548 (N_548,N_22,N_224);
and U549 (N_549,N_37,N_87);
nor U550 (N_550,N_57,N_376);
and U551 (N_551,N_56,N_11);
and U552 (N_552,N_315,N_434);
and U553 (N_553,N_16,N_266);
xor U554 (N_554,N_407,N_253);
xor U555 (N_555,N_323,N_289);
or U556 (N_556,N_304,N_329);
or U557 (N_557,N_374,N_383);
or U558 (N_558,N_364,N_215);
and U559 (N_559,N_380,N_361);
nand U560 (N_560,N_425,N_290);
and U561 (N_561,N_115,N_246);
or U562 (N_562,N_43,N_48);
or U563 (N_563,N_177,N_134);
nand U564 (N_564,N_131,N_439);
nand U565 (N_565,N_456,N_278);
and U566 (N_566,N_46,N_389);
xor U567 (N_567,N_232,N_453);
nand U568 (N_568,N_95,N_299);
or U569 (N_569,N_263,N_366);
nand U570 (N_570,N_367,N_309);
nor U571 (N_571,N_164,N_358);
nand U572 (N_572,N_88,N_494);
xnor U573 (N_573,N_277,N_359);
or U574 (N_574,N_451,N_113);
nor U575 (N_575,N_118,N_200);
nor U576 (N_576,N_350,N_229);
xnor U577 (N_577,N_422,N_39);
nand U578 (N_578,N_260,N_7);
and U579 (N_579,N_59,N_430);
or U580 (N_580,N_170,N_19);
xor U581 (N_581,N_174,N_352);
and U582 (N_582,N_3,N_261);
or U583 (N_583,N_228,N_403);
nand U584 (N_584,N_208,N_335);
nor U585 (N_585,N_445,N_271);
nor U586 (N_586,N_140,N_167);
nand U587 (N_587,N_349,N_80);
nand U588 (N_588,N_462,N_166);
nand U589 (N_589,N_198,N_138);
xnor U590 (N_590,N_188,N_438);
xnor U591 (N_591,N_457,N_338);
and U592 (N_592,N_77,N_114);
and U593 (N_593,N_402,N_178);
and U594 (N_594,N_285,N_496);
or U595 (N_595,N_373,N_307);
nand U596 (N_596,N_326,N_128);
or U597 (N_597,N_267,N_443);
nand U598 (N_598,N_372,N_317);
xnor U599 (N_599,N_479,N_110);
and U600 (N_600,N_397,N_141);
or U601 (N_601,N_35,N_417);
xnor U602 (N_602,N_256,N_204);
and U603 (N_603,N_180,N_165);
nor U604 (N_604,N_40,N_410);
nand U605 (N_605,N_201,N_26);
or U606 (N_606,N_428,N_353);
nand U607 (N_607,N_41,N_109);
and U608 (N_608,N_241,N_288);
xnor U609 (N_609,N_274,N_211);
nand U610 (N_610,N_442,N_413);
or U611 (N_611,N_139,N_210);
and U612 (N_612,N_169,N_159);
xor U613 (N_613,N_90,N_68);
nor U614 (N_614,N_319,N_18);
xor U615 (N_615,N_357,N_467);
xor U616 (N_616,N_230,N_52);
nand U617 (N_617,N_103,N_196);
and U618 (N_618,N_415,N_9);
and U619 (N_619,N_91,N_385);
and U620 (N_620,N_143,N_78);
nand U621 (N_621,N_21,N_94);
nor U622 (N_622,N_34,N_199);
nor U623 (N_623,N_404,N_472);
or U624 (N_624,N_4,N_286);
nor U625 (N_625,N_83,N_195);
or U626 (N_626,N_440,N_347);
xnor U627 (N_627,N_136,N_145);
or U628 (N_628,N_108,N_480);
nand U629 (N_629,N_470,N_30);
nand U630 (N_630,N_488,N_156);
xor U631 (N_631,N_339,N_497);
or U632 (N_632,N_296,N_8);
nand U633 (N_633,N_365,N_123);
or U634 (N_634,N_433,N_132);
nor U635 (N_635,N_86,N_291);
xor U636 (N_636,N_70,N_61);
nand U637 (N_637,N_426,N_42);
nand U638 (N_638,N_194,N_142);
nand U639 (N_639,N_391,N_236);
nand U640 (N_640,N_324,N_485);
nor U641 (N_641,N_0,N_185);
and U642 (N_642,N_119,N_222);
or U643 (N_643,N_424,N_1);
nor U644 (N_644,N_351,N_301);
nand U645 (N_645,N_454,N_247);
or U646 (N_646,N_259,N_491);
xnor U647 (N_647,N_469,N_328);
and U648 (N_648,N_36,N_206);
or U649 (N_649,N_47,N_257);
and U650 (N_650,N_431,N_477);
xnor U651 (N_651,N_125,N_302);
xnor U652 (N_652,N_65,N_388);
and U653 (N_653,N_423,N_449);
or U654 (N_654,N_314,N_155);
or U655 (N_655,N_105,N_393);
nor U656 (N_656,N_334,N_370);
nor U657 (N_657,N_310,N_158);
xnor U658 (N_658,N_416,N_356);
and U659 (N_659,N_76,N_221);
xnor U660 (N_660,N_487,N_226);
nand U661 (N_661,N_28,N_193);
or U662 (N_662,N_384,N_216);
and U663 (N_663,N_62,N_387);
xnor U664 (N_664,N_498,N_120);
or U665 (N_665,N_107,N_64);
or U666 (N_666,N_217,N_168);
xnor U667 (N_667,N_405,N_297);
or U668 (N_668,N_293,N_60);
or U669 (N_669,N_282,N_446);
or U670 (N_670,N_318,N_316);
and U671 (N_671,N_45,N_360);
nand U672 (N_672,N_332,N_458);
or U673 (N_673,N_175,N_157);
nor U674 (N_674,N_72,N_499);
or U675 (N_675,N_197,N_129);
nand U676 (N_676,N_313,N_20);
or U677 (N_677,N_148,N_460);
and U678 (N_678,N_203,N_225);
xor U679 (N_679,N_205,N_343);
or U680 (N_680,N_398,N_50);
nand U681 (N_681,N_220,N_27);
and U682 (N_682,N_162,N_320);
or U683 (N_683,N_71,N_401);
nor U684 (N_684,N_493,N_436);
xnor U685 (N_685,N_321,N_483);
and U686 (N_686,N_29,N_55);
nor U687 (N_687,N_223,N_213);
nor U688 (N_688,N_32,N_400);
and U689 (N_689,N_172,N_484);
nor U690 (N_690,N_354,N_173);
nor U691 (N_691,N_92,N_58);
nand U692 (N_692,N_84,N_465);
xnor U693 (N_693,N_283,N_306);
and U694 (N_694,N_331,N_342);
nand U695 (N_695,N_294,N_377);
and U696 (N_696,N_295,N_15);
nor U697 (N_697,N_191,N_218);
and U698 (N_698,N_396,N_250);
nand U699 (N_699,N_149,N_176);
or U700 (N_700,N_272,N_279);
xor U701 (N_701,N_146,N_10);
nor U702 (N_702,N_25,N_209);
xor U703 (N_703,N_378,N_281);
and U704 (N_704,N_459,N_284);
nor U705 (N_705,N_233,N_49);
nand U706 (N_706,N_242,N_130);
xnor U707 (N_707,N_441,N_67);
or U708 (N_708,N_184,N_305);
nand U709 (N_709,N_340,N_327);
nor U710 (N_710,N_348,N_447);
or U711 (N_711,N_238,N_235);
or U712 (N_712,N_381,N_53);
or U713 (N_713,N_116,N_249);
or U714 (N_714,N_399,N_163);
xor U715 (N_715,N_337,N_81);
xor U716 (N_716,N_476,N_38);
nand U717 (N_717,N_183,N_190);
nand U718 (N_718,N_102,N_51);
nand U719 (N_719,N_270,N_444);
xnor U720 (N_720,N_111,N_254);
or U721 (N_721,N_341,N_179);
or U722 (N_722,N_448,N_219);
xnor U723 (N_723,N_239,N_369);
xor U724 (N_724,N_355,N_411);
or U725 (N_725,N_248,N_427);
or U726 (N_726,N_276,N_435);
or U727 (N_727,N_273,N_231);
nor U728 (N_728,N_312,N_363);
nor U729 (N_729,N_379,N_437);
or U730 (N_730,N_336,N_482);
xor U731 (N_731,N_150,N_475);
xor U732 (N_732,N_275,N_368);
xnor U733 (N_733,N_214,N_386);
xnor U734 (N_734,N_414,N_450);
or U735 (N_735,N_96,N_463);
and U736 (N_736,N_17,N_481);
nor U737 (N_737,N_420,N_382);
nand U738 (N_738,N_63,N_344);
or U739 (N_739,N_13,N_473);
and U740 (N_740,N_117,N_322);
and U741 (N_741,N_362,N_492);
xor U742 (N_742,N_392,N_300);
nand U743 (N_743,N_135,N_298);
or U744 (N_744,N_152,N_412);
nand U745 (N_745,N_406,N_227);
and U746 (N_746,N_121,N_262);
or U747 (N_747,N_264,N_330);
and U748 (N_748,N_2,N_466);
nand U749 (N_749,N_73,N_14);
xor U750 (N_750,N_41,N_392);
nor U751 (N_751,N_380,N_353);
nand U752 (N_752,N_68,N_151);
nand U753 (N_753,N_293,N_379);
nand U754 (N_754,N_45,N_254);
or U755 (N_755,N_16,N_466);
nor U756 (N_756,N_294,N_135);
or U757 (N_757,N_443,N_450);
and U758 (N_758,N_135,N_76);
nor U759 (N_759,N_49,N_46);
nand U760 (N_760,N_57,N_403);
or U761 (N_761,N_474,N_159);
and U762 (N_762,N_97,N_414);
nor U763 (N_763,N_83,N_241);
or U764 (N_764,N_401,N_249);
nor U765 (N_765,N_355,N_21);
nand U766 (N_766,N_490,N_333);
or U767 (N_767,N_328,N_337);
or U768 (N_768,N_459,N_324);
or U769 (N_769,N_119,N_109);
xnor U770 (N_770,N_288,N_451);
or U771 (N_771,N_36,N_231);
nand U772 (N_772,N_14,N_76);
or U773 (N_773,N_420,N_216);
nand U774 (N_774,N_216,N_138);
xor U775 (N_775,N_271,N_165);
nand U776 (N_776,N_128,N_357);
and U777 (N_777,N_138,N_76);
xor U778 (N_778,N_15,N_242);
and U779 (N_779,N_353,N_340);
or U780 (N_780,N_342,N_426);
nand U781 (N_781,N_153,N_306);
nor U782 (N_782,N_358,N_423);
nand U783 (N_783,N_373,N_321);
and U784 (N_784,N_37,N_72);
or U785 (N_785,N_80,N_60);
or U786 (N_786,N_115,N_96);
nand U787 (N_787,N_417,N_282);
nand U788 (N_788,N_75,N_470);
or U789 (N_789,N_389,N_196);
nand U790 (N_790,N_147,N_363);
or U791 (N_791,N_310,N_115);
or U792 (N_792,N_176,N_266);
and U793 (N_793,N_164,N_36);
xor U794 (N_794,N_177,N_447);
nand U795 (N_795,N_373,N_35);
and U796 (N_796,N_403,N_273);
xor U797 (N_797,N_156,N_205);
or U798 (N_798,N_498,N_164);
or U799 (N_799,N_31,N_173);
or U800 (N_800,N_119,N_291);
nand U801 (N_801,N_158,N_239);
or U802 (N_802,N_216,N_136);
or U803 (N_803,N_192,N_245);
nor U804 (N_804,N_152,N_483);
and U805 (N_805,N_144,N_235);
nand U806 (N_806,N_197,N_432);
nor U807 (N_807,N_61,N_154);
nand U808 (N_808,N_447,N_90);
and U809 (N_809,N_155,N_393);
and U810 (N_810,N_378,N_21);
and U811 (N_811,N_148,N_383);
nand U812 (N_812,N_366,N_184);
nand U813 (N_813,N_42,N_4);
nor U814 (N_814,N_471,N_380);
xnor U815 (N_815,N_300,N_196);
or U816 (N_816,N_4,N_48);
or U817 (N_817,N_405,N_478);
or U818 (N_818,N_158,N_372);
nand U819 (N_819,N_405,N_462);
or U820 (N_820,N_72,N_490);
and U821 (N_821,N_367,N_227);
xnor U822 (N_822,N_386,N_480);
nand U823 (N_823,N_438,N_86);
xor U824 (N_824,N_382,N_368);
xor U825 (N_825,N_35,N_161);
nand U826 (N_826,N_498,N_455);
or U827 (N_827,N_313,N_344);
xor U828 (N_828,N_132,N_237);
and U829 (N_829,N_353,N_442);
xnor U830 (N_830,N_33,N_434);
nand U831 (N_831,N_7,N_352);
nand U832 (N_832,N_8,N_354);
and U833 (N_833,N_74,N_376);
and U834 (N_834,N_249,N_112);
nand U835 (N_835,N_295,N_290);
and U836 (N_836,N_319,N_39);
or U837 (N_837,N_32,N_101);
xor U838 (N_838,N_372,N_387);
or U839 (N_839,N_498,N_101);
nor U840 (N_840,N_73,N_110);
or U841 (N_841,N_450,N_449);
xor U842 (N_842,N_201,N_342);
xor U843 (N_843,N_400,N_334);
nor U844 (N_844,N_17,N_459);
xnor U845 (N_845,N_471,N_75);
nor U846 (N_846,N_431,N_107);
nor U847 (N_847,N_282,N_468);
xor U848 (N_848,N_301,N_185);
xor U849 (N_849,N_298,N_56);
or U850 (N_850,N_176,N_490);
xnor U851 (N_851,N_217,N_318);
or U852 (N_852,N_287,N_414);
and U853 (N_853,N_212,N_374);
and U854 (N_854,N_455,N_407);
nor U855 (N_855,N_137,N_130);
nand U856 (N_856,N_382,N_292);
xnor U857 (N_857,N_486,N_30);
nand U858 (N_858,N_285,N_214);
nor U859 (N_859,N_103,N_83);
nand U860 (N_860,N_239,N_43);
nor U861 (N_861,N_234,N_230);
xnor U862 (N_862,N_389,N_8);
or U863 (N_863,N_246,N_453);
xor U864 (N_864,N_92,N_238);
or U865 (N_865,N_46,N_292);
and U866 (N_866,N_48,N_234);
xor U867 (N_867,N_165,N_186);
and U868 (N_868,N_127,N_375);
or U869 (N_869,N_285,N_156);
nand U870 (N_870,N_16,N_68);
xnor U871 (N_871,N_49,N_38);
or U872 (N_872,N_94,N_87);
xor U873 (N_873,N_112,N_288);
nor U874 (N_874,N_389,N_216);
xnor U875 (N_875,N_420,N_76);
xnor U876 (N_876,N_363,N_9);
and U877 (N_877,N_200,N_279);
nor U878 (N_878,N_111,N_117);
xor U879 (N_879,N_67,N_224);
and U880 (N_880,N_160,N_103);
and U881 (N_881,N_262,N_13);
xnor U882 (N_882,N_375,N_150);
nor U883 (N_883,N_115,N_102);
nand U884 (N_884,N_340,N_149);
and U885 (N_885,N_432,N_95);
and U886 (N_886,N_23,N_18);
or U887 (N_887,N_404,N_310);
nand U888 (N_888,N_354,N_326);
xor U889 (N_889,N_424,N_180);
nor U890 (N_890,N_345,N_88);
and U891 (N_891,N_453,N_39);
nor U892 (N_892,N_426,N_9);
xor U893 (N_893,N_370,N_481);
and U894 (N_894,N_159,N_63);
nand U895 (N_895,N_495,N_244);
nor U896 (N_896,N_281,N_316);
nand U897 (N_897,N_102,N_238);
and U898 (N_898,N_459,N_240);
xor U899 (N_899,N_441,N_41);
xor U900 (N_900,N_365,N_28);
nand U901 (N_901,N_48,N_19);
and U902 (N_902,N_484,N_137);
and U903 (N_903,N_58,N_161);
or U904 (N_904,N_422,N_498);
nand U905 (N_905,N_57,N_274);
nand U906 (N_906,N_141,N_467);
or U907 (N_907,N_209,N_52);
xnor U908 (N_908,N_5,N_82);
nand U909 (N_909,N_484,N_263);
or U910 (N_910,N_36,N_6);
xor U911 (N_911,N_354,N_480);
or U912 (N_912,N_292,N_68);
nand U913 (N_913,N_474,N_411);
nand U914 (N_914,N_318,N_379);
nor U915 (N_915,N_52,N_495);
nand U916 (N_916,N_38,N_245);
or U917 (N_917,N_446,N_68);
nand U918 (N_918,N_92,N_205);
nor U919 (N_919,N_497,N_0);
nand U920 (N_920,N_287,N_350);
and U921 (N_921,N_265,N_419);
nor U922 (N_922,N_171,N_123);
nand U923 (N_923,N_382,N_358);
nor U924 (N_924,N_261,N_233);
or U925 (N_925,N_156,N_453);
xor U926 (N_926,N_140,N_367);
xor U927 (N_927,N_295,N_455);
nand U928 (N_928,N_237,N_82);
or U929 (N_929,N_458,N_498);
and U930 (N_930,N_337,N_1);
xnor U931 (N_931,N_157,N_263);
xnor U932 (N_932,N_238,N_98);
nor U933 (N_933,N_117,N_375);
nor U934 (N_934,N_238,N_413);
xnor U935 (N_935,N_418,N_354);
nand U936 (N_936,N_116,N_13);
or U937 (N_937,N_492,N_276);
xor U938 (N_938,N_55,N_413);
nand U939 (N_939,N_63,N_5);
or U940 (N_940,N_435,N_83);
xnor U941 (N_941,N_318,N_274);
nand U942 (N_942,N_467,N_60);
xnor U943 (N_943,N_90,N_444);
xnor U944 (N_944,N_365,N_440);
nand U945 (N_945,N_312,N_322);
xnor U946 (N_946,N_336,N_226);
nor U947 (N_947,N_349,N_130);
and U948 (N_948,N_39,N_79);
nand U949 (N_949,N_315,N_122);
nand U950 (N_950,N_477,N_74);
xor U951 (N_951,N_367,N_14);
or U952 (N_952,N_392,N_432);
nand U953 (N_953,N_278,N_19);
or U954 (N_954,N_304,N_12);
nand U955 (N_955,N_139,N_494);
or U956 (N_956,N_42,N_237);
or U957 (N_957,N_378,N_61);
and U958 (N_958,N_351,N_366);
and U959 (N_959,N_151,N_8);
nand U960 (N_960,N_450,N_460);
xnor U961 (N_961,N_283,N_460);
and U962 (N_962,N_468,N_108);
nand U963 (N_963,N_92,N_427);
nor U964 (N_964,N_495,N_434);
xnor U965 (N_965,N_362,N_155);
nand U966 (N_966,N_421,N_84);
and U967 (N_967,N_74,N_0);
xor U968 (N_968,N_498,N_416);
nand U969 (N_969,N_119,N_364);
nand U970 (N_970,N_188,N_355);
nand U971 (N_971,N_380,N_240);
nor U972 (N_972,N_411,N_136);
nor U973 (N_973,N_157,N_122);
or U974 (N_974,N_422,N_351);
xnor U975 (N_975,N_142,N_245);
xnor U976 (N_976,N_463,N_209);
nand U977 (N_977,N_349,N_395);
xor U978 (N_978,N_281,N_173);
or U979 (N_979,N_27,N_84);
nand U980 (N_980,N_238,N_251);
or U981 (N_981,N_297,N_258);
nand U982 (N_982,N_65,N_371);
xnor U983 (N_983,N_209,N_83);
or U984 (N_984,N_364,N_70);
nor U985 (N_985,N_489,N_42);
nor U986 (N_986,N_99,N_487);
nand U987 (N_987,N_231,N_285);
nor U988 (N_988,N_83,N_468);
nor U989 (N_989,N_93,N_355);
and U990 (N_990,N_56,N_376);
and U991 (N_991,N_207,N_429);
nor U992 (N_992,N_414,N_390);
or U993 (N_993,N_72,N_468);
and U994 (N_994,N_337,N_259);
xor U995 (N_995,N_30,N_239);
and U996 (N_996,N_54,N_318);
xnor U997 (N_997,N_25,N_177);
xnor U998 (N_998,N_218,N_82);
nor U999 (N_999,N_405,N_195);
xnor U1000 (N_1000,N_859,N_773);
nor U1001 (N_1001,N_753,N_601);
xor U1002 (N_1002,N_841,N_991);
or U1003 (N_1003,N_503,N_634);
xnor U1004 (N_1004,N_555,N_643);
and U1005 (N_1005,N_558,N_963);
nor U1006 (N_1006,N_699,N_548);
or U1007 (N_1007,N_722,N_955);
xnor U1008 (N_1008,N_587,N_563);
nand U1009 (N_1009,N_917,N_671);
or U1010 (N_1010,N_879,N_877);
and U1011 (N_1011,N_874,N_886);
nor U1012 (N_1012,N_669,N_903);
nor U1013 (N_1013,N_956,N_665);
xnor U1014 (N_1014,N_901,N_790);
and U1015 (N_1015,N_633,N_570);
nand U1016 (N_1016,N_964,N_774);
xnor U1017 (N_1017,N_935,N_615);
nor U1018 (N_1018,N_793,N_698);
xor U1019 (N_1019,N_940,N_989);
and U1020 (N_1020,N_529,N_702);
nor U1021 (N_1021,N_816,N_912);
nor U1022 (N_1022,N_937,N_673);
and U1023 (N_1023,N_830,N_664);
xor U1024 (N_1024,N_967,N_779);
or U1025 (N_1025,N_726,N_850);
xor U1026 (N_1026,N_540,N_672);
nand U1027 (N_1027,N_904,N_560);
nand U1028 (N_1028,N_678,N_688);
or U1029 (N_1029,N_791,N_693);
nor U1030 (N_1030,N_647,N_527);
nand U1031 (N_1031,N_957,N_590);
xnor U1032 (N_1032,N_719,N_677);
or U1033 (N_1033,N_938,N_889);
nor U1034 (N_1034,N_523,N_717);
nor U1035 (N_1035,N_605,N_799);
and U1036 (N_1036,N_784,N_724);
nor U1037 (N_1037,N_593,N_819);
or U1038 (N_1038,N_860,N_913);
nand U1039 (N_1039,N_676,N_679);
nor U1040 (N_1040,N_635,N_667);
nor U1041 (N_1041,N_567,N_852);
nand U1042 (N_1042,N_561,N_858);
xnor U1043 (N_1043,N_900,N_620);
and U1044 (N_1044,N_661,N_756);
or U1045 (N_1045,N_574,N_554);
and U1046 (N_1046,N_746,N_832);
and U1047 (N_1047,N_878,N_537);
nand U1048 (N_1048,N_622,N_725);
nor U1049 (N_1049,N_557,N_782);
nor U1050 (N_1050,N_776,N_599);
or U1051 (N_1051,N_847,N_608);
xnor U1052 (N_1052,N_959,N_736);
nand U1053 (N_1053,N_862,N_780);
nand U1054 (N_1054,N_972,N_979);
and U1055 (N_1055,N_546,N_990);
and U1056 (N_1056,N_500,N_777);
and U1057 (N_1057,N_640,N_769);
and U1058 (N_1058,N_604,N_969);
or U1059 (N_1059,N_517,N_807);
or U1060 (N_1060,N_943,N_525);
nor U1061 (N_1061,N_703,N_648);
or U1062 (N_1062,N_742,N_933);
nor U1063 (N_1063,N_508,N_638);
xor U1064 (N_1064,N_873,N_603);
or U1065 (N_1065,N_871,N_797);
nor U1066 (N_1066,N_962,N_765);
nand U1067 (N_1067,N_521,N_583);
nand U1068 (N_1068,N_865,N_729);
nor U1069 (N_1069,N_822,N_727);
nor U1070 (N_1070,N_785,N_761);
or U1071 (N_1071,N_654,N_749);
nand U1072 (N_1072,N_939,N_787);
or U1073 (N_1073,N_515,N_843);
xor U1074 (N_1074,N_663,N_857);
or U1075 (N_1075,N_668,N_636);
or U1076 (N_1076,N_910,N_586);
xnor U1077 (N_1077,N_612,N_792);
and U1078 (N_1078,N_660,N_994);
nand U1079 (N_1079,N_501,N_690);
nor U1080 (N_1080,N_805,N_579);
nor U1081 (N_1081,N_600,N_613);
nor U1082 (N_1082,N_571,N_524);
nor U1083 (N_1083,N_614,N_934);
nand U1084 (N_1084,N_533,N_602);
nand U1085 (N_1085,N_550,N_627);
nor U1086 (N_1086,N_844,N_752);
xnor U1087 (N_1087,N_706,N_650);
nand U1088 (N_1088,N_762,N_783);
xnor U1089 (N_1089,N_915,N_845);
nor U1090 (N_1090,N_885,N_924);
or U1091 (N_1091,N_794,N_788);
nor U1092 (N_1092,N_732,N_733);
and U1093 (N_1093,N_922,N_929);
nor U1094 (N_1094,N_894,N_639);
and U1095 (N_1095,N_998,N_800);
and U1096 (N_1096,N_547,N_584);
xor U1097 (N_1097,N_683,N_629);
nor U1098 (N_1098,N_948,N_754);
or U1099 (N_1099,N_568,N_666);
xnor U1100 (N_1100,N_812,N_597);
xor U1101 (N_1101,N_853,N_839);
nand U1102 (N_1102,N_806,N_867);
nor U1103 (N_1103,N_866,N_653);
nor U1104 (N_1104,N_512,N_897);
xnor U1105 (N_1105,N_905,N_594);
xnor U1106 (N_1106,N_846,N_573);
nor U1107 (N_1107,N_704,N_976);
or U1108 (N_1108,N_528,N_518);
xor U1109 (N_1109,N_809,N_516);
and U1110 (N_1110,N_825,N_811);
or U1111 (N_1111,N_914,N_607);
nand U1112 (N_1112,N_646,N_535);
nand U1113 (N_1113,N_623,N_823);
nor U1114 (N_1114,N_686,N_795);
and U1115 (N_1115,N_649,N_952);
nor U1116 (N_1116,N_510,N_804);
nand U1117 (N_1117,N_735,N_829);
xor U1118 (N_1118,N_684,N_896);
nor U1119 (N_1119,N_714,N_760);
xor U1120 (N_1120,N_697,N_692);
nor U1121 (N_1121,N_960,N_662);
nand U1122 (N_1122,N_808,N_999);
xnor U1123 (N_1123,N_609,N_522);
xor U1124 (N_1124,N_730,N_958);
or U1125 (N_1125,N_595,N_575);
xnor U1126 (N_1126,N_840,N_995);
nor U1127 (N_1127,N_641,N_552);
nor U1128 (N_1128,N_656,N_718);
xor U1129 (N_1129,N_580,N_659);
xnor U1130 (N_1130,N_848,N_739);
or U1131 (N_1131,N_977,N_970);
or U1132 (N_1132,N_961,N_710);
or U1133 (N_1133,N_950,N_982);
and U1134 (N_1134,N_927,N_987);
or U1135 (N_1135,N_941,N_534);
nand U1136 (N_1136,N_842,N_833);
nor U1137 (N_1137,N_888,N_854);
xor U1138 (N_1138,N_916,N_771);
xor U1139 (N_1139,N_655,N_519);
and U1140 (N_1140,N_576,N_838);
or U1141 (N_1141,N_585,N_925);
or U1142 (N_1142,N_531,N_514);
nand U1143 (N_1143,N_954,N_545);
xor U1144 (N_1144,N_930,N_868);
xor U1145 (N_1145,N_626,N_707);
and U1146 (N_1146,N_949,N_831);
nand U1147 (N_1147,N_751,N_750);
and U1148 (N_1148,N_712,N_951);
nor U1149 (N_1149,N_931,N_968);
or U1150 (N_1150,N_978,N_820);
nand U1151 (N_1151,N_919,N_887);
nand U1152 (N_1152,N_700,N_920);
or U1153 (N_1153,N_834,N_836);
xnor U1154 (N_1154,N_544,N_911);
nor U1155 (N_1155,N_705,N_694);
xor U1156 (N_1156,N_876,N_932);
xor U1157 (N_1157,N_711,N_869);
xnor U1158 (N_1158,N_974,N_606);
or U1159 (N_1159,N_723,N_542);
and U1160 (N_1160,N_892,N_658);
xor U1161 (N_1161,N_973,N_588);
nor U1162 (N_1162,N_906,N_965);
or U1163 (N_1163,N_745,N_637);
nand U1164 (N_1164,N_993,N_625);
xor U1165 (N_1165,N_875,N_505);
or U1166 (N_1166,N_996,N_682);
nor U1167 (N_1167,N_872,N_763);
xor U1168 (N_1168,N_882,N_734);
xor U1169 (N_1169,N_992,N_827);
xnor U1170 (N_1170,N_675,N_775);
nand U1171 (N_1171,N_617,N_803);
nor U1172 (N_1172,N_810,N_944);
xnor U1173 (N_1173,N_559,N_755);
xor U1174 (N_1174,N_980,N_591);
xnor U1175 (N_1175,N_926,N_764);
nor U1176 (N_1176,N_526,N_506);
or U1177 (N_1177,N_975,N_908);
or U1178 (N_1178,N_856,N_851);
nor U1179 (N_1179,N_767,N_988);
xnor U1180 (N_1180,N_511,N_578);
nor U1181 (N_1181,N_828,N_946);
and U1182 (N_1182,N_945,N_708);
and U1183 (N_1183,N_680,N_880);
nor U1184 (N_1184,N_881,N_986);
xnor U1185 (N_1185,N_981,N_624);
or U1186 (N_1186,N_824,N_596);
or U1187 (N_1187,N_520,N_566);
xnor U1188 (N_1188,N_772,N_644);
nor U1189 (N_1189,N_928,N_863);
or U1190 (N_1190,N_870,N_918);
or U1191 (N_1191,N_757,N_509);
xnor U1192 (N_1192,N_652,N_691);
nor U1193 (N_1193,N_921,N_738);
nor U1194 (N_1194,N_770,N_689);
xor U1195 (N_1195,N_815,N_695);
nor U1196 (N_1196,N_632,N_781);
or U1197 (N_1197,N_942,N_883);
nand U1198 (N_1198,N_778,N_630);
and U1199 (N_1199,N_923,N_759);
and U1200 (N_1200,N_818,N_985);
or U1201 (N_1201,N_907,N_709);
nor U1202 (N_1202,N_565,N_947);
and U1203 (N_1203,N_616,N_837);
nor U1204 (N_1204,N_551,N_543);
nand U1205 (N_1205,N_628,N_909);
and U1206 (N_1206,N_720,N_539);
nand U1207 (N_1207,N_786,N_572);
nor U1208 (N_1208,N_621,N_541);
nand U1209 (N_1209,N_696,N_670);
xor U1210 (N_1210,N_651,N_610);
or U1211 (N_1211,N_536,N_504);
nand U1212 (N_1212,N_817,N_768);
xnor U1213 (N_1213,N_619,N_891);
or U1214 (N_1214,N_744,N_814);
xor U1215 (N_1215,N_731,N_631);
or U1216 (N_1216,N_741,N_701);
or U1217 (N_1217,N_530,N_645);
or U1218 (N_1218,N_821,N_953);
xnor U1219 (N_1219,N_502,N_743);
or U1220 (N_1220,N_685,N_895);
and U1221 (N_1221,N_674,N_618);
xor U1222 (N_1222,N_716,N_581);
xnor U1223 (N_1223,N_898,N_747);
xnor U1224 (N_1224,N_549,N_532);
nor U1225 (N_1225,N_899,N_864);
nand U1226 (N_1226,N_758,N_721);
nor U1227 (N_1227,N_564,N_589);
xor U1228 (N_1228,N_681,N_893);
or U1229 (N_1229,N_592,N_798);
xor U1230 (N_1230,N_890,N_737);
nand U1231 (N_1231,N_507,N_728);
or U1232 (N_1232,N_556,N_902);
nand U1233 (N_1233,N_687,N_642);
nor U1234 (N_1234,N_611,N_983);
xor U1235 (N_1235,N_796,N_855);
xor U1236 (N_1236,N_748,N_562);
nor U1237 (N_1237,N_598,N_971);
nor U1238 (N_1238,N_936,N_997);
nor U1239 (N_1239,N_861,N_813);
or U1240 (N_1240,N_984,N_740);
nor U1241 (N_1241,N_766,N_577);
xnor U1242 (N_1242,N_966,N_582);
nor U1243 (N_1243,N_657,N_538);
nor U1244 (N_1244,N_884,N_826);
or U1245 (N_1245,N_569,N_802);
nand U1246 (N_1246,N_849,N_835);
and U1247 (N_1247,N_789,N_713);
and U1248 (N_1248,N_801,N_553);
nor U1249 (N_1249,N_715,N_513);
xor U1250 (N_1250,N_759,N_890);
nor U1251 (N_1251,N_651,N_912);
nand U1252 (N_1252,N_543,N_935);
nor U1253 (N_1253,N_807,N_983);
nand U1254 (N_1254,N_772,N_616);
xor U1255 (N_1255,N_530,N_902);
or U1256 (N_1256,N_884,N_521);
nand U1257 (N_1257,N_623,N_938);
or U1258 (N_1258,N_905,N_797);
nor U1259 (N_1259,N_737,N_638);
xor U1260 (N_1260,N_812,N_925);
nor U1261 (N_1261,N_971,N_915);
and U1262 (N_1262,N_722,N_751);
nor U1263 (N_1263,N_742,N_905);
or U1264 (N_1264,N_604,N_926);
xnor U1265 (N_1265,N_990,N_717);
nand U1266 (N_1266,N_587,N_597);
nor U1267 (N_1267,N_586,N_880);
and U1268 (N_1268,N_690,N_859);
or U1269 (N_1269,N_641,N_559);
nor U1270 (N_1270,N_557,N_762);
nor U1271 (N_1271,N_611,N_710);
nor U1272 (N_1272,N_929,N_933);
xor U1273 (N_1273,N_818,N_975);
or U1274 (N_1274,N_631,N_693);
xor U1275 (N_1275,N_837,N_550);
and U1276 (N_1276,N_706,N_771);
xor U1277 (N_1277,N_728,N_919);
nor U1278 (N_1278,N_771,N_669);
and U1279 (N_1279,N_839,N_963);
and U1280 (N_1280,N_786,N_653);
nor U1281 (N_1281,N_630,N_633);
xnor U1282 (N_1282,N_902,N_584);
nand U1283 (N_1283,N_937,N_666);
xnor U1284 (N_1284,N_786,N_837);
and U1285 (N_1285,N_776,N_633);
nor U1286 (N_1286,N_825,N_697);
nor U1287 (N_1287,N_806,N_770);
nor U1288 (N_1288,N_706,N_909);
or U1289 (N_1289,N_621,N_512);
nor U1290 (N_1290,N_742,N_879);
or U1291 (N_1291,N_584,N_608);
or U1292 (N_1292,N_939,N_609);
nand U1293 (N_1293,N_907,N_757);
or U1294 (N_1294,N_663,N_782);
xor U1295 (N_1295,N_706,N_828);
nor U1296 (N_1296,N_687,N_784);
xnor U1297 (N_1297,N_798,N_948);
or U1298 (N_1298,N_612,N_900);
nor U1299 (N_1299,N_741,N_867);
nor U1300 (N_1300,N_852,N_929);
and U1301 (N_1301,N_743,N_848);
nand U1302 (N_1302,N_851,N_967);
nand U1303 (N_1303,N_708,N_676);
xnor U1304 (N_1304,N_814,N_918);
xor U1305 (N_1305,N_996,N_680);
nor U1306 (N_1306,N_991,N_518);
xor U1307 (N_1307,N_766,N_987);
or U1308 (N_1308,N_736,N_838);
or U1309 (N_1309,N_980,N_641);
nand U1310 (N_1310,N_989,N_799);
xor U1311 (N_1311,N_531,N_840);
and U1312 (N_1312,N_577,N_993);
nor U1313 (N_1313,N_520,N_688);
and U1314 (N_1314,N_988,N_537);
and U1315 (N_1315,N_976,N_655);
xor U1316 (N_1316,N_717,N_669);
and U1317 (N_1317,N_905,N_785);
or U1318 (N_1318,N_613,N_913);
nor U1319 (N_1319,N_926,N_921);
or U1320 (N_1320,N_930,N_646);
nand U1321 (N_1321,N_579,N_751);
nand U1322 (N_1322,N_831,N_663);
nor U1323 (N_1323,N_610,N_765);
nand U1324 (N_1324,N_626,N_695);
or U1325 (N_1325,N_698,N_610);
nand U1326 (N_1326,N_645,N_876);
xor U1327 (N_1327,N_622,N_518);
nor U1328 (N_1328,N_804,N_742);
xor U1329 (N_1329,N_614,N_829);
and U1330 (N_1330,N_561,N_884);
nand U1331 (N_1331,N_836,N_970);
or U1332 (N_1332,N_831,N_572);
nand U1333 (N_1333,N_500,N_654);
or U1334 (N_1334,N_743,N_823);
nor U1335 (N_1335,N_773,N_979);
nand U1336 (N_1336,N_709,N_854);
nor U1337 (N_1337,N_696,N_506);
nand U1338 (N_1338,N_701,N_791);
and U1339 (N_1339,N_770,N_921);
or U1340 (N_1340,N_815,N_789);
xnor U1341 (N_1341,N_644,N_806);
nand U1342 (N_1342,N_601,N_644);
nor U1343 (N_1343,N_858,N_898);
nor U1344 (N_1344,N_519,N_738);
or U1345 (N_1345,N_678,N_958);
nor U1346 (N_1346,N_984,N_544);
xnor U1347 (N_1347,N_758,N_995);
xnor U1348 (N_1348,N_700,N_620);
xnor U1349 (N_1349,N_767,N_641);
xnor U1350 (N_1350,N_809,N_883);
nand U1351 (N_1351,N_524,N_718);
and U1352 (N_1352,N_743,N_969);
nor U1353 (N_1353,N_832,N_763);
and U1354 (N_1354,N_956,N_900);
xnor U1355 (N_1355,N_528,N_668);
or U1356 (N_1356,N_845,N_659);
or U1357 (N_1357,N_925,N_553);
nand U1358 (N_1358,N_688,N_604);
xnor U1359 (N_1359,N_969,N_718);
xnor U1360 (N_1360,N_864,N_546);
and U1361 (N_1361,N_712,N_943);
nor U1362 (N_1362,N_730,N_712);
and U1363 (N_1363,N_615,N_605);
nor U1364 (N_1364,N_984,N_942);
and U1365 (N_1365,N_778,N_670);
xnor U1366 (N_1366,N_892,N_581);
xnor U1367 (N_1367,N_607,N_663);
and U1368 (N_1368,N_786,N_542);
nor U1369 (N_1369,N_888,N_709);
and U1370 (N_1370,N_886,N_818);
and U1371 (N_1371,N_555,N_973);
and U1372 (N_1372,N_996,N_803);
xor U1373 (N_1373,N_740,N_795);
or U1374 (N_1374,N_608,N_579);
or U1375 (N_1375,N_638,N_642);
nand U1376 (N_1376,N_940,N_993);
nor U1377 (N_1377,N_503,N_988);
or U1378 (N_1378,N_792,N_862);
xnor U1379 (N_1379,N_860,N_959);
or U1380 (N_1380,N_640,N_908);
or U1381 (N_1381,N_540,N_808);
or U1382 (N_1382,N_638,N_527);
or U1383 (N_1383,N_930,N_797);
and U1384 (N_1384,N_841,N_549);
or U1385 (N_1385,N_593,N_598);
and U1386 (N_1386,N_595,N_594);
nand U1387 (N_1387,N_828,N_511);
nor U1388 (N_1388,N_854,N_770);
and U1389 (N_1389,N_691,N_589);
nand U1390 (N_1390,N_702,N_652);
nor U1391 (N_1391,N_835,N_986);
or U1392 (N_1392,N_777,N_888);
nor U1393 (N_1393,N_504,N_929);
nand U1394 (N_1394,N_719,N_553);
and U1395 (N_1395,N_580,N_728);
and U1396 (N_1396,N_858,N_743);
nand U1397 (N_1397,N_879,N_792);
nor U1398 (N_1398,N_849,N_888);
nor U1399 (N_1399,N_597,N_534);
nand U1400 (N_1400,N_972,N_753);
and U1401 (N_1401,N_566,N_771);
and U1402 (N_1402,N_565,N_818);
nand U1403 (N_1403,N_731,N_993);
xor U1404 (N_1404,N_530,N_882);
nand U1405 (N_1405,N_899,N_976);
nor U1406 (N_1406,N_722,N_913);
nor U1407 (N_1407,N_854,N_530);
xor U1408 (N_1408,N_661,N_827);
or U1409 (N_1409,N_630,N_640);
and U1410 (N_1410,N_580,N_958);
nor U1411 (N_1411,N_525,N_871);
xor U1412 (N_1412,N_518,N_556);
nand U1413 (N_1413,N_910,N_776);
nand U1414 (N_1414,N_644,N_627);
and U1415 (N_1415,N_900,N_756);
nand U1416 (N_1416,N_826,N_740);
and U1417 (N_1417,N_829,N_698);
nand U1418 (N_1418,N_593,N_690);
or U1419 (N_1419,N_513,N_719);
nor U1420 (N_1420,N_996,N_653);
or U1421 (N_1421,N_743,N_778);
nand U1422 (N_1422,N_887,N_600);
or U1423 (N_1423,N_842,N_506);
or U1424 (N_1424,N_990,N_789);
or U1425 (N_1425,N_821,N_752);
or U1426 (N_1426,N_966,N_749);
xnor U1427 (N_1427,N_867,N_702);
xor U1428 (N_1428,N_987,N_624);
nand U1429 (N_1429,N_821,N_852);
xnor U1430 (N_1430,N_536,N_640);
nor U1431 (N_1431,N_939,N_597);
and U1432 (N_1432,N_759,N_618);
and U1433 (N_1433,N_743,N_986);
nand U1434 (N_1434,N_771,N_752);
and U1435 (N_1435,N_736,N_847);
or U1436 (N_1436,N_884,N_754);
and U1437 (N_1437,N_781,N_898);
nand U1438 (N_1438,N_550,N_598);
and U1439 (N_1439,N_552,N_691);
xnor U1440 (N_1440,N_969,N_990);
xnor U1441 (N_1441,N_574,N_567);
or U1442 (N_1442,N_663,N_862);
or U1443 (N_1443,N_715,N_514);
nor U1444 (N_1444,N_612,N_877);
nor U1445 (N_1445,N_626,N_659);
xor U1446 (N_1446,N_652,N_848);
and U1447 (N_1447,N_950,N_805);
xnor U1448 (N_1448,N_747,N_859);
xor U1449 (N_1449,N_535,N_757);
xor U1450 (N_1450,N_849,N_996);
nand U1451 (N_1451,N_839,N_791);
nand U1452 (N_1452,N_715,N_879);
or U1453 (N_1453,N_894,N_844);
xnor U1454 (N_1454,N_752,N_976);
xor U1455 (N_1455,N_996,N_535);
or U1456 (N_1456,N_682,N_972);
nor U1457 (N_1457,N_807,N_650);
and U1458 (N_1458,N_948,N_802);
nor U1459 (N_1459,N_966,N_607);
nor U1460 (N_1460,N_819,N_908);
and U1461 (N_1461,N_664,N_686);
or U1462 (N_1462,N_956,N_908);
xor U1463 (N_1463,N_757,N_666);
xor U1464 (N_1464,N_771,N_768);
nand U1465 (N_1465,N_519,N_668);
and U1466 (N_1466,N_590,N_873);
or U1467 (N_1467,N_620,N_670);
or U1468 (N_1468,N_559,N_537);
or U1469 (N_1469,N_601,N_946);
and U1470 (N_1470,N_759,N_684);
or U1471 (N_1471,N_849,N_968);
nor U1472 (N_1472,N_794,N_983);
xnor U1473 (N_1473,N_848,N_853);
nand U1474 (N_1474,N_972,N_969);
nand U1475 (N_1475,N_903,N_723);
nor U1476 (N_1476,N_519,N_773);
nor U1477 (N_1477,N_855,N_951);
xnor U1478 (N_1478,N_879,N_898);
nor U1479 (N_1479,N_668,N_810);
or U1480 (N_1480,N_784,N_534);
xor U1481 (N_1481,N_650,N_925);
or U1482 (N_1482,N_735,N_921);
nand U1483 (N_1483,N_644,N_891);
nand U1484 (N_1484,N_863,N_631);
xnor U1485 (N_1485,N_887,N_597);
or U1486 (N_1486,N_695,N_539);
and U1487 (N_1487,N_985,N_714);
nor U1488 (N_1488,N_804,N_880);
nand U1489 (N_1489,N_787,N_916);
nand U1490 (N_1490,N_700,N_565);
or U1491 (N_1491,N_948,N_858);
nor U1492 (N_1492,N_565,N_885);
and U1493 (N_1493,N_517,N_598);
xor U1494 (N_1494,N_579,N_852);
nor U1495 (N_1495,N_617,N_844);
or U1496 (N_1496,N_670,N_526);
nand U1497 (N_1497,N_920,N_826);
xnor U1498 (N_1498,N_501,N_616);
or U1499 (N_1499,N_994,N_910);
xor U1500 (N_1500,N_1253,N_1365);
nand U1501 (N_1501,N_1068,N_1191);
xnor U1502 (N_1502,N_1203,N_1437);
or U1503 (N_1503,N_1199,N_1492);
or U1504 (N_1504,N_1081,N_1467);
nand U1505 (N_1505,N_1360,N_1497);
xor U1506 (N_1506,N_1217,N_1012);
xnor U1507 (N_1507,N_1063,N_1072);
nor U1508 (N_1508,N_1073,N_1006);
nand U1509 (N_1509,N_1168,N_1115);
or U1510 (N_1510,N_1055,N_1296);
xor U1511 (N_1511,N_1487,N_1196);
or U1512 (N_1512,N_1194,N_1209);
nand U1513 (N_1513,N_1318,N_1268);
xnor U1514 (N_1514,N_1080,N_1300);
and U1515 (N_1515,N_1283,N_1202);
xnor U1516 (N_1516,N_1198,N_1440);
nor U1517 (N_1517,N_1151,N_1161);
nand U1518 (N_1518,N_1120,N_1106);
xnor U1519 (N_1519,N_1478,N_1383);
nand U1520 (N_1520,N_1025,N_1000);
or U1521 (N_1521,N_1001,N_1225);
nor U1522 (N_1522,N_1314,N_1320);
nand U1523 (N_1523,N_1157,N_1014);
or U1524 (N_1524,N_1430,N_1394);
and U1525 (N_1525,N_1469,N_1257);
xnor U1526 (N_1526,N_1102,N_1319);
nor U1527 (N_1527,N_1446,N_1143);
nor U1528 (N_1528,N_1463,N_1295);
xnor U1529 (N_1529,N_1181,N_1219);
xnor U1530 (N_1530,N_1018,N_1003);
xnor U1531 (N_1531,N_1404,N_1036);
nand U1532 (N_1532,N_1121,N_1167);
nor U1533 (N_1533,N_1131,N_1348);
nand U1534 (N_1534,N_1359,N_1379);
nor U1535 (N_1535,N_1122,N_1316);
or U1536 (N_1536,N_1340,N_1256);
or U1537 (N_1537,N_1431,N_1236);
or U1538 (N_1538,N_1491,N_1037);
or U1539 (N_1539,N_1083,N_1206);
or U1540 (N_1540,N_1438,N_1325);
nand U1541 (N_1541,N_1347,N_1481);
nand U1542 (N_1542,N_1103,N_1165);
nand U1543 (N_1543,N_1228,N_1371);
nand U1544 (N_1544,N_1039,N_1263);
and U1545 (N_1545,N_1145,N_1368);
or U1546 (N_1546,N_1062,N_1096);
nor U1547 (N_1547,N_1237,N_1173);
nor U1548 (N_1548,N_1499,N_1141);
and U1549 (N_1549,N_1419,N_1066);
or U1550 (N_1550,N_1375,N_1222);
and U1551 (N_1551,N_1490,N_1462);
xnor U1552 (N_1552,N_1224,N_1200);
or U1553 (N_1553,N_1221,N_1321);
nor U1554 (N_1554,N_1307,N_1303);
nand U1555 (N_1555,N_1390,N_1124);
xor U1556 (N_1556,N_1464,N_1341);
xor U1557 (N_1557,N_1028,N_1337);
nand U1558 (N_1558,N_1232,N_1309);
or U1559 (N_1559,N_1429,N_1479);
nand U1560 (N_1560,N_1048,N_1097);
and U1561 (N_1561,N_1053,N_1470);
or U1562 (N_1562,N_1010,N_1249);
nor U1563 (N_1563,N_1107,N_1288);
nor U1564 (N_1564,N_1433,N_1245);
and U1565 (N_1565,N_1231,N_1241);
nor U1566 (N_1566,N_1212,N_1354);
xnor U1567 (N_1567,N_1136,N_1422);
and U1568 (N_1568,N_1054,N_1411);
xor U1569 (N_1569,N_1474,N_1074);
nand U1570 (N_1570,N_1070,N_1333);
xnor U1571 (N_1571,N_1450,N_1110);
xnor U1572 (N_1572,N_1078,N_1473);
xor U1573 (N_1573,N_1287,N_1235);
nor U1574 (N_1574,N_1112,N_1328);
nor U1575 (N_1575,N_1468,N_1108);
and U1576 (N_1576,N_1133,N_1412);
or U1577 (N_1577,N_1127,N_1410);
or U1578 (N_1578,N_1076,N_1372);
nor U1579 (N_1579,N_1452,N_1331);
or U1580 (N_1580,N_1238,N_1449);
or U1581 (N_1581,N_1436,N_1493);
or U1582 (N_1582,N_1432,N_1482);
and U1583 (N_1583,N_1192,N_1351);
or U1584 (N_1584,N_1104,N_1195);
nand U1585 (N_1585,N_1138,N_1310);
or U1586 (N_1586,N_1471,N_1069);
nand U1587 (N_1587,N_1135,N_1058);
xor U1588 (N_1588,N_1274,N_1414);
xnor U1589 (N_1589,N_1455,N_1038);
nand U1590 (N_1590,N_1182,N_1021);
nor U1591 (N_1591,N_1226,N_1046);
nor U1592 (N_1592,N_1119,N_1329);
or U1593 (N_1593,N_1160,N_1130);
or U1594 (N_1594,N_1376,N_1197);
xnor U1595 (N_1595,N_1162,N_1483);
or U1596 (N_1596,N_1211,N_1453);
or U1597 (N_1597,N_1134,N_1171);
xnor U1598 (N_1598,N_1444,N_1246);
xor U1599 (N_1599,N_1435,N_1460);
or U1600 (N_1600,N_1401,N_1396);
and U1601 (N_1601,N_1304,N_1448);
or U1602 (N_1602,N_1098,N_1045);
nand U1603 (N_1603,N_1011,N_1049);
nor U1604 (N_1604,N_1137,N_1056);
nor U1605 (N_1605,N_1311,N_1207);
or U1606 (N_1606,N_1451,N_1291);
or U1607 (N_1607,N_1034,N_1265);
xnor U1608 (N_1608,N_1132,N_1178);
and U1609 (N_1609,N_1496,N_1352);
and U1610 (N_1610,N_1156,N_1426);
nor U1611 (N_1611,N_1044,N_1125);
nand U1612 (N_1612,N_1233,N_1260);
and U1613 (N_1613,N_1230,N_1113);
nor U1614 (N_1614,N_1082,N_1442);
nand U1615 (N_1615,N_1077,N_1266);
nand U1616 (N_1616,N_1051,N_1094);
or U1617 (N_1617,N_1060,N_1363);
xnor U1618 (N_1618,N_1214,N_1189);
nor U1619 (N_1619,N_1085,N_1087);
and U1620 (N_1620,N_1179,N_1391);
nand U1621 (N_1621,N_1476,N_1382);
nor U1622 (N_1622,N_1275,N_1336);
or U1623 (N_1623,N_1445,N_1421);
nor U1624 (N_1624,N_1008,N_1213);
nand U1625 (N_1625,N_1240,N_1284);
or U1626 (N_1626,N_1064,N_1272);
xnor U1627 (N_1627,N_1163,N_1343);
and U1628 (N_1628,N_1261,N_1408);
or U1629 (N_1629,N_1251,N_1042);
or U1630 (N_1630,N_1282,N_1244);
nor U1631 (N_1631,N_1356,N_1392);
nand U1632 (N_1632,N_1158,N_1279);
and U1633 (N_1633,N_1239,N_1061);
and U1634 (N_1634,N_1201,N_1254);
xor U1635 (N_1635,N_1020,N_1031);
nor U1636 (N_1636,N_1250,N_1378);
or U1637 (N_1637,N_1218,N_1458);
nor U1638 (N_1638,N_1278,N_1465);
nand U1639 (N_1639,N_1308,N_1007);
and U1640 (N_1640,N_1398,N_1126);
nor U1641 (N_1641,N_1367,N_1317);
xnor U1642 (N_1642,N_1457,N_1393);
nor U1643 (N_1643,N_1050,N_1400);
nor U1644 (N_1644,N_1033,N_1153);
or U1645 (N_1645,N_1361,N_1243);
and U1646 (N_1646,N_1397,N_1447);
nor U1647 (N_1647,N_1403,N_1227);
nor U1648 (N_1648,N_1399,N_1323);
nand U1649 (N_1649,N_1079,N_1327);
nor U1650 (N_1650,N_1088,N_1386);
nand U1651 (N_1651,N_1334,N_1150);
and U1652 (N_1652,N_1415,N_1099);
xor U1653 (N_1653,N_1215,N_1186);
xnor U1654 (N_1654,N_1023,N_1017);
or U1655 (N_1655,N_1242,N_1461);
or U1656 (N_1656,N_1180,N_1032);
nor U1657 (N_1657,N_1148,N_1116);
or U1658 (N_1658,N_1117,N_1100);
xnor U1659 (N_1659,N_1128,N_1385);
nor U1660 (N_1660,N_1423,N_1188);
nor U1661 (N_1661,N_1208,N_1067);
and U1662 (N_1662,N_1387,N_1484);
nand U1663 (N_1663,N_1346,N_1312);
xnor U1664 (N_1664,N_1271,N_1377);
xor U1665 (N_1665,N_1280,N_1286);
or U1666 (N_1666,N_1264,N_1417);
nor U1667 (N_1667,N_1357,N_1149);
nor U1668 (N_1668,N_1190,N_1290);
and U1669 (N_1669,N_1485,N_1276);
or U1670 (N_1670,N_1258,N_1090);
or U1671 (N_1671,N_1349,N_1248);
nor U1672 (N_1672,N_1342,N_1140);
or U1673 (N_1673,N_1488,N_1364);
nor U1674 (N_1674,N_1353,N_1252);
or U1675 (N_1675,N_1294,N_1315);
nand U1676 (N_1676,N_1152,N_1184);
or U1677 (N_1677,N_1495,N_1172);
nor U1678 (N_1678,N_1105,N_1216);
and U1679 (N_1679,N_1302,N_1101);
nor U1680 (N_1680,N_1427,N_1456);
nand U1681 (N_1681,N_1166,N_1289);
or U1682 (N_1682,N_1164,N_1029);
nor U1683 (N_1683,N_1022,N_1477);
nor U1684 (N_1684,N_1380,N_1281);
or U1685 (N_1685,N_1373,N_1139);
nand U1686 (N_1686,N_1247,N_1059);
nor U1687 (N_1687,N_1093,N_1299);
and U1688 (N_1688,N_1406,N_1187);
nand U1689 (N_1689,N_1027,N_1052);
or U1690 (N_1690,N_1154,N_1009);
nor U1691 (N_1691,N_1402,N_1019);
or U1692 (N_1692,N_1220,N_1015);
and U1693 (N_1693,N_1144,N_1210);
or U1694 (N_1694,N_1147,N_1277);
nor U1695 (N_1695,N_1142,N_1185);
xnor U1696 (N_1696,N_1409,N_1259);
and U1697 (N_1697,N_1395,N_1075);
or U1698 (N_1698,N_1177,N_1267);
nor U1699 (N_1699,N_1370,N_1002);
xnor U1700 (N_1700,N_1486,N_1285);
nand U1701 (N_1701,N_1350,N_1205);
nand U1702 (N_1702,N_1326,N_1155);
nor U1703 (N_1703,N_1114,N_1109);
nand U1704 (N_1704,N_1338,N_1111);
xnor U1705 (N_1705,N_1358,N_1129);
nor U1706 (N_1706,N_1324,N_1335);
xor U1707 (N_1707,N_1384,N_1204);
or U1708 (N_1708,N_1322,N_1084);
nor U1709 (N_1709,N_1234,N_1193);
nand U1710 (N_1710,N_1418,N_1043);
or U1711 (N_1711,N_1389,N_1273);
and U1712 (N_1712,N_1494,N_1047);
xnor U1713 (N_1713,N_1293,N_1040);
xnor U1714 (N_1714,N_1089,N_1344);
nor U1715 (N_1715,N_1298,N_1086);
nand U1716 (N_1716,N_1441,N_1305);
nor U1717 (N_1717,N_1065,N_1388);
or U1718 (N_1718,N_1475,N_1005);
nand U1719 (N_1719,N_1345,N_1269);
or U1720 (N_1720,N_1374,N_1366);
xnor U1721 (N_1721,N_1013,N_1413);
xor U1722 (N_1722,N_1118,N_1057);
xor U1723 (N_1723,N_1306,N_1159);
and U1724 (N_1724,N_1175,N_1091);
xnor U1725 (N_1725,N_1416,N_1035);
nand U1726 (N_1726,N_1489,N_1439);
or U1727 (N_1727,N_1174,N_1223);
and U1728 (N_1728,N_1407,N_1169);
nor U1729 (N_1729,N_1434,N_1297);
nor U1730 (N_1730,N_1146,N_1498);
xnor U1731 (N_1731,N_1428,N_1292);
xor U1732 (N_1732,N_1092,N_1016);
and U1733 (N_1733,N_1459,N_1024);
and U1734 (N_1734,N_1041,N_1381);
and U1735 (N_1735,N_1355,N_1332);
or U1736 (N_1736,N_1026,N_1369);
or U1737 (N_1737,N_1443,N_1262);
and U1738 (N_1738,N_1095,N_1454);
nor U1739 (N_1739,N_1183,N_1472);
and U1740 (N_1740,N_1176,N_1123);
or U1741 (N_1741,N_1255,N_1480);
and U1742 (N_1742,N_1425,N_1405);
xor U1743 (N_1743,N_1362,N_1339);
xnor U1744 (N_1744,N_1330,N_1313);
and U1745 (N_1745,N_1229,N_1170);
nand U1746 (N_1746,N_1420,N_1270);
nand U1747 (N_1747,N_1466,N_1071);
nand U1748 (N_1748,N_1301,N_1424);
or U1749 (N_1749,N_1004,N_1030);
or U1750 (N_1750,N_1199,N_1461);
and U1751 (N_1751,N_1031,N_1056);
xor U1752 (N_1752,N_1048,N_1462);
and U1753 (N_1753,N_1340,N_1066);
nor U1754 (N_1754,N_1377,N_1049);
and U1755 (N_1755,N_1289,N_1069);
or U1756 (N_1756,N_1432,N_1221);
nor U1757 (N_1757,N_1153,N_1074);
xor U1758 (N_1758,N_1129,N_1231);
nor U1759 (N_1759,N_1119,N_1014);
and U1760 (N_1760,N_1120,N_1227);
and U1761 (N_1761,N_1379,N_1011);
or U1762 (N_1762,N_1064,N_1271);
or U1763 (N_1763,N_1083,N_1319);
nor U1764 (N_1764,N_1388,N_1078);
xor U1765 (N_1765,N_1082,N_1047);
nor U1766 (N_1766,N_1266,N_1476);
xnor U1767 (N_1767,N_1021,N_1237);
xor U1768 (N_1768,N_1471,N_1125);
nand U1769 (N_1769,N_1387,N_1237);
nand U1770 (N_1770,N_1182,N_1143);
nand U1771 (N_1771,N_1397,N_1136);
xor U1772 (N_1772,N_1055,N_1471);
or U1773 (N_1773,N_1463,N_1375);
or U1774 (N_1774,N_1404,N_1324);
and U1775 (N_1775,N_1232,N_1015);
nand U1776 (N_1776,N_1160,N_1073);
or U1777 (N_1777,N_1110,N_1204);
nor U1778 (N_1778,N_1076,N_1492);
xor U1779 (N_1779,N_1034,N_1085);
nand U1780 (N_1780,N_1476,N_1497);
or U1781 (N_1781,N_1299,N_1416);
or U1782 (N_1782,N_1211,N_1143);
nor U1783 (N_1783,N_1473,N_1417);
xor U1784 (N_1784,N_1283,N_1078);
nor U1785 (N_1785,N_1210,N_1023);
nand U1786 (N_1786,N_1414,N_1011);
nor U1787 (N_1787,N_1217,N_1405);
nand U1788 (N_1788,N_1312,N_1011);
and U1789 (N_1789,N_1357,N_1408);
nand U1790 (N_1790,N_1226,N_1027);
nand U1791 (N_1791,N_1287,N_1393);
or U1792 (N_1792,N_1259,N_1146);
nor U1793 (N_1793,N_1075,N_1358);
and U1794 (N_1794,N_1450,N_1314);
xnor U1795 (N_1795,N_1440,N_1315);
nor U1796 (N_1796,N_1469,N_1088);
and U1797 (N_1797,N_1077,N_1378);
nor U1798 (N_1798,N_1476,N_1136);
and U1799 (N_1799,N_1104,N_1040);
xnor U1800 (N_1800,N_1104,N_1459);
xor U1801 (N_1801,N_1107,N_1281);
nand U1802 (N_1802,N_1336,N_1243);
or U1803 (N_1803,N_1001,N_1417);
or U1804 (N_1804,N_1183,N_1062);
or U1805 (N_1805,N_1076,N_1390);
or U1806 (N_1806,N_1392,N_1455);
nor U1807 (N_1807,N_1259,N_1161);
nand U1808 (N_1808,N_1260,N_1050);
and U1809 (N_1809,N_1004,N_1431);
nand U1810 (N_1810,N_1037,N_1028);
xnor U1811 (N_1811,N_1410,N_1388);
nor U1812 (N_1812,N_1246,N_1405);
or U1813 (N_1813,N_1373,N_1133);
and U1814 (N_1814,N_1001,N_1367);
or U1815 (N_1815,N_1373,N_1218);
nor U1816 (N_1816,N_1152,N_1232);
xnor U1817 (N_1817,N_1021,N_1239);
nand U1818 (N_1818,N_1243,N_1177);
nor U1819 (N_1819,N_1380,N_1109);
and U1820 (N_1820,N_1107,N_1356);
and U1821 (N_1821,N_1409,N_1068);
or U1822 (N_1822,N_1402,N_1308);
xnor U1823 (N_1823,N_1343,N_1082);
or U1824 (N_1824,N_1018,N_1111);
nand U1825 (N_1825,N_1009,N_1104);
or U1826 (N_1826,N_1016,N_1036);
nor U1827 (N_1827,N_1464,N_1320);
and U1828 (N_1828,N_1030,N_1340);
xor U1829 (N_1829,N_1069,N_1368);
or U1830 (N_1830,N_1113,N_1442);
or U1831 (N_1831,N_1096,N_1208);
xnor U1832 (N_1832,N_1240,N_1404);
nor U1833 (N_1833,N_1439,N_1006);
xor U1834 (N_1834,N_1246,N_1335);
nand U1835 (N_1835,N_1164,N_1289);
and U1836 (N_1836,N_1107,N_1210);
xor U1837 (N_1837,N_1204,N_1066);
nor U1838 (N_1838,N_1043,N_1133);
nor U1839 (N_1839,N_1206,N_1175);
nor U1840 (N_1840,N_1055,N_1289);
or U1841 (N_1841,N_1451,N_1300);
nand U1842 (N_1842,N_1426,N_1194);
or U1843 (N_1843,N_1177,N_1025);
or U1844 (N_1844,N_1039,N_1303);
and U1845 (N_1845,N_1363,N_1346);
and U1846 (N_1846,N_1042,N_1467);
nand U1847 (N_1847,N_1014,N_1052);
xnor U1848 (N_1848,N_1127,N_1003);
nor U1849 (N_1849,N_1307,N_1245);
nand U1850 (N_1850,N_1151,N_1318);
nand U1851 (N_1851,N_1144,N_1464);
and U1852 (N_1852,N_1429,N_1394);
nand U1853 (N_1853,N_1120,N_1292);
and U1854 (N_1854,N_1433,N_1083);
nand U1855 (N_1855,N_1441,N_1232);
or U1856 (N_1856,N_1475,N_1284);
nand U1857 (N_1857,N_1340,N_1494);
nand U1858 (N_1858,N_1026,N_1011);
nor U1859 (N_1859,N_1348,N_1377);
and U1860 (N_1860,N_1417,N_1002);
and U1861 (N_1861,N_1435,N_1172);
nand U1862 (N_1862,N_1178,N_1148);
xnor U1863 (N_1863,N_1308,N_1077);
nand U1864 (N_1864,N_1214,N_1430);
nand U1865 (N_1865,N_1193,N_1375);
nor U1866 (N_1866,N_1000,N_1130);
nand U1867 (N_1867,N_1092,N_1469);
or U1868 (N_1868,N_1376,N_1073);
nor U1869 (N_1869,N_1117,N_1138);
nor U1870 (N_1870,N_1439,N_1206);
and U1871 (N_1871,N_1177,N_1006);
nor U1872 (N_1872,N_1169,N_1319);
or U1873 (N_1873,N_1197,N_1166);
nor U1874 (N_1874,N_1107,N_1151);
or U1875 (N_1875,N_1349,N_1036);
nand U1876 (N_1876,N_1177,N_1200);
and U1877 (N_1877,N_1188,N_1398);
or U1878 (N_1878,N_1020,N_1002);
and U1879 (N_1879,N_1492,N_1100);
and U1880 (N_1880,N_1341,N_1042);
nand U1881 (N_1881,N_1039,N_1196);
xor U1882 (N_1882,N_1288,N_1480);
and U1883 (N_1883,N_1499,N_1002);
xor U1884 (N_1884,N_1283,N_1088);
nor U1885 (N_1885,N_1411,N_1261);
nand U1886 (N_1886,N_1037,N_1035);
xor U1887 (N_1887,N_1493,N_1151);
nor U1888 (N_1888,N_1340,N_1245);
or U1889 (N_1889,N_1175,N_1438);
or U1890 (N_1890,N_1097,N_1256);
nand U1891 (N_1891,N_1174,N_1283);
or U1892 (N_1892,N_1031,N_1366);
nor U1893 (N_1893,N_1133,N_1361);
and U1894 (N_1894,N_1420,N_1494);
and U1895 (N_1895,N_1497,N_1081);
and U1896 (N_1896,N_1369,N_1470);
or U1897 (N_1897,N_1181,N_1354);
xnor U1898 (N_1898,N_1167,N_1126);
nor U1899 (N_1899,N_1319,N_1433);
or U1900 (N_1900,N_1348,N_1236);
nand U1901 (N_1901,N_1145,N_1242);
xor U1902 (N_1902,N_1215,N_1138);
nand U1903 (N_1903,N_1264,N_1218);
nand U1904 (N_1904,N_1016,N_1048);
and U1905 (N_1905,N_1276,N_1133);
nor U1906 (N_1906,N_1387,N_1005);
nand U1907 (N_1907,N_1197,N_1475);
nor U1908 (N_1908,N_1374,N_1112);
xor U1909 (N_1909,N_1102,N_1208);
nor U1910 (N_1910,N_1248,N_1360);
or U1911 (N_1911,N_1157,N_1266);
xor U1912 (N_1912,N_1440,N_1097);
nand U1913 (N_1913,N_1096,N_1161);
nor U1914 (N_1914,N_1227,N_1452);
or U1915 (N_1915,N_1149,N_1210);
nand U1916 (N_1916,N_1335,N_1243);
xnor U1917 (N_1917,N_1033,N_1440);
and U1918 (N_1918,N_1303,N_1129);
nand U1919 (N_1919,N_1197,N_1249);
nor U1920 (N_1920,N_1432,N_1006);
xnor U1921 (N_1921,N_1319,N_1215);
and U1922 (N_1922,N_1320,N_1027);
nor U1923 (N_1923,N_1424,N_1348);
or U1924 (N_1924,N_1370,N_1294);
nor U1925 (N_1925,N_1032,N_1293);
xnor U1926 (N_1926,N_1322,N_1056);
xnor U1927 (N_1927,N_1410,N_1120);
and U1928 (N_1928,N_1173,N_1464);
or U1929 (N_1929,N_1190,N_1309);
or U1930 (N_1930,N_1443,N_1496);
nor U1931 (N_1931,N_1429,N_1217);
xor U1932 (N_1932,N_1061,N_1440);
and U1933 (N_1933,N_1465,N_1067);
and U1934 (N_1934,N_1294,N_1154);
xnor U1935 (N_1935,N_1060,N_1400);
or U1936 (N_1936,N_1201,N_1446);
and U1937 (N_1937,N_1420,N_1058);
or U1938 (N_1938,N_1208,N_1314);
nand U1939 (N_1939,N_1311,N_1133);
and U1940 (N_1940,N_1188,N_1006);
nand U1941 (N_1941,N_1113,N_1381);
nor U1942 (N_1942,N_1431,N_1076);
and U1943 (N_1943,N_1053,N_1166);
nor U1944 (N_1944,N_1426,N_1355);
nand U1945 (N_1945,N_1362,N_1452);
or U1946 (N_1946,N_1388,N_1356);
nand U1947 (N_1947,N_1116,N_1438);
nand U1948 (N_1948,N_1093,N_1281);
or U1949 (N_1949,N_1390,N_1417);
or U1950 (N_1950,N_1145,N_1191);
nor U1951 (N_1951,N_1407,N_1456);
nand U1952 (N_1952,N_1085,N_1097);
or U1953 (N_1953,N_1047,N_1104);
and U1954 (N_1954,N_1075,N_1424);
xnor U1955 (N_1955,N_1351,N_1167);
xor U1956 (N_1956,N_1352,N_1035);
xnor U1957 (N_1957,N_1314,N_1243);
xnor U1958 (N_1958,N_1332,N_1337);
xor U1959 (N_1959,N_1265,N_1121);
xnor U1960 (N_1960,N_1201,N_1453);
nor U1961 (N_1961,N_1333,N_1145);
xor U1962 (N_1962,N_1464,N_1049);
or U1963 (N_1963,N_1474,N_1292);
and U1964 (N_1964,N_1372,N_1034);
and U1965 (N_1965,N_1100,N_1421);
xor U1966 (N_1966,N_1337,N_1009);
nor U1967 (N_1967,N_1246,N_1421);
or U1968 (N_1968,N_1436,N_1265);
or U1969 (N_1969,N_1099,N_1250);
nand U1970 (N_1970,N_1429,N_1212);
or U1971 (N_1971,N_1203,N_1088);
nor U1972 (N_1972,N_1000,N_1263);
nand U1973 (N_1973,N_1282,N_1380);
nor U1974 (N_1974,N_1280,N_1284);
nand U1975 (N_1975,N_1301,N_1280);
or U1976 (N_1976,N_1354,N_1057);
and U1977 (N_1977,N_1417,N_1150);
and U1978 (N_1978,N_1177,N_1241);
xor U1979 (N_1979,N_1056,N_1089);
nand U1980 (N_1980,N_1287,N_1448);
nand U1981 (N_1981,N_1488,N_1272);
xnor U1982 (N_1982,N_1255,N_1077);
or U1983 (N_1983,N_1073,N_1153);
nor U1984 (N_1984,N_1178,N_1043);
nand U1985 (N_1985,N_1035,N_1430);
xor U1986 (N_1986,N_1199,N_1303);
xnor U1987 (N_1987,N_1167,N_1002);
nand U1988 (N_1988,N_1256,N_1039);
or U1989 (N_1989,N_1172,N_1250);
xor U1990 (N_1990,N_1265,N_1447);
nor U1991 (N_1991,N_1475,N_1350);
xor U1992 (N_1992,N_1171,N_1236);
and U1993 (N_1993,N_1459,N_1108);
nand U1994 (N_1994,N_1132,N_1333);
and U1995 (N_1995,N_1175,N_1087);
nor U1996 (N_1996,N_1456,N_1453);
xor U1997 (N_1997,N_1298,N_1196);
and U1998 (N_1998,N_1487,N_1020);
or U1999 (N_1999,N_1008,N_1302);
nand U2000 (N_2000,N_1746,N_1676);
nand U2001 (N_2001,N_1708,N_1784);
or U2002 (N_2002,N_1909,N_1572);
nand U2003 (N_2003,N_1902,N_1817);
xor U2004 (N_2004,N_1797,N_1921);
xor U2005 (N_2005,N_1924,N_1658);
nand U2006 (N_2006,N_1701,N_1827);
xor U2007 (N_2007,N_1925,N_1699);
or U2008 (N_2008,N_1846,N_1588);
nand U2009 (N_2009,N_1770,N_1918);
xnor U2010 (N_2010,N_1691,N_1564);
xor U2011 (N_2011,N_1887,N_1839);
or U2012 (N_2012,N_1578,N_1737);
or U2013 (N_2013,N_1514,N_1653);
nor U2014 (N_2014,N_1785,N_1888);
nor U2015 (N_2015,N_1634,N_1545);
nand U2016 (N_2016,N_1940,N_1939);
and U2017 (N_2017,N_1961,N_1717);
or U2018 (N_2018,N_1875,N_1582);
nand U2019 (N_2019,N_1745,N_1769);
and U2020 (N_2020,N_1811,N_1816);
or U2021 (N_2021,N_1858,N_1738);
nor U2022 (N_2022,N_1655,N_1501);
and U2023 (N_2023,N_1793,N_1806);
nor U2024 (N_2024,N_1744,N_1788);
xnor U2025 (N_2025,N_1766,N_1830);
nand U2026 (N_2026,N_1725,N_1966);
and U2027 (N_2027,N_1824,N_1599);
or U2028 (N_2028,N_1706,N_1511);
or U2029 (N_2029,N_1563,N_1883);
and U2030 (N_2030,N_1669,N_1739);
and U2031 (N_2031,N_1664,N_1923);
xnor U2032 (N_2032,N_1568,N_1715);
nand U2033 (N_2033,N_1755,N_1507);
and U2034 (N_2034,N_1976,N_1927);
or U2035 (N_2035,N_1565,N_1642);
xnor U2036 (N_2036,N_1714,N_1576);
and U2037 (N_2037,N_1900,N_1767);
nand U2038 (N_2038,N_1533,N_1825);
and U2039 (N_2039,N_1851,N_1876);
nand U2040 (N_2040,N_1865,N_1988);
xor U2041 (N_2041,N_1983,N_1823);
nand U2042 (N_2042,N_1668,N_1581);
nor U2043 (N_2043,N_1525,N_1529);
or U2044 (N_2044,N_1638,N_1585);
or U2045 (N_2045,N_1869,N_1652);
and U2046 (N_2046,N_1898,N_1840);
nand U2047 (N_2047,N_1849,N_1882);
nor U2048 (N_2048,N_1621,N_1947);
nor U2049 (N_2049,N_1504,N_1941);
or U2050 (N_2050,N_1731,N_1712);
or U2051 (N_2051,N_1886,N_1660);
and U2052 (N_2052,N_1553,N_1765);
nand U2053 (N_2053,N_1709,N_1522);
xor U2054 (N_2054,N_1815,N_1975);
nand U2055 (N_2055,N_1508,N_1512);
or U2056 (N_2056,N_1969,N_1573);
nand U2057 (N_2057,N_1982,N_1786);
nor U2058 (N_2058,N_1977,N_1598);
xor U2059 (N_2059,N_1632,N_1594);
and U2060 (N_2060,N_1566,N_1792);
nor U2061 (N_2061,N_1832,N_1555);
nand U2062 (N_2062,N_1778,N_1633);
xnor U2063 (N_2063,N_1985,N_1844);
and U2064 (N_2064,N_1689,N_1607);
xor U2065 (N_2065,N_1644,N_1716);
and U2066 (N_2066,N_1885,N_1570);
nor U2067 (N_2067,N_1949,N_1505);
xnor U2068 (N_2068,N_1757,N_1877);
xnor U2069 (N_2069,N_1680,N_1605);
xor U2070 (N_2070,N_1659,N_1648);
or U2071 (N_2071,N_1650,N_1855);
or U2072 (N_2072,N_1773,N_1749);
and U2073 (N_2073,N_1772,N_1734);
and U2074 (N_2074,N_1908,N_1758);
nand U2075 (N_2075,N_1780,N_1932);
and U2076 (N_2076,N_1556,N_1550);
or U2077 (N_2077,N_1782,N_1736);
nor U2078 (N_2078,N_1881,N_1965);
or U2079 (N_2079,N_1804,N_1960);
and U2080 (N_2080,N_1794,N_1561);
nand U2081 (N_2081,N_1575,N_1847);
nand U2082 (N_2082,N_1623,N_1611);
and U2083 (N_2083,N_1899,N_1674);
and U2084 (N_2084,N_1904,N_1592);
nor U2085 (N_2085,N_1917,N_1748);
and U2086 (N_2086,N_1903,N_1972);
nand U2087 (N_2087,N_1548,N_1723);
nor U2088 (N_2088,N_1532,N_1558);
or U2089 (N_2089,N_1958,N_1584);
and U2090 (N_2090,N_1603,N_1610);
nand U2091 (N_2091,N_1818,N_1656);
xnor U2092 (N_2092,N_1586,N_1795);
nor U2093 (N_2093,N_1953,N_1829);
nand U2094 (N_2094,N_1624,N_1973);
xnor U2095 (N_2095,N_1537,N_1552);
nand U2096 (N_2096,N_1518,N_1579);
nand U2097 (N_2097,N_1628,N_1934);
xor U2098 (N_2098,N_1682,N_1892);
nor U2099 (N_2099,N_1720,N_1856);
nand U2100 (N_2100,N_1919,N_1989);
xnor U2101 (N_2101,N_1936,N_1681);
nor U2102 (N_2102,N_1747,N_1860);
xor U2103 (N_2103,N_1796,N_1781);
and U2104 (N_2104,N_1604,N_1678);
xnor U2105 (N_2105,N_1896,N_1554);
xor U2106 (N_2106,N_1543,N_1742);
or U2107 (N_2107,N_1893,N_1672);
nand U2108 (N_2108,N_1959,N_1713);
nor U2109 (N_2109,N_1547,N_1651);
and U2110 (N_2110,N_1948,N_1928);
or U2111 (N_2111,N_1540,N_1994);
xor U2112 (N_2112,N_1687,N_1873);
or U2113 (N_2113,N_1990,N_1690);
and U2114 (N_2114,N_1527,N_1662);
or U2115 (N_2115,N_1931,N_1724);
or U2116 (N_2116,N_1536,N_1768);
nand U2117 (N_2117,N_1673,N_1759);
xnor U2118 (N_2118,N_1967,N_1852);
and U2119 (N_2119,N_1538,N_1968);
nor U2120 (N_2120,N_1671,N_1719);
or U2121 (N_2121,N_1641,N_1562);
nor U2122 (N_2122,N_1620,N_1663);
and U2123 (N_2123,N_1841,N_1848);
and U2124 (N_2124,N_1718,N_1695);
xnor U2125 (N_2125,N_1774,N_1962);
nor U2126 (N_2126,N_1534,N_1914);
or U2127 (N_2127,N_1801,N_1912);
and U2128 (N_2128,N_1952,N_1812);
or U2129 (N_2129,N_1987,N_1643);
nand U2130 (N_2130,N_1686,N_1986);
and U2131 (N_2131,N_1991,N_1984);
or U2132 (N_2132,N_1995,N_1526);
or U2133 (N_2133,N_1910,N_1577);
and U2134 (N_2134,N_1750,N_1684);
xnor U2135 (N_2135,N_1916,N_1798);
or U2136 (N_2136,N_1626,N_1964);
and U2137 (N_2137,N_1726,N_1835);
xnor U2138 (N_2138,N_1970,N_1971);
xor U2139 (N_2139,N_1542,N_1509);
xnor U2140 (N_2140,N_1814,N_1800);
and U2141 (N_2141,N_1665,N_1837);
nor U2142 (N_2142,N_1933,N_1583);
nand U2143 (N_2143,N_1833,N_1707);
nand U2144 (N_2144,N_1506,N_1728);
or U2145 (N_2145,N_1826,N_1836);
or U2146 (N_2146,N_1627,N_1629);
or U2147 (N_2147,N_1870,N_1697);
or U2148 (N_2148,N_1807,N_1974);
xor U2149 (N_2149,N_1503,N_1649);
or U2150 (N_2150,N_1587,N_1703);
or U2151 (N_2151,N_1890,N_1571);
xnor U2152 (N_2152,N_1612,N_1645);
xnor U2153 (N_2153,N_1515,N_1791);
and U2154 (N_2154,N_1661,N_1636);
nor U2155 (N_2155,N_1838,N_1955);
nor U2156 (N_2156,N_1635,N_1820);
nand U2157 (N_2157,N_1705,N_1569);
nand U2158 (N_2158,N_1609,N_1520);
and U2159 (N_2159,N_1618,N_1999);
and U2160 (N_2160,N_1938,N_1622);
xor U2161 (N_2161,N_1859,N_1613);
xor U2162 (N_2162,N_1615,N_1625);
nor U2163 (N_2163,N_1597,N_1863);
nand U2164 (N_2164,N_1861,N_1915);
xnor U2165 (N_2165,N_1637,N_1677);
or U2166 (N_2166,N_1992,N_1884);
nand U2167 (N_2167,N_1872,N_1698);
xor U2168 (N_2168,N_1614,N_1789);
nor U2169 (N_2169,N_1721,N_1761);
nor U2170 (N_2170,N_1616,N_1907);
and U2171 (N_2171,N_1790,N_1963);
xor U2172 (N_2172,N_1601,N_1930);
nand U2173 (N_2173,N_1667,N_1831);
and U2174 (N_2174,N_1606,N_1843);
nand U2175 (N_2175,N_1654,N_1640);
or U2176 (N_2176,N_1779,N_1946);
nand U2177 (N_2177,N_1819,N_1546);
nor U2178 (N_2178,N_1805,N_1513);
nand U2179 (N_2179,N_1929,N_1600);
nand U2180 (N_2180,N_1523,N_1871);
nor U2181 (N_2181,N_1978,N_1740);
nand U2182 (N_2182,N_1980,N_1531);
xnor U2183 (N_2183,N_1775,N_1741);
nand U2184 (N_2184,N_1935,N_1864);
and U2185 (N_2185,N_1822,N_1889);
or U2186 (N_2186,N_1894,N_1942);
or U2187 (N_2187,N_1981,N_1596);
xor U2188 (N_2188,N_1866,N_1752);
xor U2189 (N_2189,N_1710,N_1679);
and U2190 (N_2190,N_1783,N_1617);
xnor U2191 (N_2191,N_1760,N_1944);
nor U2192 (N_2192,N_1862,N_1593);
xor U2193 (N_2193,N_1702,N_1762);
nand U2194 (N_2194,N_1510,N_1549);
nor U2195 (N_2195,N_1897,N_1901);
nor U2196 (N_2196,N_1521,N_1878);
xnor U2197 (N_2197,N_1693,N_1683);
and U2198 (N_2198,N_1937,N_1891);
nor U2199 (N_2199,N_1590,N_1993);
nand U2200 (N_2200,N_1979,N_1530);
xor U2201 (N_2201,N_1517,N_1813);
nor U2202 (N_2202,N_1945,N_1730);
or U2203 (N_2203,N_1675,N_1560);
nand U2204 (N_2204,N_1591,N_1722);
or U2205 (N_2205,N_1842,N_1828);
nand U2206 (N_2206,N_1764,N_1943);
or U2207 (N_2207,N_1754,N_1519);
nand U2208 (N_2208,N_1853,N_1954);
xnor U2209 (N_2209,N_1895,N_1619);
and U2210 (N_2210,N_1666,N_1763);
nand U2211 (N_2211,N_1574,N_1926);
and U2212 (N_2212,N_1580,N_1704);
and U2213 (N_2213,N_1834,N_1639);
xnor U2214 (N_2214,N_1711,N_1777);
or U2215 (N_2215,N_1729,N_1694);
nand U2216 (N_2216,N_1631,N_1559);
and U2217 (N_2217,N_1700,N_1957);
and U2218 (N_2218,N_1857,N_1913);
and U2219 (N_2219,N_1539,N_1692);
nor U2220 (N_2220,N_1595,N_1500);
nor U2221 (N_2221,N_1911,N_1850);
nand U2222 (N_2222,N_1630,N_1541);
xnor U2223 (N_2223,N_1733,N_1922);
xor U2224 (N_2224,N_1920,N_1799);
nand U2225 (N_2225,N_1776,N_1685);
nand U2226 (N_2226,N_1646,N_1551);
xnor U2227 (N_2227,N_1516,N_1802);
nand U2228 (N_2228,N_1544,N_1803);
nand U2229 (N_2229,N_1854,N_1771);
or U2230 (N_2230,N_1727,N_1753);
nand U2231 (N_2231,N_1567,N_1524);
and U2232 (N_2232,N_1528,N_1997);
and U2233 (N_2233,N_1821,N_1998);
and U2234 (N_2234,N_1845,N_1657);
nand U2235 (N_2235,N_1787,N_1906);
nand U2236 (N_2236,N_1756,N_1951);
nand U2237 (N_2237,N_1735,N_1956);
nand U2238 (N_2238,N_1557,N_1867);
nand U2239 (N_2239,N_1688,N_1502);
or U2240 (N_2240,N_1880,N_1751);
nand U2241 (N_2241,N_1535,N_1647);
nand U2242 (N_2242,N_1670,N_1743);
xor U2243 (N_2243,N_1868,N_1950);
xnor U2244 (N_2244,N_1608,N_1905);
or U2245 (N_2245,N_1589,N_1810);
or U2246 (N_2246,N_1809,N_1879);
xnor U2247 (N_2247,N_1602,N_1808);
or U2248 (N_2248,N_1874,N_1996);
nand U2249 (N_2249,N_1732,N_1696);
nor U2250 (N_2250,N_1959,N_1942);
or U2251 (N_2251,N_1971,N_1541);
nand U2252 (N_2252,N_1523,N_1601);
or U2253 (N_2253,N_1875,N_1825);
or U2254 (N_2254,N_1752,N_1578);
xor U2255 (N_2255,N_1885,N_1622);
and U2256 (N_2256,N_1623,N_1517);
nand U2257 (N_2257,N_1504,N_1935);
or U2258 (N_2258,N_1700,N_1803);
xnor U2259 (N_2259,N_1501,N_1678);
xnor U2260 (N_2260,N_1624,N_1790);
or U2261 (N_2261,N_1880,N_1646);
and U2262 (N_2262,N_1618,N_1933);
xnor U2263 (N_2263,N_1850,N_1603);
nand U2264 (N_2264,N_1636,N_1698);
nand U2265 (N_2265,N_1900,N_1734);
nor U2266 (N_2266,N_1934,N_1880);
nor U2267 (N_2267,N_1753,N_1620);
nand U2268 (N_2268,N_1560,N_1582);
and U2269 (N_2269,N_1737,N_1692);
or U2270 (N_2270,N_1680,N_1946);
xor U2271 (N_2271,N_1988,N_1727);
xor U2272 (N_2272,N_1844,N_1934);
nand U2273 (N_2273,N_1686,N_1922);
xnor U2274 (N_2274,N_1563,N_1937);
nand U2275 (N_2275,N_1657,N_1887);
or U2276 (N_2276,N_1637,N_1993);
or U2277 (N_2277,N_1697,N_1509);
nand U2278 (N_2278,N_1642,N_1755);
xnor U2279 (N_2279,N_1780,N_1573);
or U2280 (N_2280,N_1734,N_1717);
or U2281 (N_2281,N_1748,N_1551);
or U2282 (N_2282,N_1876,N_1937);
nor U2283 (N_2283,N_1718,N_1640);
or U2284 (N_2284,N_1821,N_1635);
nand U2285 (N_2285,N_1865,N_1620);
nand U2286 (N_2286,N_1745,N_1652);
nor U2287 (N_2287,N_1777,N_1703);
nand U2288 (N_2288,N_1725,N_1610);
and U2289 (N_2289,N_1685,N_1640);
nor U2290 (N_2290,N_1689,N_1927);
nand U2291 (N_2291,N_1778,N_1880);
nand U2292 (N_2292,N_1711,N_1793);
and U2293 (N_2293,N_1539,N_1812);
and U2294 (N_2294,N_1575,N_1770);
nor U2295 (N_2295,N_1878,N_1770);
xnor U2296 (N_2296,N_1989,N_1888);
nor U2297 (N_2297,N_1837,N_1636);
nand U2298 (N_2298,N_1595,N_1733);
or U2299 (N_2299,N_1638,N_1751);
nor U2300 (N_2300,N_1618,N_1711);
nor U2301 (N_2301,N_1962,N_1599);
nor U2302 (N_2302,N_1534,N_1632);
xnor U2303 (N_2303,N_1946,N_1578);
nand U2304 (N_2304,N_1953,N_1910);
nand U2305 (N_2305,N_1858,N_1562);
or U2306 (N_2306,N_1911,N_1569);
nand U2307 (N_2307,N_1739,N_1542);
xnor U2308 (N_2308,N_1585,N_1562);
and U2309 (N_2309,N_1701,N_1523);
xnor U2310 (N_2310,N_1537,N_1953);
nand U2311 (N_2311,N_1822,N_1655);
and U2312 (N_2312,N_1884,N_1837);
nor U2313 (N_2313,N_1527,N_1757);
nand U2314 (N_2314,N_1564,N_1993);
or U2315 (N_2315,N_1523,N_1712);
xnor U2316 (N_2316,N_1584,N_1534);
nor U2317 (N_2317,N_1672,N_1602);
and U2318 (N_2318,N_1612,N_1549);
nor U2319 (N_2319,N_1789,N_1610);
and U2320 (N_2320,N_1836,N_1518);
xor U2321 (N_2321,N_1940,N_1852);
xor U2322 (N_2322,N_1933,N_1837);
xnor U2323 (N_2323,N_1610,N_1507);
or U2324 (N_2324,N_1860,N_1674);
xnor U2325 (N_2325,N_1840,N_1663);
nor U2326 (N_2326,N_1863,N_1531);
or U2327 (N_2327,N_1520,N_1894);
and U2328 (N_2328,N_1649,N_1952);
or U2329 (N_2329,N_1551,N_1776);
xor U2330 (N_2330,N_1827,N_1651);
xnor U2331 (N_2331,N_1819,N_1868);
or U2332 (N_2332,N_1967,N_1958);
nor U2333 (N_2333,N_1741,N_1590);
or U2334 (N_2334,N_1843,N_1785);
or U2335 (N_2335,N_1521,N_1586);
and U2336 (N_2336,N_1695,N_1760);
or U2337 (N_2337,N_1583,N_1651);
or U2338 (N_2338,N_1695,N_1750);
nor U2339 (N_2339,N_1602,N_1614);
xor U2340 (N_2340,N_1584,N_1920);
and U2341 (N_2341,N_1592,N_1996);
and U2342 (N_2342,N_1680,N_1696);
nor U2343 (N_2343,N_1731,N_1644);
nand U2344 (N_2344,N_1636,N_1712);
and U2345 (N_2345,N_1620,N_1607);
or U2346 (N_2346,N_1676,N_1895);
and U2347 (N_2347,N_1648,N_1779);
nor U2348 (N_2348,N_1722,N_1661);
nand U2349 (N_2349,N_1740,N_1840);
xor U2350 (N_2350,N_1532,N_1526);
and U2351 (N_2351,N_1553,N_1851);
nand U2352 (N_2352,N_1693,N_1679);
nand U2353 (N_2353,N_1778,N_1799);
or U2354 (N_2354,N_1932,N_1985);
nor U2355 (N_2355,N_1942,N_1714);
and U2356 (N_2356,N_1784,N_1801);
and U2357 (N_2357,N_1988,N_1979);
or U2358 (N_2358,N_1657,N_1753);
nor U2359 (N_2359,N_1697,N_1761);
and U2360 (N_2360,N_1680,N_1937);
xor U2361 (N_2361,N_1512,N_1831);
or U2362 (N_2362,N_1682,N_1582);
or U2363 (N_2363,N_1994,N_1884);
xor U2364 (N_2364,N_1546,N_1960);
xnor U2365 (N_2365,N_1832,N_1784);
nor U2366 (N_2366,N_1546,N_1582);
nand U2367 (N_2367,N_1966,N_1624);
nor U2368 (N_2368,N_1688,N_1739);
xnor U2369 (N_2369,N_1772,N_1547);
nand U2370 (N_2370,N_1606,N_1687);
nor U2371 (N_2371,N_1566,N_1788);
nand U2372 (N_2372,N_1696,N_1827);
and U2373 (N_2373,N_1692,N_1954);
xor U2374 (N_2374,N_1615,N_1850);
nor U2375 (N_2375,N_1996,N_1739);
or U2376 (N_2376,N_1672,N_1836);
nand U2377 (N_2377,N_1626,N_1771);
nand U2378 (N_2378,N_1728,N_1958);
or U2379 (N_2379,N_1730,N_1708);
xnor U2380 (N_2380,N_1891,N_1749);
and U2381 (N_2381,N_1792,N_1597);
nand U2382 (N_2382,N_1689,N_1989);
and U2383 (N_2383,N_1917,N_1654);
nor U2384 (N_2384,N_1664,N_1931);
or U2385 (N_2385,N_1676,N_1520);
xor U2386 (N_2386,N_1696,N_1840);
nor U2387 (N_2387,N_1736,N_1653);
xor U2388 (N_2388,N_1524,N_1758);
xnor U2389 (N_2389,N_1502,N_1574);
or U2390 (N_2390,N_1749,N_1689);
and U2391 (N_2391,N_1802,N_1529);
and U2392 (N_2392,N_1571,N_1994);
xnor U2393 (N_2393,N_1783,N_1682);
nand U2394 (N_2394,N_1838,N_1878);
nand U2395 (N_2395,N_1588,N_1786);
or U2396 (N_2396,N_1981,N_1632);
xnor U2397 (N_2397,N_1741,N_1640);
nand U2398 (N_2398,N_1552,N_1957);
xnor U2399 (N_2399,N_1527,N_1942);
nor U2400 (N_2400,N_1825,N_1859);
nor U2401 (N_2401,N_1661,N_1662);
nor U2402 (N_2402,N_1629,N_1630);
or U2403 (N_2403,N_1985,N_1647);
nor U2404 (N_2404,N_1723,N_1936);
nand U2405 (N_2405,N_1679,N_1786);
nor U2406 (N_2406,N_1764,N_1658);
nand U2407 (N_2407,N_1711,N_1891);
or U2408 (N_2408,N_1963,N_1658);
nand U2409 (N_2409,N_1958,N_1814);
xor U2410 (N_2410,N_1629,N_1718);
or U2411 (N_2411,N_1636,N_1758);
and U2412 (N_2412,N_1681,N_1750);
or U2413 (N_2413,N_1911,N_1515);
xnor U2414 (N_2414,N_1613,N_1741);
nor U2415 (N_2415,N_1766,N_1815);
nor U2416 (N_2416,N_1956,N_1877);
nor U2417 (N_2417,N_1669,N_1755);
xnor U2418 (N_2418,N_1786,N_1874);
or U2419 (N_2419,N_1702,N_1530);
and U2420 (N_2420,N_1832,N_1868);
and U2421 (N_2421,N_1672,N_1645);
nor U2422 (N_2422,N_1654,N_1673);
and U2423 (N_2423,N_1827,N_1513);
nand U2424 (N_2424,N_1559,N_1755);
and U2425 (N_2425,N_1747,N_1995);
xor U2426 (N_2426,N_1963,N_1884);
and U2427 (N_2427,N_1984,N_1553);
and U2428 (N_2428,N_1851,N_1836);
xor U2429 (N_2429,N_1509,N_1692);
and U2430 (N_2430,N_1614,N_1879);
nor U2431 (N_2431,N_1707,N_1943);
xnor U2432 (N_2432,N_1537,N_1868);
and U2433 (N_2433,N_1607,N_1683);
nor U2434 (N_2434,N_1980,N_1659);
nand U2435 (N_2435,N_1587,N_1621);
and U2436 (N_2436,N_1693,N_1913);
or U2437 (N_2437,N_1522,N_1638);
or U2438 (N_2438,N_1921,N_1820);
and U2439 (N_2439,N_1832,N_1880);
xnor U2440 (N_2440,N_1832,N_1872);
and U2441 (N_2441,N_1635,N_1584);
or U2442 (N_2442,N_1643,N_1962);
xnor U2443 (N_2443,N_1791,N_1855);
nor U2444 (N_2444,N_1634,N_1758);
nand U2445 (N_2445,N_1703,N_1537);
nor U2446 (N_2446,N_1756,N_1862);
nand U2447 (N_2447,N_1895,N_1767);
xor U2448 (N_2448,N_1895,N_1772);
or U2449 (N_2449,N_1734,N_1766);
nor U2450 (N_2450,N_1670,N_1720);
and U2451 (N_2451,N_1607,N_1742);
nand U2452 (N_2452,N_1632,N_1743);
and U2453 (N_2453,N_1540,N_1943);
xnor U2454 (N_2454,N_1641,N_1665);
or U2455 (N_2455,N_1822,N_1800);
xor U2456 (N_2456,N_1656,N_1692);
or U2457 (N_2457,N_1673,N_1884);
nor U2458 (N_2458,N_1985,N_1560);
nand U2459 (N_2459,N_1707,N_1727);
or U2460 (N_2460,N_1545,N_1773);
and U2461 (N_2461,N_1575,N_1938);
nand U2462 (N_2462,N_1785,N_1995);
xor U2463 (N_2463,N_1875,N_1532);
nor U2464 (N_2464,N_1735,N_1955);
or U2465 (N_2465,N_1605,N_1726);
or U2466 (N_2466,N_1919,N_1808);
and U2467 (N_2467,N_1602,N_1676);
nor U2468 (N_2468,N_1990,N_1915);
nor U2469 (N_2469,N_1552,N_1909);
xor U2470 (N_2470,N_1985,N_1824);
and U2471 (N_2471,N_1670,N_1813);
and U2472 (N_2472,N_1619,N_1780);
or U2473 (N_2473,N_1550,N_1646);
xnor U2474 (N_2474,N_1818,N_1921);
and U2475 (N_2475,N_1826,N_1574);
xor U2476 (N_2476,N_1525,N_1870);
and U2477 (N_2477,N_1821,N_1527);
nand U2478 (N_2478,N_1840,N_1601);
nor U2479 (N_2479,N_1514,N_1790);
and U2480 (N_2480,N_1711,N_1736);
nand U2481 (N_2481,N_1712,N_1836);
nor U2482 (N_2482,N_1590,N_1651);
nor U2483 (N_2483,N_1861,N_1504);
nor U2484 (N_2484,N_1923,N_1885);
and U2485 (N_2485,N_1980,N_1752);
or U2486 (N_2486,N_1631,N_1580);
and U2487 (N_2487,N_1588,N_1716);
and U2488 (N_2488,N_1911,N_1968);
and U2489 (N_2489,N_1579,N_1546);
nand U2490 (N_2490,N_1998,N_1632);
xor U2491 (N_2491,N_1909,N_1738);
nand U2492 (N_2492,N_1829,N_1868);
xnor U2493 (N_2493,N_1927,N_1515);
and U2494 (N_2494,N_1522,N_1601);
and U2495 (N_2495,N_1762,N_1562);
nor U2496 (N_2496,N_1823,N_1531);
nor U2497 (N_2497,N_1583,N_1895);
xnor U2498 (N_2498,N_1984,N_1847);
xor U2499 (N_2499,N_1568,N_1806);
nor U2500 (N_2500,N_2307,N_2313);
nor U2501 (N_2501,N_2454,N_2168);
xnor U2502 (N_2502,N_2211,N_2170);
nor U2503 (N_2503,N_2256,N_2364);
nor U2504 (N_2504,N_2300,N_2347);
nand U2505 (N_2505,N_2016,N_2284);
or U2506 (N_2506,N_2000,N_2132);
nor U2507 (N_2507,N_2065,N_2370);
and U2508 (N_2508,N_2298,N_2182);
nor U2509 (N_2509,N_2362,N_2352);
xnor U2510 (N_2510,N_2475,N_2048);
or U2511 (N_2511,N_2176,N_2494);
nor U2512 (N_2512,N_2009,N_2416);
and U2513 (N_2513,N_2237,N_2202);
or U2514 (N_2514,N_2442,N_2072);
xor U2515 (N_2515,N_2154,N_2261);
and U2516 (N_2516,N_2389,N_2192);
nand U2517 (N_2517,N_2451,N_2367);
or U2518 (N_2518,N_2265,N_2255);
and U2519 (N_2519,N_2226,N_2366);
or U2520 (N_2520,N_2477,N_2338);
nand U2521 (N_2521,N_2495,N_2167);
xnor U2522 (N_2522,N_2243,N_2474);
or U2523 (N_2523,N_2463,N_2396);
nor U2524 (N_2524,N_2342,N_2281);
nor U2525 (N_2525,N_2283,N_2285);
or U2526 (N_2526,N_2008,N_2238);
nand U2527 (N_2527,N_2398,N_2058);
and U2528 (N_2528,N_2275,N_2128);
or U2529 (N_2529,N_2091,N_2252);
xnor U2530 (N_2530,N_2085,N_2411);
and U2531 (N_2531,N_2024,N_2186);
nor U2532 (N_2532,N_2376,N_2172);
and U2533 (N_2533,N_2457,N_2053);
or U2534 (N_2534,N_2253,N_2310);
xor U2535 (N_2535,N_2086,N_2328);
nor U2536 (N_2536,N_2138,N_2049);
xnor U2537 (N_2537,N_2054,N_2026);
or U2538 (N_2538,N_2305,N_2287);
or U2539 (N_2539,N_2007,N_2493);
and U2540 (N_2540,N_2302,N_2316);
or U2541 (N_2541,N_2120,N_2260);
nor U2542 (N_2542,N_2344,N_2365);
or U2543 (N_2543,N_2384,N_2435);
nor U2544 (N_2544,N_2066,N_2239);
nor U2545 (N_2545,N_2481,N_2188);
nor U2546 (N_2546,N_2062,N_2277);
xnor U2547 (N_2547,N_2415,N_2464);
xor U2548 (N_2548,N_2232,N_2381);
or U2549 (N_2549,N_2423,N_2038);
and U2550 (N_2550,N_2087,N_2198);
and U2551 (N_2551,N_2079,N_2269);
nor U2552 (N_2552,N_2019,N_2482);
nor U2553 (N_2553,N_2222,N_2057);
nand U2554 (N_2554,N_2459,N_2109);
nor U2555 (N_2555,N_2174,N_2356);
and U2556 (N_2556,N_2273,N_2040);
nor U2557 (N_2557,N_2304,N_2225);
or U2558 (N_2558,N_2361,N_2075);
nand U2559 (N_2559,N_2246,N_2044);
or U2560 (N_2560,N_2006,N_2125);
xnor U2561 (N_2561,N_2490,N_2478);
or U2562 (N_2562,N_2324,N_2144);
nor U2563 (N_2563,N_2380,N_2249);
or U2564 (N_2564,N_2343,N_2122);
nand U2565 (N_2565,N_2462,N_2374);
xnor U2566 (N_2566,N_2259,N_2034);
xor U2567 (N_2567,N_2220,N_2404);
nor U2568 (N_2568,N_2254,N_2156);
and U2569 (N_2569,N_2378,N_2081);
xor U2570 (N_2570,N_2201,N_2326);
or U2571 (N_2571,N_2403,N_2311);
or U2572 (N_2572,N_2372,N_2020);
or U2573 (N_2573,N_2089,N_2064);
xor U2574 (N_2574,N_2409,N_2166);
or U2575 (N_2575,N_2045,N_2337);
and U2576 (N_2576,N_2179,N_2397);
xnor U2577 (N_2577,N_2074,N_2441);
nand U2578 (N_2578,N_2090,N_2180);
and U2579 (N_2579,N_2102,N_2427);
xnor U2580 (N_2580,N_2197,N_2418);
xnor U2581 (N_2581,N_2194,N_2270);
nand U2582 (N_2582,N_2061,N_2139);
or U2583 (N_2583,N_2185,N_2327);
nor U2584 (N_2584,N_2046,N_2425);
xor U2585 (N_2585,N_2027,N_2401);
or U2586 (N_2586,N_2227,N_2395);
nand U2587 (N_2587,N_2322,N_2083);
nand U2588 (N_2588,N_2465,N_2199);
nor U2589 (N_2589,N_2035,N_2468);
xor U2590 (N_2590,N_2453,N_2334);
and U2591 (N_2591,N_2108,N_2244);
or U2592 (N_2592,N_2496,N_2150);
or U2593 (N_2593,N_2208,N_2306);
xor U2594 (N_2594,N_2455,N_2101);
nor U2595 (N_2595,N_2210,N_2025);
or U2596 (N_2596,N_2400,N_2349);
nor U2597 (N_2597,N_2206,N_2052);
or U2598 (N_2598,N_2391,N_2345);
xnor U2599 (N_2599,N_2013,N_2258);
xor U2600 (N_2600,N_2437,N_2164);
or U2601 (N_2601,N_2426,N_2088);
and U2602 (N_2602,N_2387,N_2432);
nand U2603 (N_2603,N_2183,N_2360);
xor U2604 (N_2604,N_2195,N_2375);
xnor U2605 (N_2605,N_2330,N_2077);
nor U2606 (N_2606,N_2341,N_2290);
nand U2607 (N_2607,N_2155,N_2143);
nor U2608 (N_2608,N_2385,N_2325);
xnor U2609 (N_2609,N_2317,N_2279);
nor U2610 (N_2610,N_2377,N_2333);
and U2611 (N_2611,N_2012,N_2294);
nor U2612 (N_2612,N_2022,N_2363);
xor U2613 (N_2613,N_2408,N_2039);
xor U2614 (N_2614,N_2359,N_2178);
nor U2615 (N_2615,N_2340,N_2036);
xnor U2616 (N_2616,N_2469,N_2422);
nor U2617 (N_2617,N_2131,N_2191);
nor U2618 (N_2618,N_2297,N_2233);
and U2619 (N_2619,N_2114,N_2096);
or U2620 (N_2620,N_2230,N_2419);
or U2621 (N_2621,N_2082,N_2456);
xor U2622 (N_2622,N_2399,N_2460);
or U2623 (N_2623,N_2461,N_2486);
nor U2624 (N_2624,N_2219,N_2388);
or U2625 (N_2625,N_2187,N_2073);
xor U2626 (N_2626,N_2485,N_2162);
xnor U2627 (N_2627,N_2234,N_2315);
and U2628 (N_2628,N_2030,N_2293);
or U2629 (N_2629,N_2371,N_2173);
or U2630 (N_2630,N_2355,N_2257);
nand U2631 (N_2631,N_2177,N_2029);
or U2632 (N_2632,N_2130,N_2115);
nand U2633 (N_2633,N_2386,N_2149);
or U2634 (N_2634,N_2228,N_2031);
nand U2635 (N_2635,N_2193,N_2446);
and U2636 (N_2636,N_2161,N_2003);
nand U2637 (N_2637,N_2402,N_2248);
or U2638 (N_2638,N_2134,N_2165);
or U2639 (N_2639,N_2353,N_2414);
or U2640 (N_2640,N_2288,N_2190);
xnor U2641 (N_2641,N_2487,N_2434);
xor U2642 (N_2642,N_2189,N_2145);
xnor U2643 (N_2643,N_2392,N_2480);
or U2644 (N_2644,N_2421,N_2080);
and U2645 (N_2645,N_2171,N_2280);
xnor U2646 (N_2646,N_2471,N_2267);
or U2647 (N_2647,N_2215,N_2436);
or U2648 (N_2648,N_2470,N_2428);
nand U2649 (N_2649,N_2406,N_2489);
xnor U2650 (N_2650,N_2444,N_2107);
xor U2651 (N_2651,N_2430,N_2231);
and U2652 (N_2652,N_2032,N_2136);
or U2653 (N_2653,N_2263,N_2323);
or U2654 (N_2654,N_2318,N_2303);
nand U2655 (N_2655,N_2407,N_2092);
and U2656 (N_2656,N_2289,N_2240);
and U2657 (N_2657,N_2214,N_2157);
or U2658 (N_2658,N_2339,N_2181);
or U2659 (N_2659,N_2160,N_2296);
nand U2660 (N_2660,N_2110,N_2466);
and U2661 (N_2661,N_2041,N_2119);
or U2662 (N_2662,N_2060,N_2314);
nand U2663 (N_2663,N_2169,N_2247);
nand U2664 (N_2664,N_2123,N_2412);
nand U2665 (N_2665,N_2264,N_2135);
nor U2666 (N_2666,N_2076,N_2213);
nand U2667 (N_2667,N_2438,N_2033);
or U2668 (N_2668,N_2229,N_2368);
and U2669 (N_2669,N_2382,N_2433);
or U2670 (N_2670,N_2320,N_2440);
xor U2671 (N_2671,N_2209,N_2319);
nor U2672 (N_2672,N_2014,N_2393);
nand U2673 (N_2673,N_2274,N_2004);
nand U2674 (N_2674,N_2093,N_2429);
xnor U2675 (N_2675,N_2152,N_2050);
xor U2676 (N_2676,N_2126,N_2499);
or U2677 (N_2677,N_2413,N_2498);
nand U2678 (N_2678,N_2002,N_2309);
or U2679 (N_2679,N_2443,N_2017);
xnor U2680 (N_2680,N_2484,N_2373);
xor U2681 (N_2681,N_2369,N_2301);
nand U2682 (N_2682,N_2175,N_2278);
nor U2683 (N_2683,N_2291,N_2070);
nor U2684 (N_2684,N_2184,N_2104);
or U2685 (N_2685,N_2133,N_2335);
xnor U2686 (N_2686,N_2223,N_2106);
nor U2687 (N_2687,N_2063,N_2351);
nor U2688 (N_2688,N_2268,N_2148);
and U2689 (N_2689,N_2023,N_2312);
and U2690 (N_2690,N_2121,N_2488);
or U2691 (N_2691,N_2336,N_2221);
xnor U2692 (N_2692,N_2417,N_2483);
nor U2693 (N_2693,N_2151,N_2276);
and U2694 (N_2694,N_2078,N_2216);
nand U2695 (N_2695,N_2479,N_2129);
nand U2696 (N_2696,N_2118,N_2051);
nor U2697 (N_2697,N_2207,N_2147);
nand U2698 (N_2698,N_2218,N_2266);
xnor U2699 (N_2699,N_2105,N_2021);
nand U2700 (N_2700,N_2212,N_2405);
and U2701 (N_2701,N_2067,N_2042);
or U2702 (N_2702,N_2292,N_2011);
nor U2703 (N_2703,N_2410,N_2431);
nand U2704 (N_2704,N_2037,N_2449);
xor U2705 (N_2705,N_2069,N_2439);
nor U2706 (N_2706,N_2295,N_2491);
nand U2707 (N_2707,N_2354,N_2472);
nor U2708 (N_2708,N_2346,N_2348);
nand U2709 (N_2709,N_2163,N_2332);
nor U2710 (N_2710,N_2497,N_2241);
xor U2711 (N_2711,N_2245,N_2250);
nor U2712 (N_2712,N_2424,N_2116);
nor U2713 (N_2713,N_2055,N_2084);
and U2714 (N_2714,N_2282,N_2350);
nand U2715 (N_2715,N_2094,N_2321);
and U2716 (N_2716,N_2196,N_2331);
xor U2717 (N_2717,N_2420,N_2095);
xor U2718 (N_2718,N_2271,N_2127);
nor U2719 (N_2719,N_2358,N_2113);
or U2720 (N_2720,N_2200,N_2390);
or U2721 (N_2721,N_2111,N_2262);
or U2722 (N_2722,N_2142,N_2203);
nor U2723 (N_2723,N_2100,N_2047);
and U2724 (N_2724,N_2492,N_2236);
nor U2725 (N_2725,N_2137,N_2001);
or U2726 (N_2726,N_2272,N_2447);
or U2727 (N_2727,N_2224,N_2010);
nor U2728 (N_2728,N_2098,N_2379);
or U2729 (N_2729,N_2242,N_2357);
nand U2730 (N_2730,N_2467,N_2028);
xnor U2731 (N_2731,N_2286,N_2056);
nor U2732 (N_2732,N_2251,N_2205);
nand U2733 (N_2733,N_2124,N_2099);
nor U2734 (N_2734,N_2043,N_2097);
nand U2735 (N_2735,N_2068,N_2448);
xnor U2736 (N_2736,N_2217,N_2140);
and U2737 (N_2737,N_2005,N_2473);
nand U2738 (N_2738,N_2158,N_2146);
nor U2739 (N_2739,N_2383,N_2117);
nor U2740 (N_2740,N_2015,N_2059);
xor U2741 (N_2741,N_2071,N_2141);
and U2742 (N_2742,N_2103,N_2394);
and U2743 (N_2743,N_2153,N_2204);
xnor U2744 (N_2744,N_2445,N_2329);
xor U2745 (N_2745,N_2458,N_2112);
xnor U2746 (N_2746,N_2235,N_2452);
or U2747 (N_2747,N_2308,N_2018);
xor U2748 (N_2748,N_2299,N_2476);
and U2749 (N_2749,N_2450,N_2159);
nor U2750 (N_2750,N_2057,N_2178);
or U2751 (N_2751,N_2179,N_2335);
nand U2752 (N_2752,N_2232,N_2466);
nand U2753 (N_2753,N_2332,N_2467);
nor U2754 (N_2754,N_2113,N_2319);
nor U2755 (N_2755,N_2006,N_2386);
and U2756 (N_2756,N_2163,N_2325);
nand U2757 (N_2757,N_2107,N_2457);
nand U2758 (N_2758,N_2185,N_2042);
or U2759 (N_2759,N_2145,N_2457);
nor U2760 (N_2760,N_2369,N_2248);
and U2761 (N_2761,N_2446,N_2363);
nor U2762 (N_2762,N_2083,N_2167);
or U2763 (N_2763,N_2473,N_2137);
nor U2764 (N_2764,N_2376,N_2315);
nor U2765 (N_2765,N_2444,N_2285);
nand U2766 (N_2766,N_2456,N_2145);
nor U2767 (N_2767,N_2039,N_2401);
xor U2768 (N_2768,N_2140,N_2019);
xor U2769 (N_2769,N_2195,N_2284);
and U2770 (N_2770,N_2100,N_2092);
or U2771 (N_2771,N_2118,N_2386);
xor U2772 (N_2772,N_2033,N_2228);
nor U2773 (N_2773,N_2168,N_2396);
nand U2774 (N_2774,N_2100,N_2314);
nand U2775 (N_2775,N_2401,N_2298);
or U2776 (N_2776,N_2157,N_2360);
or U2777 (N_2777,N_2481,N_2024);
nand U2778 (N_2778,N_2411,N_2406);
and U2779 (N_2779,N_2455,N_2430);
nor U2780 (N_2780,N_2175,N_2150);
xnor U2781 (N_2781,N_2069,N_2491);
nor U2782 (N_2782,N_2427,N_2208);
and U2783 (N_2783,N_2142,N_2164);
and U2784 (N_2784,N_2137,N_2046);
or U2785 (N_2785,N_2070,N_2024);
xnor U2786 (N_2786,N_2120,N_2272);
or U2787 (N_2787,N_2439,N_2477);
nand U2788 (N_2788,N_2478,N_2200);
or U2789 (N_2789,N_2173,N_2000);
nor U2790 (N_2790,N_2031,N_2265);
and U2791 (N_2791,N_2331,N_2008);
and U2792 (N_2792,N_2228,N_2495);
nor U2793 (N_2793,N_2255,N_2178);
xor U2794 (N_2794,N_2395,N_2164);
and U2795 (N_2795,N_2482,N_2165);
xnor U2796 (N_2796,N_2313,N_2054);
or U2797 (N_2797,N_2099,N_2054);
xnor U2798 (N_2798,N_2277,N_2005);
and U2799 (N_2799,N_2001,N_2319);
nor U2800 (N_2800,N_2121,N_2487);
and U2801 (N_2801,N_2300,N_2271);
xor U2802 (N_2802,N_2488,N_2193);
xnor U2803 (N_2803,N_2117,N_2171);
and U2804 (N_2804,N_2248,N_2327);
nand U2805 (N_2805,N_2392,N_2251);
xor U2806 (N_2806,N_2222,N_2219);
nand U2807 (N_2807,N_2488,N_2406);
xor U2808 (N_2808,N_2066,N_2443);
xor U2809 (N_2809,N_2342,N_2348);
nor U2810 (N_2810,N_2215,N_2101);
or U2811 (N_2811,N_2200,N_2042);
or U2812 (N_2812,N_2169,N_2439);
nand U2813 (N_2813,N_2092,N_2061);
or U2814 (N_2814,N_2116,N_2015);
nor U2815 (N_2815,N_2070,N_2297);
or U2816 (N_2816,N_2323,N_2314);
and U2817 (N_2817,N_2048,N_2013);
nand U2818 (N_2818,N_2254,N_2342);
xor U2819 (N_2819,N_2241,N_2159);
and U2820 (N_2820,N_2156,N_2245);
nand U2821 (N_2821,N_2071,N_2208);
and U2822 (N_2822,N_2407,N_2281);
nand U2823 (N_2823,N_2352,N_2408);
nor U2824 (N_2824,N_2487,N_2294);
or U2825 (N_2825,N_2372,N_2311);
or U2826 (N_2826,N_2250,N_2282);
xnor U2827 (N_2827,N_2164,N_2221);
and U2828 (N_2828,N_2148,N_2231);
or U2829 (N_2829,N_2098,N_2481);
and U2830 (N_2830,N_2179,N_2262);
and U2831 (N_2831,N_2042,N_2347);
or U2832 (N_2832,N_2055,N_2112);
or U2833 (N_2833,N_2281,N_2390);
and U2834 (N_2834,N_2100,N_2084);
nor U2835 (N_2835,N_2427,N_2295);
nand U2836 (N_2836,N_2497,N_2350);
xor U2837 (N_2837,N_2025,N_2058);
nand U2838 (N_2838,N_2089,N_2429);
nor U2839 (N_2839,N_2059,N_2070);
nand U2840 (N_2840,N_2354,N_2080);
and U2841 (N_2841,N_2482,N_2091);
xor U2842 (N_2842,N_2047,N_2140);
xor U2843 (N_2843,N_2371,N_2355);
nand U2844 (N_2844,N_2182,N_2161);
xor U2845 (N_2845,N_2367,N_2340);
nor U2846 (N_2846,N_2088,N_2342);
xor U2847 (N_2847,N_2060,N_2137);
or U2848 (N_2848,N_2465,N_2042);
and U2849 (N_2849,N_2208,N_2343);
nor U2850 (N_2850,N_2352,N_2219);
and U2851 (N_2851,N_2273,N_2022);
or U2852 (N_2852,N_2299,N_2195);
and U2853 (N_2853,N_2478,N_2259);
and U2854 (N_2854,N_2437,N_2371);
or U2855 (N_2855,N_2134,N_2253);
or U2856 (N_2856,N_2400,N_2078);
xnor U2857 (N_2857,N_2411,N_2347);
nand U2858 (N_2858,N_2102,N_2303);
xor U2859 (N_2859,N_2330,N_2179);
nand U2860 (N_2860,N_2454,N_2096);
and U2861 (N_2861,N_2211,N_2201);
nor U2862 (N_2862,N_2118,N_2183);
and U2863 (N_2863,N_2238,N_2176);
and U2864 (N_2864,N_2029,N_2195);
or U2865 (N_2865,N_2094,N_2402);
nor U2866 (N_2866,N_2054,N_2308);
or U2867 (N_2867,N_2348,N_2270);
or U2868 (N_2868,N_2055,N_2178);
or U2869 (N_2869,N_2266,N_2484);
or U2870 (N_2870,N_2003,N_2415);
xor U2871 (N_2871,N_2023,N_2055);
xnor U2872 (N_2872,N_2321,N_2273);
nand U2873 (N_2873,N_2455,N_2154);
nor U2874 (N_2874,N_2028,N_2181);
nor U2875 (N_2875,N_2284,N_2313);
xnor U2876 (N_2876,N_2080,N_2470);
xor U2877 (N_2877,N_2111,N_2243);
or U2878 (N_2878,N_2177,N_2392);
and U2879 (N_2879,N_2345,N_2475);
xor U2880 (N_2880,N_2214,N_2291);
xnor U2881 (N_2881,N_2021,N_2497);
nor U2882 (N_2882,N_2494,N_2354);
or U2883 (N_2883,N_2403,N_2238);
or U2884 (N_2884,N_2194,N_2163);
and U2885 (N_2885,N_2257,N_2236);
nor U2886 (N_2886,N_2080,N_2033);
xnor U2887 (N_2887,N_2148,N_2238);
xnor U2888 (N_2888,N_2369,N_2472);
nor U2889 (N_2889,N_2326,N_2444);
nand U2890 (N_2890,N_2378,N_2050);
or U2891 (N_2891,N_2499,N_2164);
or U2892 (N_2892,N_2369,N_2304);
or U2893 (N_2893,N_2344,N_2101);
or U2894 (N_2894,N_2465,N_2043);
xnor U2895 (N_2895,N_2323,N_2461);
xnor U2896 (N_2896,N_2232,N_2017);
nor U2897 (N_2897,N_2024,N_2161);
xnor U2898 (N_2898,N_2206,N_2424);
and U2899 (N_2899,N_2465,N_2141);
xnor U2900 (N_2900,N_2265,N_2206);
xnor U2901 (N_2901,N_2475,N_2422);
nor U2902 (N_2902,N_2451,N_2038);
nand U2903 (N_2903,N_2278,N_2028);
nor U2904 (N_2904,N_2196,N_2241);
and U2905 (N_2905,N_2051,N_2129);
nor U2906 (N_2906,N_2016,N_2000);
xor U2907 (N_2907,N_2499,N_2034);
xor U2908 (N_2908,N_2208,N_2256);
nor U2909 (N_2909,N_2450,N_2142);
nand U2910 (N_2910,N_2116,N_2386);
and U2911 (N_2911,N_2043,N_2254);
or U2912 (N_2912,N_2117,N_2060);
nor U2913 (N_2913,N_2305,N_2200);
nor U2914 (N_2914,N_2021,N_2441);
nand U2915 (N_2915,N_2449,N_2162);
and U2916 (N_2916,N_2214,N_2196);
xnor U2917 (N_2917,N_2052,N_2333);
xor U2918 (N_2918,N_2376,N_2464);
nor U2919 (N_2919,N_2378,N_2426);
and U2920 (N_2920,N_2285,N_2385);
or U2921 (N_2921,N_2411,N_2134);
nor U2922 (N_2922,N_2259,N_2301);
and U2923 (N_2923,N_2409,N_2456);
nor U2924 (N_2924,N_2302,N_2044);
or U2925 (N_2925,N_2265,N_2300);
xor U2926 (N_2926,N_2243,N_2379);
xnor U2927 (N_2927,N_2136,N_2301);
and U2928 (N_2928,N_2036,N_2338);
and U2929 (N_2929,N_2386,N_2469);
nor U2930 (N_2930,N_2461,N_2290);
xnor U2931 (N_2931,N_2426,N_2050);
and U2932 (N_2932,N_2188,N_2409);
or U2933 (N_2933,N_2259,N_2226);
and U2934 (N_2934,N_2257,N_2386);
or U2935 (N_2935,N_2353,N_2235);
xnor U2936 (N_2936,N_2323,N_2075);
nor U2937 (N_2937,N_2406,N_2273);
or U2938 (N_2938,N_2399,N_2176);
or U2939 (N_2939,N_2069,N_2477);
or U2940 (N_2940,N_2286,N_2308);
nand U2941 (N_2941,N_2005,N_2482);
xor U2942 (N_2942,N_2497,N_2189);
nor U2943 (N_2943,N_2463,N_2186);
or U2944 (N_2944,N_2399,N_2223);
nor U2945 (N_2945,N_2017,N_2207);
or U2946 (N_2946,N_2361,N_2056);
xnor U2947 (N_2947,N_2290,N_2441);
nor U2948 (N_2948,N_2193,N_2111);
and U2949 (N_2949,N_2352,N_2357);
or U2950 (N_2950,N_2392,N_2174);
or U2951 (N_2951,N_2155,N_2056);
or U2952 (N_2952,N_2458,N_2420);
xnor U2953 (N_2953,N_2222,N_2210);
nor U2954 (N_2954,N_2388,N_2241);
xnor U2955 (N_2955,N_2474,N_2323);
xnor U2956 (N_2956,N_2376,N_2228);
xor U2957 (N_2957,N_2410,N_2348);
nor U2958 (N_2958,N_2474,N_2331);
xor U2959 (N_2959,N_2123,N_2307);
xor U2960 (N_2960,N_2358,N_2181);
or U2961 (N_2961,N_2418,N_2117);
xor U2962 (N_2962,N_2104,N_2294);
or U2963 (N_2963,N_2467,N_2380);
nand U2964 (N_2964,N_2218,N_2455);
nor U2965 (N_2965,N_2042,N_2120);
nor U2966 (N_2966,N_2142,N_2028);
xnor U2967 (N_2967,N_2280,N_2174);
and U2968 (N_2968,N_2328,N_2288);
nand U2969 (N_2969,N_2414,N_2320);
nand U2970 (N_2970,N_2467,N_2382);
or U2971 (N_2971,N_2094,N_2267);
xor U2972 (N_2972,N_2302,N_2461);
or U2973 (N_2973,N_2332,N_2442);
nor U2974 (N_2974,N_2277,N_2263);
xnor U2975 (N_2975,N_2219,N_2008);
nor U2976 (N_2976,N_2167,N_2194);
or U2977 (N_2977,N_2076,N_2429);
and U2978 (N_2978,N_2099,N_2138);
or U2979 (N_2979,N_2337,N_2193);
and U2980 (N_2980,N_2284,N_2122);
or U2981 (N_2981,N_2104,N_2108);
xnor U2982 (N_2982,N_2035,N_2093);
or U2983 (N_2983,N_2226,N_2146);
and U2984 (N_2984,N_2293,N_2034);
xnor U2985 (N_2985,N_2085,N_2294);
nor U2986 (N_2986,N_2101,N_2353);
and U2987 (N_2987,N_2322,N_2310);
nor U2988 (N_2988,N_2499,N_2016);
nor U2989 (N_2989,N_2074,N_2096);
nor U2990 (N_2990,N_2342,N_2169);
xnor U2991 (N_2991,N_2106,N_2382);
and U2992 (N_2992,N_2032,N_2015);
or U2993 (N_2993,N_2087,N_2234);
nand U2994 (N_2994,N_2366,N_2168);
or U2995 (N_2995,N_2180,N_2371);
nor U2996 (N_2996,N_2302,N_2262);
or U2997 (N_2997,N_2066,N_2017);
nor U2998 (N_2998,N_2264,N_2017);
nand U2999 (N_2999,N_2316,N_2076);
nor U3000 (N_3000,N_2644,N_2777);
or U3001 (N_3001,N_2517,N_2625);
nor U3002 (N_3002,N_2804,N_2505);
nand U3003 (N_3003,N_2569,N_2978);
or U3004 (N_3004,N_2530,N_2573);
nor U3005 (N_3005,N_2768,N_2692);
nor U3006 (N_3006,N_2633,N_2997);
nand U3007 (N_3007,N_2657,N_2595);
xnor U3008 (N_3008,N_2811,N_2765);
and U3009 (N_3009,N_2709,N_2776);
xnor U3010 (N_3010,N_2626,N_2553);
xnor U3011 (N_3011,N_2965,N_2749);
and U3012 (N_3012,N_2945,N_2634);
xor U3013 (N_3013,N_2724,N_2981);
nor U3014 (N_3014,N_2693,N_2576);
and U3015 (N_3015,N_2786,N_2887);
nand U3016 (N_3016,N_2800,N_2868);
or U3017 (N_3017,N_2881,N_2852);
nand U3018 (N_3018,N_2829,N_2900);
nor U3019 (N_3019,N_2734,N_2739);
xnor U3020 (N_3020,N_2884,N_2820);
nand U3021 (N_3021,N_2919,N_2585);
nand U3022 (N_3022,N_2617,N_2509);
nor U3023 (N_3023,N_2688,N_2527);
and U3024 (N_3024,N_2694,N_2774);
or U3025 (N_3025,N_2912,N_2841);
and U3026 (N_3026,N_2977,N_2715);
nor U3027 (N_3027,N_2669,N_2629);
xor U3028 (N_3028,N_2973,N_2848);
nand U3029 (N_3029,N_2771,N_2551);
nand U3030 (N_3030,N_2850,N_2647);
or U3031 (N_3031,N_2787,N_2728);
nand U3032 (N_3032,N_2955,N_2914);
and U3033 (N_3033,N_2649,N_2807);
nor U3034 (N_3034,N_2612,N_2825);
nand U3035 (N_3035,N_2792,N_2526);
and U3036 (N_3036,N_2913,N_2990);
nand U3037 (N_3037,N_2580,N_2630);
nand U3038 (N_3038,N_2520,N_2677);
nand U3039 (N_3039,N_2872,N_2631);
or U3040 (N_3040,N_2966,N_2687);
xnor U3041 (N_3041,N_2581,N_2718);
nor U3042 (N_3042,N_2579,N_2860);
nand U3043 (N_3043,N_2938,N_2871);
and U3044 (N_3044,N_2598,N_2703);
nand U3045 (N_3045,N_2643,N_2952);
nand U3046 (N_3046,N_2590,N_2722);
nor U3047 (N_3047,N_2500,N_2970);
or U3048 (N_3048,N_2753,N_2655);
xnor U3049 (N_3049,N_2660,N_2839);
and U3050 (N_3050,N_2568,N_2866);
nand U3051 (N_3051,N_2911,N_2802);
or U3052 (N_3052,N_2556,N_2983);
or U3053 (N_3053,N_2897,N_2591);
and U3054 (N_3054,N_2759,N_2535);
or U3055 (N_3055,N_2902,N_2817);
xnor U3056 (N_3056,N_2691,N_2925);
nand U3057 (N_3057,N_2684,N_2957);
xor U3058 (N_3058,N_2732,N_2798);
nor U3059 (N_3059,N_2958,N_2922);
or U3060 (N_3060,N_2570,N_2609);
and U3061 (N_3061,N_2908,N_2877);
and U3062 (N_3062,N_2931,N_2658);
nor U3063 (N_3063,N_2894,N_2823);
nor U3064 (N_3064,N_2795,N_2755);
xnor U3065 (N_3065,N_2775,N_2843);
xor U3066 (N_3066,N_2700,N_2679);
nand U3067 (N_3067,N_2803,N_2648);
nand U3068 (N_3068,N_2704,N_2519);
nor U3069 (N_3069,N_2555,N_2758);
nand U3070 (N_3070,N_2858,N_2623);
nand U3071 (N_3071,N_2599,N_2670);
nor U3072 (N_3072,N_2501,N_2636);
or U3073 (N_3073,N_2559,N_2948);
xnor U3074 (N_3074,N_2707,N_2906);
xor U3075 (N_3075,N_2793,N_2600);
xnor U3076 (N_3076,N_2762,N_2743);
xnor U3077 (N_3077,N_2515,N_2571);
nor U3078 (N_3078,N_2550,N_2790);
nor U3079 (N_3079,N_2674,N_2893);
nand U3080 (N_3080,N_2514,N_2750);
xor U3081 (N_3081,N_2689,N_2988);
nand U3082 (N_3082,N_2933,N_2961);
nor U3083 (N_3083,N_2661,N_2747);
and U3084 (N_3084,N_2865,N_2620);
nor U3085 (N_3085,N_2540,N_2699);
or U3086 (N_3086,N_2736,N_2766);
nand U3087 (N_3087,N_2979,N_2932);
nand U3088 (N_3088,N_2849,N_2903);
xnor U3089 (N_3089,N_2830,N_2876);
and U3090 (N_3090,N_2896,N_2974);
xor U3091 (N_3091,N_2522,N_2992);
xnor U3092 (N_3092,N_2980,N_2589);
nand U3093 (N_3093,N_2744,N_2534);
or U3094 (N_3094,N_2951,N_2929);
or U3095 (N_3095,N_2822,N_2667);
or U3096 (N_3096,N_2878,N_2873);
nor U3097 (N_3097,N_2563,N_2676);
or U3098 (N_3098,N_2883,N_2835);
and U3099 (N_3099,N_2603,N_2627);
nor U3100 (N_3100,N_2761,N_2711);
nor U3101 (N_3101,N_2574,N_2921);
or U3102 (N_3102,N_2808,N_2543);
xnor U3103 (N_3103,N_2721,N_2898);
nor U3104 (N_3104,N_2927,N_2828);
nand U3105 (N_3105,N_2837,N_2564);
nand U3106 (N_3106,N_2751,N_2546);
nand U3107 (N_3107,N_2549,N_2935);
or U3108 (N_3108,N_2583,N_2597);
or U3109 (N_3109,N_2943,N_2991);
nor U3110 (N_3110,N_2586,N_2614);
nand U3111 (N_3111,N_2842,N_2740);
and U3112 (N_3112,N_2696,N_2741);
nor U3113 (N_3113,N_2662,N_2999);
nand U3114 (N_3114,N_2639,N_2710);
or U3115 (N_3115,N_2757,N_2924);
and U3116 (N_3116,N_2596,N_2818);
nor U3117 (N_3117,N_2557,N_2838);
nor U3118 (N_3118,N_2545,N_2554);
xnor U3119 (N_3119,N_2953,N_2746);
nor U3120 (N_3120,N_2941,N_2544);
nand U3121 (N_3121,N_2909,N_2760);
nand U3122 (N_3122,N_2816,N_2552);
and U3123 (N_3123,N_2613,N_2770);
nand U3124 (N_3124,N_2652,N_2806);
xor U3125 (N_3125,N_2604,N_2507);
or U3126 (N_3126,N_2588,N_2930);
xnor U3127 (N_3127,N_2752,N_2976);
and U3128 (N_3128,N_2989,N_2745);
and U3129 (N_3129,N_2510,N_2869);
and U3130 (N_3130,N_2946,N_2767);
nand U3131 (N_3131,N_2528,N_2809);
or U3132 (N_3132,N_2685,N_2686);
nand U3133 (N_3133,N_2713,N_2610);
xor U3134 (N_3134,N_2511,N_2773);
nor U3135 (N_3135,N_2531,N_2650);
xor U3136 (N_3136,N_2797,N_2738);
nor U3137 (N_3137,N_2547,N_2791);
and U3138 (N_3138,N_2857,N_2731);
xnor U3139 (N_3139,N_2836,N_2907);
nor U3140 (N_3140,N_2889,N_2833);
xnor U3141 (N_3141,N_2780,N_2541);
or U3142 (N_3142,N_2993,N_2725);
and U3143 (N_3143,N_2592,N_2533);
xor U3144 (N_3144,N_2844,N_2910);
nor U3145 (N_3145,N_2769,N_2706);
or U3146 (N_3146,N_2875,N_2892);
nand U3147 (N_3147,N_2882,N_2819);
or U3148 (N_3148,N_2512,N_2834);
or U3149 (N_3149,N_2895,N_2575);
or U3150 (N_3150,N_2779,N_2923);
or U3151 (N_3151,N_2645,N_2523);
or U3152 (N_3152,N_2611,N_2672);
nand U3153 (N_3153,N_2680,N_2944);
and U3154 (N_3154,N_2756,N_2683);
nor U3155 (N_3155,N_2789,N_2864);
xor U3156 (N_3156,N_2840,N_2524);
xor U3157 (N_3157,N_2954,N_2862);
nand U3158 (N_3158,N_2577,N_2561);
or U3159 (N_3159,N_2947,N_2607);
xnor U3160 (N_3160,N_2995,N_2717);
or U3161 (N_3161,N_2937,N_2730);
nor U3162 (N_3162,N_2506,N_2879);
nand U3163 (N_3163,N_2542,N_2987);
nor U3164 (N_3164,N_2861,N_2982);
xnor U3165 (N_3165,N_2619,N_2827);
nor U3166 (N_3166,N_2681,N_2601);
nor U3167 (N_3167,N_2608,N_2962);
nand U3168 (N_3168,N_2521,N_2801);
nand U3169 (N_3169,N_2621,N_2967);
and U3170 (N_3170,N_2796,N_2504);
nand U3171 (N_3171,N_2939,N_2984);
nor U3172 (N_3172,N_2959,N_2641);
xnor U3173 (N_3173,N_2794,N_2782);
or U3174 (N_3174,N_2664,N_2513);
nand U3175 (N_3175,N_2847,N_2508);
nor U3176 (N_3176,N_2863,N_2783);
xnor U3177 (N_3177,N_2714,N_2737);
and U3178 (N_3178,N_2594,N_2697);
and U3179 (N_3179,N_2905,N_2821);
or U3180 (N_3180,N_2870,N_2815);
xnor U3181 (N_3181,N_2651,N_2781);
nand U3182 (N_3182,N_2587,N_2695);
nor U3183 (N_3183,N_2605,N_2845);
xnor U3184 (N_3184,N_2727,N_2719);
and U3185 (N_3185,N_2940,N_2560);
and U3186 (N_3186,N_2867,N_2874);
nand U3187 (N_3187,N_2969,N_2936);
xor U3188 (N_3188,N_2723,N_2538);
nand U3189 (N_3189,N_2890,N_2671);
nor U3190 (N_3190,N_2562,N_2615);
nand U3191 (N_3191,N_2733,N_2772);
and U3192 (N_3192,N_2566,N_2885);
xor U3193 (N_3193,N_2754,N_2656);
nand U3194 (N_3194,N_2826,N_2799);
nand U3195 (N_3195,N_2539,N_2659);
or U3196 (N_3196,N_2701,N_2891);
and U3197 (N_3197,N_2788,N_2675);
and U3198 (N_3198,N_2996,N_2926);
nand U3199 (N_3199,N_2690,N_2968);
or U3200 (N_3200,N_2646,N_2628);
xor U3201 (N_3201,N_2637,N_2720);
or U3202 (N_3202,N_2853,N_2904);
or U3203 (N_3203,N_2582,N_2934);
nor U3204 (N_3204,N_2854,N_2640);
or U3205 (N_3205,N_2712,N_2888);
xor U3206 (N_3206,N_2666,N_2972);
nand U3207 (N_3207,N_2994,N_2813);
or U3208 (N_3208,N_2502,N_2537);
xor U3209 (N_3209,N_2529,N_2729);
or U3210 (N_3210,N_2812,N_2971);
and U3211 (N_3211,N_2763,N_2824);
and U3212 (N_3212,N_2602,N_2856);
nor U3213 (N_3213,N_2949,N_2964);
or U3214 (N_3214,N_2920,N_2654);
and U3215 (N_3215,N_2682,N_2899);
or U3216 (N_3216,N_2525,N_2831);
or U3217 (N_3217,N_2632,N_2678);
or U3218 (N_3218,N_2916,N_2986);
or U3219 (N_3219,N_2518,N_2859);
or U3220 (N_3220,N_2572,N_2653);
and U3221 (N_3221,N_2901,N_2846);
nand U3222 (N_3222,N_2668,N_2764);
and U3223 (N_3223,N_2698,N_2503);
nand U3224 (N_3224,N_2702,N_2998);
or U3225 (N_3225,N_2622,N_2624);
nand U3226 (N_3226,N_2942,N_2716);
xor U3227 (N_3227,N_2532,N_2810);
nand U3228 (N_3228,N_2880,N_2778);
or U3229 (N_3229,N_2814,N_2805);
and U3230 (N_3230,N_2950,N_2638);
nor U3231 (N_3231,N_2708,N_2917);
nor U3232 (N_3232,N_2663,N_2673);
nand U3233 (N_3233,N_2616,N_2726);
nand U3234 (N_3234,N_2928,N_2536);
nand U3235 (N_3235,N_2963,N_2665);
nand U3236 (N_3236,N_2618,N_2548);
xnor U3237 (N_3237,N_2584,N_2516);
nor U3238 (N_3238,N_2567,N_2985);
or U3239 (N_3239,N_2960,N_2855);
nor U3240 (N_3240,N_2558,N_2851);
nor U3241 (N_3241,N_2735,N_2565);
xnor U3242 (N_3242,N_2784,N_2956);
xor U3243 (N_3243,N_2886,N_2593);
or U3244 (N_3244,N_2642,N_2832);
or U3245 (N_3245,N_2606,N_2785);
and U3246 (N_3246,N_2635,N_2742);
nand U3247 (N_3247,N_2915,N_2918);
xnor U3248 (N_3248,N_2748,N_2578);
xnor U3249 (N_3249,N_2705,N_2975);
xor U3250 (N_3250,N_2684,N_2961);
xnor U3251 (N_3251,N_2616,N_2628);
nor U3252 (N_3252,N_2933,N_2872);
or U3253 (N_3253,N_2849,N_2527);
xnor U3254 (N_3254,N_2827,N_2815);
and U3255 (N_3255,N_2819,N_2612);
nand U3256 (N_3256,N_2528,N_2566);
nor U3257 (N_3257,N_2527,N_2968);
nor U3258 (N_3258,N_2736,N_2825);
nand U3259 (N_3259,N_2984,N_2714);
nor U3260 (N_3260,N_2936,N_2689);
nand U3261 (N_3261,N_2762,N_2652);
nand U3262 (N_3262,N_2510,N_2604);
and U3263 (N_3263,N_2986,N_2640);
nor U3264 (N_3264,N_2991,N_2522);
and U3265 (N_3265,N_2716,N_2558);
and U3266 (N_3266,N_2512,N_2795);
xor U3267 (N_3267,N_2946,N_2864);
nand U3268 (N_3268,N_2789,N_2727);
or U3269 (N_3269,N_2805,N_2812);
or U3270 (N_3270,N_2912,N_2635);
xnor U3271 (N_3271,N_2544,N_2688);
xor U3272 (N_3272,N_2971,N_2928);
or U3273 (N_3273,N_2718,N_2770);
or U3274 (N_3274,N_2618,N_2506);
nand U3275 (N_3275,N_2548,N_2512);
nor U3276 (N_3276,N_2833,N_2644);
or U3277 (N_3277,N_2811,N_2540);
or U3278 (N_3278,N_2507,N_2686);
nor U3279 (N_3279,N_2756,N_2534);
xnor U3280 (N_3280,N_2833,N_2968);
or U3281 (N_3281,N_2519,N_2911);
or U3282 (N_3282,N_2563,N_2599);
nor U3283 (N_3283,N_2770,N_2989);
or U3284 (N_3284,N_2687,N_2837);
and U3285 (N_3285,N_2982,N_2806);
or U3286 (N_3286,N_2508,N_2945);
or U3287 (N_3287,N_2621,N_2576);
and U3288 (N_3288,N_2884,N_2769);
and U3289 (N_3289,N_2917,N_2572);
and U3290 (N_3290,N_2817,N_2620);
xor U3291 (N_3291,N_2963,N_2649);
and U3292 (N_3292,N_2546,N_2998);
and U3293 (N_3293,N_2735,N_2864);
xnor U3294 (N_3294,N_2862,N_2936);
and U3295 (N_3295,N_2886,N_2585);
nor U3296 (N_3296,N_2862,N_2839);
nand U3297 (N_3297,N_2541,N_2507);
nand U3298 (N_3298,N_2506,N_2617);
xnor U3299 (N_3299,N_2977,N_2564);
nor U3300 (N_3300,N_2902,N_2709);
or U3301 (N_3301,N_2615,N_2577);
nor U3302 (N_3302,N_2824,N_2896);
nand U3303 (N_3303,N_2882,N_2778);
or U3304 (N_3304,N_2843,N_2771);
nand U3305 (N_3305,N_2894,N_2547);
nor U3306 (N_3306,N_2799,N_2504);
or U3307 (N_3307,N_2706,N_2753);
nand U3308 (N_3308,N_2778,N_2839);
and U3309 (N_3309,N_2987,N_2564);
or U3310 (N_3310,N_2738,N_2516);
nor U3311 (N_3311,N_2677,N_2551);
nand U3312 (N_3312,N_2500,N_2860);
or U3313 (N_3313,N_2551,N_2858);
nor U3314 (N_3314,N_2814,N_2501);
and U3315 (N_3315,N_2594,N_2785);
nand U3316 (N_3316,N_2929,N_2515);
xnor U3317 (N_3317,N_2859,N_2830);
and U3318 (N_3318,N_2710,N_2874);
xnor U3319 (N_3319,N_2543,N_2611);
nor U3320 (N_3320,N_2568,N_2877);
nand U3321 (N_3321,N_2578,N_2682);
nand U3322 (N_3322,N_2979,N_2672);
nand U3323 (N_3323,N_2932,N_2920);
and U3324 (N_3324,N_2510,N_2990);
and U3325 (N_3325,N_2736,N_2550);
and U3326 (N_3326,N_2640,N_2683);
nor U3327 (N_3327,N_2887,N_2803);
nor U3328 (N_3328,N_2686,N_2540);
and U3329 (N_3329,N_2506,N_2589);
nand U3330 (N_3330,N_2554,N_2594);
and U3331 (N_3331,N_2714,N_2578);
nor U3332 (N_3332,N_2854,N_2694);
or U3333 (N_3333,N_2745,N_2904);
nor U3334 (N_3334,N_2956,N_2501);
and U3335 (N_3335,N_2607,N_2855);
nor U3336 (N_3336,N_2678,N_2537);
or U3337 (N_3337,N_2583,N_2752);
xnor U3338 (N_3338,N_2948,N_2679);
and U3339 (N_3339,N_2900,N_2907);
and U3340 (N_3340,N_2802,N_2861);
and U3341 (N_3341,N_2607,N_2586);
or U3342 (N_3342,N_2682,N_2577);
xnor U3343 (N_3343,N_2794,N_2888);
or U3344 (N_3344,N_2995,N_2633);
or U3345 (N_3345,N_2868,N_2678);
or U3346 (N_3346,N_2874,N_2881);
xor U3347 (N_3347,N_2626,N_2798);
nand U3348 (N_3348,N_2754,N_2775);
xnor U3349 (N_3349,N_2518,N_2578);
or U3350 (N_3350,N_2762,N_2672);
or U3351 (N_3351,N_2925,N_2705);
xor U3352 (N_3352,N_2813,N_2636);
or U3353 (N_3353,N_2535,N_2800);
nand U3354 (N_3354,N_2509,N_2924);
xor U3355 (N_3355,N_2586,N_2760);
nor U3356 (N_3356,N_2812,N_2883);
xnor U3357 (N_3357,N_2638,N_2769);
and U3358 (N_3358,N_2948,N_2606);
xnor U3359 (N_3359,N_2751,N_2574);
or U3360 (N_3360,N_2549,N_2633);
or U3361 (N_3361,N_2871,N_2933);
xnor U3362 (N_3362,N_2519,N_2503);
or U3363 (N_3363,N_2553,N_2564);
nor U3364 (N_3364,N_2733,N_2775);
and U3365 (N_3365,N_2628,N_2930);
nand U3366 (N_3366,N_2517,N_2662);
nand U3367 (N_3367,N_2718,N_2902);
xor U3368 (N_3368,N_2642,N_2914);
and U3369 (N_3369,N_2758,N_2594);
nor U3370 (N_3370,N_2707,N_2594);
nand U3371 (N_3371,N_2665,N_2924);
nand U3372 (N_3372,N_2948,N_2538);
xor U3373 (N_3373,N_2843,N_2779);
nand U3374 (N_3374,N_2906,N_2911);
nand U3375 (N_3375,N_2967,N_2534);
nand U3376 (N_3376,N_2531,N_2945);
nor U3377 (N_3377,N_2676,N_2677);
nor U3378 (N_3378,N_2814,N_2779);
or U3379 (N_3379,N_2587,N_2502);
or U3380 (N_3380,N_2694,N_2925);
nand U3381 (N_3381,N_2605,N_2926);
nand U3382 (N_3382,N_2636,N_2760);
or U3383 (N_3383,N_2859,N_2832);
nor U3384 (N_3384,N_2633,N_2564);
xor U3385 (N_3385,N_2690,N_2916);
xor U3386 (N_3386,N_2514,N_2804);
nand U3387 (N_3387,N_2612,N_2968);
xor U3388 (N_3388,N_2703,N_2937);
xor U3389 (N_3389,N_2828,N_2537);
nand U3390 (N_3390,N_2916,N_2595);
nor U3391 (N_3391,N_2701,N_2776);
nand U3392 (N_3392,N_2951,N_2717);
and U3393 (N_3393,N_2775,N_2640);
nand U3394 (N_3394,N_2767,N_2980);
and U3395 (N_3395,N_2811,N_2590);
xor U3396 (N_3396,N_2652,N_2569);
nand U3397 (N_3397,N_2608,N_2896);
nor U3398 (N_3398,N_2689,N_2637);
xor U3399 (N_3399,N_2650,N_2643);
or U3400 (N_3400,N_2522,N_2940);
nand U3401 (N_3401,N_2643,N_2661);
or U3402 (N_3402,N_2624,N_2890);
xnor U3403 (N_3403,N_2610,N_2598);
and U3404 (N_3404,N_2533,N_2750);
or U3405 (N_3405,N_2737,N_2557);
or U3406 (N_3406,N_2781,N_2634);
and U3407 (N_3407,N_2911,N_2728);
and U3408 (N_3408,N_2701,N_2868);
and U3409 (N_3409,N_2623,N_2819);
nand U3410 (N_3410,N_2911,N_2625);
and U3411 (N_3411,N_2746,N_2910);
nand U3412 (N_3412,N_2811,N_2893);
xnor U3413 (N_3413,N_2715,N_2901);
and U3414 (N_3414,N_2775,N_2540);
nor U3415 (N_3415,N_2574,N_2703);
or U3416 (N_3416,N_2867,N_2595);
and U3417 (N_3417,N_2738,N_2994);
nand U3418 (N_3418,N_2646,N_2909);
xor U3419 (N_3419,N_2819,N_2974);
nor U3420 (N_3420,N_2604,N_2838);
nand U3421 (N_3421,N_2554,N_2531);
nand U3422 (N_3422,N_2743,N_2786);
xnor U3423 (N_3423,N_2851,N_2973);
nor U3424 (N_3424,N_2529,N_2877);
nand U3425 (N_3425,N_2879,N_2821);
nor U3426 (N_3426,N_2590,N_2544);
and U3427 (N_3427,N_2551,N_2764);
nor U3428 (N_3428,N_2931,N_2994);
and U3429 (N_3429,N_2617,N_2751);
or U3430 (N_3430,N_2500,N_2692);
and U3431 (N_3431,N_2784,N_2840);
or U3432 (N_3432,N_2896,N_2966);
nor U3433 (N_3433,N_2639,N_2610);
and U3434 (N_3434,N_2671,N_2985);
xor U3435 (N_3435,N_2714,N_2716);
and U3436 (N_3436,N_2844,N_2917);
and U3437 (N_3437,N_2608,N_2651);
and U3438 (N_3438,N_2907,N_2593);
or U3439 (N_3439,N_2890,N_2759);
nor U3440 (N_3440,N_2980,N_2930);
nor U3441 (N_3441,N_2753,N_2896);
nor U3442 (N_3442,N_2574,N_2722);
and U3443 (N_3443,N_2686,N_2819);
nand U3444 (N_3444,N_2934,N_2722);
xor U3445 (N_3445,N_2821,N_2622);
and U3446 (N_3446,N_2994,N_2923);
and U3447 (N_3447,N_2950,N_2645);
or U3448 (N_3448,N_2735,N_2832);
nor U3449 (N_3449,N_2845,N_2604);
and U3450 (N_3450,N_2824,N_2735);
and U3451 (N_3451,N_2593,N_2990);
xor U3452 (N_3452,N_2637,N_2997);
nand U3453 (N_3453,N_2933,N_2652);
nor U3454 (N_3454,N_2559,N_2669);
xor U3455 (N_3455,N_2732,N_2769);
and U3456 (N_3456,N_2782,N_2832);
or U3457 (N_3457,N_2757,N_2945);
xnor U3458 (N_3458,N_2977,N_2706);
nor U3459 (N_3459,N_2794,N_2799);
nor U3460 (N_3460,N_2756,N_2518);
nand U3461 (N_3461,N_2815,N_2940);
nand U3462 (N_3462,N_2903,N_2526);
or U3463 (N_3463,N_2535,N_2785);
xor U3464 (N_3464,N_2927,N_2633);
xnor U3465 (N_3465,N_2744,N_2985);
and U3466 (N_3466,N_2662,N_2564);
nand U3467 (N_3467,N_2958,N_2845);
or U3468 (N_3468,N_2818,N_2714);
or U3469 (N_3469,N_2713,N_2878);
xor U3470 (N_3470,N_2553,N_2901);
and U3471 (N_3471,N_2913,N_2663);
nand U3472 (N_3472,N_2929,N_2717);
nor U3473 (N_3473,N_2778,N_2700);
nand U3474 (N_3474,N_2638,N_2796);
xnor U3475 (N_3475,N_2934,N_2988);
nor U3476 (N_3476,N_2589,N_2755);
nor U3477 (N_3477,N_2512,N_2757);
or U3478 (N_3478,N_2513,N_2812);
and U3479 (N_3479,N_2582,N_2681);
or U3480 (N_3480,N_2890,N_2567);
xnor U3481 (N_3481,N_2946,N_2827);
nor U3482 (N_3482,N_2515,N_2844);
nand U3483 (N_3483,N_2955,N_2613);
and U3484 (N_3484,N_2604,N_2950);
nor U3485 (N_3485,N_2585,N_2751);
nor U3486 (N_3486,N_2694,N_2735);
nor U3487 (N_3487,N_2565,N_2502);
nor U3488 (N_3488,N_2662,N_2840);
nand U3489 (N_3489,N_2594,N_2913);
and U3490 (N_3490,N_2798,N_2938);
or U3491 (N_3491,N_2783,N_2714);
nor U3492 (N_3492,N_2642,N_2908);
or U3493 (N_3493,N_2677,N_2932);
and U3494 (N_3494,N_2637,N_2977);
nor U3495 (N_3495,N_2945,N_2635);
nand U3496 (N_3496,N_2786,N_2594);
xor U3497 (N_3497,N_2652,N_2727);
or U3498 (N_3498,N_2502,N_2880);
or U3499 (N_3499,N_2590,N_2626);
nor U3500 (N_3500,N_3077,N_3062);
nand U3501 (N_3501,N_3485,N_3020);
xor U3502 (N_3502,N_3185,N_3309);
nand U3503 (N_3503,N_3172,N_3432);
and U3504 (N_3504,N_3425,N_3001);
xnor U3505 (N_3505,N_3434,N_3035);
xor U3506 (N_3506,N_3312,N_3021);
nor U3507 (N_3507,N_3481,N_3064);
and U3508 (N_3508,N_3043,N_3073);
and U3509 (N_3509,N_3294,N_3359);
or U3510 (N_3510,N_3013,N_3322);
xnor U3511 (N_3511,N_3166,N_3347);
xnor U3512 (N_3512,N_3007,N_3205);
xnor U3513 (N_3513,N_3125,N_3213);
and U3514 (N_3514,N_3230,N_3232);
and U3515 (N_3515,N_3228,N_3423);
or U3516 (N_3516,N_3149,N_3463);
and U3517 (N_3517,N_3492,N_3006);
or U3518 (N_3518,N_3300,N_3250);
or U3519 (N_3519,N_3406,N_3473);
and U3520 (N_3520,N_3333,N_3157);
nor U3521 (N_3521,N_3163,N_3272);
nand U3522 (N_3522,N_3118,N_3199);
nor U3523 (N_3523,N_3459,N_3256);
or U3524 (N_3524,N_3382,N_3072);
nor U3525 (N_3525,N_3321,N_3109);
xor U3526 (N_3526,N_3115,N_3107);
xor U3527 (N_3527,N_3191,N_3193);
xnor U3528 (N_3528,N_3451,N_3048);
nand U3529 (N_3529,N_3237,N_3045);
and U3530 (N_3530,N_3236,N_3344);
nor U3531 (N_3531,N_3208,N_3132);
nor U3532 (N_3532,N_3354,N_3489);
xnor U3533 (N_3533,N_3366,N_3116);
xor U3534 (N_3534,N_3084,N_3245);
xnor U3535 (N_3535,N_3260,N_3327);
nor U3536 (N_3536,N_3337,N_3097);
and U3537 (N_3537,N_3170,N_3197);
or U3538 (N_3538,N_3217,N_3202);
nor U3539 (N_3539,N_3352,N_3470);
or U3540 (N_3540,N_3238,N_3144);
and U3541 (N_3541,N_3449,N_3285);
and U3542 (N_3542,N_3355,N_3464);
xor U3543 (N_3543,N_3324,N_3437);
nor U3544 (N_3544,N_3117,N_3283);
xnor U3545 (N_3545,N_3365,N_3036);
and U3546 (N_3546,N_3046,N_3054);
xor U3547 (N_3547,N_3000,N_3494);
xor U3548 (N_3548,N_3016,N_3305);
xor U3549 (N_3549,N_3303,N_3334);
and U3550 (N_3550,N_3094,N_3204);
nand U3551 (N_3551,N_3279,N_3291);
nor U3552 (N_3552,N_3152,N_3075);
or U3553 (N_3553,N_3474,N_3251);
nand U3554 (N_3554,N_3158,N_3289);
nand U3555 (N_3555,N_3402,N_3362);
or U3556 (N_3556,N_3393,N_3058);
nor U3557 (N_3557,N_3374,N_3074);
and U3558 (N_3558,N_3477,N_3031);
and U3559 (N_3559,N_3153,N_3141);
or U3560 (N_3560,N_3188,N_3219);
nand U3561 (N_3561,N_3379,N_3468);
nor U3562 (N_3562,N_3318,N_3323);
nor U3563 (N_3563,N_3056,N_3039);
xnor U3564 (N_3564,N_3241,N_3346);
or U3565 (N_3565,N_3174,N_3326);
and U3566 (N_3566,N_3395,N_3435);
nand U3567 (N_3567,N_3431,N_3348);
nand U3568 (N_3568,N_3335,N_3308);
nor U3569 (N_3569,N_3438,N_3079);
nor U3570 (N_3570,N_3415,N_3055);
and U3571 (N_3571,N_3159,N_3288);
and U3572 (N_3572,N_3221,N_3223);
and U3573 (N_3573,N_3028,N_3088);
or U3574 (N_3574,N_3037,N_3201);
xnor U3575 (N_3575,N_3195,N_3310);
xnor U3576 (N_3576,N_3194,N_3081);
and U3577 (N_3577,N_3102,N_3375);
nor U3578 (N_3578,N_3212,N_3218);
nand U3579 (N_3579,N_3082,N_3178);
and U3580 (N_3580,N_3340,N_3063);
nand U3581 (N_3581,N_3397,N_3248);
nand U3582 (N_3582,N_3286,N_3096);
and U3583 (N_3583,N_3461,N_3014);
xnor U3584 (N_3584,N_3325,N_3413);
or U3585 (N_3585,N_3167,N_3025);
nor U3586 (N_3586,N_3436,N_3122);
xor U3587 (N_3587,N_3311,N_3295);
nand U3588 (N_3588,N_3076,N_3069);
xnor U3589 (N_3589,N_3380,N_3403);
nor U3590 (N_3590,N_3343,N_3098);
xnor U3591 (N_3591,N_3146,N_3095);
nand U3592 (N_3592,N_3239,N_3426);
nor U3593 (N_3593,N_3130,N_3314);
or U3594 (N_3594,N_3227,N_3086);
nor U3595 (N_3595,N_3244,N_3261);
or U3596 (N_3596,N_3008,N_3377);
or U3597 (N_3597,N_3392,N_3255);
or U3598 (N_3598,N_3078,N_3369);
or U3599 (N_3599,N_3089,N_3487);
and U3600 (N_3600,N_3262,N_3042);
or U3601 (N_3601,N_3259,N_3113);
xnor U3602 (N_3602,N_3090,N_3421);
nand U3603 (N_3603,N_3498,N_3067);
nand U3604 (N_3604,N_3383,N_3091);
nor U3605 (N_3605,N_3401,N_3015);
xor U3606 (N_3606,N_3371,N_3472);
nor U3607 (N_3607,N_3004,N_3277);
nor U3608 (N_3608,N_3411,N_3271);
or U3609 (N_3609,N_3351,N_3247);
nand U3610 (N_3610,N_3111,N_3475);
nor U3611 (N_3611,N_3229,N_3356);
xnor U3612 (N_3612,N_3011,N_3243);
nand U3613 (N_3613,N_3126,N_3386);
and U3614 (N_3614,N_3302,N_3336);
nor U3615 (N_3615,N_3137,N_3496);
or U3616 (N_3616,N_3452,N_3206);
nor U3617 (N_3617,N_3161,N_3427);
or U3618 (N_3618,N_3190,N_3198);
nand U3619 (N_3619,N_3129,N_3160);
nand U3620 (N_3620,N_3209,N_3136);
xnor U3621 (N_3621,N_3495,N_3032);
nor U3622 (N_3622,N_3071,N_3417);
xor U3623 (N_3623,N_3368,N_3215);
and U3624 (N_3624,N_3155,N_3430);
nand U3625 (N_3625,N_3350,N_3026);
nand U3626 (N_3626,N_3278,N_3376);
xnor U3627 (N_3627,N_3499,N_3273);
nor U3628 (N_3628,N_3292,N_3252);
or U3629 (N_3629,N_3372,N_3328);
nor U3630 (N_3630,N_3341,N_3342);
nand U3631 (N_3631,N_3154,N_3164);
nand U3632 (N_3632,N_3070,N_3454);
nand U3633 (N_3633,N_3460,N_3304);
and U3634 (N_3634,N_3287,N_3384);
nor U3635 (N_3635,N_3225,N_3192);
nand U3636 (N_3636,N_3038,N_3106);
and U3637 (N_3637,N_3447,N_3444);
or U3638 (N_3638,N_3274,N_3398);
nor U3639 (N_3639,N_3246,N_3400);
xnor U3640 (N_3640,N_3222,N_3133);
nor U3641 (N_3641,N_3234,N_3316);
or U3642 (N_3642,N_3009,N_3183);
nand U3643 (N_3643,N_3265,N_3490);
nor U3644 (N_3644,N_3023,N_3235);
xor U3645 (N_3645,N_3105,N_3150);
and U3646 (N_3646,N_3266,N_3066);
nand U3647 (N_3647,N_3207,N_3173);
and U3648 (N_3648,N_3442,N_3177);
or U3649 (N_3649,N_3012,N_3339);
nor U3650 (N_3650,N_3297,N_3405);
xor U3651 (N_3651,N_3301,N_3242);
or U3652 (N_3652,N_3491,N_3162);
xnor U3653 (N_3653,N_3329,N_3019);
or U3654 (N_3654,N_3493,N_3175);
or U3655 (N_3655,N_3138,N_3299);
nand U3656 (N_3656,N_3214,N_3093);
nand U3657 (N_3657,N_3226,N_3358);
and U3658 (N_3658,N_3044,N_3453);
xor U3659 (N_3659,N_3134,N_3349);
xnor U3660 (N_3660,N_3186,N_3257);
xor U3661 (N_3661,N_3361,N_3331);
and U3662 (N_3662,N_3387,N_3254);
nor U3663 (N_3663,N_3357,N_3414);
xor U3664 (N_3664,N_3378,N_3433);
xor U3665 (N_3665,N_3180,N_3099);
and U3666 (N_3666,N_3267,N_3418);
nor U3667 (N_3667,N_3410,N_3027);
xnor U3668 (N_3668,N_3142,N_3441);
xor U3669 (N_3669,N_3263,N_3030);
nor U3670 (N_3670,N_3282,N_3087);
or U3671 (N_3671,N_3168,N_3047);
and U3672 (N_3672,N_3385,N_3497);
xnor U3673 (N_3673,N_3345,N_3332);
or U3674 (N_3674,N_3184,N_3367);
or U3675 (N_3675,N_3315,N_3484);
or U3676 (N_3676,N_3196,N_3049);
nor U3677 (N_3677,N_3145,N_3462);
and U3678 (N_3678,N_3258,N_3440);
or U3679 (N_3679,N_3253,N_3085);
xnor U3680 (N_3680,N_3276,N_3059);
or U3681 (N_3681,N_3017,N_3060);
or U3682 (N_3682,N_3083,N_3156);
nor U3683 (N_3683,N_3370,N_3317);
and U3684 (N_3684,N_3033,N_3293);
or U3685 (N_3685,N_3419,N_3306);
nor U3686 (N_3686,N_3388,N_3373);
and U3687 (N_3687,N_3139,N_3108);
xor U3688 (N_3688,N_3050,N_3381);
and U3689 (N_3689,N_3429,N_3466);
and U3690 (N_3690,N_3284,N_3412);
nor U3691 (N_3691,N_3231,N_3068);
xnor U3692 (N_3692,N_3439,N_3456);
nor U3693 (N_3693,N_3220,N_3280);
xor U3694 (N_3694,N_3135,N_3101);
xnor U3695 (N_3695,N_3147,N_3005);
xor U3696 (N_3696,N_3364,N_3320);
and U3697 (N_3697,N_3034,N_3269);
xor U3698 (N_3698,N_3128,N_3446);
nor U3699 (N_3699,N_3457,N_3471);
or U3700 (N_3700,N_3171,N_3458);
and U3701 (N_3701,N_3298,N_3399);
nor U3702 (N_3702,N_3053,N_3169);
or U3703 (N_3703,N_3482,N_3182);
xnor U3704 (N_3704,N_3022,N_3396);
nand U3705 (N_3705,N_3103,N_3124);
or U3706 (N_3706,N_3408,N_3181);
or U3707 (N_3707,N_3420,N_3151);
xnor U3708 (N_3708,N_3313,N_3448);
nor U3709 (N_3709,N_3469,N_3216);
or U3710 (N_3710,N_3424,N_3203);
and U3711 (N_3711,N_3330,N_3140);
xnor U3712 (N_3712,N_3065,N_3428);
and U3713 (N_3713,N_3479,N_3409);
xnor U3714 (N_3714,N_3394,N_3176);
and U3715 (N_3715,N_3391,N_3003);
nand U3716 (N_3716,N_3120,N_3480);
or U3717 (N_3717,N_3040,N_3467);
nor U3718 (N_3718,N_3143,N_3240);
xnor U3719 (N_3719,N_3264,N_3057);
or U3720 (N_3720,N_3390,N_3029);
nand U3721 (N_3721,N_3363,N_3131);
nor U3722 (N_3722,N_3112,N_3478);
xor U3723 (N_3723,N_3224,N_3445);
nor U3724 (N_3724,N_3148,N_3407);
nor U3725 (N_3725,N_3052,N_3307);
nor U3726 (N_3726,N_3486,N_3002);
xor U3727 (N_3727,N_3092,N_3443);
nand U3728 (N_3728,N_3114,N_3483);
xor U3729 (N_3729,N_3249,N_3121);
nor U3730 (N_3730,N_3123,N_3100);
or U3731 (N_3731,N_3465,N_3281);
and U3732 (N_3732,N_3275,N_3189);
or U3733 (N_3733,N_3422,N_3450);
nand U3734 (N_3734,N_3290,N_3187);
or U3735 (N_3735,N_3051,N_3389);
and U3736 (N_3736,N_3455,N_3080);
nand U3737 (N_3737,N_3268,N_3110);
or U3738 (N_3738,N_3270,N_3296);
nor U3739 (N_3739,N_3338,N_3200);
xnor U3740 (N_3740,N_3010,N_3319);
or U3741 (N_3741,N_3061,N_3024);
nand U3742 (N_3742,N_3404,N_3476);
and U3743 (N_3743,N_3360,N_3416);
nor U3744 (N_3744,N_3488,N_3127);
and U3745 (N_3745,N_3211,N_3119);
and U3746 (N_3746,N_3104,N_3165);
and U3747 (N_3747,N_3018,N_3233);
or U3748 (N_3748,N_3041,N_3179);
and U3749 (N_3749,N_3353,N_3210);
or U3750 (N_3750,N_3119,N_3057);
xnor U3751 (N_3751,N_3242,N_3166);
and U3752 (N_3752,N_3073,N_3356);
or U3753 (N_3753,N_3154,N_3045);
or U3754 (N_3754,N_3105,N_3318);
or U3755 (N_3755,N_3244,N_3169);
xnor U3756 (N_3756,N_3457,N_3396);
or U3757 (N_3757,N_3021,N_3150);
and U3758 (N_3758,N_3301,N_3041);
nor U3759 (N_3759,N_3066,N_3238);
nor U3760 (N_3760,N_3019,N_3154);
or U3761 (N_3761,N_3415,N_3234);
and U3762 (N_3762,N_3041,N_3346);
or U3763 (N_3763,N_3126,N_3012);
nor U3764 (N_3764,N_3292,N_3058);
nor U3765 (N_3765,N_3098,N_3042);
nor U3766 (N_3766,N_3009,N_3479);
and U3767 (N_3767,N_3294,N_3103);
xor U3768 (N_3768,N_3269,N_3498);
nor U3769 (N_3769,N_3008,N_3068);
or U3770 (N_3770,N_3023,N_3362);
xor U3771 (N_3771,N_3457,N_3164);
and U3772 (N_3772,N_3375,N_3221);
xor U3773 (N_3773,N_3446,N_3068);
xor U3774 (N_3774,N_3171,N_3204);
nand U3775 (N_3775,N_3301,N_3262);
and U3776 (N_3776,N_3263,N_3035);
nor U3777 (N_3777,N_3253,N_3040);
nor U3778 (N_3778,N_3166,N_3100);
and U3779 (N_3779,N_3307,N_3433);
xnor U3780 (N_3780,N_3496,N_3353);
nor U3781 (N_3781,N_3459,N_3029);
and U3782 (N_3782,N_3019,N_3457);
xor U3783 (N_3783,N_3056,N_3127);
nor U3784 (N_3784,N_3445,N_3337);
and U3785 (N_3785,N_3070,N_3049);
nand U3786 (N_3786,N_3015,N_3407);
and U3787 (N_3787,N_3299,N_3408);
and U3788 (N_3788,N_3016,N_3062);
and U3789 (N_3789,N_3319,N_3015);
nor U3790 (N_3790,N_3308,N_3253);
or U3791 (N_3791,N_3480,N_3059);
nand U3792 (N_3792,N_3422,N_3101);
or U3793 (N_3793,N_3018,N_3340);
and U3794 (N_3794,N_3269,N_3264);
and U3795 (N_3795,N_3305,N_3252);
xnor U3796 (N_3796,N_3376,N_3486);
or U3797 (N_3797,N_3306,N_3149);
or U3798 (N_3798,N_3003,N_3364);
and U3799 (N_3799,N_3159,N_3293);
nor U3800 (N_3800,N_3034,N_3294);
or U3801 (N_3801,N_3261,N_3487);
or U3802 (N_3802,N_3055,N_3137);
nand U3803 (N_3803,N_3162,N_3347);
and U3804 (N_3804,N_3426,N_3110);
nand U3805 (N_3805,N_3165,N_3384);
and U3806 (N_3806,N_3046,N_3156);
xnor U3807 (N_3807,N_3032,N_3253);
and U3808 (N_3808,N_3324,N_3090);
nand U3809 (N_3809,N_3443,N_3378);
nand U3810 (N_3810,N_3068,N_3434);
or U3811 (N_3811,N_3311,N_3455);
xnor U3812 (N_3812,N_3352,N_3395);
nor U3813 (N_3813,N_3120,N_3425);
or U3814 (N_3814,N_3006,N_3281);
xnor U3815 (N_3815,N_3335,N_3376);
xor U3816 (N_3816,N_3004,N_3328);
or U3817 (N_3817,N_3412,N_3455);
xor U3818 (N_3818,N_3256,N_3233);
nand U3819 (N_3819,N_3092,N_3097);
and U3820 (N_3820,N_3444,N_3146);
nand U3821 (N_3821,N_3427,N_3293);
and U3822 (N_3822,N_3118,N_3223);
nand U3823 (N_3823,N_3111,N_3224);
nor U3824 (N_3824,N_3218,N_3214);
nor U3825 (N_3825,N_3407,N_3362);
xor U3826 (N_3826,N_3153,N_3103);
xnor U3827 (N_3827,N_3216,N_3410);
xnor U3828 (N_3828,N_3381,N_3479);
nor U3829 (N_3829,N_3405,N_3343);
nor U3830 (N_3830,N_3264,N_3205);
xnor U3831 (N_3831,N_3416,N_3194);
xor U3832 (N_3832,N_3066,N_3120);
xor U3833 (N_3833,N_3333,N_3210);
nand U3834 (N_3834,N_3041,N_3078);
xnor U3835 (N_3835,N_3187,N_3031);
and U3836 (N_3836,N_3024,N_3169);
or U3837 (N_3837,N_3442,N_3352);
and U3838 (N_3838,N_3031,N_3275);
nor U3839 (N_3839,N_3448,N_3328);
or U3840 (N_3840,N_3296,N_3308);
or U3841 (N_3841,N_3394,N_3253);
or U3842 (N_3842,N_3488,N_3182);
or U3843 (N_3843,N_3339,N_3006);
nor U3844 (N_3844,N_3160,N_3315);
and U3845 (N_3845,N_3073,N_3089);
or U3846 (N_3846,N_3369,N_3116);
or U3847 (N_3847,N_3278,N_3035);
nor U3848 (N_3848,N_3114,N_3039);
nand U3849 (N_3849,N_3100,N_3410);
nand U3850 (N_3850,N_3371,N_3179);
and U3851 (N_3851,N_3353,N_3228);
xor U3852 (N_3852,N_3031,N_3200);
nand U3853 (N_3853,N_3330,N_3403);
or U3854 (N_3854,N_3147,N_3131);
nor U3855 (N_3855,N_3233,N_3279);
nand U3856 (N_3856,N_3070,N_3123);
xnor U3857 (N_3857,N_3381,N_3104);
nand U3858 (N_3858,N_3132,N_3111);
nand U3859 (N_3859,N_3313,N_3210);
nor U3860 (N_3860,N_3026,N_3223);
and U3861 (N_3861,N_3139,N_3441);
or U3862 (N_3862,N_3381,N_3436);
nand U3863 (N_3863,N_3099,N_3332);
or U3864 (N_3864,N_3251,N_3440);
xnor U3865 (N_3865,N_3335,N_3439);
or U3866 (N_3866,N_3430,N_3336);
xor U3867 (N_3867,N_3123,N_3187);
or U3868 (N_3868,N_3450,N_3211);
nor U3869 (N_3869,N_3357,N_3101);
nand U3870 (N_3870,N_3125,N_3463);
nand U3871 (N_3871,N_3353,N_3124);
or U3872 (N_3872,N_3283,N_3131);
and U3873 (N_3873,N_3234,N_3097);
nand U3874 (N_3874,N_3361,N_3422);
nor U3875 (N_3875,N_3160,N_3224);
nand U3876 (N_3876,N_3036,N_3127);
nor U3877 (N_3877,N_3364,N_3396);
or U3878 (N_3878,N_3287,N_3045);
or U3879 (N_3879,N_3211,N_3453);
or U3880 (N_3880,N_3035,N_3119);
xor U3881 (N_3881,N_3286,N_3038);
xor U3882 (N_3882,N_3270,N_3004);
xnor U3883 (N_3883,N_3011,N_3228);
or U3884 (N_3884,N_3176,N_3400);
nand U3885 (N_3885,N_3077,N_3333);
or U3886 (N_3886,N_3452,N_3073);
and U3887 (N_3887,N_3136,N_3212);
nor U3888 (N_3888,N_3003,N_3257);
nor U3889 (N_3889,N_3144,N_3374);
nand U3890 (N_3890,N_3305,N_3275);
and U3891 (N_3891,N_3147,N_3251);
nor U3892 (N_3892,N_3182,N_3163);
xnor U3893 (N_3893,N_3389,N_3306);
and U3894 (N_3894,N_3010,N_3485);
nand U3895 (N_3895,N_3228,N_3471);
and U3896 (N_3896,N_3485,N_3139);
nor U3897 (N_3897,N_3011,N_3203);
nand U3898 (N_3898,N_3433,N_3011);
or U3899 (N_3899,N_3081,N_3488);
nand U3900 (N_3900,N_3225,N_3337);
or U3901 (N_3901,N_3378,N_3406);
nor U3902 (N_3902,N_3201,N_3465);
xor U3903 (N_3903,N_3426,N_3309);
or U3904 (N_3904,N_3222,N_3048);
nor U3905 (N_3905,N_3484,N_3331);
or U3906 (N_3906,N_3361,N_3239);
xnor U3907 (N_3907,N_3023,N_3020);
xor U3908 (N_3908,N_3374,N_3010);
nand U3909 (N_3909,N_3261,N_3181);
or U3910 (N_3910,N_3483,N_3216);
and U3911 (N_3911,N_3438,N_3138);
nor U3912 (N_3912,N_3424,N_3011);
xor U3913 (N_3913,N_3044,N_3067);
xor U3914 (N_3914,N_3434,N_3232);
nand U3915 (N_3915,N_3097,N_3057);
nand U3916 (N_3916,N_3193,N_3218);
nor U3917 (N_3917,N_3420,N_3208);
or U3918 (N_3918,N_3266,N_3481);
and U3919 (N_3919,N_3463,N_3270);
xor U3920 (N_3920,N_3287,N_3376);
and U3921 (N_3921,N_3319,N_3380);
or U3922 (N_3922,N_3239,N_3079);
nor U3923 (N_3923,N_3131,N_3340);
and U3924 (N_3924,N_3348,N_3352);
nand U3925 (N_3925,N_3378,N_3485);
xor U3926 (N_3926,N_3244,N_3083);
and U3927 (N_3927,N_3456,N_3341);
or U3928 (N_3928,N_3292,N_3340);
and U3929 (N_3929,N_3126,N_3023);
xnor U3930 (N_3930,N_3480,N_3263);
nand U3931 (N_3931,N_3266,N_3408);
or U3932 (N_3932,N_3307,N_3442);
xnor U3933 (N_3933,N_3288,N_3371);
or U3934 (N_3934,N_3361,N_3207);
and U3935 (N_3935,N_3477,N_3418);
xor U3936 (N_3936,N_3497,N_3300);
and U3937 (N_3937,N_3319,N_3007);
and U3938 (N_3938,N_3218,N_3172);
nand U3939 (N_3939,N_3197,N_3123);
and U3940 (N_3940,N_3401,N_3210);
xnor U3941 (N_3941,N_3417,N_3360);
or U3942 (N_3942,N_3421,N_3108);
nand U3943 (N_3943,N_3161,N_3127);
and U3944 (N_3944,N_3290,N_3055);
or U3945 (N_3945,N_3078,N_3429);
xor U3946 (N_3946,N_3332,N_3014);
or U3947 (N_3947,N_3004,N_3183);
and U3948 (N_3948,N_3284,N_3323);
nor U3949 (N_3949,N_3368,N_3127);
nand U3950 (N_3950,N_3374,N_3418);
or U3951 (N_3951,N_3326,N_3243);
nor U3952 (N_3952,N_3163,N_3248);
and U3953 (N_3953,N_3295,N_3240);
nand U3954 (N_3954,N_3496,N_3393);
xor U3955 (N_3955,N_3452,N_3287);
nand U3956 (N_3956,N_3143,N_3321);
xor U3957 (N_3957,N_3200,N_3394);
xnor U3958 (N_3958,N_3129,N_3005);
and U3959 (N_3959,N_3476,N_3040);
nand U3960 (N_3960,N_3084,N_3221);
or U3961 (N_3961,N_3088,N_3150);
xor U3962 (N_3962,N_3215,N_3378);
and U3963 (N_3963,N_3383,N_3273);
xor U3964 (N_3964,N_3299,N_3083);
and U3965 (N_3965,N_3457,N_3392);
nor U3966 (N_3966,N_3204,N_3035);
xor U3967 (N_3967,N_3386,N_3141);
xnor U3968 (N_3968,N_3252,N_3014);
and U3969 (N_3969,N_3175,N_3159);
and U3970 (N_3970,N_3413,N_3362);
or U3971 (N_3971,N_3487,N_3399);
and U3972 (N_3972,N_3193,N_3123);
or U3973 (N_3973,N_3193,N_3249);
nand U3974 (N_3974,N_3336,N_3444);
nand U3975 (N_3975,N_3008,N_3481);
nand U3976 (N_3976,N_3215,N_3454);
or U3977 (N_3977,N_3311,N_3478);
nand U3978 (N_3978,N_3196,N_3279);
nand U3979 (N_3979,N_3135,N_3028);
nand U3980 (N_3980,N_3458,N_3424);
nor U3981 (N_3981,N_3155,N_3471);
xor U3982 (N_3982,N_3105,N_3457);
nor U3983 (N_3983,N_3223,N_3455);
nor U3984 (N_3984,N_3482,N_3032);
or U3985 (N_3985,N_3398,N_3071);
and U3986 (N_3986,N_3373,N_3249);
nor U3987 (N_3987,N_3127,N_3042);
xor U3988 (N_3988,N_3452,N_3375);
and U3989 (N_3989,N_3129,N_3376);
or U3990 (N_3990,N_3344,N_3086);
or U3991 (N_3991,N_3492,N_3430);
nor U3992 (N_3992,N_3329,N_3239);
or U3993 (N_3993,N_3496,N_3155);
or U3994 (N_3994,N_3094,N_3244);
xnor U3995 (N_3995,N_3135,N_3232);
nor U3996 (N_3996,N_3371,N_3172);
nand U3997 (N_3997,N_3214,N_3113);
or U3998 (N_3998,N_3386,N_3199);
nand U3999 (N_3999,N_3226,N_3144);
nand U4000 (N_4000,N_3775,N_3789);
and U4001 (N_4001,N_3574,N_3701);
and U4002 (N_4002,N_3704,N_3793);
or U4003 (N_4003,N_3761,N_3950);
xnor U4004 (N_4004,N_3845,N_3999);
and U4005 (N_4005,N_3519,N_3549);
nor U4006 (N_4006,N_3912,N_3843);
xor U4007 (N_4007,N_3740,N_3550);
or U4008 (N_4008,N_3933,N_3865);
nand U4009 (N_4009,N_3997,N_3665);
or U4010 (N_4010,N_3504,N_3615);
and U4011 (N_4011,N_3828,N_3813);
and U4012 (N_4012,N_3600,N_3962);
or U4013 (N_4013,N_3895,N_3893);
nor U4014 (N_4014,N_3899,N_3710);
and U4015 (N_4015,N_3898,N_3564);
nand U4016 (N_4016,N_3544,N_3526);
or U4017 (N_4017,N_3919,N_3726);
xor U4018 (N_4018,N_3973,N_3667);
xor U4019 (N_4019,N_3802,N_3623);
and U4020 (N_4020,N_3513,N_3786);
nand U4021 (N_4021,N_3599,N_3931);
nor U4022 (N_4022,N_3588,N_3668);
xnor U4023 (N_4023,N_3800,N_3760);
nor U4024 (N_4024,N_3986,N_3712);
nor U4025 (N_4025,N_3993,N_3757);
nand U4026 (N_4026,N_3691,N_3830);
nor U4027 (N_4027,N_3706,N_3971);
and U4028 (N_4028,N_3792,N_3988);
nand U4029 (N_4029,N_3685,N_3984);
and U4030 (N_4030,N_3774,N_3658);
and U4031 (N_4031,N_3829,N_3539);
or U4032 (N_4032,N_3769,N_3812);
xnor U4033 (N_4033,N_3578,N_3776);
or U4034 (N_4034,N_3814,N_3671);
xor U4035 (N_4035,N_3705,N_3683);
and U4036 (N_4036,N_3916,N_3906);
and U4037 (N_4037,N_3958,N_3889);
xor U4038 (N_4038,N_3690,N_3503);
nor U4039 (N_4039,N_3649,N_3921);
and U4040 (N_4040,N_3815,N_3888);
nand U4041 (N_4041,N_3556,N_3720);
or U4042 (N_4042,N_3577,N_3585);
nand U4043 (N_4043,N_3531,N_3907);
xnor U4044 (N_4044,N_3863,N_3532);
and U4045 (N_4045,N_3927,N_3978);
nor U4046 (N_4046,N_3651,N_3887);
and U4047 (N_4047,N_3542,N_3969);
and U4048 (N_4048,N_3631,N_3902);
nor U4049 (N_4049,N_3954,N_3892);
or U4050 (N_4050,N_3590,N_3678);
nand U4051 (N_4051,N_3976,N_3809);
nand U4052 (N_4052,N_3963,N_3537);
and U4053 (N_4053,N_3557,N_3834);
and U4054 (N_4054,N_3891,N_3900);
nor U4055 (N_4055,N_3525,N_3764);
nand U4056 (N_4056,N_3729,N_3838);
xnor U4057 (N_4057,N_3894,N_3995);
nor U4058 (N_4058,N_3872,N_3570);
xor U4059 (N_4059,N_3832,N_3553);
nand U4060 (N_4060,N_3536,N_3647);
or U4061 (N_4061,N_3998,N_3979);
and U4062 (N_4062,N_3660,N_3929);
nand U4063 (N_4063,N_3846,N_3604);
nand U4064 (N_4064,N_3853,N_3591);
nor U4065 (N_4065,N_3538,N_3878);
or U4066 (N_4066,N_3696,N_3836);
or U4067 (N_4067,N_3505,N_3896);
xor U4068 (N_4068,N_3567,N_3662);
or U4069 (N_4069,N_3733,N_3635);
nand U4070 (N_4070,N_3746,N_3805);
and U4071 (N_4071,N_3956,N_3871);
nor U4072 (N_4072,N_3583,N_3960);
nand U4073 (N_4073,N_3653,N_3937);
xnor U4074 (N_4074,N_3822,N_3932);
xor U4075 (N_4075,N_3571,N_3890);
nor U4076 (N_4076,N_3692,N_3796);
nand U4077 (N_4077,N_3780,N_3918);
or U4078 (N_4078,N_3881,N_3844);
and U4079 (N_4079,N_3713,N_3753);
and U4080 (N_4080,N_3940,N_3610);
or U4081 (N_4081,N_3632,N_3755);
or U4082 (N_4082,N_3679,N_3548);
and U4083 (N_4083,N_3695,N_3811);
nand U4084 (N_4084,N_3731,N_3910);
nand U4085 (N_4085,N_3687,N_3595);
and U4086 (N_4086,N_3861,N_3628);
nor U4087 (N_4087,N_3707,N_3598);
and U4088 (N_4088,N_3512,N_3520);
and U4089 (N_4089,N_3914,N_3763);
and U4090 (N_4090,N_3586,N_3752);
or U4091 (N_4091,N_3930,N_3742);
and U4092 (N_4092,N_3938,N_3766);
and U4093 (N_4093,N_3990,N_3642);
xnor U4094 (N_4094,N_3747,N_3873);
nand U4095 (N_4095,N_3573,N_3510);
and U4096 (N_4096,N_3854,N_3566);
nand U4097 (N_4097,N_3529,N_3939);
and U4098 (N_4098,N_3735,N_3905);
and U4099 (N_4099,N_3522,N_3677);
nor U4100 (N_4100,N_3517,N_3945);
nor U4101 (N_4101,N_3655,N_3778);
or U4102 (N_4102,N_3868,N_3736);
xnor U4103 (N_4103,N_3797,N_3622);
and U4104 (N_4104,N_3975,N_3739);
or U4105 (N_4105,N_3597,N_3639);
and U4106 (N_4106,N_3967,N_3611);
and U4107 (N_4107,N_3850,N_3772);
or U4108 (N_4108,N_3546,N_3580);
xor U4109 (N_4109,N_3547,N_3527);
nand U4110 (N_4110,N_3782,N_3637);
nand U4111 (N_4111,N_3788,N_3502);
and U4112 (N_4112,N_3727,N_3841);
or U4113 (N_4113,N_3784,N_3652);
and U4114 (N_4114,N_3922,N_3987);
nor U4115 (N_4115,N_3816,N_3605);
xor U4116 (N_4116,N_3565,N_3661);
nand U4117 (N_4117,N_3837,N_3749);
and U4118 (N_4118,N_3882,N_3773);
nor U4119 (N_4119,N_3709,N_3810);
xnor U4120 (N_4120,N_3614,N_3911);
or U4121 (N_4121,N_3982,N_3768);
xor U4122 (N_4122,N_3646,N_3582);
nor U4123 (N_4123,N_3901,N_3756);
and U4124 (N_4124,N_3924,N_3869);
nor U4125 (N_4125,N_3804,N_3974);
nor U4126 (N_4126,N_3762,N_3823);
nor U4127 (N_4127,N_3783,N_3636);
nor U4128 (N_4128,N_3886,N_3857);
and U4129 (N_4129,N_3721,N_3750);
and U4130 (N_4130,N_3554,N_3920);
xnor U4131 (N_4131,N_3790,N_3851);
xor U4132 (N_4132,N_3877,N_3684);
or U4133 (N_4133,N_3942,N_3584);
nor U4134 (N_4134,N_3926,N_3657);
nand U4135 (N_4135,N_3983,N_3759);
xnor U4136 (N_4136,N_3659,N_3785);
or U4137 (N_4137,N_3620,N_3618);
or U4138 (N_4138,N_3608,N_3957);
nand U4139 (N_4139,N_3880,N_3514);
and U4140 (N_4140,N_3533,N_3501);
or U4141 (N_4141,N_3612,N_3737);
nor U4142 (N_4142,N_3825,N_3540);
nor U4143 (N_4143,N_3745,N_3682);
nand U4144 (N_4144,N_3860,N_3650);
or U4145 (N_4145,N_3708,N_3643);
or U4146 (N_4146,N_3627,N_3791);
nand U4147 (N_4147,N_3603,N_3725);
and U4148 (N_4148,N_3619,N_3609);
nor U4149 (N_4149,N_3594,N_3732);
and U4150 (N_4150,N_3511,N_3852);
xnor U4151 (N_4151,N_3738,N_3915);
and U4152 (N_4152,N_3728,N_3961);
nor U4153 (N_4153,N_3601,N_3833);
and U4154 (N_4154,N_3716,N_3876);
nor U4155 (N_4155,N_3848,N_3644);
nand U4156 (N_4156,N_3944,N_3581);
and U4157 (N_4157,N_3593,N_3719);
nand U4158 (N_4158,N_3913,N_3941);
and U4159 (N_4159,N_3909,N_3681);
xor U4160 (N_4160,N_3903,N_3858);
or U4161 (N_4161,N_3528,N_3779);
xnor U4162 (N_4162,N_3686,N_3640);
nand U4163 (N_4163,N_3697,N_3748);
or U4164 (N_4164,N_3641,N_3630);
xor U4165 (N_4165,N_3718,N_3568);
or U4166 (N_4166,N_3981,N_3934);
and U4167 (N_4167,N_3569,N_3948);
nor U4168 (N_4168,N_3664,N_3508);
xor U4169 (N_4169,N_3606,N_3558);
nor U4170 (N_4170,N_3827,N_3625);
and U4171 (N_4171,N_3806,N_3935);
or U4172 (N_4172,N_3607,N_3803);
or U4173 (N_4173,N_3648,N_3840);
nor U4174 (N_4174,N_3777,N_3572);
or U4175 (N_4175,N_3798,N_3801);
xnor U4176 (N_4176,N_3817,N_3980);
nand U4177 (N_4177,N_3953,N_3855);
or U4178 (N_4178,N_3885,N_3771);
nand U4179 (N_4179,N_3949,N_3579);
or U4180 (N_4180,N_3821,N_3613);
and U4181 (N_4181,N_3518,N_3835);
nand U4182 (N_4182,N_3964,N_3996);
nand U4183 (N_4183,N_3589,N_3543);
and U4184 (N_4184,N_3820,N_3879);
nor U4185 (N_4185,N_3730,N_3500);
or U4186 (N_4186,N_3856,N_3634);
xor U4187 (N_4187,N_3535,N_3952);
nand U4188 (N_4188,N_3521,N_3758);
or U4189 (N_4189,N_3884,N_3951);
xor U4190 (N_4190,N_3781,N_3754);
nand U4191 (N_4191,N_3819,N_3663);
or U4192 (N_4192,N_3711,N_3917);
or U4193 (N_4193,N_3616,N_3698);
or U4194 (N_4194,N_3559,N_3562);
nor U4195 (N_4195,N_3859,N_3847);
or U4196 (N_4196,N_3770,N_3626);
nor U4197 (N_4197,N_3946,N_3693);
nand U4198 (N_4198,N_3509,N_3734);
nand U4199 (N_4199,N_3507,N_3966);
or U4200 (N_4200,N_3875,N_3994);
and U4201 (N_4201,N_3824,N_3575);
xor U4202 (N_4202,N_3751,N_3831);
and U4203 (N_4203,N_3767,N_3743);
nor U4204 (N_4204,N_3638,N_3675);
and U4205 (N_4205,N_3723,N_3702);
nand U4206 (N_4206,N_3670,N_3959);
or U4207 (N_4207,N_3596,N_3965);
nor U4208 (N_4208,N_3674,N_3799);
nand U4209 (N_4209,N_3936,N_3807);
nor U4210 (N_4210,N_3794,N_3666);
and U4211 (N_4211,N_3883,N_3870);
and U4212 (N_4212,N_3842,N_3688);
and U4213 (N_4213,N_3699,N_3560);
and U4214 (N_4214,N_3795,N_3724);
and U4215 (N_4215,N_3587,N_3977);
or U4216 (N_4216,N_3516,N_3592);
and U4217 (N_4217,N_3867,N_3633);
nand U4218 (N_4218,N_3862,N_3629);
nor U4219 (N_4219,N_3617,N_3694);
nor U4220 (N_4220,N_3530,N_3656);
nor U4221 (N_4221,N_3808,N_3555);
or U4222 (N_4222,N_3897,N_3992);
nor U4223 (N_4223,N_3839,N_3714);
and U4224 (N_4224,N_3700,N_3654);
xnor U4225 (N_4225,N_3904,N_3703);
and U4226 (N_4226,N_3506,N_3715);
xor U4227 (N_4227,N_3645,N_3561);
xnor U4228 (N_4228,N_3722,N_3524);
and U4229 (N_4229,N_3908,N_3947);
and U4230 (N_4230,N_3943,N_3744);
or U4231 (N_4231,N_3576,N_3989);
nor U4232 (N_4232,N_3968,N_3563);
xnor U4233 (N_4233,N_3874,N_3669);
xnor U4234 (N_4234,N_3923,N_3673);
or U4235 (N_4235,N_3545,N_3925);
xnor U4236 (N_4236,N_3864,N_3972);
nand U4237 (N_4237,N_3717,N_3866);
nor U4238 (N_4238,N_3534,N_3787);
nor U4239 (N_4239,N_3741,N_3689);
or U4240 (N_4240,N_3985,N_3818);
and U4241 (N_4241,N_3765,N_3541);
xnor U4242 (N_4242,N_3680,N_3849);
xor U4243 (N_4243,N_3602,N_3676);
nor U4244 (N_4244,N_3955,N_3928);
and U4245 (N_4245,N_3552,N_3826);
and U4246 (N_4246,N_3551,N_3970);
nand U4247 (N_4247,N_3621,N_3515);
nor U4248 (N_4248,N_3991,N_3624);
nand U4249 (N_4249,N_3523,N_3672);
and U4250 (N_4250,N_3635,N_3798);
nor U4251 (N_4251,N_3871,N_3918);
xor U4252 (N_4252,N_3903,N_3521);
nor U4253 (N_4253,N_3822,N_3757);
nor U4254 (N_4254,N_3857,N_3939);
nor U4255 (N_4255,N_3723,N_3758);
and U4256 (N_4256,N_3504,N_3941);
xor U4257 (N_4257,N_3683,N_3527);
xor U4258 (N_4258,N_3950,N_3990);
nand U4259 (N_4259,N_3561,N_3662);
nand U4260 (N_4260,N_3525,N_3856);
or U4261 (N_4261,N_3635,N_3769);
or U4262 (N_4262,N_3974,N_3655);
and U4263 (N_4263,N_3755,N_3816);
and U4264 (N_4264,N_3764,N_3726);
xnor U4265 (N_4265,N_3676,N_3554);
xnor U4266 (N_4266,N_3884,N_3964);
nor U4267 (N_4267,N_3726,N_3745);
and U4268 (N_4268,N_3635,N_3744);
or U4269 (N_4269,N_3785,N_3884);
nand U4270 (N_4270,N_3859,N_3965);
nor U4271 (N_4271,N_3561,N_3569);
and U4272 (N_4272,N_3659,N_3594);
and U4273 (N_4273,N_3771,N_3689);
xnor U4274 (N_4274,N_3824,N_3967);
nor U4275 (N_4275,N_3975,N_3979);
nor U4276 (N_4276,N_3808,N_3568);
nor U4277 (N_4277,N_3823,N_3500);
and U4278 (N_4278,N_3660,N_3882);
nand U4279 (N_4279,N_3692,N_3915);
or U4280 (N_4280,N_3798,N_3628);
or U4281 (N_4281,N_3960,N_3589);
and U4282 (N_4282,N_3571,N_3670);
nor U4283 (N_4283,N_3795,N_3654);
or U4284 (N_4284,N_3586,N_3843);
and U4285 (N_4285,N_3776,N_3716);
nand U4286 (N_4286,N_3703,N_3722);
or U4287 (N_4287,N_3584,N_3674);
nor U4288 (N_4288,N_3800,N_3593);
nand U4289 (N_4289,N_3556,N_3788);
or U4290 (N_4290,N_3918,N_3526);
nand U4291 (N_4291,N_3770,N_3528);
or U4292 (N_4292,N_3665,N_3577);
or U4293 (N_4293,N_3565,N_3703);
or U4294 (N_4294,N_3666,N_3935);
xnor U4295 (N_4295,N_3700,N_3935);
xor U4296 (N_4296,N_3560,N_3847);
nand U4297 (N_4297,N_3690,N_3954);
or U4298 (N_4298,N_3713,N_3606);
nor U4299 (N_4299,N_3787,N_3899);
nand U4300 (N_4300,N_3613,N_3522);
xor U4301 (N_4301,N_3715,N_3545);
nand U4302 (N_4302,N_3780,N_3531);
or U4303 (N_4303,N_3597,N_3771);
nor U4304 (N_4304,N_3912,N_3898);
nor U4305 (N_4305,N_3917,N_3934);
nand U4306 (N_4306,N_3637,N_3821);
and U4307 (N_4307,N_3752,N_3714);
xor U4308 (N_4308,N_3676,N_3927);
or U4309 (N_4309,N_3961,N_3812);
nor U4310 (N_4310,N_3711,N_3977);
or U4311 (N_4311,N_3893,N_3707);
xnor U4312 (N_4312,N_3707,N_3953);
nor U4313 (N_4313,N_3891,N_3629);
nor U4314 (N_4314,N_3889,N_3909);
xor U4315 (N_4315,N_3765,N_3568);
or U4316 (N_4316,N_3869,N_3796);
nor U4317 (N_4317,N_3579,N_3500);
and U4318 (N_4318,N_3631,N_3789);
xnor U4319 (N_4319,N_3836,N_3733);
or U4320 (N_4320,N_3936,N_3529);
nand U4321 (N_4321,N_3823,N_3758);
nand U4322 (N_4322,N_3731,N_3502);
nand U4323 (N_4323,N_3993,N_3771);
and U4324 (N_4324,N_3838,N_3959);
nor U4325 (N_4325,N_3812,N_3931);
or U4326 (N_4326,N_3870,N_3844);
nor U4327 (N_4327,N_3856,N_3526);
xnor U4328 (N_4328,N_3799,N_3817);
and U4329 (N_4329,N_3752,N_3781);
or U4330 (N_4330,N_3559,N_3548);
and U4331 (N_4331,N_3604,N_3944);
and U4332 (N_4332,N_3830,N_3966);
nor U4333 (N_4333,N_3819,N_3662);
and U4334 (N_4334,N_3974,N_3648);
and U4335 (N_4335,N_3852,N_3810);
and U4336 (N_4336,N_3661,N_3636);
and U4337 (N_4337,N_3878,N_3644);
xnor U4338 (N_4338,N_3793,N_3766);
xnor U4339 (N_4339,N_3997,N_3722);
nand U4340 (N_4340,N_3817,N_3660);
nor U4341 (N_4341,N_3754,N_3626);
or U4342 (N_4342,N_3580,N_3679);
nand U4343 (N_4343,N_3905,N_3677);
nor U4344 (N_4344,N_3668,N_3889);
or U4345 (N_4345,N_3553,N_3978);
and U4346 (N_4346,N_3752,N_3918);
nand U4347 (N_4347,N_3895,N_3905);
xor U4348 (N_4348,N_3753,N_3729);
nor U4349 (N_4349,N_3832,N_3651);
nor U4350 (N_4350,N_3841,N_3902);
or U4351 (N_4351,N_3817,N_3935);
and U4352 (N_4352,N_3913,N_3519);
and U4353 (N_4353,N_3809,N_3587);
nand U4354 (N_4354,N_3639,N_3548);
xor U4355 (N_4355,N_3672,N_3928);
nand U4356 (N_4356,N_3970,N_3516);
xnor U4357 (N_4357,N_3583,N_3829);
or U4358 (N_4358,N_3894,N_3988);
nand U4359 (N_4359,N_3912,N_3944);
xor U4360 (N_4360,N_3878,N_3558);
and U4361 (N_4361,N_3827,N_3667);
nor U4362 (N_4362,N_3962,N_3621);
and U4363 (N_4363,N_3950,N_3957);
nand U4364 (N_4364,N_3636,N_3599);
nand U4365 (N_4365,N_3921,N_3769);
nor U4366 (N_4366,N_3888,N_3754);
or U4367 (N_4367,N_3910,N_3933);
nand U4368 (N_4368,N_3785,N_3787);
nand U4369 (N_4369,N_3634,N_3501);
and U4370 (N_4370,N_3612,N_3907);
nor U4371 (N_4371,N_3698,N_3542);
and U4372 (N_4372,N_3695,N_3682);
nand U4373 (N_4373,N_3800,N_3757);
xor U4374 (N_4374,N_3648,N_3897);
and U4375 (N_4375,N_3573,N_3762);
xnor U4376 (N_4376,N_3647,N_3563);
and U4377 (N_4377,N_3934,N_3928);
and U4378 (N_4378,N_3789,N_3843);
and U4379 (N_4379,N_3664,N_3996);
xor U4380 (N_4380,N_3890,N_3993);
or U4381 (N_4381,N_3803,N_3820);
xnor U4382 (N_4382,N_3574,N_3594);
xnor U4383 (N_4383,N_3952,N_3775);
xor U4384 (N_4384,N_3909,N_3928);
or U4385 (N_4385,N_3992,N_3913);
or U4386 (N_4386,N_3719,N_3675);
and U4387 (N_4387,N_3727,N_3700);
xor U4388 (N_4388,N_3533,N_3612);
nor U4389 (N_4389,N_3811,N_3622);
xor U4390 (N_4390,N_3838,N_3580);
nor U4391 (N_4391,N_3981,N_3612);
nand U4392 (N_4392,N_3659,N_3799);
or U4393 (N_4393,N_3725,N_3596);
xnor U4394 (N_4394,N_3803,N_3927);
xor U4395 (N_4395,N_3566,N_3659);
nand U4396 (N_4396,N_3802,N_3804);
nand U4397 (N_4397,N_3854,N_3515);
xor U4398 (N_4398,N_3625,N_3963);
or U4399 (N_4399,N_3522,N_3614);
nor U4400 (N_4400,N_3648,N_3822);
nand U4401 (N_4401,N_3516,N_3864);
nand U4402 (N_4402,N_3611,N_3951);
nand U4403 (N_4403,N_3706,N_3560);
nor U4404 (N_4404,N_3940,N_3545);
nand U4405 (N_4405,N_3626,N_3528);
xnor U4406 (N_4406,N_3648,N_3784);
nor U4407 (N_4407,N_3584,N_3995);
nand U4408 (N_4408,N_3967,N_3578);
xor U4409 (N_4409,N_3672,N_3706);
and U4410 (N_4410,N_3513,N_3796);
nand U4411 (N_4411,N_3560,N_3948);
nand U4412 (N_4412,N_3544,N_3647);
or U4413 (N_4413,N_3564,N_3933);
xnor U4414 (N_4414,N_3889,N_3552);
or U4415 (N_4415,N_3751,N_3665);
or U4416 (N_4416,N_3569,N_3936);
and U4417 (N_4417,N_3579,N_3613);
nor U4418 (N_4418,N_3742,N_3790);
xor U4419 (N_4419,N_3648,N_3935);
nor U4420 (N_4420,N_3782,N_3828);
nor U4421 (N_4421,N_3890,N_3808);
nor U4422 (N_4422,N_3927,N_3832);
or U4423 (N_4423,N_3679,N_3915);
or U4424 (N_4424,N_3554,N_3848);
or U4425 (N_4425,N_3709,N_3550);
or U4426 (N_4426,N_3703,N_3879);
and U4427 (N_4427,N_3655,N_3645);
or U4428 (N_4428,N_3854,N_3766);
nand U4429 (N_4429,N_3834,N_3859);
nor U4430 (N_4430,N_3630,N_3779);
and U4431 (N_4431,N_3808,N_3943);
and U4432 (N_4432,N_3639,N_3865);
or U4433 (N_4433,N_3813,N_3940);
nor U4434 (N_4434,N_3907,N_3953);
nor U4435 (N_4435,N_3595,N_3790);
xor U4436 (N_4436,N_3869,N_3870);
nor U4437 (N_4437,N_3816,N_3766);
or U4438 (N_4438,N_3652,N_3692);
and U4439 (N_4439,N_3782,N_3717);
or U4440 (N_4440,N_3706,N_3553);
nor U4441 (N_4441,N_3768,N_3939);
nand U4442 (N_4442,N_3831,N_3746);
nor U4443 (N_4443,N_3877,N_3695);
or U4444 (N_4444,N_3677,N_3850);
and U4445 (N_4445,N_3734,N_3524);
xor U4446 (N_4446,N_3526,N_3542);
and U4447 (N_4447,N_3706,N_3615);
and U4448 (N_4448,N_3897,N_3623);
nor U4449 (N_4449,N_3510,N_3803);
nand U4450 (N_4450,N_3740,N_3908);
or U4451 (N_4451,N_3857,N_3605);
or U4452 (N_4452,N_3702,N_3846);
and U4453 (N_4453,N_3614,N_3509);
nand U4454 (N_4454,N_3579,N_3618);
xor U4455 (N_4455,N_3871,N_3910);
or U4456 (N_4456,N_3743,N_3733);
nor U4457 (N_4457,N_3703,N_3724);
nor U4458 (N_4458,N_3812,N_3504);
nand U4459 (N_4459,N_3633,N_3708);
nand U4460 (N_4460,N_3585,N_3596);
or U4461 (N_4461,N_3944,N_3504);
nor U4462 (N_4462,N_3993,N_3901);
xnor U4463 (N_4463,N_3732,N_3517);
nor U4464 (N_4464,N_3544,N_3778);
xor U4465 (N_4465,N_3715,N_3741);
nand U4466 (N_4466,N_3869,N_3553);
xor U4467 (N_4467,N_3762,N_3686);
and U4468 (N_4468,N_3898,N_3600);
and U4469 (N_4469,N_3631,N_3767);
nand U4470 (N_4470,N_3549,N_3766);
or U4471 (N_4471,N_3992,N_3534);
nor U4472 (N_4472,N_3943,N_3964);
and U4473 (N_4473,N_3558,N_3910);
or U4474 (N_4474,N_3743,N_3996);
and U4475 (N_4475,N_3848,N_3624);
nand U4476 (N_4476,N_3684,N_3638);
xnor U4477 (N_4477,N_3633,N_3715);
nor U4478 (N_4478,N_3786,N_3632);
nor U4479 (N_4479,N_3649,N_3784);
nor U4480 (N_4480,N_3794,N_3945);
xnor U4481 (N_4481,N_3753,N_3925);
or U4482 (N_4482,N_3610,N_3816);
and U4483 (N_4483,N_3789,N_3999);
nor U4484 (N_4484,N_3588,N_3651);
nor U4485 (N_4485,N_3877,N_3937);
and U4486 (N_4486,N_3793,N_3727);
xor U4487 (N_4487,N_3722,N_3689);
xnor U4488 (N_4488,N_3540,N_3828);
and U4489 (N_4489,N_3772,N_3910);
and U4490 (N_4490,N_3754,N_3766);
nor U4491 (N_4491,N_3575,N_3741);
nand U4492 (N_4492,N_3513,N_3991);
xor U4493 (N_4493,N_3512,N_3655);
xnor U4494 (N_4494,N_3804,N_3787);
nand U4495 (N_4495,N_3637,N_3783);
or U4496 (N_4496,N_3587,N_3904);
nor U4497 (N_4497,N_3836,N_3762);
or U4498 (N_4498,N_3725,N_3867);
and U4499 (N_4499,N_3875,N_3714);
xor U4500 (N_4500,N_4343,N_4029);
xnor U4501 (N_4501,N_4072,N_4196);
and U4502 (N_4502,N_4168,N_4437);
or U4503 (N_4503,N_4497,N_4372);
and U4504 (N_4504,N_4291,N_4172);
or U4505 (N_4505,N_4231,N_4084);
and U4506 (N_4506,N_4401,N_4462);
nor U4507 (N_4507,N_4298,N_4346);
nor U4508 (N_4508,N_4481,N_4390);
and U4509 (N_4509,N_4123,N_4446);
nor U4510 (N_4510,N_4178,N_4070);
nand U4511 (N_4511,N_4017,N_4167);
nor U4512 (N_4512,N_4096,N_4485);
xor U4513 (N_4513,N_4301,N_4465);
xnor U4514 (N_4514,N_4133,N_4169);
or U4515 (N_4515,N_4214,N_4281);
or U4516 (N_4516,N_4366,N_4182);
xor U4517 (N_4517,N_4382,N_4201);
and U4518 (N_4518,N_4073,N_4449);
and U4519 (N_4519,N_4140,N_4049);
nand U4520 (N_4520,N_4012,N_4216);
xor U4521 (N_4521,N_4408,N_4082);
or U4522 (N_4522,N_4160,N_4180);
and U4523 (N_4523,N_4286,N_4130);
nor U4524 (N_4524,N_4177,N_4021);
nor U4525 (N_4525,N_4268,N_4228);
nor U4526 (N_4526,N_4314,N_4024);
xor U4527 (N_4527,N_4126,N_4436);
nor U4528 (N_4528,N_4238,N_4006);
nor U4529 (N_4529,N_4312,N_4109);
or U4530 (N_4530,N_4056,N_4272);
nand U4531 (N_4531,N_4174,N_4233);
and U4532 (N_4532,N_4015,N_4152);
nand U4533 (N_4533,N_4118,N_4209);
or U4534 (N_4534,N_4440,N_4198);
or U4535 (N_4535,N_4147,N_4033);
nor U4536 (N_4536,N_4184,N_4326);
nand U4537 (N_4537,N_4205,N_4125);
nor U4538 (N_4538,N_4302,N_4373);
nor U4539 (N_4539,N_4371,N_4085);
xor U4540 (N_4540,N_4392,N_4411);
nand U4541 (N_4541,N_4441,N_4075);
xnor U4542 (N_4542,N_4406,N_4034);
and U4543 (N_4543,N_4478,N_4250);
and U4544 (N_4544,N_4052,N_4031);
and U4545 (N_4545,N_4234,N_4431);
nor U4546 (N_4546,N_4428,N_4489);
or U4547 (N_4547,N_4087,N_4270);
xnor U4548 (N_4548,N_4499,N_4287);
nor U4549 (N_4549,N_4313,N_4309);
or U4550 (N_4550,N_4337,N_4300);
xnor U4551 (N_4551,N_4193,N_4142);
or U4552 (N_4552,N_4484,N_4289);
nor U4553 (N_4553,N_4374,N_4399);
xnor U4554 (N_4554,N_4212,N_4414);
nand U4555 (N_4555,N_4018,N_4044);
and U4556 (N_4556,N_4068,N_4080);
nand U4557 (N_4557,N_4252,N_4240);
xor U4558 (N_4558,N_4486,N_4099);
and U4559 (N_4559,N_4002,N_4463);
xnor U4560 (N_4560,N_4013,N_4415);
xor U4561 (N_4561,N_4375,N_4492);
xnor U4562 (N_4562,N_4304,N_4121);
nor U4563 (N_4563,N_4016,N_4466);
xnor U4564 (N_4564,N_4349,N_4139);
xnor U4565 (N_4565,N_4435,N_4190);
nand U4566 (N_4566,N_4275,N_4329);
xor U4567 (N_4567,N_4144,N_4066);
or U4568 (N_4568,N_4387,N_4135);
nor U4569 (N_4569,N_4469,N_4071);
xor U4570 (N_4570,N_4239,N_4086);
nor U4571 (N_4571,N_4091,N_4226);
xnor U4572 (N_4572,N_4053,N_4036);
nand U4573 (N_4573,N_4004,N_4307);
nor U4574 (N_4574,N_4403,N_4256);
xor U4575 (N_4575,N_4368,N_4297);
nand U4576 (N_4576,N_4379,N_4093);
or U4577 (N_4577,N_4124,N_4494);
nand U4578 (N_4578,N_4249,N_4248);
and U4579 (N_4579,N_4391,N_4227);
nand U4580 (N_4580,N_4456,N_4438);
xnor U4581 (N_4581,N_4305,N_4432);
xor U4582 (N_4582,N_4241,N_4213);
and U4583 (N_4583,N_4159,N_4251);
nor U4584 (N_4584,N_4204,N_4400);
xor U4585 (N_4585,N_4030,N_4100);
nor U4586 (N_4586,N_4477,N_4038);
nor U4587 (N_4587,N_4405,N_4311);
xor U4588 (N_4588,N_4334,N_4255);
nand U4589 (N_4589,N_4335,N_4430);
nor U4590 (N_4590,N_4330,N_4158);
or U4591 (N_4591,N_4134,N_4293);
nand U4592 (N_4592,N_4254,N_4377);
nor U4593 (N_4593,N_4257,N_4079);
xor U4594 (N_4594,N_4218,N_4151);
or U4595 (N_4595,N_4258,N_4360);
nor U4596 (N_4596,N_4129,N_4211);
nand U4597 (N_4597,N_4473,N_4064);
nor U4598 (N_4598,N_4023,N_4197);
xor U4599 (N_4599,N_4454,N_4367);
nand U4600 (N_4600,N_4331,N_4319);
xor U4601 (N_4601,N_4402,N_4057);
nor U4602 (N_4602,N_4146,N_4332);
xnor U4603 (N_4603,N_4318,N_4153);
nand U4604 (N_4604,N_4127,N_4076);
nor U4605 (N_4605,N_4232,N_4010);
or U4606 (N_4606,N_4092,N_4181);
or U4607 (N_4607,N_4183,N_4058);
nand U4608 (N_4608,N_4427,N_4242);
and U4609 (N_4609,N_4060,N_4453);
or U4610 (N_4610,N_4210,N_4026);
nor U4611 (N_4611,N_4221,N_4244);
xnor U4612 (N_4612,N_4479,N_4219);
and U4613 (N_4613,N_4264,N_4294);
xnor U4614 (N_4614,N_4316,N_4179);
nand U4615 (N_4615,N_4008,N_4320);
and U4616 (N_4616,N_4136,N_4116);
or U4617 (N_4617,N_4295,N_4199);
xor U4618 (N_4618,N_4452,N_4107);
xnor U4619 (N_4619,N_4222,N_4460);
or U4620 (N_4620,N_4342,N_4194);
nor U4621 (N_4621,N_4102,N_4202);
or U4622 (N_4622,N_4235,N_4271);
or U4623 (N_4623,N_4288,N_4020);
or U4624 (N_4624,N_4132,N_4365);
nor U4625 (N_4625,N_4154,N_4112);
xnor U4626 (N_4626,N_4354,N_4385);
nor U4627 (N_4627,N_4447,N_4325);
xnor U4628 (N_4628,N_4105,N_4110);
xor U4629 (N_4629,N_4364,N_4310);
nand U4630 (N_4630,N_4393,N_4128);
nand U4631 (N_4631,N_4333,N_4065);
and U4632 (N_4632,N_4359,N_4276);
xnor U4633 (N_4633,N_4472,N_4458);
nand U4634 (N_4634,N_4088,N_4009);
or U4635 (N_4635,N_4166,N_4412);
xor U4636 (N_4636,N_4113,N_4383);
or U4637 (N_4637,N_4117,N_4223);
nand U4638 (N_4638,N_4323,N_4046);
and U4639 (N_4639,N_4176,N_4426);
nand U4640 (N_4640,N_4439,N_4470);
nor U4641 (N_4641,N_4274,N_4344);
nor U4642 (N_4642,N_4069,N_4370);
and U4643 (N_4643,N_4050,N_4047);
or U4644 (N_4644,N_4421,N_4014);
or U4645 (N_4645,N_4119,N_4413);
or U4646 (N_4646,N_4417,N_4163);
and U4647 (N_4647,N_4040,N_4145);
xnor U4648 (N_4648,N_4042,N_4292);
xor U4649 (N_4649,N_4001,N_4137);
or U4650 (N_4650,N_4407,N_4488);
xnor U4651 (N_4651,N_4077,N_4162);
nand U4652 (N_4652,N_4103,N_4434);
and U4653 (N_4653,N_4063,N_4098);
or U4654 (N_4654,N_4220,N_4404);
xor U4655 (N_4655,N_4369,N_4165);
or U4656 (N_4656,N_4003,N_4261);
nor U4657 (N_4657,N_4253,N_4224);
nor U4658 (N_4658,N_4457,N_4245);
nand U4659 (N_4659,N_4269,N_4043);
nor U4660 (N_4660,N_4025,N_4280);
or U4661 (N_4661,N_4381,N_4173);
xor U4662 (N_4662,N_4247,N_4496);
nand U4663 (N_4663,N_4445,N_4206);
or U4664 (N_4664,N_4120,N_4186);
nand U4665 (N_4665,N_4322,N_4464);
nand U4666 (N_4666,N_4416,N_4078);
xor U4667 (N_4667,N_4161,N_4187);
nand U4668 (N_4668,N_4094,N_4171);
xnor U4669 (N_4669,N_4266,N_4083);
and U4670 (N_4670,N_4035,N_4418);
nor U4671 (N_4671,N_4263,N_4095);
nand U4672 (N_4672,N_4315,N_4471);
nor U4673 (N_4673,N_4422,N_4455);
xnor U4674 (N_4674,N_4000,N_4101);
xor U4675 (N_4675,N_4007,N_4037);
and U4676 (N_4676,N_4027,N_4157);
nand U4677 (N_4677,N_4350,N_4237);
xnor U4678 (N_4678,N_4389,N_4362);
xor U4679 (N_4679,N_4185,N_4208);
and U4680 (N_4680,N_4356,N_4019);
and U4681 (N_4681,N_4217,N_4459);
and U4682 (N_4682,N_4156,N_4131);
nor U4683 (N_4683,N_4476,N_4122);
and U4684 (N_4684,N_4376,N_4041);
or U4685 (N_4685,N_4203,N_4262);
nor U4686 (N_4686,N_4398,N_4150);
and U4687 (N_4687,N_4351,N_4032);
nand U4688 (N_4688,N_4143,N_4424);
or U4689 (N_4689,N_4207,N_4353);
xor U4690 (N_4690,N_4423,N_4409);
xnor U4691 (N_4691,N_4149,N_4429);
xor U4692 (N_4692,N_4467,N_4059);
xnor U4693 (N_4693,N_4442,N_4106);
xor U4694 (N_4694,N_4191,N_4277);
and U4695 (N_4695,N_4396,N_4074);
or U4696 (N_4696,N_4028,N_4327);
and U4697 (N_4697,N_4420,N_4444);
and U4698 (N_4698,N_4114,N_4200);
and U4699 (N_4699,N_4011,N_4067);
or U4700 (N_4700,N_4483,N_4246);
xor U4701 (N_4701,N_4243,N_4081);
nor U4702 (N_4702,N_4498,N_4317);
xnor U4703 (N_4703,N_4051,N_4055);
nand U4704 (N_4704,N_4397,N_4045);
or U4705 (N_4705,N_4491,N_4259);
nor U4706 (N_4706,N_4284,N_4474);
xnor U4707 (N_4707,N_4111,N_4090);
xor U4708 (N_4708,N_4410,N_4303);
nor U4709 (N_4709,N_4482,N_4361);
or U4710 (N_4710,N_4089,N_4290);
xor U4711 (N_4711,N_4054,N_4490);
nor U4712 (N_4712,N_4339,N_4148);
nor U4713 (N_4713,N_4062,N_4357);
and U4714 (N_4714,N_4475,N_4388);
nand U4715 (N_4715,N_4338,N_4487);
nor U4716 (N_4716,N_4495,N_4225);
xor U4717 (N_4717,N_4285,N_4425);
xor U4718 (N_4718,N_4321,N_4433);
nand U4719 (N_4719,N_4355,N_4155);
or U4720 (N_4720,N_4451,N_4363);
and U4721 (N_4721,N_4039,N_4005);
xnor U4722 (N_4722,N_4341,N_4308);
xnor U4723 (N_4723,N_4347,N_4282);
or U4724 (N_4724,N_4448,N_4022);
and U4725 (N_4725,N_4279,N_4278);
and U4726 (N_4726,N_4443,N_4358);
nor U4727 (N_4727,N_4192,N_4419);
and U4728 (N_4728,N_4189,N_4141);
and U4729 (N_4729,N_4493,N_4306);
or U4730 (N_4730,N_4097,N_4195);
nor U4731 (N_4731,N_4273,N_4384);
and U4732 (N_4732,N_4215,N_4115);
nand U4733 (N_4733,N_4104,N_4188);
xnor U4734 (N_4734,N_4061,N_4378);
or U4735 (N_4735,N_4352,N_4267);
xor U4736 (N_4736,N_4386,N_4138);
nand U4737 (N_4737,N_4345,N_4229);
and U4738 (N_4738,N_4299,N_4380);
or U4739 (N_4739,N_4164,N_4348);
and U4740 (N_4740,N_4328,N_4450);
xnor U4741 (N_4741,N_4260,N_4175);
nor U4742 (N_4742,N_4230,N_4394);
nor U4743 (N_4743,N_4324,N_4480);
nor U4744 (N_4744,N_4340,N_4283);
nand U4745 (N_4745,N_4236,N_4048);
or U4746 (N_4746,N_4108,N_4395);
xnor U4747 (N_4747,N_4468,N_4461);
nor U4748 (N_4748,N_4170,N_4265);
nor U4749 (N_4749,N_4336,N_4296);
or U4750 (N_4750,N_4255,N_4150);
nor U4751 (N_4751,N_4234,N_4150);
or U4752 (N_4752,N_4253,N_4110);
nor U4753 (N_4753,N_4402,N_4415);
nor U4754 (N_4754,N_4268,N_4492);
nand U4755 (N_4755,N_4463,N_4392);
or U4756 (N_4756,N_4141,N_4462);
nand U4757 (N_4757,N_4234,N_4220);
nor U4758 (N_4758,N_4426,N_4343);
nand U4759 (N_4759,N_4383,N_4205);
nand U4760 (N_4760,N_4009,N_4345);
nor U4761 (N_4761,N_4434,N_4305);
nand U4762 (N_4762,N_4108,N_4319);
nor U4763 (N_4763,N_4202,N_4412);
nand U4764 (N_4764,N_4497,N_4124);
nor U4765 (N_4765,N_4476,N_4181);
or U4766 (N_4766,N_4489,N_4242);
and U4767 (N_4767,N_4404,N_4357);
nor U4768 (N_4768,N_4413,N_4028);
and U4769 (N_4769,N_4353,N_4185);
or U4770 (N_4770,N_4125,N_4498);
xnor U4771 (N_4771,N_4304,N_4407);
xor U4772 (N_4772,N_4418,N_4112);
xnor U4773 (N_4773,N_4010,N_4270);
and U4774 (N_4774,N_4020,N_4129);
and U4775 (N_4775,N_4183,N_4052);
nand U4776 (N_4776,N_4160,N_4498);
or U4777 (N_4777,N_4096,N_4262);
nand U4778 (N_4778,N_4425,N_4300);
or U4779 (N_4779,N_4448,N_4085);
and U4780 (N_4780,N_4155,N_4318);
and U4781 (N_4781,N_4405,N_4453);
and U4782 (N_4782,N_4262,N_4234);
and U4783 (N_4783,N_4371,N_4275);
xor U4784 (N_4784,N_4180,N_4257);
and U4785 (N_4785,N_4336,N_4240);
and U4786 (N_4786,N_4144,N_4322);
xnor U4787 (N_4787,N_4061,N_4212);
nor U4788 (N_4788,N_4182,N_4300);
and U4789 (N_4789,N_4248,N_4340);
nor U4790 (N_4790,N_4260,N_4010);
nand U4791 (N_4791,N_4072,N_4458);
nor U4792 (N_4792,N_4055,N_4444);
or U4793 (N_4793,N_4380,N_4381);
and U4794 (N_4794,N_4380,N_4466);
or U4795 (N_4795,N_4159,N_4452);
xor U4796 (N_4796,N_4445,N_4226);
or U4797 (N_4797,N_4150,N_4304);
nand U4798 (N_4798,N_4246,N_4031);
or U4799 (N_4799,N_4280,N_4104);
or U4800 (N_4800,N_4090,N_4179);
or U4801 (N_4801,N_4244,N_4367);
nand U4802 (N_4802,N_4350,N_4157);
nor U4803 (N_4803,N_4384,N_4228);
xor U4804 (N_4804,N_4474,N_4022);
nand U4805 (N_4805,N_4206,N_4365);
xor U4806 (N_4806,N_4199,N_4108);
and U4807 (N_4807,N_4413,N_4272);
nor U4808 (N_4808,N_4272,N_4293);
and U4809 (N_4809,N_4385,N_4229);
nand U4810 (N_4810,N_4459,N_4051);
nor U4811 (N_4811,N_4387,N_4471);
nand U4812 (N_4812,N_4185,N_4398);
xnor U4813 (N_4813,N_4041,N_4055);
and U4814 (N_4814,N_4338,N_4339);
or U4815 (N_4815,N_4183,N_4015);
xor U4816 (N_4816,N_4445,N_4027);
nor U4817 (N_4817,N_4456,N_4296);
nor U4818 (N_4818,N_4037,N_4341);
nand U4819 (N_4819,N_4033,N_4362);
xnor U4820 (N_4820,N_4260,N_4380);
xnor U4821 (N_4821,N_4118,N_4370);
nand U4822 (N_4822,N_4415,N_4041);
nand U4823 (N_4823,N_4311,N_4468);
nor U4824 (N_4824,N_4467,N_4041);
nor U4825 (N_4825,N_4361,N_4212);
and U4826 (N_4826,N_4324,N_4342);
xnor U4827 (N_4827,N_4208,N_4299);
or U4828 (N_4828,N_4050,N_4208);
nor U4829 (N_4829,N_4208,N_4304);
and U4830 (N_4830,N_4457,N_4092);
nor U4831 (N_4831,N_4449,N_4433);
and U4832 (N_4832,N_4188,N_4204);
or U4833 (N_4833,N_4413,N_4072);
or U4834 (N_4834,N_4045,N_4139);
nand U4835 (N_4835,N_4277,N_4403);
and U4836 (N_4836,N_4240,N_4155);
or U4837 (N_4837,N_4301,N_4047);
or U4838 (N_4838,N_4155,N_4010);
nor U4839 (N_4839,N_4381,N_4458);
and U4840 (N_4840,N_4428,N_4372);
nand U4841 (N_4841,N_4252,N_4344);
or U4842 (N_4842,N_4474,N_4338);
nand U4843 (N_4843,N_4173,N_4114);
or U4844 (N_4844,N_4399,N_4411);
and U4845 (N_4845,N_4214,N_4288);
or U4846 (N_4846,N_4311,N_4258);
nor U4847 (N_4847,N_4228,N_4159);
xor U4848 (N_4848,N_4386,N_4369);
nor U4849 (N_4849,N_4495,N_4388);
or U4850 (N_4850,N_4451,N_4347);
nand U4851 (N_4851,N_4406,N_4440);
and U4852 (N_4852,N_4156,N_4388);
or U4853 (N_4853,N_4113,N_4406);
nand U4854 (N_4854,N_4240,N_4193);
or U4855 (N_4855,N_4139,N_4160);
or U4856 (N_4856,N_4279,N_4219);
nand U4857 (N_4857,N_4020,N_4257);
xnor U4858 (N_4858,N_4145,N_4407);
nand U4859 (N_4859,N_4095,N_4245);
or U4860 (N_4860,N_4184,N_4177);
nor U4861 (N_4861,N_4490,N_4442);
or U4862 (N_4862,N_4262,N_4114);
nor U4863 (N_4863,N_4207,N_4209);
xnor U4864 (N_4864,N_4007,N_4275);
nand U4865 (N_4865,N_4481,N_4098);
or U4866 (N_4866,N_4238,N_4246);
nand U4867 (N_4867,N_4268,N_4447);
nor U4868 (N_4868,N_4000,N_4191);
and U4869 (N_4869,N_4003,N_4100);
or U4870 (N_4870,N_4311,N_4413);
xnor U4871 (N_4871,N_4063,N_4435);
nand U4872 (N_4872,N_4478,N_4066);
nor U4873 (N_4873,N_4001,N_4010);
and U4874 (N_4874,N_4010,N_4011);
xor U4875 (N_4875,N_4330,N_4177);
nor U4876 (N_4876,N_4031,N_4245);
nand U4877 (N_4877,N_4355,N_4046);
nand U4878 (N_4878,N_4460,N_4406);
and U4879 (N_4879,N_4191,N_4267);
or U4880 (N_4880,N_4129,N_4297);
or U4881 (N_4881,N_4235,N_4076);
xnor U4882 (N_4882,N_4253,N_4171);
and U4883 (N_4883,N_4032,N_4293);
nand U4884 (N_4884,N_4360,N_4352);
xor U4885 (N_4885,N_4011,N_4480);
or U4886 (N_4886,N_4200,N_4357);
or U4887 (N_4887,N_4282,N_4467);
xnor U4888 (N_4888,N_4028,N_4080);
nand U4889 (N_4889,N_4157,N_4272);
xnor U4890 (N_4890,N_4477,N_4075);
and U4891 (N_4891,N_4260,N_4053);
nor U4892 (N_4892,N_4122,N_4447);
nand U4893 (N_4893,N_4409,N_4316);
or U4894 (N_4894,N_4176,N_4381);
nand U4895 (N_4895,N_4159,N_4047);
xnor U4896 (N_4896,N_4122,N_4220);
xnor U4897 (N_4897,N_4064,N_4113);
xor U4898 (N_4898,N_4315,N_4229);
nor U4899 (N_4899,N_4424,N_4227);
or U4900 (N_4900,N_4107,N_4458);
and U4901 (N_4901,N_4431,N_4025);
and U4902 (N_4902,N_4226,N_4099);
nor U4903 (N_4903,N_4039,N_4476);
xor U4904 (N_4904,N_4483,N_4275);
or U4905 (N_4905,N_4252,N_4169);
xor U4906 (N_4906,N_4310,N_4376);
xor U4907 (N_4907,N_4040,N_4292);
or U4908 (N_4908,N_4015,N_4139);
nand U4909 (N_4909,N_4302,N_4063);
or U4910 (N_4910,N_4327,N_4121);
nor U4911 (N_4911,N_4009,N_4272);
nand U4912 (N_4912,N_4339,N_4076);
or U4913 (N_4913,N_4377,N_4040);
or U4914 (N_4914,N_4109,N_4161);
nand U4915 (N_4915,N_4160,N_4269);
nor U4916 (N_4916,N_4130,N_4251);
nor U4917 (N_4917,N_4463,N_4480);
and U4918 (N_4918,N_4270,N_4083);
and U4919 (N_4919,N_4487,N_4171);
nor U4920 (N_4920,N_4369,N_4112);
and U4921 (N_4921,N_4030,N_4072);
nand U4922 (N_4922,N_4365,N_4457);
xor U4923 (N_4923,N_4347,N_4226);
or U4924 (N_4924,N_4111,N_4297);
nand U4925 (N_4925,N_4310,N_4351);
nor U4926 (N_4926,N_4156,N_4061);
or U4927 (N_4927,N_4206,N_4355);
and U4928 (N_4928,N_4138,N_4233);
and U4929 (N_4929,N_4038,N_4180);
and U4930 (N_4930,N_4333,N_4329);
nor U4931 (N_4931,N_4001,N_4330);
and U4932 (N_4932,N_4332,N_4468);
nand U4933 (N_4933,N_4291,N_4038);
nand U4934 (N_4934,N_4258,N_4126);
xnor U4935 (N_4935,N_4259,N_4056);
and U4936 (N_4936,N_4050,N_4427);
and U4937 (N_4937,N_4489,N_4184);
or U4938 (N_4938,N_4216,N_4011);
or U4939 (N_4939,N_4053,N_4377);
and U4940 (N_4940,N_4315,N_4425);
and U4941 (N_4941,N_4068,N_4181);
nand U4942 (N_4942,N_4339,N_4441);
and U4943 (N_4943,N_4366,N_4056);
and U4944 (N_4944,N_4382,N_4448);
nand U4945 (N_4945,N_4343,N_4011);
nand U4946 (N_4946,N_4310,N_4381);
or U4947 (N_4947,N_4311,N_4172);
nor U4948 (N_4948,N_4203,N_4197);
nand U4949 (N_4949,N_4470,N_4310);
nand U4950 (N_4950,N_4445,N_4362);
or U4951 (N_4951,N_4298,N_4011);
nor U4952 (N_4952,N_4274,N_4127);
or U4953 (N_4953,N_4294,N_4412);
nand U4954 (N_4954,N_4261,N_4343);
or U4955 (N_4955,N_4083,N_4427);
xor U4956 (N_4956,N_4367,N_4394);
xor U4957 (N_4957,N_4156,N_4367);
and U4958 (N_4958,N_4333,N_4366);
nor U4959 (N_4959,N_4189,N_4207);
xnor U4960 (N_4960,N_4262,N_4073);
or U4961 (N_4961,N_4474,N_4092);
or U4962 (N_4962,N_4276,N_4451);
nor U4963 (N_4963,N_4445,N_4114);
and U4964 (N_4964,N_4315,N_4396);
and U4965 (N_4965,N_4016,N_4006);
xnor U4966 (N_4966,N_4141,N_4264);
xnor U4967 (N_4967,N_4193,N_4339);
nand U4968 (N_4968,N_4174,N_4235);
and U4969 (N_4969,N_4235,N_4479);
nand U4970 (N_4970,N_4155,N_4287);
nor U4971 (N_4971,N_4471,N_4266);
or U4972 (N_4972,N_4074,N_4413);
xnor U4973 (N_4973,N_4339,N_4135);
and U4974 (N_4974,N_4084,N_4105);
and U4975 (N_4975,N_4490,N_4214);
and U4976 (N_4976,N_4433,N_4411);
nor U4977 (N_4977,N_4449,N_4023);
xnor U4978 (N_4978,N_4149,N_4217);
and U4979 (N_4979,N_4421,N_4131);
nor U4980 (N_4980,N_4032,N_4105);
nor U4981 (N_4981,N_4349,N_4404);
xor U4982 (N_4982,N_4140,N_4151);
and U4983 (N_4983,N_4347,N_4103);
nand U4984 (N_4984,N_4245,N_4187);
and U4985 (N_4985,N_4383,N_4286);
and U4986 (N_4986,N_4287,N_4070);
or U4987 (N_4987,N_4011,N_4238);
nand U4988 (N_4988,N_4424,N_4399);
nand U4989 (N_4989,N_4470,N_4215);
nor U4990 (N_4990,N_4091,N_4491);
nand U4991 (N_4991,N_4183,N_4218);
and U4992 (N_4992,N_4119,N_4198);
nor U4993 (N_4993,N_4498,N_4113);
xnor U4994 (N_4994,N_4338,N_4108);
nor U4995 (N_4995,N_4331,N_4378);
nand U4996 (N_4996,N_4187,N_4160);
and U4997 (N_4997,N_4229,N_4182);
nand U4998 (N_4998,N_4263,N_4437);
xor U4999 (N_4999,N_4428,N_4087);
xor U5000 (N_5000,N_4611,N_4658);
or U5001 (N_5001,N_4656,N_4731);
or U5002 (N_5002,N_4872,N_4883);
nand U5003 (N_5003,N_4616,N_4913);
nor U5004 (N_5004,N_4782,N_4725);
xor U5005 (N_5005,N_4528,N_4794);
nor U5006 (N_5006,N_4818,N_4605);
or U5007 (N_5007,N_4539,N_4683);
nand U5008 (N_5008,N_4881,N_4576);
xnor U5009 (N_5009,N_4541,N_4737);
nor U5010 (N_5010,N_4892,N_4595);
or U5011 (N_5011,N_4633,N_4618);
nor U5012 (N_5012,N_4695,N_4841);
nor U5013 (N_5013,N_4889,N_4918);
nand U5014 (N_5014,N_4977,N_4817);
or U5015 (N_5015,N_4857,N_4899);
xnor U5016 (N_5016,N_4575,N_4993);
nand U5017 (N_5017,N_4902,N_4740);
or U5018 (N_5018,N_4885,N_4769);
nand U5019 (N_5019,N_4504,N_4578);
nor U5020 (N_5020,N_4719,N_4558);
or U5021 (N_5021,N_4743,N_4998);
xnor U5022 (N_5022,N_4523,N_4583);
nand U5023 (N_5023,N_4750,N_4777);
nand U5024 (N_5024,N_4861,N_4820);
nor U5025 (N_5025,N_4712,N_4568);
nor U5026 (N_5026,N_4636,N_4515);
nor U5027 (N_5027,N_4707,N_4659);
nor U5028 (N_5028,N_4943,N_4842);
nand U5029 (N_5029,N_4718,N_4500);
xor U5030 (N_5030,N_4845,N_4688);
xnor U5031 (N_5031,N_4631,N_4660);
nand U5032 (N_5032,N_4796,N_4952);
nand U5033 (N_5033,N_4798,N_4766);
and U5034 (N_5034,N_4713,N_4741);
and U5035 (N_5035,N_4704,N_4646);
nand U5036 (N_5036,N_4623,N_4738);
or U5037 (N_5037,N_4942,N_4839);
or U5038 (N_5038,N_4599,N_4870);
nor U5039 (N_5039,N_4744,N_4603);
nand U5040 (N_5040,N_4856,N_4774);
nand U5041 (N_5041,N_4989,N_4812);
nor U5042 (N_5042,N_4877,N_4642);
xnor U5043 (N_5043,N_4852,N_4672);
xnor U5044 (N_5044,N_4544,N_4874);
nor U5045 (N_5045,N_4914,N_4823);
nor U5046 (N_5046,N_4795,N_4722);
nand U5047 (N_5047,N_4621,N_4501);
xnor U5048 (N_5048,N_4982,N_4530);
nor U5049 (N_5049,N_4521,N_4570);
and U5050 (N_5050,N_4553,N_4598);
or U5051 (N_5051,N_4994,N_4939);
xor U5052 (N_5052,N_4807,N_4559);
xnor U5053 (N_5053,N_4723,N_4549);
or U5054 (N_5054,N_4664,N_4630);
nor U5055 (N_5055,N_4536,N_4752);
nand U5056 (N_5056,N_4730,N_4832);
xnor U5057 (N_5057,N_4567,N_4503);
or U5058 (N_5058,N_4887,N_4655);
xor U5059 (N_5059,N_4555,N_4937);
nand U5060 (N_5060,N_4975,N_4565);
nor U5061 (N_5061,N_4510,N_4542);
or U5062 (N_5062,N_4779,N_4844);
and U5063 (N_5063,N_4591,N_4692);
and U5064 (N_5064,N_4703,N_4518);
nand U5065 (N_5065,N_4974,N_4619);
nor U5066 (N_5066,N_4825,N_4635);
nand U5067 (N_5067,N_4678,N_4761);
and U5068 (N_5068,N_4984,N_4961);
xor U5069 (N_5069,N_4965,N_4920);
nand U5070 (N_5070,N_4606,N_4934);
xnor U5071 (N_5071,N_4677,N_4617);
nor U5072 (N_5072,N_4764,N_4679);
or U5073 (N_5073,N_4905,N_4579);
and U5074 (N_5074,N_4944,N_4900);
and U5075 (N_5075,N_4760,N_4991);
nor U5076 (N_5076,N_4751,N_4897);
nand U5077 (N_5077,N_4732,N_4529);
nor U5078 (N_5078,N_4724,N_4551);
nand U5079 (N_5079,N_4929,N_4850);
nand U5080 (N_5080,N_4608,N_4875);
nor U5081 (N_5081,N_4627,N_4871);
and U5082 (N_5082,N_4600,N_4868);
xor U5083 (N_5083,N_4907,N_4711);
nor U5084 (N_5084,N_4853,N_4728);
nor U5085 (N_5085,N_4860,N_4886);
or U5086 (N_5086,N_4609,N_4690);
xnor U5087 (N_5087,N_4505,N_4949);
nor U5088 (N_5088,N_4569,N_4550);
nand U5089 (N_5089,N_4957,N_4896);
xnor U5090 (N_5090,N_4936,N_4654);
or U5091 (N_5091,N_4562,N_4894);
or U5092 (N_5092,N_4727,N_4950);
nand U5093 (N_5093,N_4921,N_4590);
or U5094 (N_5094,N_4806,N_4509);
and U5095 (N_5095,N_4720,N_4978);
or U5096 (N_5096,N_4815,N_4780);
or U5097 (N_5097,N_4849,N_4945);
nor U5098 (N_5098,N_4987,N_4924);
xnor U5099 (N_5099,N_4746,N_4891);
nor U5100 (N_5100,N_4747,N_4869);
xnor U5101 (N_5101,N_4745,N_4502);
xor U5102 (N_5102,N_4548,N_4773);
xor U5103 (N_5103,N_4916,N_4833);
nor U5104 (N_5104,N_4564,N_4634);
nand U5105 (N_5105,N_4863,N_4985);
nand U5106 (N_5106,N_4647,N_4622);
or U5107 (N_5107,N_4666,N_4753);
nand U5108 (N_5108,N_4763,N_4824);
nor U5109 (N_5109,N_4802,N_4652);
nor U5110 (N_5110,N_4847,N_4915);
nor U5111 (N_5111,N_4601,N_4586);
and U5112 (N_5112,N_4992,N_4888);
or U5113 (N_5113,N_4697,N_4629);
and U5114 (N_5114,N_4657,N_4685);
xor U5115 (N_5115,N_4514,N_4653);
and U5116 (N_5116,N_4986,N_4959);
or U5117 (N_5117,N_4814,N_4827);
nor U5118 (N_5118,N_4733,N_4904);
xnor U5119 (N_5119,N_4717,N_4917);
and U5120 (N_5120,N_4637,N_4572);
or U5121 (N_5121,N_4864,N_4604);
and U5122 (N_5122,N_4848,N_4787);
nor U5123 (N_5123,N_4947,N_4701);
nor U5124 (N_5124,N_4674,N_4784);
nor U5125 (N_5125,N_4808,N_4736);
nor U5126 (N_5126,N_4726,N_4835);
nand U5127 (N_5127,N_4734,N_4557);
nand U5128 (N_5128,N_4791,N_4826);
nand U5129 (N_5129,N_4762,N_4997);
nand U5130 (N_5130,N_4522,N_4527);
nand U5131 (N_5131,N_4585,N_4926);
and U5132 (N_5132,N_4946,N_4615);
xnor U5133 (N_5133,N_4644,N_4571);
nor U5134 (N_5134,N_4865,N_4516);
and U5135 (N_5135,N_4925,N_4940);
or U5136 (N_5136,N_4963,N_4687);
nand U5137 (N_5137,N_4577,N_4938);
or U5138 (N_5138,N_4797,N_4996);
and U5139 (N_5139,N_4547,N_4866);
and U5140 (N_5140,N_4691,N_4922);
xor U5141 (N_5141,N_4563,N_4816);
or U5142 (N_5142,N_4840,N_4748);
nand U5143 (N_5143,N_4681,N_4649);
nand U5144 (N_5144,N_4513,N_4771);
and U5145 (N_5145,N_4596,N_4698);
nand U5146 (N_5146,N_4830,N_4846);
and U5147 (N_5147,N_4828,N_4667);
and U5148 (N_5148,N_4638,N_4742);
nand U5149 (N_5149,N_4783,N_4676);
nor U5150 (N_5150,N_4620,N_4593);
xor U5151 (N_5151,N_4931,N_4836);
nor U5152 (N_5152,N_4757,N_4966);
nand U5153 (N_5153,N_4976,N_4507);
and U5154 (N_5154,N_4535,N_4715);
nand U5155 (N_5155,N_4822,N_4858);
nor U5156 (N_5156,N_4967,N_4765);
and U5157 (N_5157,N_4511,N_4910);
and U5158 (N_5158,N_4906,N_4767);
xnor U5159 (N_5159,N_4813,N_4506);
nand U5160 (N_5160,N_4758,N_4867);
and U5161 (N_5161,N_4809,N_4556);
nor U5162 (N_5162,N_4930,N_4702);
nand U5163 (N_5163,N_4793,N_4612);
and U5164 (N_5164,N_4970,N_4641);
and U5165 (N_5165,N_4948,N_4661);
or U5166 (N_5166,N_4573,N_4895);
and U5167 (N_5167,N_4545,N_4995);
or U5168 (N_5168,N_4680,N_4626);
nor U5169 (N_5169,N_4554,N_4819);
nand U5170 (N_5170,N_4706,N_4954);
xor U5171 (N_5171,N_4588,N_4582);
xor U5172 (N_5172,N_4756,N_4941);
and U5173 (N_5173,N_4537,N_4625);
nor U5174 (N_5174,N_4508,N_4810);
nor U5175 (N_5175,N_4804,N_4768);
nor U5176 (N_5176,N_4632,N_4968);
nand U5177 (N_5177,N_4911,N_4580);
xnor U5178 (N_5178,N_4800,N_4581);
xor U5179 (N_5179,N_4643,N_4855);
nand U5180 (N_5180,N_4532,N_4898);
nor U5181 (N_5181,N_4546,N_4755);
nand U5182 (N_5182,N_4587,N_4831);
nor U5183 (N_5183,N_4524,N_4973);
or U5184 (N_5184,N_4584,N_4958);
or U5185 (N_5185,N_4955,N_4531);
and U5186 (N_5186,N_4935,N_4517);
nor U5187 (N_5187,N_4933,N_4597);
and U5188 (N_5188,N_4801,N_4684);
nand U5189 (N_5189,N_4811,N_4624);
nor U5190 (N_5190,N_4613,N_4754);
nand U5191 (N_5191,N_4526,N_4893);
xnor U5192 (N_5192,N_4971,N_4969);
or U5193 (N_5193,N_4951,N_4979);
and U5194 (N_5194,N_4749,N_4790);
and U5195 (N_5195,N_4566,N_4928);
nand U5196 (N_5196,N_4650,N_4829);
or U5197 (N_5197,N_4610,N_4834);
nor U5198 (N_5198,N_4614,N_4540);
and U5199 (N_5199,N_4699,N_4909);
nor U5200 (N_5200,N_4901,N_4882);
and U5201 (N_5201,N_4594,N_4772);
and U5202 (N_5202,N_4923,N_4561);
nand U5203 (N_5203,N_4639,N_4805);
nand U5204 (N_5204,N_4686,N_4781);
or U5205 (N_5205,N_4775,N_4983);
or U5206 (N_5206,N_4729,N_4803);
or U5207 (N_5207,N_4838,N_4689);
nor U5208 (N_5208,N_4714,N_4880);
and U5209 (N_5209,N_4520,N_4721);
and U5210 (N_5210,N_4759,N_4962);
or U5211 (N_5211,N_4876,N_4675);
nor U5212 (N_5212,N_4552,N_4873);
or U5213 (N_5213,N_4673,N_4776);
or U5214 (N_5214,N_4533,N_4932);
or U5215 (N_5215,N_4927,N_4980);
nand U5216 (N_5216,N_4543,N_4696);
xnor U5217 (N_5217,N_4651,N_4878);
xnor U5218 (N_5218,N_4648,N_4972);
xor U5219 (N_5219,N_4525,N_4890);
or U5220 (N_5220,N_4710,N_4964);
or U5221 (N_5221,N_4859,N_4669);
nand U5222 (N_5222,N_4693,N_4988);
nand U5223 (N_5223,N_4960,N_4792);
and U5224 (N_5224,N_4709,N_4862);
nand U5225 (N_5225,N_4519,N_4837);
or U5226 (N_5226,N_4999,N_4682);
and U5227 (N_5227,N_4645,N_4879);
xnor U5228 (N_5228,N_4854,N_4602);
and U5229 (N_5229,N_4700,N_4534);
nor U5230 (N_5230,N_4739,N_4786);
nor U5231 (N_5231,N_4694,N_4851);
nor U5232 (N_5232,N_4785,N_4908);
or U5233 (N_5233,N_4663,N_4884);
nor U5234 (N_5234,N_4990,N_4640);
xnor U5235 (N_5235,N_4981,N_4607);
nor U5236 (N_5236,N_4799,N_4708);
nor U5237 (N_5237,N_4560,N_4770);
xor U5238 (N_5238,N_4670,N_4668);
nand U5239 (N_5239,N_4705,N_4716);
nor U5240 (N_5240,N_4789,N_4671);
xnor U5241 (N_5241,N_4778,N_4592);
xor U5242 (N_5242,N_4843,N_4821);
nor U5243 (N_5243,N_4574,N_4665);
xnor U5244 (N_5244,N_4788,N_4919);
nand U5245 (N_5245,N_4912,N_4956);
xor U5246 (N_5246,N_4538,N_4953);
and U5247 (N_5247,N_4589,N_4628);
and U5248 (N_5248,N_4662,N_4903);
and U5249 (N_5249,N_4735,N_4512);
nand U5250 (N_5250,N_4657,N_4970);
nand U5251 (N_5251,N_4790,N_4939);
nand U5252 (N_5252,N_4593,N_4687);
or U5253 (N_5253,N_4896,N_4698);
or U5254 (N_5254,N_4785,N_4682);
nor U5255 (N_5255,N_4821,N_4744);
and U5256 (N_5256,N_4771,N_4698);
xnor U5257 (N_5257,N_4923,N_4683);
xnor U5258 (N_5258,N_4908,N_4988);
or U5259 (N_5259,N_4776,N_4945);
and U5260 (N_5260,N_4533,N_4514);
nand U5261 (N_5261,N_4501,N_4750);
nand U5262 (N_5262,N_4753,N_4745);
nand U5263 (N_5263,N_4899,N_4867);
and U5264 (N_5264,N_4834,N_4578);
xor U5265 (N_5265,N_4800,N_4708);
and U5266 (N_5266,N_4735,N_4700);
nor U5267 (N_5267,N_4958,N_4734);
nor U5268 (N_5268,N_4942,N_4869);
or U5269 (N_5269,N_4722,N_4510);
nor U5270 (N_5270,N_4897,N_4724);
nor U5271 (N_5271,N_4795,N_4695);
nor U5272 (N_5272,N_4823,N_4638);
and U5273 (N_5273,N_4853,N_4714);
nor U5274 (N_5274,N_4694,N_4624);
xnor U5275 (N_5275,N_4991,N_4744);
xor U5276 (N_5276,N_4706,N_4753);
nor U5277 (N_5277,N_4777,N_4839);
xor U5278 (N_5278,N_4943,N_4590);
nor U5279 (N_5279,N_4543,N_4921);
nand U5280 (N_5280,N_4979,N_4506);
nand U5281 (N_5281,N_4850,N_4935);
or U5282 (N_5282,N_4693,N_4898);
or U5283 (N_5283,N_4509,N_4788);
xor U5284 (N_5284,N_4616,N_4954);
xor U5285 (N_5285,N_4689,N_4766);
nor U5286 (N_5286,N_4953,N_4505);
and U5287 (N_5287,N_4900,N_4511);
or U5288 (N_5288,N_4834,N_4660);
and U5289 (N_5289,N_4773,N_4966);
or U5290 (N_5290,N_4999,N_4843);
and U5291 (N_5291,N_4827,N_4900);
nor U5292 (N_5292,N_4644,N_4808);
and U5293 (N_5293,N_4685,N_4659);
and U5294 (N_5294,N_4722,N_4951);
and U5295 (N_5295,N_4977,N_4553);
or U5296 (N_5296,N_4693,N_4744);
nor U5297 (N_5297,N_4861,N_4598);
xor U5298 (N_5298,N_4568,N_4696);
or U5299 (N_5299,N_4866,N_4743);
nor U5300 (N_5300,N_4863,N_4778);
nor U5301 (N_5301,N_4980,N_4747);
xor U5302 (N_5302,N_4803,N_4776);
or U5303 (N_5303,N_4954,N_4516);
and U5304 (N_5304,N_4998,N_4832);
xor U5305 (N_5305,N_4673,N_4803);
xor U5306 (N_5306,N_4638,N_4910);
nand U5307 (N_5307,N_4793,N_4527);
and U5308 (N_5308,N_4819,N_4618);
nor U5309 (N_5309,N_4520,N_4828);
or U5310 (N_5310,N_4861,N_4910);
xnor U5311 (N_5311,N_4987,N_4909);
xnor U5312 (N_5312,N_4811,N_4521);
xnor U5313 (N_5313,N_4962,N_4978);
and U5314 (N_5314,N_4539,N_4525);
or U5315 (N_5315,N_4740,N_4916);
nor U5316 (N_5316,N_4962,N_4579);
or U5317 (N_5317,N_4794,N_4959);
xor U5318 (N_5318,N_4983,N_4955);
nor U5319 (N_5319,N_4783,N_4749);
and U5320 (N_5320,N_4880,N_4840);
nor U5321 (N_5321,N_4891,N_4973);
nor U5322 (N_5322,N_4951,N_4807);
xor U5323 (N_5323,N_4638,N_4547);
nand U5324 (N_5324,N_4652,N_4633);
xnor U5325 (N_5325,N_4856,N_4867);
or U5326 (N_5326,N_4754,N_4506);
nor U5327 (N_5327,N_4938,N_4967);
and U5328 (N_5328,N_4722,N_4995);
nand U5329 (N_5329,N_4731,N_4691);
nand U5330 (N_5330,N_4524,N_4848);
nor U5331 (N_5331,N_4532,N_4618);
nor U5332 (N_5332,N_4511,N_4860);
and U5333 (N_5333,N_4524,N_4855);
or U5334 (N_5334,N_4879,N_4527);
or U5335 (N_5335,N_4568,N_4987);
nor U5336 (N_5336,N_4837,N_4797);
and U5337 (N_5337,N_4837,N_4743);
xnor U5338 (N_5338,N_4550,N_4957);
nor U5339 (N_5339,N_4907,N_4729);
or U5340 (N_5340,N_4575,N_4823);
nand U5341 (N_5341,N_4740,N_4797);
xnor U5342 (N_5342,N_4534,N_4978);
nand U5343 (N_5343,N_4619,N_4621);
or U5344 (N_5344,N_4972,N_4673);
nand U5345 (N_5345,N_4836,N_4898);
nand U5346 (N_5346,N_4635,N_4643);
and U5347 (N_5347,N_4980,N_4717);
nor U5348 (N_5348,N_4565,N_4893);
and U5349 (N_5349,N_4560,N_4870);
nand U5350 (N_5350,N_4601,N_4950);
xnor U5351 (N_5351,N_4776,N_4634);
or U5352 (N_5352,N_4607,N_4738);
and U5353 (N_5353,N_4568,N_4861);
nand U5354 (N_5354,N_4811,N_4531);
xnor U5355 (N_5355,N_4713,N_4789);
xnor U5356 (N_5356,N_4989,N_4923);
nor U5357 (N_5357,N_4959,N_4784);
or U5358 (N_5358,N_4893,N_4968);
or U5359 (N_5359,N_4881,N_4770);
or U5360 (N_5360,N_4863,N_4687);
nand U5361 (N_5361,N_4979,N_4678);
nand U5362 (N_5362,N_4899,N_4803);
xnor U5363 (N_5363,N_4649,N_4785);
nand U5364 (N_5364,N_4823,N_4951);
xor U5365 (N_5365,N_4886,N_4545);
or U5366 (N_5366,N_4802,N_4775);
nor U5367 (N_5367,N_4674,N_4927);
xor U5368 (N_5368,N_4797,N_4677);
and U5369 (N_5369,N_4962,N_4530);
nor U5370 (N_5370,N_4909,N_4765);
xor U5371 (N_5371,N_4938,N_4764);
or U5372 (N_5372,N_4644,N_4721);
and U5373 (N_5373,N_4860,N_4938);
nand U5374 (N_5374,N_4984,N_4828);
xor U5375 (N_5375,N_4648,N_4893);
and U5376 (N_5376,N_4818,N_4923);
and U5377 (N_5377,N_4902,N_4694);
nand U5378 (N_5378,N_4887,N_4926);
or U5379 (N_5379,N_4993,N_4983);
and U5380 (N_5380,N_4893,N_4840);
or U5381 (N_5381,N_4515,N_4977);
or U5382 (N_5382,N_4553,N_4943);
xnor U5383 (N_5383,N_4933,N_4609);
xnor U5384 (N_5384,N_4694,N_4653);
and U5385 (N_5385,N_4831,N_4999);
nor U5386 (N_5386,N_4636,N_4919);
nor U5387 (N_5387,N_4535,N_4829);
or U5388 (N_5388,N_4895,N_4922);
and U5389 (N_5389,N_4911,N_4895);
xnor U5390 (N_5390,N_4702,N_4959);
and U5391 (N_5391,N_4931,N_4723);
nand U5392 (N_5392,N_4965,N_4977);
and U5393 (N_5393,N_4714,N_4652);
nor U5394 (N_5394,N_4839,N_4935);
or U5395 (N_5395,N_4666,N_4544);
xor U5396 (N_5396,N_4551,N_4637);
and U5397 (N_5397,N_4981,N_4794);
nor U5398 (N_5398,N_4710,N_4903);
nor U5399 (N_5399,N_4757,N_4951);
nand U5400 (N_5400,N_4627,N_4901);
and U5401 (N_5401,N_4879,N_4726);
and U5402 (N_5402,N_4803,N_4502);
and U5403 (N_5403,N_4582,N_4953);
nand U5404 (N_5404,N_4590,N_4727);
xor U5405 (N_5405,N_4931,N_4562);
xor U5406 (N_5406,N_4506,N_4513);
or U5407 (N_5407,N_4525,N_4699);
nand U5408 (N_5408,N_4969,N_4878);
nand U5409 (N_5409,N_4705,N_4736);
or U5410 (N_5410,N_4685,N_4631);
or U5411 (N_5411,N_4796,N_4769);
nand U5412 (N_5412,N_4546,N_4887);
or U5413 (N_5413,N_4742,N_4795);
or U5414 (N_5414,N_4812,N_4851);
or U5415 (N_5415,N_4771,N_4820);
nand U5416 (N_5416,N_4656,N_4684);
nor U5417 (N_5417,N_4948,N_4906);
xnor U5418 (N_5418,N_4803,N_4954);
and U5419 (N_5419,N_4623,N_4871);
or U5420 (N_5420,N_4870,N_4935);
nand U5421 (N_5421,N_4524,N_4925);
nor U5422 (N_5422,N_4961,N_4966);
and U5423 (N_5423,N_4623,N_4632);
nand U5424 (N_5424,N_4643,N_4791);
nand U5425 (N_5425,N_4895,N_4519);
or U5426 (N_5426,N_4892,N_4570);
xor U5427 (N_5427,N_4688,N_4884);
and U5428 (N_5428,N_4994,N_4585);
xnor U5429 (N_5429,N_4873,N_4527);
xor U5430 (N_5430,N_4646,N_4616);
and U5431 (N_5431,N_4873,N_4623);
nor U5432 (N_5432,N_4874,N_4623);
or U5433 (N_5433,N_4745,N_4552);
and U5434 (N_5434,N_4723,N_4814);
xor U5435 (N_5435,N_4549,N_4926);
or U5436 (N_5436,N_4552,N_4543);
nor U5437 (N_5437,N_4610,N_4741);
or U5438 (N_5438,N_4762,N_4917);
nor U5439 (N_5439,N_4591,N_4884);
and U5440 (N_5440,N_4646,N_4822);
xor U5441 (N_5441,N_4983,N_4776);
xnor U5442 (N_5442,N_4793,N_4861);
nand U5443 (N_5443,N_4742,N_4915);
and U5444 (N_5444,N_4664,N_4773);
or U5445 (N_5445,N_4816,N_4621);
xor U5446 (N_5446,N_4648,N_4813);
xor U5447 (N_5447,N_4980,N_4864);
or U5448 (N_5448,N_4901,N_4831);
nor U5449 (N_5449,N_4821,N_4735);
nor U5450 (N_5450,N_4590,N_4689);
or U5451 (N_5451,N_4621,N_4989);
and U5452 (N_5452,N_4589,N_4654);
nor U5453 (N_5453,N_4731,N_4790);
and U5454 (N_5454,N_4786,N_4957);
nand U5455 (N_5455,N_4892,N_4646);
or U5456 (N_5456,N_4699,N_4824);
and U5457 (N_5457,N_4972,N_4860);
and U5458 (N_5458,N_4623,N_4856);
and U5459 (N_5459,N_4786,N_4995);
nand U5460 (N_5460,N_4765,N_4816);
and U5461 (N_5461,N_4874,N_4780);
and U5462 (N_5462,N_4730,N_4838);
and U5463 (N_5463,N_4587,N_4636);
nor U5464 (N_5464,N_4938,N_4631);
or U5465 (N_5465,N_4786,N_4531);
or U5466 (N_5466,N_4587,N_4737);
or U5467 (N_5467,N_4836,N_4595);
xor U5468 (N_5468,N_4997,N_4907);
nand U5469 (N_5469,N_4597,N_4526);
nand U5470 (N_5470,N_4756,N_4839);
xor U5471 (N_5471,N_4743,N_4843);
xor U5472 (N_5472,N_4766,N_4822);
nor U5473 (N_5473,N_4885,N_4703);
nand U5474 (N_5474,N_4693,N_4662);
or U5475 (N_5475,N_4728,N_4543);
nor U5476 (N_5476,N_4648,N_4888);
nor U5477 (N_5477,N_4873,N_4984);
nor U5478 (N_5478,N_4961,N_4776);
or U5479 (N_5479,N_4953,N_4769);
nor U5480 (N_5480,N_4985,N_4514);
nand U5481 (N_5481,N_4528,N_4520);
xor U5482 (N_5482,N_4727,N_4872);
xor U5483 (N_5483,N_4756,N_4994);
nor U5484 (N_5484,N_4562,N_4910);
xor U5485 (N_5485,N_4820,N_4785);
xnor U5486 (N_5486,N_4770,N_4664);
nor U5487 (N_5487,N_4808,N_4890);
or U5488 (N_5488,N_4655,N_4786);
nor U5489 (N_5489,N_4861,N_4742);
xor U5490 (N_5490,N_4876,N_4804);
and U5491 (N_5491,N_4669,N_4977);
nand U5492 (N_5492,N_4841,N_4776);
or U5493 (N_5493,N_4722,N_4668);
and U5494 (N_5494,N_4547,N_4895);
and U5495 (N_5495,N_4918,N_4948);
nand U5496 (N_5496,N_4833,N_4683);
nor U5497 (N_5497,N_4682,N_4522);
or U5498 (N_5498,N_4935,N_4925);
xnor U5499 (N_5499,N_4776,N_4807);
or U5500 (N_5500,N_5347,N_5326);
nand U5501 (N_5501,N_5272,N_5041);
xor U5502 (N_5502,N_5410,N_5091);
and U5503 (N_5503,N_5423,N_5336);
nor U5504 (N_5504,N_5366,N_5044);
or U5505 (N_5505,N_5493,N_5032);
or U5506 (N_5506,N_5431,N_5169);
and U5507 (N_5507,N_5452,N_5327);
xor U5508 (N_5508,N_5024,N_5198);
nand U5509 (N_5509,N_5181,N_5102);
and U5510 (N_5510,N_5385,N_5241);
nand U5511 (N_5511,N_5222,N_5252);
and U5512 (N_5512,N_5417,N_5116);
nor U5513 (N_5513,N_5176,N_5226);
or U5514 (N_5514,N_5060,N_5473);
nand U5515 (N_5515,N_5190,N_5085);
nand U5516 (N_5516,N_5031,N_5063);
nand U5517 (N_5517,N_5273,N_5158);
or U5518 (N_5518,N_5195,N_5406);
or U5519 (N_5519,N_5334,N_5426);
or U5520 (N_5520,N_5332,N_5098);
or U5521 (N_5521,N_5090,N_5320);
nor U5522 (N_5522,N_5046,N_5216);
xnor U5523 (N_5523,N_5424,N_5300);
xnor U5524 (N_5524,N_5125,N_5382);
or U5525 (N_5525,N_5022,N_5053);
and U5526 (N_5526,N_5271,N_5159);
nor U5527 (N_5527,N_5244,N_5330);
or U5528 (N_5528,N_5391,N_5435);
or U5529 (N_5529,N_5135,N_5077);
or U5530 (N_5530,N_5317,N_5064);
nor U5531 (N_5531,N_5008,N_5472);
nand U5532 (N_5532,N_5021,N_5062);
or U5533 (N_5533,N_5051,N_5066);
or U5534 (N_5534,N_5365,N_5175);
nand U5535 (N_5535,N_5476,N_5335);
or U5536 (N_5536,N_5166,N_5362);
and U5537 (N_5537,N_5274,N_5034);
xnor U5538 (N_5538,N_5133,N_5261);
and U5539 (N_5539,N_5318,N_5432);
or U5540 (N_5540,N_5170,N_5314);
nand U5541 (N_5541,N_5210,N_5356);
and U5542 (N_5542,N_5402,N_5427);
and U5543 (N_5543,N_5388,N_5136);
xnor U5544 (N_5544,N_5396,N_5011);
xor U5545 (N_5545,N_5023,N_5143);
or U5546 (N_5546,N_5313,N_5139);
xnor U5547 (N_5547,N_5351,N_5392);
xnor U5548 (N_5548,N_5304,N_5411);
nand U5549 (N_5549,N_5324,N_5217);
and U5550 (N_5550,N_5377,N_5269);
nand U5551 (N_5551,N_5279,N_5033);
nand U5552 (N_5552,N_5214,N_5122);
nand U5553 (N_5553,N_5444,N_5087);
nor U5554 (N_5554,N_5455,N_5393);
xnor U5555 (N_5555,N_5134,N_5132);
or U5556 (N_5556,N_5345,N_5038);
xnor U5557 (N_5557,N_5479,N_5086);
or U5558 (N_5558,N_5164,N_5243);
nor U5559 (N_5559,N_5291,N_5121);
xnor U5560 (N_5560,N_5384,N_5364);
xnor U5561 (N_5561,N_5020,N_5311);
nor U5562 (N_5562,N_5454,N_5144);
nand U5563 (N_5563,N_5386,N_5154);
nor U5564 (N_5564,N_5376,N_5110);
and U5565 (N_5565,N_5497,N_5453);
nor U5566 (N_5566,N_5319,N_5468);
nor U5567 (N_5567,N_5178,N_5138);
nand U5568 (N_5568,N_5446,N_5367);
or U5569 (N_5569,N_5416,N_5074);
or U5570 (N_5570,N_5076,N_5151);
and U5571 (N_5571,N_5192,N_5496);
nand U5572 (N_5572,N_5147,N_5407);
xor U5573 (N_5573,N_5389,N_5254);
and U5574 (N_5574,N_5232,N_5073);
or U5575 (N_5575,N_5089,N_5039);
nand U5576 (N_5576,N_5126,N_5301);
nor U5577 (N_5577,N_5184,N_5413);
nor U5578 (N_5578,N_5266,N_5149);
and U5579 (N_5579,N_5310,N_5280);
or U5580 (N_5580,N_5483,N_5030);
and U5581 (N_5581,N_5474,N_5270);
nand U5582 (N_5582,N_5227,N_5489);
or U5583 (N_5583,N_5357,N_5234);
or U5584 (N_5584,N_5460,N_5448);
nand U5585 (N_5585,N_5208,N_5119);
nand U5586 (N_5586,N_5302,N_5199);
nand U5587 (N_5587,N_5415,N_5428);
and U5588 (N_5588,N_5488,N_5399);
xor U5589 (N_5589,N_5188,N_5442);
or U5590 (N_5590,N_5200,N_5451);
xor U5591 (N_5591,N_5436,N_5128);
nand U5592 (N_5592,N_5145,N_5215);
xnor U5593 (N_5593,N_5464,N_5204);
and U5594 (N_5594,N_5485,N_5095);
xor U5595 (N_5595,N_5109,N_5012);
xor U5596 (N_5596,N_5056,N_5323);
xnor U5597 (N_5597,N_5219,N_5420);
or U5598 (N_5598,N_5113,N_5398);
or U5599 (N_5599,N_5306,N_5209);
nor U5600 (N_5600,N_5434,N_5194);
nand U5601 (N_5601,N_5054,N_5425);
xor U5602 (N_5602,N_5189,N_5440);
or U5603 (N_5603,N_5287,N_5106);
nor U5604 (N_5604,N_5043,N_5185);
and U5605 (N_5605,N_5491,N_5341);
xor U5606 (N_5606,N_5490,N_5017);
nand U5607 (N_5607,N_5156,N_5340);
nor U5608 (N_5608,N_5183,N_5288);
nand U5609 (N_5609,N_5167,N_5492);
and U5610 (N_5610,N_5006,N_5371);
and U5611 (N_5611,N_5463,N_5299);
xor U5612 (N_5612,N_5173,N_5289);
or U5613 (N_5613,N_5224,N_5403);
nand U5614 (N_5614,N_5025,N_5267);
nor U5615 (N_5615,N_5005,N_5001);
nor U5616 (N_5616,N_5029,N_5478);
xor U5617 (N_5617,N_5482,N_5450);
nand U5618 (N_5618,N_5157,N_5142);
or U5619 (N_5619,N_5187,N_5048);
and U5620 (N_5620,N_5329,N_5177);
xnor U5621 (N_5621,N_5223,N_5408);
nand U5622 (N_5622,N_5247,N_5305);
nand U5623 (N_5623,N_5103,N_5160);
and U5624 (N_5624,N_5118,N_5211);
and U5625 (N_5625,N_5007,N_5100);
or U5626 (N_5626,N_5284,N_5239);
or U5627 (N_5627,N_5081,N_5421);
nor U5628 (N_5628,N_5148,N_5262);
and U5629 (N_5629,N_5179,N_5096);
nor U5630 (N_5630,N_5229,N_5378);
xor U5631 (N_5631,N_5484,N_5027);
nor U5632 (N_5632,N_5242,N_5141);
nor U5633 (N_5633,N_5225,N_5111);
or U5634 (N_5634,N_5088,N_5000);
xor U5635 (N_5635,N_5083,N_5315);
nand U5636 (N_5636,N_5487,N_5220);
xnor U5637 (N_5637,N_5494,N_5236);
nand U5638 (N_5638,N_5230,N_5297);
xor U5639 (N_5639,N_5369,N_5438);
nand U5640 (N_5640,N_5316,N_5035);
xor U5641 (N_5641,N_5061,N_5155);
or U5642 (N_5642,N_5124,N_5354);
or U5643 (N_5643,N_5481,N_5248);
xnor U5644 (N_5644,N_5449,N_5397);
nor U5645 (N_5645,N_5268,N_5312);
or U5646 (N_5646,N_5099,N_5245);
nand U5647 (N_5647,N_5338,N_5499);
nand U5648 (N_5648,N_5146,N_5470);
nand U5649 (N_5649,N_5174,N_5105);
or U5650 (N_5650,N_5249,N_5298);
xnor U5651 (N_5651,N_5040,N_5441);
xnor U5652 (N_5652,N_5309,N_5419);
xnor U5653 (N_5653,N_5107,N_5221);
and U5654 (N_5654,N_5331,N_5094);
xor U5655 (N_5655,N_5387,N_5457);
and U5656 (N_5656,N_5072,N_5079);
nand U5657 (N_5657,N_5127,N_5153);
nor U5658 (N_5658,N_5395,N_5131);
nor U5659 (N_5659,N_5171,N_5019);
and U5660 (N_5660,N_5276,N_5193);
xnor U5661 (N_5661,N_5429,N_5228);
or U5662 (N_5662,N_5295,N_5028);
and U5663 (N_5663,N_5477,N_5161);
or U5664 (N_5664,N_5333,N_5152);
or U5665 (N_5665,N_5137,N_5165);
nand U5666 (N_5666,N_5069,N_5070);
or U5667 (N_5667,N_5401,N_5058);
nor U5668 (N_5668,N_5277,N_5379);
xor U5669 (N_5669,N_5359,N_5250);
or U5670 (N_5670,N_5466,N_5114);
nand U5671 (N_5671,N_5003,N_5002);
nor U5672 (N_5672,N_5337,N_5071);
nand U5673 (N_5673,N_5349,N_5462);
xnor U5674 (N_5674,N_5253,N_5237);
nor U5675 (N_5675,N_5405,N_5016);
or U5676 (N_5676,N_5263,N_5358);
and U5677 (N_5677,N_5258,N_5037);
or U5678 (N_5678,N_5422,N_5456);
nor U5679 (N_5679,N_5049,N_5256);
xnor U5680 (N_5680,N_5394,N_5055);
or U5681 (N_5681,N_5368,N_5196);
or U5682 (N_5682,N_5197,N_5057);
nand U5683 (N_5683,N_5260,N_5259);
xnor U5684 (N_5684,N_5308,N_5380);
nand U5685 (N_5685,N_5212,N_5129);
or U5686 (N_5686,N_5445,N_5495);
nand U5687 (N_5687,N_5350,N_5443);
or U5688 (N_5688,N_5162,N_5293);
nand U5689 (N_5689,N_5026,N_5172);
nand U5690 (N_5690,N_5010,N_5205);
nand U5691 (N_5691,N_5339,N_5059);
and U5692 (N_5692,N_5409,N_5264);
xnor U5693 (N_5693,N_5251,N_5104);
or U5694 (N_5694,N_5286,N_5383);
and U5695 (N_5695,N_5290,N_5275);
nor U5696 (N_5696,N_5203,N_5437);
xnor U5697 (N_5697,N_5123,N_5285);
nand U5698 (N_5698,N_5303,N_5404);
or U5699 (N_5699,N_5467,N_5322);
xor U5700 (N_5700,N_5082,N_5292);
and U5701 (N_5701,N_5238,N_5014);
and U5702 (N_5702,N_5186,N_5112);
or U5703 (N_5703,N_5414,N_5080);
xor U5704 (N_5704,N_5042,N_5370);
xnor U5705 (N_5705,N_5018,N_5231);
and U5706 (N_5706,N_5321,N_5108);
or U5707 (N_5707,N_5004,N_5343);
nor U5708 (N_5708,N_5328,N_5180);
or U5709 (N_5709,N_5418,N_5400);
nor U5710 (N_5710,N_5355,N_5045);
and U5711 (N_5711,N_5361,N_5353);
or U5712 (N_5712,N_5430,N_5342);
nand U5713 (N_5713,N_5218,N_5480);
nor U5714 (N_5714,N_5207,N_5465);
nor U5715 (N_5715,N_5078,N_5201);
nor U5716 (N_5716,N_5294,N_5412);
nand U5717 (N_5717,N_5240,N_5191);
and U5718 (N_5718,N_5101,N_5013);
xnor U5719 (N_5719,N_5352,N_5381);
and U5720 (N_5720,N_5296,N_5498);
and U5721 (N_5721,N_5447,N_5439);
xnor U5722 (N_5722,N_5117,N_5283);
or U5723 (N_5723,N_5475,N_5307);
xnor U5724 (N_5724,N_5206,N_5140);
xor U5725 (N_5725,N_5233,N_5325);
and U5726 (N_5726,N_5246,N_5068);
nor U5727 (N_5727,N_5150,N_5459);
nor U5728 (N_5728,N_5075,N_5346);
nor U5729 (N_5729,N_5363,N_5213);
or U5730 (N_5730,N_5265,N_5015);
nand U5731 (N_5731,N_5458,N_5278);
or U5732 (N_5732,N_5130,N_5050);
nand U5733 (N_5733,N_5168,N_5255);
and U5734 (N_5734,N_5052,N_5390);
xnor U5735 (N_5735,N_5084,N_5486);
and U5736 (N_5736,N_5433,N_5461);
xor U5737 (N_5737,N_5374,N_5065);
nor U5738 (N_5738,N_5036,N_5469);
or U5739 (N_5739,N_5348,N_5182);
nor U5740 (N_5740,N_5163,N_5092);
and U5741 (N_5741,N_5471,N_5344);
and U5742 (N_5742,N_5372,N_5257);
nor U5743 (N_5743,N_5115,N_5120);
nand U5744 (N_5744,N_5067,N_5097);
or U5745 (N_5745,N_5047,N_5235);
nand U5746 (N_5746,N_5009,N_5282);
and U5747 (N_5747,N_5375,N_5360);
nand U5748 (N_5748,N_5093,N_5202);
and U5749 (N_5749,N_5373,N_5281);
nor U5750 (N_5750,N_5301,N_5079);
nor U5751 (N_5751,N_5387,N_5403);
nand U5752 (N_5752,N_5367,N_5098);
nand U5753 (N_5753,N_5478,N_5091);
and U5754 (N_5754,N_5056,N_5063);
or U5755 (N_5755,N_5085,N_5107);
or U5756 (N_5756,N_5247,N_5076);
nand U5757 (N_5757,N_5373,N_5411);
nand U5758 (N_5758,N_5487,N_5410);
and U5759 (N_5759,N_5147,N_5341);
nand U5760 (N_5760,N_5066,N_5235);
xnor U5761 (N_5761,N_5077,N_5018);
or U5762 (N_5762,N_5006,N_5142);
nand U5763 (N_5763,N_5170,N_5302);
and U5764 (N_5764,N_5203,N_5059);
nand U5765 (N_5765,N_5187,N_5405);
and U5766 (N_5766,N_5127,N_5035);
xor U5767 (N_5767,N_5077,N_5218);
nand U5768 (N_5768,N_5303,N_5362);
and U5769 (N_5769,N_5469,N_5493);
and U5770 (N_5770,N_5263,N_5078);
xor U5771 (N_5771,N_5360,N_5002);
and U5772 (N_5772,N_5245,N_5355);
and U5773 (N_5773,N_5442,N_5006);
xor U5774 (N_5774,N_5021,N_5222);
xnor U5775 (N_5775,N_5462,N_5030);
or U5776 (N_5776,N_5020,N_5291);
or U5777 (N_5777,N_5331,N_5249);
and U5778 (N_5778,N_5161,N_5077);
xnor U5779 (N_5779,N_5175,N_5071);
and U5780 (N_5780,N_5135,N_5299);
nand U5781 (N_5781,N_5118,N_5004);
nor U5782 (N_5782,N_5186,N_5373);
nor U5783 (N_5783,N_5247,N_5472);
nor U5784 (N_5784,N_5077,N_5497);
nor U5785 (N_5785,N_5182,N_5491);
and U5786 (N_5786,N_5381,N_5285);
xnor U5787 (N_5787,N_5019,N_5219);
xnor U5788 (N_5788,N_5431,N_5349);
xor U5789 (N_5789,N_5281,N_5382);
nand U5790 (N_5790,N_5157,N_5222);
or U5791 (N_5791,N_5148,N_5028);
or U5792 (N_5792,N_5018,N_5189);
nor U5793 (N_5793,N_5421,N_5429);
nor U5794 (N_5794,N_5192,N_5374);
nor U5795 (N_5795,N_5115,N_5490);
nor U5796 (N_5796,N_5030,N_5167);
nor U5797 (N_5797,N_5046,N_5149);
or U5798 (N_5798,N_5163,N_5198);
xor U5799 (N_5799,N_5275,N_5177);
xnor U5800 (N_5800,N_5380,N_5144);
nand U5801 (N_5801,N_5300,N_5233);
or U5802 (N_5802,N_5223,N_5139);
or U5803 (N_5803,N_5048,N_5237);
xor U5804 (N_5804,N_5236,N_5212);
nor U5805 (N_5805,N_5405,N_5066);
nand U5806 (N_5806,N_5120,N_5098);
and U5807 (N_5807,N_5056,N_5055);
nand U5808 (N_5808,N_5227,N_5268);
xor U5809 (N_5809,N_5229,N_5364);
nor U5810 (N_5810,N_5005,N_5179);
or U5811 (N_5811,N_5365,N_5047);
nand U5812 (N_5812,N_5448,N_5323);
xor U5813 (N_5813,N_5295,N_5177);
and U5814 (N_5814,N_5239,N_5290);
nand U5815 (N_5815,N_5175,N_5310);
nand U5816 (N_5816,N_5034,N_5002);
or U5817 (N_5817,N_5134,N_5332);
or U5818 (N_5818,N_5149,N_5446);
nor U5819 (N_5819,N_5089,N_5178);
or U5820 (N_5820,N_5198,N_5058);
nand U5821 (N_5821,N_5061,N_5100);
nor U5822 (N_5822,N_5497,N_5285);
nor U5823 (N_5823,N_5020,N_5226);
and U5824 (N_5824,N_5442,N_5097);
or U5825 (N_5825,N_5352,N_5150);
or U5826 (N_5826,N_5205,N_5044);
and U5827 (N_5827,N_5172,N_5370);
xor U5828 (N_5828,N_5303,N_5413);
or U5829 (N_5829,N_5487,N_5070);
and U5830 (N_5830,N_5432,N_5240);
or U5831 (N_5831,N_5359,N_5135);
xor U5832 (N_5832,N_5447,N_5098);
nor U5833 (N_5833,N_5130,N_5177);
xnor U5834 (N_5834,N_5173,N_5170);
nand U5835 (N_5835,N_5279,N_5179);
nand U5836 (N_5836,N_5241,N_5358);
nand U5837 (N_5837,N_5355,N_5459);
nor U5838 (N_5838,N_5153,N_5256);
xnor U5839 (N_5839,N_5481,N_5147);
nor U5840 (N_5840,N_5458,N_5098);
or U5841 (N_5841,N_5159,N_5182);
xnor U5842 (N_5842,N_5253,N_5034);
and U5843 (N_5843,N_5288,N_5370);
nor U5844 (N_5844,N_5489,N_5478);
xnor U5845 (N_5845,N_5092,N_5110);
or U5846 (N_5846,N_5382,N_5261);
and U5847 (N_5847,N_5260,N_5111);
and U5848 (N_5848,N_5012,N_5492);
or U5849 (N_5849,N_5489,N_5050);
and U5850 (N_5850,N_5364,N_5095);
xnor U5851 (N_5851,N_5197,N_5040);
or U5852 (N_5852,N_5352,N_5084);
nand U5853 (N_5853,N_5372,N_5464);
and U5854 (N_5854,N_5198,N_5226);
nand U5855 (N_5855,N_5150,N_5409);
or U5856 (N_5856,N_5320,N_5110);
nand U5857 (N_5857,N_5464,N_5487);
or U5858 (N_5858,N_5064,N_5310);
and U5859 (N_5859,N_5119,N_5228);
nor U5860 (N_5860,N_5429,N_5216);
xor U5861 (N_5861,N_5069,N_5291);
xor U5862 (N_5862,N_5430,N_5042);
nor U5863 (N_5863,N_5024,N_5426);
nor U5864 (N_5864,N_5472,N_5309);
or U5865 (N_5865,N_5280,N_5403);
xor U5866 (N_5866,N_5460,N_5085);
and U5867 (N_5867,N_5262,N_5477);
and U5868 (N_5868,N_5254,N_5111);
nor U5869 (N_5869,N_5236,N_5154);
nand U5870 (N_5870,N_5211,N_5181);
xor U5871 (N_5871,N_5345,N_5230);
nor U5872 (N_5872,N_5150,N_5470);
or U5873 (N_5873,N_5217,N_5368);
xnor U5874 (N_5874,N_5149,N_5468);
xnor U5875 (N_5875,N_5249,N_5434);
nand U5876 (N_5876,N_5106,N_5380);
nand U5877 (N_5877,N_5254,N_5313);
xor U5878 (N_5878,N_5051,N_5421);
and U5879 (N_5879,N_5499,N_5311);
nand U5880 (N_5880,N_5143,N_5154);
nand U5881 (N_5881,N_5249,N_5010);
and U5882 (N_5882,N_5247,N_5185);
or U5883 (N_5883,N_5044,N_5093);
and U5884 (N_5884,N_5147,N_5279);
nand U5885 (N_5885,N_5107,N_5429);
nor U5886 (N_5886,N_5336,N_5065);
nand U5887 (N_5887,N_5392,N_5339);
and U5888 (N_5888,N_5382,N_5499);
and U5889 (N_5889,N_5103,N_5071);
or U5890 (N_5890,N_5070,N_5037);
or U5891 (N_5891,N_5202,N_5240);
nor U5892 (N_5892,N_5092,N_5141);
and U5893 (N_5893,N_5394,N_5309);
nand U5894 (N_5894,N_5031,N_5109);
or U5895 (N_5895,N_5109,N_5039);
xor U5896 (N_5896,N_5223,N_5258);
nor U5897 (N_5897,N_5143,N_5315);
nor U5898 (N_5898,N_5405,N_5363);
nand U5899 (N_5899,N_5495,N_5231);
and U5900 (N_5900,N_5253,N_5369);
nand U5901 (N_5901,N_5118,N_5061);
nor U5902 (N_5902,N_5013,N_5422);
nor U5903 (N_5903,N_5068,N_5228);
and U5904 (N_5904,N_5470,N_5220);
or U5905 (N_5905,N_5188,N_5032);
or U5906 (N_5906,N_5161,N_5162);
nand U5907 (N_5907,N_5047,N_5155);
or U5908 (N_5908,N_5385,N_5218);
and U5909 (N_5909,N_5175,N_5156);
and U5910 (N_5910,N_5449,N_5280);
nor U5911 (N_5911,N_5197,N_5465);
xnor U5912 (N_5912,N_5412,N_5378);
nor U5913 (N_5913,N_5287,N_5200);
nor U5914 (N_5914,N_5239,N_5258);
xor U5915 (N_5915,N_5232,N_5149);
or U5916 (N_5916,N_5367,N_5176);
and U5917 (N_5917,N_5476,N_5040);
or U5918 (N_5918,N_5252,N_5375);
or U5919 (N_5919,N_5168,N_5293);
or U5920 (N_5920,N_5365,N_5129);
nand U5921 (N_5921,N_5498,N_5271);
or U5922 (N_5922,N_5413,N_5132);
or U5923 (N_5923,N_5065,N_5254);
nand U5924 (N_5924,N_5379,N_5387);
nor U5925 (N_5925,N_5122,N_5165);
or U5926 (N_5926,N_5182,N_5034);
xor U5927 (N_5927,N_5195,N_5317);
xnor U5928 (N_5928,N_5312,N_5117);
nand U5929 (N_5929,N_5466,N_5359);
xor U5930 (N_5930,N_5398,N_5250);
or U5931 (N_5931,N_5136,N_5391);
xor U5932 (N_5932,N_5269,N_5492);
or U5933 (N_5933,N_5202,N_5025);
or U5934 (N_5934,N_5053,N_5123);
and U5935 (N_5935,N_5123,N_5404);
xor U5936 (N_5936,N_5176,N_5127);
or U5937 (N_5937,N_5452,N_5409);
nor U5938 (N_5938,N_5299,N_5143);
xor U5939 (N_5939,N_5399,N_5425);
or U5940 (N_5940,N_5302,N_5165);
and U5941 (N_5941,N_5378,N_5196);
xor U5942 (N_5942,N_5406,N_5011);
nor U5943 (N_5943,N_5203,N_5172);
nand U5944 (N_5944,N_5020,N_5147);
and U5945 (N_5945,N_5429,N_5094);
and U5946 (N_5946,N_5264,N_5391);
nor U5947 (N_5947,N_5385,N_5416);
or U5948 (N_5948,N_5353,N_5461);
or U5949 (N_5949,N_5064,N_5011);
nand U5950 (N_5950,N_5157,N_5172);
and U5951 (N_5951,N_5004,N_5060);
nor U5952 (N_5952,N_5402,N_5471);
nand U5953 (N_5953,N_5394,N_5139);
or U5954 (N_5954,N_5074,N_5238);
and U5955 (N_5955,N_5134,N_5043);
or U5956 (N_5956,N_5046,N_5191);
nor U5957 (N_5957,N_5427,N_5428);
xor U5958 (N_5958,N_5363,N_5218);
nor U5959 (N_5959,N_5159,N_5254);
nor U5960 (N_5960,N_5133,N_5449);
or U5961 (N_5961,N_5211,N_5371);
xor U5962 (N_5962,N_5016,N_5045);
and U5963 (N_5963,N_5359,N_5042);
nand U5964 (N_5964,N_5230,N_5323);
nor U5965 (N_5965,N_5347,N_5394);
or U5966 (N_5966,N_5074,N_5452);
and U5967 (N_5967,N_5477,N_5273);
and U5968 (N_5968,N_5297,N_5449);
nand U5969 (N_5969,N_5135,N_5056);
or U5970 (N_5970,N_5416,N_5400);
xnor U5971 (N_5971,N_5457,N_5136);
nor U5972 (N_5972,N_5211,N_5293);
xnor U5973 (N_5973,N_5306,N_5494);
nand U5974 (N_5974,N_5074,N_5262);
xnor U5975 (N_5975,N_5168,N_5037);
nor U5976 (N_5976,N_5106,N_5401);
xor U5977 (N_5977,N_5277,N_5417);
and U5978 (N_5978,N_5132,N_5350);
nand U5979 (N_5979,N_5274,N_5268);
nand U5980 (N_5980,N_5401,N_5034);
nand U5981 (N_5981,N_5075,N_5162);
nand U5982 (N_5982,N_5208,N_5270);
or U5983 (N_5983,N_5053,N_5361);
and U5984 (N_5984,N_5252,N_5030);
nor U5985 (N_5985,N_5377,N_5270);
or U5986 (N_5986,N_5050,N_5358);
and U5987 (N_5987,N_5480,N_5002);
and U5988 (N_5988,N_5052,N_5440);
nor U5989 (N_5989,N_5156,N_5420);
nand U5990 (N_5990,N_5060,N_5128);
or U5991 (N_5991,N_5148,N_5130);
or U5992 (N_5992,N_5373,N_5237);
nor U5993 (N_5993,N_5060,N_5255);
and U5994 (N_5994,N_5016,N_5415);
and U5995 (N_5995,N_5211,N_5006);
xnor U5996 (N_5996,N_5265,N_5197);
xor U5997 (N_5997,N_5427,N_5192);
nand U5998 (N_5998,N_5462,N_5174);
xor U5999 (N_5999,N_5306,N_5345);
or U6000 (N_6000,N_5754,N_5873);
nor U6001 (N_6001,N_5811,N_5631);
xor U6002 (N_6002,N_5720,N_5749);
or U6003 (N_6003,N_5905,N_5939);
or U6004 (N_6004,N_5763,N_5746);
or U6005 (N_6005,N_5551,N_5675);
xnor U6006 (N_6006,N_5888,N_5825);
and U6007 (N_6007,N_5724,N_5819);
nor U6008 (N_6008,N_5598,N_5542);
xor U6009 (N_6009,N_5883,N_5773);
xnor U6010 (N_6010,N_5771,N_5816);
xor U6011 (N_6011,N_5574,N_5823);
nand U6012 (N_6012,N_5988,N_5790);
nand U6013 (N_6013,N_5989,N_5959);
nand U6014 (N_6014,N_5945,N_5686);
and U6015 (N_6015,N_5616,N_5697);
and U6016 (N_6016,N_5795,N_5668);
xnor U6017 (N_6017,N_5858,N_5878);
nor U6018 (N_6018,N_5608,N_5926);
or U6019 (N_6019,N_5728,N_5798);
nor U6020 (N_6020,N_5534,N_5700);
nand U6021 (N_6021,N_5956,N_5914);
nor U6022 (N_6022,N_5953,N_5979);
xnor U6023 (N_6023,N_5894,N_5593);
nor U6024 (N_6024,N_5557,N_5850);
nand U6025 (N_6025,N_5931,N_5703);
nor U6026 (N_6026,N_5961,N_5709);
nor U6027 (N_6027,N_5937,N_5846);
xor U6028 (N_6028,N_5607,N_5717);
nor U6029 (N_6029,N_5929,N_5652);
xnor U6030 (N_6030,N_5814,N_5995);
nand U6031 (N_6031,N_5853,N_5576);
nor U6032 (N_6032,N_5788,N_5716);
and U6033 (N_6033,N_5884,N_5969);
xnor U6034 (N_6034,N_5752,N_5662);
xnor U6035 (N_6035,N_5781,N_5568);
nand U6036 (N_6036,N_5789,N_5810);
and U6037 (N_6037,N_5513,N_5676);
nand U6038 (N_6038,N_5733,N_5645);
and U6039 (N_6039,N_5832,N_5923);
xor U6040 (N_6040,N_5635,N_5644);
or U6041 (N_6041,N_5550,N_5751);
xnor U6042 (N_6042,N_5809,N_5669);
and U6043 (N_6043,N_5680,N_5651);
and U6044 (N_6044,N_5708,N_5572);
xor U6045 (N_6045,N_5687,N_5666);
xor U6046 (N_6046,N_5737,N_5583);
xor U6047 (N_6047,N_5802,N_5739);
nor U6048 (N_6048,N_5590,N_5515);
and U6049 (N_6049,N_5615,N_5711);
nand U6050 (N_6050,N_5978,N_5529);
and U6051 (N_6051,N_5786,N_5831);
or U6052 (N_6052,N_5672,N_5560);
nor U6053 (N_6053,N_5817,N_5868);
and U6054 (N_6054,N_5648,N_5877);
nor U6055 (N_6055,N_5656,N_5958);
and U6056 (N_6056,N_5533,N_5954);
nor U6057 (N_6057,N_5587,N_5628);
nand U6058 (N_6058,N_5854,N_5876);
xor U6059 (N_6059,N_5775,N_5862);
nand U6060 (N_6060,N_5913,N_5869);
or U6061 (N_6061,N_5928,N_5500);
xor U6062 (N_6062,N_5804,N_5655);
nor U6063 (N_6063,N_5801,N_5595);
nand U6064 (N_6064,N_5930,N_5856);
nor U6065 (N_6065,N_5911,N_5982);
or U6066 (N_6066,N_5813,N_5743);
xor U6067 (N_6067,N_5774,N_5627);
nor U6068 (N_6068,N_5924,N_5904);
or U6069 (N_6069,N_5630,N_5829);
nand U6070 (N_6070,N_5507,N_5636);
and U6071 (N_6071,N_5867,N_5667);
and U6072 (N_6072,N_5599,N_5742);
xor U6073 (N_6073,N_5646,N_5714);
or U6074 (N_6074,N_5957,N_5796);
and U6075 (N_6075,N_5983,N_5808);
and U6076 (N_6076,N_5509,N_5664);
xor U6077 (N_6077,N_5552,N_5812);
nor U6078 (N_6078,N_5562,N_5890);
xnor U6079 (N_6079,N_5575,N_5670);
and U6080 (N_6080,N_5891,N_5759);
nor U6081 (N_6081,N_5898,N_5866);
or U6082 (N_6082,N_5779,N_5525);
nor U6083 (N_6083,N_5641,N_5882);
xnor U6084 (N_6084,N_5698,N_5885);
xnor U6085 (N_6085,N_5776,N_5673);
xnor U6086 (N_6086,N_5987,N_5519);
nor U6087 (N_6087,N_5643,N_5942);
and U6088 (N_6088,N_5538,N_5563);
xor U6089 (N_6089,N_5691,N_5745);
and U6090 (N_6090,N_5503,N_5985);
or U6091 (N_6091,N_5906,N_5506);
and U6092 (N_6092,N_5947,N_5976);
or U6093 (N_6093,N_5847,N_5710);
nor U6094 (N_6094,N_5613,N_5824);
xnor U6095 (N_6095,N_5870,N_5603);
nor U6096 (N_6096,N_5696,N_5962);
nor U6097 (N_6097,N_5921,N_5879);
and U6098 (N_6098,N_5718,N_5740);
xor U6099 (N_6099,N_5963,N_5578);
nor U6100 (N_6100,N_5665,N_5586);
xor U6101 (N_6101,N_5860,N_5543);
xor U6102 (N_6102,N_5642,N_5677);
nor U6103 (N_6103,N_5756,N_5640);
and U6104 (N_6104,N_5863,N_5830);
nor U6105 (N_6105,N_5734,N_5951);
or U6106 (N_6106,N_5654,N_5547);
or U6107 (N_6107,N_5907,N_5851);
nor U6108 (N_6108,N_5544,N_5561);
nor U6109 (N_6109,N_5925,N_5764);
nor U6110 (N_6110,N_5567,N_5597);
and U6111 (N_6111,N_5539,N_5683);
nand U6112 (N_6112,N_5875,N_5622);
nor U6113 (N_6113,N_5981,N_5571);
xnor U6114 (N_6114,N_5614,N_5548);
nor U6115 (N_6115,N_5527,N_5712);
and U6116 (N_6116,N_5502,N_5611);
nor U6117 (N_6117,N_5653,N_5573);
xor U6118 (N_6118,N_5944,N_5532);
xor U6119 (N_6119,N_5591,N_5726);
nor U6120 (N_6120,N_5606,N_5577);
and U6121 (N_6121,N_5649,N_5909);
nand U6122 (N_6122,N_5835,N_5514);
and U6123 (N_6123,N_5735,N_5834);
and U6124 (N_6124,N_5657,N_5900);
xor U6125 (N_6125,N_5689,N_5715);
nor U6126 (N_6126,N_5650,N_5960);
and U6127 (N_6127,N_5827,N_5933);
and U6128 (N_6128,N_5528,N_5970);
or U6129 (N_6129,N_5510,N_5865);
or U6130 (N_6130,N_5535,N_5619);
or U6131 (N_6131,N_5524,N_5968);
nor U6132 (N_6132,N_5950,N_5936);
and U6133 (N_6133,N_5915,N_5920);
nor U6134 (N_6134,N_5517,N_5895);
and U6135 (N_6135,N_5661,N_5620);
and U6136 (N_6136,N_5741,N_5792);
nand U6137 (N_6137,N_5537,N_5545);
and U6138 (N_6138,N_5946,N_5855);
xnor U6139 (N_6139,N_5778,N_5838);
or U6140 (N_6140,N_5852,N_5549);
and U6141 (N_6141,N_5901,N_5755);
nand U6142 (N_6142,N_5526,N_5772);
or U6143 (N_6143,N_5807,N_5585);
nand U6144 (N_6144,N_5727,N_5617);
and U6145 (N_6145,N_5848,N_5972);
nor U6146 (N_6146,N_5967,N_5618);
nand U6147 (N_6147,N_5899,N_5986);
nor U6148 (N_6148,N_5629,N_5659);
and U6149 (N_6149,N_5584,N_5553);
xor U6150 (N_6150,N_5623,N_5688);
and U6151 (N_6151,N_5569,N_5540);
or U6152 (N_6152,N_5769,N_5588);
xor U6153 (N_6153,N_5766,N_5999);
and U6154 (N_6154,N_5821,N_5601);
nand U6155 (N_6155,N_5935,N_5511);
nand U6156 (N_6156,N_5632,N_5843);
nor U6157 (N_6157,N_5828,N_5785);
xor U6158 (N_6158,N_5522,N_5952);
and U6159 (N_6159,N_5530,N_5671);
nand U6160 (N_6160,N_5881,N_5818);
and U6161 (N_6161,N_5508,N_5554);
and U6162 (N_6162,N_5721,N_5908);
and U6163 (N_6163,N_5993,N_5658);
or U6164 (N_6164,N_5991,N_5621);
nand U6165 (N_6165,N_5546,N_5753);
and U6166 (N_6166,N_5725,N_5580);
and U6167 (N_6167,N_5520,N_5797);
nor U6168 (N_6168,N_5767,N_5886);
nand U6169 (N_6169,N_5592,N_5762);
nor U6170 (N_6170,N_5722,N_5996);
xnor U6171 (N_6171,N_5941,N_5761);
nor U6172 (N_6172,N_5992,N_5682);
xnor U6173 (N_6173,N_5780,N_5731);
nand U6174 (N_6174,N_5610,N_5845);
or U6175 (N_6175,N_5965,N_5706);
and U6176 (N_6176,N_5889,N_5699);
xnor U6177 (N_6177,N_5744,N_5501);
nand U6178 (N_6178,N_5581,N_5600);
or U6179 (N_6179,N_5674,N_5541);
nor U6180 (N_6180,N_5555,N_5815);
or U6181 (N_6181,N_5777,N_5663);
or U6182 (N_6182,N_5949,N_5512);
nor U6183 (N_6183,N_5861,N_5932);
xor U6184 (N_6184,N_5748,N_5806);
and U6185 (N_6185,N_5782,N_5565);
nor U6186 (N_6186,N_5826,N_5910);
nand U6187 (N_6187,N_5589,N_5694);
nor U6188 (N_6188,N_5605,N_5799);
or U6189 (N_6189,N_5844,N_5768);
xor U6190 (N_6190,N_5975,N_5912);
nand U6191 (N_6191,N_5602,N_5922);
nor U6192 (N_6192,N_5880,N_5940);
xnor U6193 (N_6193,N_5730,N_5504);
nand U6194 (N_6194,N_5903,N_5842);
or U6195 (N_6195,N_5893,N_5897);
xnor U6196 (N_6196,N_5707,N_5998);
nand U6197 (N_6197,N_5558,N_5916);
and U6198 (N_6198,N_5892,N_5849);
or U6199 (N_6199,N_5784,N_5966);
nand U6200 (N_6200,N_5639,N_5971);
nor U6201 (N_6201,N_5990,N_5692);
nor U6202 (N_6202,N_5918,N_5679);
and U6203 (N_6203,N_5633,N_5864);
nand U6204 (N_6204,N_5582,N_5841);
and U6205 (N_6205,N_5836,N_5723);
nor U6206 (N_6206,N_5750,N_5704);
xnor U6207 (N_6207,N_5833,N_5997);
or U6208 (N_6208,N_5518,N_5738);
nand U6209 (N_6209,N_5757,N_5839);
nor U6210 (N_6210,N_5747,N_5713);
or U6211 (N_6211,N_5678,N_5660);
nand U6212 (N_6212,N_5857,N_5579);
nand U6213 (N_6213,N_5917,N_5943);
nand U6214 (N_6214,N_5690,N_5758);
xor U6215 (N_6215,N_5736,N_5612);
nor U6216 (N_6216,N_5685,N_5566);
or U6217 (N_6217,N_5559,N_5505);
nor U6218 (N_6218,N_5637,N_5787);
or U6219 (N_6219,N_5556,N_5596);
nand U6220 (N_6220,N_5770,N_5783);
xnor U6221 (N_6221,N_5594,N_5570);
or U6222 (N_6222,N_5874,N_5695);
or U6223 (N_6223,N_5980,N_5872);
nor U6224 (N_6224,N_5794,N_5805);
xnor U6225 (N_6225,N_5919,N_5984);
nand U6226 (N_6226,N_5701,N_5729);
and U6227 (N_6227,N_5822,N_5803);
nor U6228 (N_6228,N_5760,N_5604);
and U6229 (N_6229,N_5955,N_5732);
xnor U6230 (N_6230,N_5793,N_5887);
or U6231 (N_6231,N_5948,N_5902);
xor U6232 (N_6232,N_5624,N_5840);
nand U6233 (N_6233,N_5681,N_5938);
xnor U6234 (N_6234,N_5837,N_5964);
xor U6235 (N_6235,N_5820,N_5536);
or U6236 (N_6236,N_5521,N_5974);
nor U6237 (N_6237,N_5871,N_5647);
nand U6238 (N_6238,N_5934,N_5896);
xnor U6239 (N_6239,N_5927,N_5977);
and U6240 (N_6240,N_5859,N_5625);
nand U6241 (N_6241,N_5531,N_5973);
xor U6242 (N_6242,N_5791,N_5638);
and U6243 (N_6243,N_5719,N_5800);
nand U6244 (N_6244,N_5994,N_5705);
nor U6245 (N_6245,N_5634,N_5693);
xor U6246 (N_6246,N_5702,N_5523);
nand U6247 (N_6247,N_5684,N_5516);
nand U6248 (N_6248,N_5765,N_5564);
nor U6249 (N_6249,N_5609,N_5626);
nor U6250 (N_6250,N_5775,N_5630);
or U6251 (N_6251,N_5522,N_5556);
and U6252 (N_6252,N_5685,N_5705);
or U6253 (N_6253,N_5566,N_5931);
or U6254 (N_6254,N_5563,N_5801);
nor U6255 (N_6255,N_5790,N_5552);
nor U6256 (N_6256,N_5954,N_5893);
or U6257 (N_6257,N_5903,N_5617);
xnor U6258 (N_6258,N_5670,N_5788);
xnor U6259 (N_6259,N_5996,N_5543);
nand U6260 (N_6260,N_5882,N_5973);
or U6261 (N_6261,N_5557,N_5512);
nor U6262 (N_6262,N_5770,N_5873);
or U6263 (N_6263,N_5522,N_5963);
or U6264 (N_6264,N_5585,N_5759);
or U6265 (N_6265,N_5583,N_5594);
or U6266 (N_6266,N_5517,N_5731);
nand U6267 (N_6267,N_5919,N_5676);
or U6268 (N_6268,N_5917,N_5914);
and U6269 (N_6269,N_5850,N_5919);
and U6270 (N_6270,N_5828,N_5986);
xor U6271 (N_6271,N_5749,N_5890);
nand U6272 (N_6272,N_5842,N_5592);
or U6273 (N_6273,N_5711,N_5827);
or U6274 (N_6274,N_5649,N_5989);
or U6275 (N_6275,N_5686,N_5680);
and U6276 (N_6276,N_5844,N_5877);
nand U6277 (N_6277,N_5909,N_5832);
nor U6278 (N_6278,N_5768,N_5789);
and U6279 (N_6279,N_5837,N_5876);
nor U6280 (N_6280,N_5680,N_5522);
nand U6281 (N_6281,N_5945,N_5578);
xnor U6282 (N_6282,N_5682,N_5790);
or U6283 (N_6283,N_5971,N_5724);
nand U6284 (N_6284,N_5664,N_5697);
or U6285 (N_6285,N_5785,N_5512);
nor U6286 (N_6286,N_5728,N_5846);
and U6287 (N_6287,N_5691,N_5613);
xnor U6288 (N_6288,N_5775,N_5677);
and U6289 (N_6289,N_5824,N_5540);
nor U6290 (N_6290,N_5842,N_5548);
xor U6291 (N_6291,N_5525,N_5724);
xor U6292 (N_6292,N_5595,N_5735);
nand U6293 (N_6293,N_5755,N_5599);
and U6294 (N_6294,N_5685,N_5922);
or U6295 (N_6295,N_5589,N_5826);
nand U6296 (N_6296,N_5540,N_5649);
nand U6297 (N_6297,N_5751,N_5523);
or U6298 (N_6298,N_5740,N_5649);
or U6299 (N_6299,N_5536,N_5766);
nand U6300 (N_6300,N_5828,N_5923);
xor U6301 (N_6301,N_5668,N_5904);
nand U6302 (N_6302,N_5715,N_5567);
nand U6303 (N_6303,N_5998,N_5619);
and U6304 (N_6304,N_5774,N_5970);
nand U6305 (N_6305,N_5768,N_5653);
nand U6306 (N_6306,N_5650,N_5928);
and U6307 (N_6307,N_5887,N_5670);
nand U6308 (N_6308,N_5636,N_5558);
or U6309 (N_6309,N_5994,N_5795);
or U6310 (N_6310,N_5908,N_5652);
nand U6311 (N_6311,N_5913,N_5505);
and U6312 (N_6312,N_5729,N_5798);
nor U6313 (N_6313,N_5917,N_5990);
or U6314 (N_6314,N_5565,N_5915);
and U6315 (N_6315,N_5840,N_5555);
and U6316 (N_6316,N_5912,N_5965);
or U6317 (N_6317,N_5858,N_5928);
nor U6318 (N_6318,N_5756,N_5810);
and U6319 (N_6319,N_5570,N_5688);
nand U6320 (N_6320,N_5733,N_5608);
xor U6321 (N_6321,N_5510,N_5623);
or U6322 (N_6322,N_5648,N_5984);
xnor U6323 (N_6323,N_5649,N_5534);
nor U6324 (N_6324,N_5777,N_5879);
nand U6325 (N_6325,N_5842,N_5661);
or U6326 (N_6326,N_5507,N_5897);
xor U6327 (N_6327,N_5796,N_5991);
nand U6328 (N_6328,N_5528,N_5564);
and U6329 (N_6329,N_5563,N_5647);
or U6330 (N_6330,N_5985,N_5870);
or U6331 (N_6331,N_5961,N_5562);
nand U6332 (N_6332,N_5768,N_5953);
nor U6333 (N_6333,N_5747,N_5799);
or U6334 (N_6334,N_5691,N_5521);
or U6335 (N_6335,N_5627,N_5673);
nand U6336 (N_6336,N_5615,N_5502);
and U6337 (N_6337,N_5765,N_5648);
or U6338 (N_6338,N_5846,N_5768);
and U6339 (N_6339,N_5542,N_5512);
nor U6340 (N_6340,N_5608,N_5977);
and U6341 (N_6341,N_5558,N_5737);
or U6342 (N_6342,N_5744,N_5968);
nand U6343 (N_6343,N_5800,N_5551);
xnor U6344 (N_6344,N_5954,N_5505);
xor U6345 (N_6345,N_5644,N_5830);
and U6346 (N_6346,N_5583,N_5577);
and U6347 (N_6347,N_5548,N_5970);
nand U6348 (N_6348,N_5873,N_5512);
xnor U6349 (N_6349,N_5584,N_5891);
nor U6350 (N_6350,N_5704,N_5916);
and U6351 (N_6351,N_5658,N_5740);
xor U6352 (N_6352,N_5710,N_5539);
xor U6353 (N_6353,N_5640,N_5522);
nand U6354 (N_6354,N_5648,N_5706);
nand U6355 (N_6355,N_5809,N_5689);
nor U6356 (N_6356,N_5974,N_5918);
or U6357 (N_6357,N_5530,N_5604);
or U6358 (N_6358,N_5586,N_5568);
and U6359 (N_6359,N_5784,N_5677);
and U6360 (N_6360,N_5689,N_5601);
nor U6361 (N_6361,N_5679,N_5814);
and U6362 (N_6362,N_5893,N_5542);
or U6363 (N_6363,N_5655,N_5629);
and U6364 (N_6364,N_5653,N_5980);
nand U6365 (N_6365,N_5632,N_5583);
or U6366 (N_6366,N_5518,N_5983);
xor U6367 (N_6367,N_5915,N_5732);
or U6368 (N_6368,N_5919,N_5736);
nand U6369 (N_6369,N_5707,N_5501);
xor U6370 (N_6370,N_5991,N_5650);
or U6371 (N_6371,N_5598,N_5895);
nand U6372 (N_6372,N_5963,N_5705);
or U6373 (N_6373,N_5520,N_5917);
xnor U6374 (N_6374,N_5885,N_5793);
nand U6375 (N_6375,N_5777,N_5505);
nand U6376 (N_6376,N_5706,N_5788);
and U6377 (N_6377,N_5892,N_5907);
or U6378 (N_6378,N_5807,N_5824);
and U6379 (N_6379,N_5628,N_5755);
and U6380 (N_6380,N_5663,N_5653);
nor U6381 (N_6381,N_5975,N_5618);
nand U6382 (N_6382,N_5755,N_5705);
nand U6383 (N_6383,N_5682,N_5656);
and U6384 (N_6384,N_5785,N_5765);
nor U6385 (N_6385,N_5859,N_5795);
xor U6386 (N_6386,N_5790,N_5962);
nand U6387 (N_6387,N_5726,N_5684);
nand U6388 (N_6388,N_5583,N_5753);
nand U6389 (N_6389,N_5521,N_5577);
and U6390 (N_6390,N_5598,N_5722);
and U6391 (N_6391,N_5772,N_5876);
nor U6392 (N_6392,N_5834,N_5507);
xor U6393 (N_6393,N_5697,N_5699);
and U6394 (N_6394,N_5627,N_5803);
xor U6395 (N_6395,N_5791,N_5916);
nor U6396 (N_6396,N_5536,N_5638);
nand U6397 (N_6397,N_5691,N_5697);
nor U6398 (N_6398,N_5867,N_5906);
and U6399 (N_6399,N_5534,N_5869);
or U6400 (N_6400,N_5712,N_5894);
nand U6401 (N_6401,N_5872,N_5895);
and U6402 (N_6402,N_5843,N_5971);
nand U6403 (N_6403,N_5539,N_5964);
nor U6404 (N_6404,N_5707,N_5945);
xor U6405 (N_6405,N_5830,N_5678);
and U6406 (N_6406,N_5812,N_5934);
nand U6407 (N_6407,N_5688,N_5705);
xor U6408 (N_6408,N_5584,N_5718);
xor U6409 (N_6409,N_5618,N_5667);
or U6410 (N_6410,N_5926,N_5693);
nand U6411 (N_6411,N_5510,N_5796);
nor U6412 (N_6412,N_5841,N_5904);
nor U6413 (N_6413,N_5663,N_5645);
xnor U6414 (N_6414,N_5701,N_5534);
and U6415 (N_6415,N_5542,N_5572);
xnor U6416 (N_6416,N_5669,N_5802);
and U6417 (N_6417,N_5662,N_5720);
xor U6418 (N_6418,N_5931,N_5777);
xnor U6419 (N_6419,N_5505,N_5610);
xnor U6420 (N_6420,N_5611,N_5670);
nand U6421 (N_6421,N_5627,N_5823);
and U6422 (N_6422,N_5926,N_5990);
or U6423 (N_6423,N_5964,N_5995);
and U6424 (N_6424,N_5943,N_5744);
nand U6425 (N_6425,N_5629,N_5796);
xnor U6426 (N_6426,N_5651,N_5976);
and U6427 (N_6427,N_5903,N_5551);
nor U6428 (N_6428,N_5678,N_5895);
nand U6429 (N_6429,N_5953,N_5806);
and U6430 (N_6430,N_5781,N_5747);
nand U6431 (N_6431,N_5993,N_5765);
nand U6432 (N_6432,N_5794,N_5834);
nor U6433 (N_6433,N_5861,N_5798);
xnor U6434 (N_6434,N_5928,N_5535);
and U6435 (N_6435,N_5711,N_5685);
xor U6436 (N_6436,N_5645,N_5564);
and U6437 (N_6437,N_5611,N_5666);
or U6438 (N_6438,N_5673,N_5781);
xor U6439 (N_6439,N_5864,N_5646);
and U6440 (N_6440,N_5902,N_5989);
nand U6441 (N_6441,N_5927,N_5737);
nand U6442 (N_6442,N_5754,N_5922);
nand U6443 (N_6443,N_5882,N_5601);
nand U6444 (N_6444,N_5887,N_5775);
or U6445 (N_6445,N_5946,N_5977);
xor U6446 (N_6446,N_5662,N_5524);
nand U6447 (N_6447,N_5734,N_5597);
nor U6448 (N_6448,N_5508,N_5641);
xnor U6449 (N_6449,N_5996,N_5612);
nand U6450 (N_6450,N_5719,N_5784);
or U6451 (N_6451,N_5615,N_5862);
nand U6452 (N_6452,N_5701,N_5781);
or U6453 (N_6453,N_5710,N_5868);
and U6454 (N_6454,N_5605,N_5881);
and U6455 (N_6455,N_5502,N_5889);
or U6456 (N_6456,N_5562,N_5566);
and U6457 (N_6457,N_5731,N_5670);
nor U6458 (N_6458,N_5730,N_5814);
nand U6459 (N_6459,N_5609,N_5970);
or U6460 (N_6460,N_5574,N_5623);
or U6461 (N_6461,N_5589,N_5558);
nand U6462 (N_6462,N_5684,N_5686);
nand U6463 (N_6463,N_5650,N_5893);
nor U6464 (N_6464,N_5768,N_5976);
xnor U6465 (N_6465,N_5850,N_5601);
and U6466 (N_6466,N_5876,N_5677);
and U6467 (N_6467,N_5717,N_5790);
nor U6468 (N_6468,N_5895,N_5868);
nor U6469 (N_6469,N_5966,N_5926);
nand U6470 (N_6470,N_5670,N_5952);
nor U6471 (N_6471,N_5768,N_5799);
or U6472 (N_6472,N_5863,N_5571);
and U6473 (N_6473,N_5880,N_5635);
or U6474 (N_6474,N_5503,N_5662);
nand U6475 (N_6475,N_5992,N_5885);
and U6476 (N_6476,N_5508,N_5948);
or U6477 (N_6477,N_5834,N_5702);
and U6478 (N_6478,N_5802,N_5936);
or U6479 (N_6479,N_5885,N_5638);
xor U6480 (N_6480,N_5689,N_5883);
nor U6481 (N_6481,N_5550,N_5907);
nor U6482 (N_6482,N_5637,N_5727);
nand U6483 (N_6483,N_5842,N_5588);
or U6484 (N_6484,N_5876,N_5781);
nor U6485 (N_6485,N_5752,N_5975);
and U6486 (N_6486,N_5984,N_5947);
and U6487 (N_6487,N_5665,N_5836);
nand U6488 (N_6488,N_5848,N_5720);
nand U6489 (N_6489,N_5561,N_5504);
nand U6490 (N_6490,N_5807,N_5935);
nor U6491 (N_6491,N_5576,N_5670);
xor U6492 (N_6492,N_5686,N_5947);
xnor U6493 (N_6493,N_5514,N_5501);
or U6494 (N_6494,N_5626,N_5749);
xor U6495 (N_6495,N_5721,N_5508);
and U6496 (N_6496,N_5916,N_5909);
and U6497 (N_6497,N_5570,N_5603);
and U6498 (N_6498,N_5724,N_5735);
and U6499 (N_6499,N_5629,N_5616);
nand U6500 (N_6500,N_6148,N_6351);
xor U6501 (N_6501,N_6265,N_6444);
xor U6502 (N_6502,N_6258,N_6389);
or U6503 (N_6503,N_6217,N_6467);
and U6504 (N_6504,N_6150,N_6303);
xor U6505 (N_6505,N_6417,N_6474);
xor U6506 (N_6506,N_6005,N_6322);
nor U6507 (N_6507,N_6455,N_6093);
nand U6508 (N_6508,N_6026,N_6177);
and U6509 (N_6509,N_6229,N_6075);
xnor U6510 (N_6510,N_6050,N_6200);
nor U6511 (N_6511,N_6245,N_6252);
nand U6512 (N_6512,N_6375,N_6097);
and U6513 (N_6513,N_6248,N_6065);
xor U6514 (N_6514,N_6007,N_6418);
nor U6515 (N_6515,N_6355,N_6391);
xor U6516 (N_6516,N_6460,N_6191);
nand U6517 (N_6517,N_6227,N_6164);
or U6518 (N_6518,N_6115,N_6190);
xnor U6519 (N_6519,N_6379,N_6036);
nand U6520 (N_6520,N_6221,N_6222);
nor U6521 (N_6521,N_6223,N_6102);
nand U6522 (N_6522,N_6293,N_6399);
and U6523 (N_6523,N_6316,N_6071);
nor U6524 (N_6524,N_6041,N_6342);
xor U6525 (N_6525,N_6407,N_6367);
nand U6526 (N_6526,N_6319,N_6084);
xnor U6527 (N_6527,N_6108,N_6347);
xor U6528 (N_6528,N_6186,N_6392);
or U6529 (N_6529,N_6061,N_6482);
or U6530 (N_6530,N_6213,N_6263);
and U6531 (N_6531,N_6219,N_6178);
and U6532 (N_6532,N_6143,N_6487);
or U6533 (N_6533,N_6353,N_6453);
or U6534 (N_6534,N_6497,N_6088);
nor U6535 (N_6535,N_6017,N_6475);
xor U6536 (N_6536,N_6476,N_6411);
nor U6537 (N_6537,N_6030,N_6096);
and U6538 (N_6538,N_6390,N_6276);
nor U6539 (N_6539,N_6449,N_6033);
nand U6540 (N_6540,N_6037,N_6433);
nand U6541 (N_6541,N_6197,N_6428);
nor U6542 (N_6542,N_6042,N_6090);
or U6543 (N_6543,N_6127,N_6193);
nand U6544 (N_6544,N_6462,N_6220);
nor U6545 (N_6545,N_6268,N_6204);
and U6546 (N_6546,N_6404,N_6354);
nor U6547 (N_6547,N_6114,N_6098);
nor U6548 (N_6548,N_6381,N_6032);
and U6549 (N_6549,N_6110,N_6142);
nor U6550 (N_6550,N_6169,N_6066);
nand U6551 (N_6551,N_6400,N_6332);
or U6552 (N_6552,N_6287,N_6124);
nor U6553 (N_6553,N_6470,N_6405);
and U6554 (N_6554,N_6130,N_6483);
xnor U6555 (N_6555,N_6089,N_6380);
nor U6556 (N_6556,N_6166,N_6402);
or U6557 (N_6557,N_6410,N_6473);
nand U6558 (N_6558,N_6225,N_6207);
and U6559 (N_6559,N_6313,N_6366);
nand U6560 (N_6560,N_6239,N_6168);
and U6561 (N_6561,N_6255,N_6120);
or U6562 (N_6562,N_6145,N_6215);
nand U6563 (N_6563,N_6495,N_6446);
and U6564 (N_6564,N_6237,N_6009);
and U6565 (N_6565,N_6294,N_6363);
or U6566 (N_6566,N_6490,N_6049);
and U6567 (N_6567,N_6011,N_6288);
and U6568 (N_6568,N_6173,N_6365);
or U6569 (N_6569,N_6430,N_6253);
xor U6570 (N_6570,N_6279,N_6264);
nand U6571 (N_6571,N_6137,N_6373);
xnor U6572 (N_6572,N_6330,N_6095);
and U6573 (N_6573,N_6002,N_6238);
xor U6574 (N_6574,N_6496,N_6395);
xor U6575 (N_6575,N_6072,N_6165);
nor U6576 (N_6576,N_6329,N_6052);
nand U6577 (N_6577,N_6208,N_6458);
or U6578 (N_6578,N_6396,N_6284);
nor U6579 (N_6579,N_6249,N_6443);
xor U6580 (N_6580,N_6292,N_6076);
or U6581 (N_6581,N_6337,N_6004);
and U6582 (N_6582,N_6015,N_6226);
and U6583 (N_6583,N_6266,N_6104);
nor U6584 (N_6584,N_6256,N_6231);
and U6585 (N_6585,N_6172,N_6014);
and U6586 (N_6586,N_6118,N_6179);
or U6587 (N_6587,N_6408,N_6484);
xor U6588 (N_6588,N_6212,N_6086);
or U6589 (N_6589,N_6491,N_6358);
or U6590 (N_6590,N_6331,N_6016);
or U6591 (N_6591,N_6485,N_6370);
and U6592 (N_6592,N_6300,N_6421);
nand U6593 (N_6593,N_6304,N_6176);
nor U6594 (N_6594,N_6480,N_6243);
nor U6595 (N_6595,N_6378,N_6278);
nand U6596 (N_6596,N_6439,N_6461);
nand U6597 (N_6597,N_6286,N_6318);
nor U6598 (N_6598,N_6478,N_6083);
or U6599 (N_6599,N_6393,N_6105);
nand U6600 (N_6600,N_6295,N_6413);
and U6601 (N_6601,N_6498,N_6234);
nand U6602 (N_6602,N_6270,N_6335);
and U6603 (N_6603,N_6369,N_6385);
or U6604 (N_6604,N_6203,N_6113);
nand U6605 (N_6605,N_6472,N_6021);
nand U6606 (N_6606,N_6438,N_6181);
nand U6607 (N_6607,N_6261,N_6306);
nand U6608 (N_6608,N_6448,N_6028);
xnor U6609 (N_6609,N_6151,N_6336);
or U6610 (N_6610,N_6383,N_6019);
nand U6611 (N_6611,N_6057,N_6103);
nand U6612 (N_6612,N_6338,N_6274);
xor U6613 (N_6613,N_6250,N_6465);
and U6614 (N_6614,N_6003,N_6459);
nor U6615 (N_6615,N_6339,N_6324);
nor U6616 (N_6616,N_6427,N_6183);
or U6617 (N_6617,N_6236,N_6131);
nand U6618 (N_6618,N_6180,N_6326);
and U6619 (N_6619,N_6348,N_6488);
xor U6620 (N_6620,N_6209,N_6139);
xnor U6621 (N_6621,N_6122,N_6006);
xnor U6622 (N_6622,N_6437,N_6155);
or U6623 (N_6623,N_6244,N_6346);
and U6624 (N_6624,N_6377,N_6479);
xnor U6625 (N_6625,N_6285,N_6423);
or U6626 (N_6626,N_6386,N_6281);
and U6627 (N_6627,N_6419,N_6382);
and U6628 (N_6628,N_6357,N_6368);
and U6629 (N_6629,N_6218,N_6315);
nand U6630 (N_6630,N_6046,N_6040);
nand U6631 (N_6631,N_6328,N_6175);
nor U6632 (N_6632,N_6327,N_6343);
or U6633 (N_6633,N_6080,N_6211);
nor U6634 (N_6634,N_6224,N_6299);
nand U6635 (N_6635,N_6436,N_6384);
nor U6636 (N_6636,N_6305,N_6492);
and U6637 (N_6637,N_6262,N_6424);
nand U6638 (N_6638,N_6310,N_6152);
xnor U6639 (N_6639,N_6260,N_6128);
nand U6640 (N_6640,N_6356,N_6109);
xor U6641 (N_6641,N_6309,N_6056);
and U6642 (N_6642,N_6493,N_6149);
nor U6643 (N_6643,N_6070,N_6422);
or U6644 (N_6644,N_6297,N_6352);
nand U6645 (N_6645,N_6350,N_6162);
xor U6646 (N_6646,N_6325,N_6282);
and U6647 (N_6647,N_6311,N_6362);
nand U6648 (N_6648,N_6060,N_6216);
nand U6649 (N_6649,N_6018,N_6147);
and U6650 (N_6650,N_6290,N_6135);
nand U6651 (N_6651,N_6298,N_6468);
nor U6652 (N_6652,N_6447,N_6100);
xor U6653 (N_6653,N_6000,N_6029);
or U6654 (N_6654,N_6425,N_6398);
and U6655 (N_6655,N_6160,N_6321);
nor U6656 (N_6656,N_6451,N_6273);
nor U6657 (N_6657,N_6232,N_6235);
nor U6658 (N_6658,N_6129,N_6012);
nor U6659 (N_6659,N_6107,N_6055);
or U6660 (N_6660,N_6241,N_6196);
or U6661 (N_6661,N_6132,N_6140);
nor U6662 (N_6662,N_6457,N_6374);
nand U6663 (N_6663,N_6494,N_6116);
nor U6664 (N_6664,N_6117,N_6091);
nand U6665 (N_6665,N_6133,N_6008);
nor U6666 (N_6666,N_6141,N_6254);
nand U6667 (N_6667,N_6340,N_6189);
and U6668 (N_6668,N_6302,N_6240);
nor U6669 (N_6669,N_6228,N_6138);
xor U6670 (N_6670,N_6397,N_6442);
or U6671 (N_6671,N_6053,N_6077);
or U6672 (N_6672,N_6202,N_6199);
xnor U6673 (N_6673,N_6047,N_6412);
and U6674 (N_6674,N_6043,N_6210);
or U6675 (N_6675,N_6456,N_6187);
or U6676 (N_6676,N_6062,N_6296);
nand U6677 (N_6677,N_6074,N_6068);
nor U6678 (N_6678,N_6185,N_6415);
xor U6679 (N_6679,N_6058,N_6073);
and U6680 (N_6680,N_6136,N_6432);
xnor U6681 (N_6681,N_6092,N_6291);
xor U6682 (N_6682,N_6440,N_6161);
nor U6683 (N_6683,N_6201,N_6333);
nand U6684 (N_6684,N_6275,N_6101);
nand U6685 (N_6685,N_6174,N_6349);
nand U6686 (N_6686,N_6431,N_6010);
nor U6687 (N_6687,N_6360,N_6403);
xor U6688 (N_6688,N_6167,N_6481);
xor U6689 (N_6689,N_6361,N_6409);
nor U6690 (N_6690,N_6289,N_6020);
nand U6691 (N_6691,N_6054,N_6125);
nor U6692 (N_6692,N_6198,N_6163);
nand U6693 (N_6693,N_6454,N_6022);
xor U6694 (N_6694,N_6230,N_6341);
and U6695 (N_6695,N_6045,N_6119);
nor U6696 (N_6696,N_6394,N_6039);
or U6697 (N_6697,N_6182,N_6111);
or U6698 (N_6698,N_6123,N_6477);
or U6699 (N_6699,N_6320,N_6445);
xnor U6700 (N_6700,N_6112,N_6401);
nor U6701 (N_6701,N_6246,N_6450);
or U6702 (N_6702,N_6001,N_6038);
or U6703 (N_6703,N_6051,N_6027);
xor U6704 (N_6704,N_6146,N_6486);
xnor U6705 (N_6705,N_6023,N_6079);
and U6706 (N_6706,N_6171,N_6069);
and U6707 (N_6707,N_6156,N_6469);
and U6708 (N_6708,N_6452,N_6188);
nor U6709 (N_6709,N_6206,N_6371);
xnor U6710 (N_6710,N_6144,N_6416);
or U6711 (N_6711,N_6087,N_6471);
xor U6712 (N_6712,N_6434,N_6426);
xnor U6713 (N_6713,N_6345,N_6194);
and U6714 (N_6714,N_6184,N_6099);
or U6715 (N_6715,N_6158,N_6134);
nand U6716 (N_6716,N_6233,N_6205);
nand U6717 (N_6717,N_6344,N_6376);
nor U6718 (N_6718,N_6435,N_6242);
xnor U6719 (N_6719,N_6153,N_6359);
or U6720 (N_6720,N_6489,N_6271);
xnor U6721 (N_6721,N_6251,N_6121);
nor U6722 (N_6722,N_6406,N_6272);
nor U6723 (N_6723,N_6214,N_6283);
nand U6724 (N_6724,N_6024,N_6280);
and U6725 (N_6725,N_6308,N_6429);
nor U6726 (N_6726,N_6126,N_6388);
nor U6727 (N_6727,N_6466,N_6067);
nor U6728 (N_6728,N_6269,N_6301);
nor U6729 (N_6729,N_6034,N_6048);
xor U6730 (N_6730,N_6044,N_6307);
xnor U6731 (N_6731,N_6170,N_6463);
nor U6732 (N_6732,N_6157,N_6013);
xnor U6733 (N_6733,N_6094,N_6025);
or U6734 (N_6734,N_6078,N_6247);
and U6735 (N_6735,N_6192,N_6195);
nor U6736 (N_6736,N_6499,N_6031);
or U6737 (N_6737,N_6035,N_6372);
nor U6738 (N_6738,N_6159,N_6064);
and U6739 (N_6739,N_6464,N_6106);
nand U6740 (N_6740,N_6257,N_6323);
or U6741 (N_6741,N_6334,N_6317);
or U6742 (N_6742,N_6420,N_6441);
or U6743 (N_6743,N_6387,N_6312);
or U6744 (N_6744,N_6085,N_6277);
xnor U6745 (N_6745,N_6082,N_6314);
xnor U6746 (N_6746,N_6259,N_6364);
and U6747 (N_6747,N_6414,N_6059);
xor U6748 (N_6748,N_6063,N_6154);
nor U6749 (N_6749,N_6267,N_6081);
or U6750 (N_6750,N_6151,N_6143);
nor U6751 (N_6751,N_6430,N_6472);
nand U6752 (N_6752,N_6389,N_6298);
and U6753 (N_6753,N_6180,N_6268);
nor U6754 (N_6754,N_6202,N_6484);
and U6755 (N_6755,N_6317,N_6498);
and U6756 (N_6756,N_6292,N_6449);
or U6757 (N_6757,N_6426,N_6414);
or U6758 (N_6758,N_6353,N_6297);
xor U6759 (N_6759,N_6176,N_6109);
xnor U6760 (N_6760,N_6214,N_6381);
or U6761 (N_6761,N_6288,N_6358);
nand U6762 (N_6762,N_6130,N_6016);
xor U6763 (N_6763,N_6169,N_6305);
nor U6764 (N_6764,N_6077,N_6282);
nand U6765 (N_6765,N_6031,N_6289);
nand U6766 (N_6766,N_6457,N_6294);
or U6767 (N_6767,N_6088,N_6384);
nand U6768 (N_6768,N_6340,N_6164);
nand U6769 (N_6769,N_6253,N_6294);
xor U6770 (N_6770,N_6441,N_6414);
nand U6771 (N_6771,N_6290,N_6049);
or U6772 (N_6772,N_6009,N_6151);
nand U6773 (N_6773,N_6289,N_6382);
nand U6774 (N_6774,N_6042,N_6404);
or U6775 (N_6775,N_6321,N_6251);
nor U6776 (N_6776,N_6171,N_6211);
and U6777 (N_6777,N_6420,N_6134);
nand U6778 (N_6778,N_6421,N_6194);
and U6779 (N_6779,N_6085,N_6366);
and U6780 (N_6780,N_6009,N_6128);
and U6781 (N_6781,N_6410,N_6353);
xnor U6782 (N_6782,N_6085,N_6144);
nor U6783 (N_6783,N_6219,N_6193);
and U6784 (N_6784,N_6214,N_6195);
or U6785 (N_6785,N_6478,N_6130);
nor U6786 (N_6786,N_6273,N_6042);
xor U6787 (N_6787,N_6024,N_6026);
xnor U6788 (N_6788,N_6284,N_6420);
nor U6789 (N_6789,N_6386,N_6046);
or U6790 (N_6790,N_6284,N_6345);
and U6791 (N_6791,N_6005,N_6393);
nor U6792 (N_6792,N_6492,N_6182);
nand U6793 (N_6793,N_6037,N_6305);
nor U6794 (N_6794,N_6270,N_6443);
nand U6795 (N_6795,N_6119,N_6261);
or U6796 (N_6796,N_6493,N_6073);
nor U6797 (N_6797,N_6161,N_6384);
nor U6798 (N_6798,N_6308,N_6033);
nor U6799 (N_6799,N_6350,N_6466);
nor U6800 (N_6800,N_6131,N_6289);
nand U6801 (N_6801,N_6231,N_6068);
or U6802 (N_6802,N_6033,N_6361);
nor U6803 (N_6803,N_6111,N_6411);
nand U6804 (N_6804,N_6498,N_6000);
nor U6805 (N_6805,N_6271,N_6095);
xor U6806 (N_6806,N_6210,N_6202);
xnor U6807 (N_6807,N_6106,N_6204);
and U6808 (N_6808,N_6061,N_6248);
or U6809 (N_6809,N_6233,N_6132);
or U6810 (N_6810,N_6138,N_6183);
nand U6811 (N_6811,N_6371,N_6254);
and U6812 (N_6812,N_6230,N_6153);
and U6813 (N_6813,N_6019,N_6332);
xnor U6814 (N_6814,N_6147,N_6062);
and U6815 (N_6815,N_6421,N_6457);
or U6816 (N_6816,N_6316,N_6058);
nand U6817 (N_6817,N_6227,N_6112);
and U6818 (N_6818,N_6424,N_6055);
or U6819 (N_6819,N_6307,N_6009);
and U6820 (N_6820,N_6151,N_6459);
nand U6821 (N_6821,N_6451,N_6403);
or U6822 (N_6822,N_6491,N_6308);
and U6823 (N_6823,N_6432,N_6034);
nor U6824 (N_6824,N_6061,N_6352);
nor U6825 (N_6825,N_6140,N_6011);
nand U6826 (N_6826,N_6167,N_6166);
or U6827 (N_6827,N_6298,N_6101);
or U6828 (N_6828,N_6009,N_6065);
or U6829 (N_6829,N_6456,N_6123);
or U6830 (N_6830,N_6343,N_6152);
xnor U6831 (N_6831,N_6105,N_6404);
or U6832 (N_6832,N_6278,N_6144);
nor U6833 (N_6833,N_6091,N_6278);
nand U6834 (N_6834,N_6408,N_6132);
nand U6835 (N_6835,N_6332,N_6447);
nor U6836 (N_6836,N_6231,N_6455);
or U6837 (N_6837,N_6152,N_6132);
xnor U6838 (N_6838,N_6113,N_6460);
and U6839 (N_6839,N_6240,N_6164);
and U6840 (N_6840,N_6130,N_6112);
and U6841 (N_6841,N_6416,N_6419);
or U6842 (N_6842,N_6068,N_6146);
or U6843 (N_6843,N_6318,N_6254);
xor U6844 (N_6844,N_6471,N_6113);
xor U6845 (N_6845,N_6438,N_6468);
nor U6846 (N_6846,N_6231,N_6108);
nor U6847 (N_6847,N_6166,N_6397);
xor U6848 (N_6848,N_6468,N_6010);
and U6849 (N_6849,N_6292,N_6497);
nor U6850 (N_6850,N_6355,N_6157);
nand U6851 (N_6851,N_6322,N_6307);
or U6852 (N_6852,N_6458,N_6014);
and U6853 (N_6853,N_6021,N_6263);
and U6854 (N_6854,N_6225,N_6413);
and U6855 (N_6855,N_6246,N_6167);
nand U6856 (N_6856,N_6190,N_6246);
nand U6857 (N_6857,N_6340,N_6348);
and U6858 (N_6858,N_6049,N_6144);
xnor U6859 (N_6859,N_6371,N_6311);
xor U6860 (N_6860,N_6208,N_6283);
or U6861 (N_6861,N_6382,N_6108);
nand U6862 (N_6862,N_6469,N_6060);
or U6863 (N_6863,N_6019,N_6099);
nand U6864 (N_6864,N_6460,N_6346);
xor U6865 (N_6865,N_6166,N_6015);
xor U6866 (N_6866,N_6034,N_6212);
xnor U6867 (N_6867,N_6115,N_6278);
and U6868 (N_6868,N_6362,N_6384);
nor U6869 (N_6869,N_6366,N_6287);
nor U6870 (N_6870,N_6479,N_6032);
xnor U6871 (N_6871,N_6035,N_6271);
or U6872 (N_6872,N_6400,N_6263);
or U6873 (N_6873,N_6247,N_6129);
xnor U6874 (N_6874,N_6293,N_6046);
or U6875 (N_6875,N_6377,N_6171);
nor U6876 (N_6876,N_6385,N_6177);
or U6877 (N_6877,N_6448,N_6361);
xor U6878 (N_6878,N_6058,N_6389);
xnor U6879 (N_6879,N_6272,N_6409);
xnor U6880 (N_6880,N_6240,N_6439);
nor U6881 (N_6881,N_6171,N_6174);
nor U6882 (N_6882,N_6471,N_6103);
or U6883 (N_6883,N_6448,N_6014);
and U6884 (N_6884,N_6048,N_6397);
nand U6885 (N_6885,N_6378,N_6439);
nand U6886 (N_6886,N_6133,N_6099);
and U6887 (N_6887,N_6041,N_6137);
nand U6888 (N_6888,N_6228,N_6447);
nor U6889 (N_6889,N_6082,N_6401);
or U6890 (N_6890,N_6289,N_6137);
xor U6891 (N_6891,N_6469,N_6187);
nor U6892 (N_6892,N_6354,N_6124);
xnor U6893 (N_6893,N_6363,N_6498);
nand U6894 (N_6894,N_6340,N_6476);
nand U6895 (N_6895,N_6177,N_6070);
nor U6896 (N_6896,N_6116,N_6087);
or U6897 (N_6897,N_6347,N_6354);
xnor U6898 (N_6898,N_6139,N_6466);
nor U6899 (N_6899,N_6491,N_6259);
nand U6900 (N_6900,N_6111,N_6484);
xnor U6901 (N_6901,N_6301,N_6008);
and U6902 (N_6902,N_6360,N_6140);
and U6903 (N_6903,N_6188,N_6306);
or U6904 (N_6904,N_6483,N_6017);
and U6905 (N_6905,N_6366,N_6166);
or U6906 (N_6906,N_6465,N_6449);
or U6907 (N_6907,N_6260,N_6116);
xnor U6908 (N_6908,N_6424,N_6052);
or U6909 (N_6909,N_6115,N_6145);
or U6910 (N_6910,N_6330,N_6127);
or U6911 (N_6911,N_6378,N_6090);
nor U6912 (N_6912,N_6262,N_6082);
xor U6913 (N_6913,N_6471,N_6116);
nand U6914 (N_6914,N_6207,N_6491);
or U6915 (N_6915,N_6047,N_6333);
or U6916 (N_6916,N_6490,N_6093);
nor U6917 (N_6917,N_6221,N_6258);
xnor U6918 (N_6918,N_6344,N_6225);
or U6919 (N_6919,N_6139,N_6245);
and U6920 (N_6920,N_6106,N_6097);
nand U6921 (N_6921,N_6138,N_6355);
nor U6922 (N_6922,N_6457,N_6082);
or U6923 (N_6923,N_6099,N_6410);
nor U6924 (N_6924,N_6373,N_6091);
nand U6925 (N_6925,N_6437,N_6311);
nand U6926 (N_6926,N_6284,N_6045);
xor U6927 (N_6927,N_6227,N_6426);
and U6928 (N_6928,N_6490,N_6128);
or U6929 (N_6929,N_6027,N_6427);
xor U6930 (N_6930,N_6376,N_6054);
nand U6931 (N_6931,N_6031,N_6376);
nand U6932 (N_6932,N_6276,N_6286);
or U6933 (N_6933,N_6462,N_6399);
or U6934 (N_6934,N_6413,N_6066);
and U6935 (N_6935,N_6389,N_6379);
nand U6936 (N_6936,N_6381,N_6112);
xnor U6937 (N_6937,N_6245,N_6207);
xor U6938 (N_6938,N_6107,N_6404);
xnor U6939 (N_6939,N_6457,N_6186);
or U6940 (N_6940,N_6260,N_6498);
nand U6941 (N_6941,N_6471,N_6042);
nand U6942 (N_6942,N_6025,N_6313);
or U6943 (N_6943,N_6339,N_6184);
nor U6944 (N_6944,N_6197,N_6144);
and U6945 (N_6945,N_6063,N_6319);
xnor U6946 (N_6946,N_6404,N_6014);
nor U6947 (N_6947,N_6447,N_6044);
nand U6948 (N_6948,N_6023,N_6412);
or U6949 (N_6949,N_6445,N_6004);
nand U6950 (N_6950,N_6023,N_6375);
xor U6951 (N_6951,N_6041,N_6328);
nand U6952 (N_6952,N_6472,N_6404);
xnor U6953 (N_6953,N_6331,N_6137);
xor U6954 (N_6954,N_6097,N_6060);
or U6955 (N_6955,N_6252,N_6071);
or U6956 (N_6956,N_6130,N_6073);
or U6957 (N_6957,N_6299,N_6121);
nand U6958 (N_6958,N_6302,N_6126);
nand U6959 (N_6959,N_6053,N_6489);
and U6960 (N_6960,N_6494,N_6227);
or U6961 (N_6961,N_6227,N_6296);
or U6962 (N_6962,N_6369,N_6485);
and U6963 (N_6963,N_6485,N_6128);
and U6964 (N_6964,N_6305,N_6429);
nor U6965 (N_6965,N_6388,N_6072);
xnor U6966 (N_6966,N_6476,N_6179);
nand U6967 (N_6967,N_6263,N_6487);
xor U6968 (N_6968,N_6346,N_6005);
nand U6969 (N_6969,N_6150,N_6286);
or U6970 (N_6970,N_6030,N_6298);
nor U6971 (N_6971,N_6060,N_6262);
and U6972 (N_6972,N_6013,N_6179);
or U6973 (N_6973,N_6310,N_6008);
and U6974 (N_6974,N_6061,N_6234);
xor U6975 (N_6975,N_6476,N_6178);
or U6976 (N_6976,N_6469,N_6033);
and U6977 (N_6977,N_6336,N_6142);
or U6978 (N_6978,N_6304,N_6147);
nor U6979 (N_6979,N_6461,N_6186);
or U6980 (N_6980,N_6369,N_6219);
nand U6981 (N_6981,N_6446,N_6488);
and U6982 (N_6982,N_6364,N_6141);
xnor U6983 (N_6983,N_6185,N_6364);
nor U6984 (N_6984,N_6370,N_6450);
nand U6985 (N_6985,N_6244,N_6353);
xor U6986 (N_6986,N_6392,N_6126);
or U6987 (N_6987,N_6027,N_6103);
nand U6988 (N_6988,N_6404,N_6296);
or U6989 (N_6989,N_6463,N_6462);
or U6990 (N_6990,N_6435,N_6236);
and U6991 (N_6991,N_6402,N_6134);
nand U6992 (N_6992,N_6301,N_6001);
or U6993 (N_6993,N_6334,N_6115);
or U6994 (N_6994,N_6069,N_6119);
and U6995 (N_6995,N_6075,N_6200);
and U6996 (N_6996,N_6226,N_6140);
nor U6997 (N_6997,N_6343,N_6232);
xor U6998 (N_6998,N_6320,N_6425);
nand U6999 (N_6999,N_6248,N_6252);
nand U7000 (N_7000,N_6760,N_6854);
or U7001 (N_7001,N_6720,N_6953);
or U7002 (N_7002,N_6729,N_6727);
nor U7003 (N_7003,N_6748,N_6965);
nor U7004 (N_7004,N_6690,N_6895);
nand U7005 (N_7005,N_6933,N_6691);
and U7006 (N_7006,N_6809,N_6635);
xnor U7007 (N_7007,N_6581,N_6761);
or U7008 (N_7008,N_6559,N_6592);
and U7009 (N_7009,N_6700,N_6603);
nor U7010 (N_7010,N_6697,N_6715);
nand U7011 (N_7011,N_6949,N_6689);
and U7012 (N_7012,N_6679,N_6529);
nand U7013 (N_7013,N_6756,N_6923);
and U7014 (N_7014,N_6580,N_6627);
and U7015 (N_7015,N_6901,N_6537);
xor U7016 (N_7016,N_6911,N_6544);
nand U7017 (N_7017,N_6740,N_6978);
nand U7018 (N_7018,N_6710,N_6881);
nor U7019 (N_7019,N_6833,N_6902);
and U7020 (N_7020,N_6670,N_6738);
and U7021 (N_7021,N_6565,N_6775);
nor U7022 (N_7022,N_6822,N_6730);
or U7023 (N_7023,N_6878,N_6557);
and U7024 (N_7024,N_6575,N_6677);
nand U7025 (N_7025,N_6708,N_6747);
or U7026 (N_7026,N_6594,N_6617);
nand U7027 (N_7027,N_6863,N_6905);
nor U7028 (N_7028,N_6610,N_6801);
xor U7029 (N_7029,N_6543,N_6716);
nand U7030 (N_7030,N_6922,N_6515);
or U7031 (N_7031,N_6717,N_6947);
xor U7032 (N_7032,N_6969,N_6852);
nand U7033 (N_7033,N_6526,N_6850);
and U7034 (N_7034,N_6551,N_6624);
and U7035 (N_7035,N_6958,N_6796);
or U7036 (N_7036,N_6636,N_6893);
nand U7037 (N_7037,N_6799,N_6827);
and U7038 (N_7038,N_6577,N_6997);
nor U7039 (N_7039,N_6582,N_6899);
or U7040 (N_7040,N_6642,N_6841);
or U7041 (N_7041,N_6814,N_6973);
nor U7042 (N_7042,N_6566,N_6888);
nor U7043 (N_7043,N_6563,N_6510);
nor U7044 (N_7044,N_6558,N_6797);
xnor U7045 (N_7045,N_6573,N_6767);
and U7046 (N_7046,N_6678,N_6823);
nor U7047 (N_7047,N_6737,N_6979);
nor U7048 (N_7048,N_6793,N_6994);
xnor U7049 (N_7049,N_6591,N_6751);
and U7050 (N_7050,N_6641,N_6638);
xnor U7051 (N_7051,N_6886,N_6934);
nor U7052 (N_7052,N_6671,N_6988);
nor U7053 (N_7053,N_6987,N_6507);
xnor U7054 (N_7054,N_6567,N_6866);
xnor U7055 (N_7055,N_6948,N_6877);
nand U7056 (N_7056,N_6693,N_6906);
and U7057 (N_7057,N_6935,N_6532);
and U7058 (N_7058,N_6658,N_6839);
and U7059 (N_7059,N_6889,N_6601);
nand U7060 (N_7060,N_6649,N_6726);
xor U7061 (N_7061,N_6596,N_6625);
nand U7062 (N_7062,N_6910,N_6813);
and U7063 (N_7063,N_6882,N_6876);
xor U7064 (N_7064,N_6540,N_6849);
and U7065 (N_7065,N_6908,N_6640);
and U7066 (N_7066,N_6611,N_6860);
nand U7067 (N_7067,N_6622,N_6890);
and U7068 (N_7068,N_6916,N_6811);
or U7069 (N_7069,N_6946,N_6976);
and U7070 (N_7070,N_6986,N_6840);
or U7071 (N_7071,N_6778,N_6975);
nand U7072 (N_7072,N_6518,N_6776);
or U7073 (N_7073,N_6912,N_6696);
nand U7074 (N_7074,N_6541,N_6629);
nand U7075 (N_7075,N_6735,N_6616);
nor U7076 (N_7076,N_6817,N_6921);
or U7077 (N_7077,N_6909,N_6780);
or U7078 (N_7078,N_6755,N_6673);
nor U7079 (N_7079,N_6523,N_6661);
nor U7080 (N_7080,N_6539,N_6856);
or U7081 (N_7081,N_6746,N_6790);
nand U7082 (N_7082,N_6545,N_6682);
nand U7083 (N_7083,N_6648,N_6514);
or U7084 (N_7084,N_6578,N_6571);
or U7085 (N_7085,N_6504,N_6595);
or U7086 (N_7086,N_6651,N_6762);
xor U7087 (N_7087,N_6675,N_6590);
xor U7088 (N_7088,N_6961,N_6832);
xor U7089 (N_7089,N_6552,N_6844);
xnor U7090 (N_7090,N_6692,N_6728);
xnor U7091 (N_7091,N_6546,N_6859);
and U7092 (N_7092,N_6868,N_6531);
xnor U7093 (N_7093,N_6954,N_6894);
nor U7094 (N_7094,N_6875,N_6530);
xor U7095 (N_7095,N_6614,N_6957);
nand U7096 (N_7096,N_6956,N_6588);
nand U7097 (N_7097,N_6794,N_6574);
nand U7098 (N_7098,N_6904,N_6597);
nand U7099 (N_7099,N_6655,N_6572);
nand U7100 (N_7100,N_6681,N_6535);
nand U7101 (N_7101,N_6712,N_6533);
or U7102 (N_7102,N_6970,N_6645);
and U7103 (N_7103,N_6963,N_6869);
xor U7104 (N_7104,N_6966,N_6960);
or U7105 (N_7105,N_6699,N_6656);
xor U7106 (N_7106,N_6620,N_6952);
nand U7107 (N_7107,N_6950,N_6806);
xor U7108 (N_7108,N_6607,N_6634);
xnor U7109 (N_7109,N_6538,N_6672);
or U7110 (N_7110,N_6884,N_6632);
nand U7111 (N_7111,N_6847,N_6600);
nand U7112 (N_7112,N_6802,N_6937);
xnor U7113 (N_7113,N_6785,N_6550);
or U7114 (N_7114,N_6944,N_6606);
nand U7115 (N_7115,N_6722,N_6668);
xor U7116 (N_7116,N_6913,N_6808);
nand U7117 (N_7117,N_6825,N_6613);
xor U7118 (N_7118,N_6653,N_6993);
nor U7119 (N_7119,N_6773,N_6804);
and U7120 (N_7120,N_6818,N_6660);
xor U7121 (N_7121,N_6664,N_6500);
nand U7122 (N_7122,N_6665,N_6974);
or U7123 (N_7123,N_6967,N_6917);
or U7124 (N_7124,N_6501,N_6983);
nor U7125 (N_7125,N_6652,N_6851);
xor U7126 (N_7126,N_6891,N_6765);
or U7127 (N_7127,N_6907,N_6705);
and U7128 (N_7128,N_6807,N_6867);
xnor U7129 (N_7129,N_6945,N_6900);
and U7130 (N_7130,N_6619,N_6879);
or U7131 (N_7131,N_6734,N_6980);
nor U7132 (N_7132,N_6770,N_6828);
xor U7133 (N_7133,N_6897,N_6824);
nor U7134 (N_7134,N_6742,N_6659);
nand U7135 (N_7135,N_6861,N_6512);
and U7136 (N_7136,N_6731,N_6657);
nor U7137 (N_7137,N_6528,N_6522);
and U7138 (N_7138,N_6815,N_6609);
nor U7139 (N_7139,N_6995,N_6676);
nor U7140 (N_7140,N_6812,N_6569);
and U7141 (N_7141,N_6741,N_6783);
or U7142 (N_7142,N_6930,N_6749);
nand U7143 (N_7143,N_6633,N_6576);
and U7144 (N_7144,N_6752,N_6745);
nor U7145 (N_7145,N_6714,N_6766);
nor U7146 (N_7146,N_6598,N_6647);
nand U7147 (N_7147,N_6803,N_6626);
xor U7148 (N_7148,N_6618,N_6781);
or U7149 (N_7149,N_6939,N_6685);
nand U7150 (N_7150,N_6709,N_6768);
xor U7151 (N_7151,N_6608,N_6789);
nor U7152 (N_7152,N_6556,N_6848);
nor U7153 (N_7153,N_6962,N_6846);
nand U7154 (N_7154,N_6564,N_6758);
or U7155 (N_7155,N_6943,N_6643);
xnor U7156 (N_7156,N_6985,N_6732);
nor U7157 (N_7157,N_6542,N_6777);
xnor U7158 (N_7158,N_6570,N_6586);
and U7159 (N_7159,N_6703,N_6555);
xor U7160 (N_7160,N_6662,N_6628);
nand U7161 (N_7161,N_6991,N_6516);
nor U7162 (N_7162,N_6724,N_6694);
nor U7163 (N_7163,N_6631,N_6654);
or U7164 (N_7164,N_6560,N_6666);
or U7165 (N_7165,N_6830,N_6887);
and U7166 (N_7166,N_6981,N_6800);
nor U7167 (N_7167,N_6561,N_6896);
xor U7168 (N_7168,N_6562,N_6763);
xnor U7169 (N_7169,N_6733,N_6698);
or U7170 (N_7170,N_6585,N_6880);
nor U7171 (N_7171,N_6502,N_6810);
xor U7172 (N_7172,N_6513,N_6924);
xor U7173 (N_7173,N_6621,N_6999);
or U7174 (N_7174,N_6547,N_6713);
xnor U7175 (N_7175,N_6787,N_6680);
xnor U7176 (N_7176,N_6862,N_6707);
nor U7177 (N_7177,N_6831,N_6858);
and U7178 (N_7178,N_6989,N_6990);
and U7179 (N_7179,N_6864,N_6927);
or U7180 (N_7180,N_6926,N_6554);
nor U7181 (N_7181,N_6898,N_6834);
or U7182 (N_7182,N_6721,N_6941);
nand U7183 (N_7183,N_6764,N_6805);
or U7184 (N_7184,N_6589,N_6769);
nor U7185 (N_7185,N_6644,N_6826);
nand U7186 (N_7186,N_6599,N_6968);
xor U7187 (N_7187,N_6593,N_6838);
nor U7188 (N_7188,N_6548,N_6669);
or U7189 (N_7189,N_6524,N_6754);
nand U7190 (N_7190,N_6646,N_6885);
and U7191 (N_7191,N_6929,N_6959);
and U7192 (N_7192,N_6798,N_6719);
xnor U7193 (N_7193,N_6931,N_6744);
nor U7194 (N_7194,N_6568,N_6736);
or U7195 (N_7195,N_6503,N_6883);
nand U7196 (N_7196,N_6602,N_6955);
xnor U7197 (N_7197,N_6753,N_6845);
nand U7198 (N_7198,N_6505,N_6871);
xnor U7199 (N_7199,N_6938,N_6820);
or U7200 (N_7200,N_6639,N_6772);
nand U7201 (N_7201,N_6704,N_6982);
nor U7202 (N_7202,N_6816,N_6992);
nand U7203 (N_7203,N_6612,N_6914);
nor U7204 (N_7204,N_6795,N_6873);
nand U7205 (N_7205,N_6527,N_6759);
xor U7206 (N_7206,N_6872,N_6821);
nand U7207 (N_7207,N_6604,N_6553);
and U7208 (N_7208,N_6792,N_6837);
xnor U7209 (N_7209,N_6637,N_6774);
nand U7210 (N_7210,N_6951,N_6791);
nand U7211 (N_7211,N_6743,N_6865);
nor U7212 (N_7212,N_6757,N_6701);
and U7213 (N_7213,N_6525,N_6725);
and U7214 (N_7214,N_6788,N_6605);
and U7215 (N_7215,N_6684,N_6892);
nor U7216 (N_7216,N_6920,N_6579);
xor U7217 (N_7217,N_6819,N_6786);
or U7218 (N_7218,N_6857,N_6519);
nand U7219 (N_7219,N_6936,N_6686);
xnor U7220 (N_7220,N_6750,N_6506);
and U7221 (N_7221,N_6509,N_6843);
nand U7222 (N_7222,N_6964,N_6663);
nand U7223 (N_7223,N_6919,N_6903);
and U7224 (N_7224,N_6855,N_6771);
and U7225 (N_7225,N_6695,N_6998);
xor U7226 (N_7226,N_6842,N_6549);
and U7227 (N_7227,N_6711,N_6942);
and U7228 (N_7228,N_6784,N_6702);
xnor U7229 (N_7229,N_6674,N_6996);
xnor U7230 (N_7230,N_6932,N_6940);
nand U7231 (N_7231,N_6683,N_6874);
and U7232 (N_7232,N_6971,N_6984);
and U7233 (N_7233,N_6623,N_6667);
xnor U7234 (N_7234,N_6521,N_6915);
xnor U7235 (N_7235,N_6853,N_6918);
and U7236 (N_7236,N_6782,N_6511);
nor U7237 (N_7237,N_6587,N_6520);
and U7238 (N_7238,N_6536,N_6584);
nor U7239 (N_7239,N_6650,N_6517);
and U7240 (N_7240,N_6836,N_6583);
or U7241 (N_7241,N_6835,N_6829);
or U7242 (N_7242,N_6688,N_6687);
nor U7243 (N_7243,N_6870,N_6718);
nand U7244 (N_7244,N_6972,N_6534);
xor U7245 (N_7245,N_6928,N_6925);
xnor U7246 (N_7246,N_6630,N_6779);
nand U7247 (N_7247,N_6723,N_6977);
or U7248 (N_7248,N_6615,N_6739);
xor U7249 (N_7249,N_6706,N_6508);
nor U7250 (N_7250,N_6912,N_6734);
nand U7251 (N_7251,N_6632,N_6811);
xor U7252 (N_7252,N_6653,N_6726);
xnor U7253 (N_7253,N_6737,N_6746);
nand U7254 (N_7254,N_6541,N_6993);
xnor U7255 (N_7255,N_6635,N_6897);
xnor U7256 (N_7256,N_6991,N_6593);
or U7257 (N_7257,N_6837,N_6731);
or U7258 (N_7258,N_6892,N_6999);
nand U7259 (N_7259,N_6595,N_6862);
nand U7260 (N_7260,N_6745,N_6896);
and U7261 (N_7261,N_6544,N_6718);
and U7262 (N_7262,N_6751,N_6682);
nand U7263 (N_7263,N_6657,N_6966);
and U7264 (N_7264,N_6614,N_6589);
nand U7265 (N_7265,N_6687,N_6831);
xor U7266 (N_7266,N_6770,N_6889);
and U7267 (N_7267,N_6521,N_6841);
nand U7268 (N_7268,N_6905,N_6903);
nor U7269 (N_7269,N_6568,N_6939);
nor U7270 (N_7270,N_6850,N_6905);
or U7271 (N_7271,N_6891,N_6561);
and U7272 (N_7272,N_6719,N_6855);
or U7273 (N_7273,N_6980,N_6609);
or U7274 (N_7274,N_6891,N_6552);
xnor U7275 (N_7275,N_6515,N_6914);
nand U7276 (N_7276,N_6730,N_6748);
xor U7277 (N_7277,N_6504,N_6536);
and U7278 (N_7278,N_6819,N_6790);
nand U7279 (N_7279,N_6750,N_6501);
nor U7280 (N_7280,N_6798,N_6636);
or U7281 (N_7281,N_6641,N_6978);
or U7282 (N_7282,N_6787,N_6912);
or U7283 (N_7283,N_6677,N_6753);
xnor U7284 (N_7284,N_6563,N_6964);
nor U7285 (N_7285,N_6588,N_6697);
and U7286 (N_7286,N_6648,N_6704);
xnor U7287 (N_7287,N_6936,N_6811);
or U7288 (N_7288,N_6527,N_6760);
or U7289 (N_7289,N_6800,N_6524);
nand U7290 (N_7290,N_6566,N_6545);
and U7291 (N_7291,N_6999,N_6544);
and U7292 (N_7292,N_6931,N_6641);
xor U7293 (N_7293,N_6923,N_6758);
and U7294 (N_7294,N_6618,N_6613);
nor U7295 (N_7295,N_6640,N_6792);
and U7296 (N_7296,N_6960,N_6672);
xor U7297 (N_7297,N_6683,N_6628);
nor U7298 (N_7298,N_6934,N_6520);
or U7299 (N_7299,N_6874,N_6703);
and U7300 (N_7300,N_6908,N_6887);
xor U7301 (N_7301,N_6757,N_6673);
and U7302 (N_7302,N_6848,N_6963);
and U7303 (N_7303,N_6543,N_6774);
and U7304 (N_7304,N_6936,N_6712);
and U7305 (N_7305,N_6545,N_6915);
xnor U7306 (N_7306,N_6586,N_6779);
nor U7307 (N_7307,N_6703,N_6623);
or U7308 (N_7308,N_6820,N_6861);
nor U7309 (N_7309,N_6847,N_6666);
xnor U7310 (N_7310,N_6502,N_6873);
xnor U7311 (N_7311,N_6773,N_6989);
nor U7312 (N_7312,N_6522,N_6526);
nor U7313 (N_7313,N_6892,N_6564);
nand U7314 (N_7314,N_6929,N_6886);
xnor U7315 (N_7315,N_6780,N_6659);
nand U7316 (N_7316,N_6888,N_6917);
xor U7317 (N_7317,N_6541,N_6536);
nand U7318 (N_7318,N_6722,N_6931);
or U7319 (N_7319,N_6615,N_6994);
nand U7320 (N_7320,N_6961,N_6555);
and U7321 (N_7321,N_6816,N_6921);
nand U7322 (N_7322,N_6648,N_6991);
or U7323 (N_7323,N_6963,N_6763);
or U7324 (N_7324,N_6934,N_6698);
xor U7325 (N_7325,N_6920,N_6795);
nand U7326 (N_7326,N_6574,N_6917);
nand U7327 (N_7327,N_6786,N_6723);
nor U7328 (N_7328,N_6535,N_6671);
or U7329 (N_7329,N_6941,N_6854);
nor U7330 (N_7330,N_6816,N_6769);
or U7331 (N_7331,N_6745,N_6633);
and U7332 (N_7332,N_6535,N_6884);
nor U7333 (N_7333,N_6535,N_6502);
xnor U7334 (N_7334,N_6934,N_6969);
nand U7335 (N_7335,N_6650,N_6866);
nand U7336 (N_7336,N_6799,N_6531);
xnor U7337 (N_7337,N_6556,N_6513);
nand U7338 (N_7338,N_6536,N_6961);
and U7339 (N_7339,N_6507,N_6961);
and U7340 (N_7340,N_6711,N_6998);
nor U7341 (N_7341,N_6962,N_6786);
xor U7342 (N_7342,N_6896,N_6514);
nand U7343 (N_7343,N_6595,N_6583);
or U7344 (N_7344,N_6881,N_6714);
nor U7345 (N_7345,N_6619,N_6649);
and U7346 (N_7346,N_6571,N_6641);
nand U7347 (N_7347,N_6636,N_6652);
or U7348 (N_7348,N_6928,N_6529);
nor U7349 (N_7349,N_6551,N_6517);
nand U7350 (N_7350,N_6605,N_6738);
or U7351 (N_7351,N_6569,N_6558);
or U7352 (N_7352,N_6982,N_6680);
xor U7353 (N_7353,N_6701,N_6912);
nand U7354 (N_7354,N_6649,N_6797);
or U7355 (N_7355,N_6566,N_6861);
nor U7356 (N_7356,N_6635,N_6719);
and U7357 (N_7357,N_6885,N_6888);
nor U7358 (N_7358,N_6610,N_6999);
xnor U7359 (N_7359,N_6927,N_6784);
nor U7360 (N_7360,N_6966,N_6760);
nand U7361 (N_7361,N_6927,N_6509);
nor U7362 (N_7362,N_6594,N_6985);
xor U7363 (N_7363,N_6551,N_6594);
and U7364 (N_7364,N_6911,N_6771);
and U7365 (N_7365,N_6668,N_6700);
nand U7366 (N_7366,N_6691,N_6584);
and U7367 (N_7367,N_6764,N_6644);
or U7368 (N_7368,N_6639,N_6641);
xnor U7369 (N_7369,N_6551,N_6576);
nand U7370 (N_7370,N_6766,N_6571);
and U7371 (N_7371,N_6659,N_6797);
and U7372 (N_7372,N_6758,N_6788);
xor U7373 (N_7373,N_6604,N_6593);
nor U7374 (N_7374,N_6643,N_6751);
xnor U7375 (N_7375,N_6652,N_6515);
and U7376 (N_7376,N_6914,N_6845);
and U7377 (N_7377,N_6824,N_6719);
nand U7378 (N_7378,N_6732,N_6904);
xor U7379 (N_7379,N_6832,N_6555);
nand U7380 (N_7380,N_6711,N_6639);
nand U7381 (N_7381,N_6597,N_6755);
and U7382 (N_7382,N_6608,N_6899);
xnor U7383 (N_7383,N_6581,N_6838);
or U7384 (N_7384,N_6768,N_6626);
xnor U7385 (N_7385,N_6822,N_6736);
or U7386 (N_7386,N_6937,N_6975);
nor U7387 (N_7387,N_6905,N_6656);
nand U7388 (N_7388,N_6592,N_6552);
nand U7389 (N_7389,N_6967,N_6803);
and U7390 (N_7390,N_6995,N_6880);
nand U7391 (N_7391,N_6822,N_6857);
xnor U7392 (N_7392,N_6604,N_6900);
nand U7393 (N_7393,N_6854,N_6732);
or U7394 (N_7394,N_6814,N_6529);
nor U7395 (N_7395,N_6737,N_6940);
xnor U7396 (N_7396,N_6838,N_6709);
nand U7397 (N_7397,N_6629,N_6968);
or U7398 (N_7398,N_6821,N_6512);
or U7399 (N_7399,N_6775,N_6858);
xnor U7400 (N_7400,N_6535,N_6666);
xnor U7401 (N_7401,N_6696,N_6773);
or U7402 (N_7402,N_6707,N_6793);
xor U7403 (N_7403,N_6597,N_6516);
and U7404 (N_7404,N_6592,N_6625);
and U7405 (N_7405,N_6719,N_6602);
and U7406 (N_7406,N_6665,N_6835);
or U7407 (N_7407,N_6633,N_6596);
xnor U7408 (N_7408,N_6953,N_6769);
nor U7409 (N_7409,N_6774,N_6945);
nand U7410 (N_7410,N_6942,N_6917);
xnor U7411 (N_7411,N_6561,N_6804);
nor U7412 (N_7412,N_6728,N_6868);
and U7413 (N_7413,N_6528,N_6637);
and U7414 (N_7414,N_6942,N_6854);
or U7415 (N_7415,N_6600,N_6690);
and U7416 (N_7416,N_6871,N_6658);
xor U7417 (N_7417,N_6842,N_6662);
xor U7418 (N_7418,N_6519,N_6745);
nand U7419 (N_7419,N_6571,N_6558);
nand U7420 (N_7420,N_6898,N_6675);
or U7421 (N_7421,N_6946,N_6582);
and U7422 (N_7422,N_6515,N_6629);
nand U7423 (N_7423,N_6831,N_6656);
nor U7424 (N_7424,N_6948,N_6919);
and U7425 (N_7425,N_6951,N_6620);
or U7426 (N_7426,N_6906,N_6645);
nand U7427 (N_7427,N_6522,N_6562);
xnor U7428 (N_7428,N_6912,N_6816);
nor U7429 (N_7429,N_6846,N_6590);
and U7430 (N_7430,N_6620,N_6963);
nor U7431 (N_7431,N_6546,N_6545);
and U7432 (N_7432,N_6717,N_6900);
nor U7433 (N_7433,N_6791,N_6540);
nor U7434 (N_7434,N_6787,N_6525);
and U7435 (N_7435,N_6759,N_6850);
and U7436 (N_7436,N_6860,N_6980);
and U7437 (N_7437,N_6863,N_6918);
nor U7438 (N_7438,N_6618,N_6643);
xor U7439 (N_7439,N_6658,N_6586);
nor U7440 (N_7440,N_6687,N_6790);
or U7441 (N_7441,N_6898,N_6539);
nor U7442 (N_7442,N_6981,N_6795);
and U7443 (N_7443,N_6830,N_6816);
or U7444 (N_7444,N_6762,N_6732);
xor U7445 (N_7445,N_6677,N_6862);
and U7446 (N_7446,N_6594,N_6847);
nand U7447 (N_7447,N_6901,N_6720);
or U7448 (N_7448,N_6740,N_6644);
nor U7449 (N_7449,N_6999,N_6617);
nor U7450 (N_7450,N_6611,N_6729);
and U7451 (N_7451,N_6891,N_6933);
and U7452 (N_7452,N_6974,N_6593);
nor U7453 (N_7453,N_6705,N_6831);
nand U7454 (N_7454,N_6841,N_6895);
and U7455 (N_7455,N_6699,N_6953);
nor U7456 (N_7456,N_6998,N_6651);
nor U7457 (N_7457,N_6847,N_6746);
or U7458 (N_7458,N_6776,N_6968);
xor U7459 (N_7459,N_6532,N_6713);
xnor U7460 (N_7460,N_6674,N_6743);
nor U7461 (N_7461,N_6996,N_6842);
nand U7462 (N_7462,N_6788,N_6675);
nand U7463 (N_7463,N_6998,N_6550);
and U7464 (N_7464,N_6768,N_6967);
nor U7465 (N_7465,N_6647,N_6608);
and U7466 (N_7466,N_6884,N_6798);
nor U7467 (N_7467,N_6572,N_6992);
or U7468 (N_7468,N_6686,N_6724);
xnor U7469 (N_7469,N_6992,N_6882);
or U7470 (N_7470,N_6745,N_6948);
xnor U7471 (N_7471,N_6967,N_6903);
xnor U7472 (N_7472,N_6745,N_6783);
xnor U7473 (N_7473,N_6611,N_6936);
nand U7474 (N_7474,N_6683,N_6999);
and U7475 (N_7475,N_6663,N_6981);
or U7476 (N_7476,N_6692,N_6992);
or U7477 (N_7477,N_6599,N_6950);
nor U7478 (N_7478,N_6964,N_6723);
xnor U7479 (N_7479,N_6650,N_6596);
xor U7480 (N_7480,N_6529,N_6643);
nand U7481 (N_7481,N_6963,N_6966);
nor U7482 (N_7482,N_6832,N_6940);
nand U7483 (N_7483,N_6965,N_6632);
xnor U7484 (N_7484,N_6792,N_6908);
nor U7485 (N_7485,N_6900,N_6757);
and U7486 (N_7486,N_6768,N_6753);
xor U7487 (N_7487,N_6972,N_6630);
and U7488 (N_7488,N_6860,N_6519);
or U7489 (N_7489,N_6946,N_6573);
or U7490 (N_7490,N_6620,N_6536);
and U7491 (N_7491,N_6581,N_6527);
and U7492 (N_7492,N_6939,N_6612);
or U7493 (N_7493,N_6666,N_6737);
xnor U7494 (N_7494,N_6617,N_6692);
and U7495 (N_7495,N_6886,N_6880);
or U7496 (N_7496,N_6762,N_6777);
nor U7497 (N_7497,N_6734,N_6781);
nor U7498 (N_7498,N_6817,N_6878);
nand U7499 (N_7499,N_6949,N_6641);
nand U7500 (N_7500,N_7407,N_7354);
and U7501 (N_7501,N_7272,N_7220);
and U7502 (N_7502,N_7203,N_7015);
xnor U7503 (N_7503,N_7329,N_7419);
xnor U7504 (N_7504,N_7165,N_7382);
xnor U7505 (N_7505,N_7294,N_7484);
xnor U7506 (N_7506,N_7136,N_7411);
or U7507 (N_7507,N_7172,N_7247);
nand U7508 (N_7508,N_7207,N_7129);
and U7509 (N_7509,N_7389,N_7492);
nor U7510 (N_7510,N_7016,N_7280);
xor U7511 (N_7511,N_7221,N_7415);
xor U7512 (N_7512,N_7087,N_7008);
xor U7513 (N_7513,N_7326,N_7195);
or U7514 (N_7514,N_7343,N_7350);
xor U7515 (N_7515,N_7310,N_7019);
nor U7516 (N_7516,N_7024,N_7298);
nand U7517 (N_7517,N_7145,N_7338);
xor U7518 (N_7518,N_7096,N_7238);
or U7519 (N_7519,N_7159,N_7370);
nor U7520 (N_7520,N_7134,N_7114);
nor U7521 (N_7521,N_7327,N_7355);
or U7522 (N_7522,N_7292,N_7251);
or U7523 (N_7523,N_7451,N_7192);
and U7524 (N_7524,N_7112,N_7356);
and U7525 (N_7525,N_7498,N_7284);
and U7526 (N_7526,N_7265,N_7325);
nor U7527 (N_7527,N_7275,N_7150);
nand U7528 (N_7528,N_7068,N_7462);
and U7529 (N_7529,N_7149,N_7035);
nand U7530 (N_7530,N_7119,N_7315);
xnor U7531 (N_7531,N_7128,N_7433);
nor U7532 (N_7532,N_7281,N_7100);
and U7533 (N_7533,N_7291,N_7362);
nand U7534 (N_7534,N_7347,N_7293);
nor U7535 (N_7535,N_7188,N_7465);
and U7536 (N_7536,N_7029,N_7250);
nor U7537 (N_7537,N_7001,N_7122);
nand U7538 (N_7538,N_7233,N_7160);
xnor U7539 (N_7539,N_7330,N_7146);
nor U7540 (N_7540,N_7286,N_7263);
nand U7541 (N_7541,N_7390,N_7060);
nor U7542 (N_7542,N_7197,N_7053);
nand U7543 (N_7543,N_7471,N_7425);
nand U7544 (N_7544,N_7467,N_7475);
nor U7545 (N_7545,N_7032,N_7083);
and U7546 (N_7546,N_7398,N_7490);
xnor U7547 (N_7547,N_7456,N_7086);
nand U7548 (N_7548,N_7311,N_7124);
and U7549 (N_7549,N_7174,N_7092);
and U7550 (N_7550,N_7191,N_7052);
nand U7551 (N_7551,N_7358,N_7206);
nand U7552 (N_7552,N_7385,N_7455);
and U7553 (N_7553,N_7241,N_7156);
or U7554 (N_7554,N_7464,N_7460);
nor U7555 (N_7555,N_7094,N_7065);
or U7556 (N_7556,N_7349,N_7219);
nand U7557 (N_7557,N_7255,N_7289);
or U7558 (N_7558,N_7374,N_7082);
xor U7559 (N_7559,N_7055,N_7260);
xnor U7560 (N_7560,N_7023,N_7266);
or U7561 (N_7561,N_7007,N_7231);
nand U7562 (N_7562,N_7163,N_7333);
and U7563 (N_7563,N_7063,N_7208);
xor U7564 (N_7564,N_7057,N_7239);
nand U7565 (N_7565,N_7453,N_7256);
nand U7566 (N_7566,N_7090,N_7274);
nor U7567 (N_7567,N_7416,N_7491);
xnor U7568 (N_7568,N_7116,N_7170);
xnor U7569 (N_7569,N_7177,N_7393);
nor U7570 (N_7570,N_7067,N_7249);
xor U7571 (N_7571,N_7078,N_7152);
or U7572 (N_7572,N_7366,N_7230);
and U7573 (N_7573,N_7200,N_7039);
and U7574 (N_7574,N_7401,N_7080);
nand U7575 (N_7575,N_7345,N_7364);
or U7576 (N_7576,N_7320,N_7316);
or U7577 (N_7577,N_7406,N_7106);
and U7578 (N_7578,N_7384,N_7095);
and U7579 (N_7579,N_7269,N_7157);
nor U7580 (N_7580,N_7353,N_7395);
nor U7581 (N_7581,N_7357,N_7105);
xnor U7582 (N_7582,N_7414,N_7481);
xor U7583 (N_7583,N_7000,N_7193);
nor U7584 (N_7584,N_7210,N_7113);
or U7585 (N_7585,N_7161,N_7006);
xnor U7586 (N_7586,N_7312,N_7089);
or U7587 (N_7587,N_7304,N_7405);
or U7588 (N_7588,N_7287,N_7378);
xnor U7589 (N_7589,N_7391,N_7137);
xnor U7590 (N_7590,N_7229,N_7380);
and U7591 (N_7591,N_7010,N_7253);
nor U7592 (N_7592,N_7457,N_7302);
and U7593 (N_7593,N_7369,N_7199);
nand U7594 (N_7594,N_7427,N_7102);
or U7595 (N_7595,N_7386,N_7336);
nand U7596 (N_7596,N_7025,N_7158);
nor U7597 (N_7597,N_7109,N_7012);
nor U7598 (N_7598,N_7301,N_7037);
xor U7599 (N_7599,N_7098,N_7004);
and U7600 (N_7600,N_7468,N_7139);
xnor U7601 (N_7601,N_7348,N_7365);
nand U7602 (N_7602,N_7189,N_7056);
or U7603 (N_7603,N_7176,N_7043);
or U7604 (N_7604,N_7283,N_7215);
and U7605 (N_7605,N_7408,N_7021);
and U7606 (N_7606,N_7248,N_7088);
and U7607 (N_7607,N_7066,N_7036);
or U7608 (N_7608,N_7166,N_7496);
and U7609 (N_7609,N_7171,N_7482);
or U7610 (N_7610,N_7448,N_7246);
nand U7611 (N_7611,N_7198,N_7243);
and U7612 (N_7612,N_7091,N_7334);
xnor U7613 (N_7613,N_7031,N_7225);
xnor U7614 (N_7614,N_7264,N_7423);
or U7615 (N_7615,N_7050,N_7131);
or U7616 (N_7616,N_7309,N_7242);
nor U7617 (N_7617,N_7073,N_7232);
xnor U7618 (N_7618,N_7072,N_7376);
or U7619 (N_7619,N_7279,N_7125);
and U7620 (N_7620,N_7173,N_7144);
xor U7621 (N_7621,N_7108,N_7235);
xnor U7622 (N_7622,N_7034,N_7194);
nand U7623 (N_7623,N_7142,N_7313);
xnor U7624 (N_7624,N_7305,N_7214);
or U7625 (N_7625,N_7442,N_7169);
or U7626 (N_7626,N_7138,N_7318);
xor U7627 (N_7627,N_7300,N_7352);
or U7628 (N_7628,N_7201,N_7420);
nand U7629 (N_7629,N_7101,N_7441);
and U7630 (N_7630,N_7271,N_7216);
xor U7631 (N_7631,N_7017,N_7440);
nor U7632 (N_7632,N_7314,N_7217);
or U7633 (N_7633,N_7470,N_7099);
and U7634 (N_7634,N_7324,N_7209);
nor U7635 (N_7635,N_7093,N_7267);
nand U7636 (N_7636,N_7426,N_7054);
and U7637 (N_7637,N_7028,N_7466);
and U7638 (N_7638,N_7273,N_7104);
nand U7639 (N_7639,N_7205,N_7282);
nor U7640 (N_7640,N_7046,N_7003);
xnor U7641 (N_7641,N_7436,N_7047);
nand U7642 (N_7642,N_7444,N_7022);
nand U7643 (N_7643,N_7387,N_7458);
nand U7644 (N_7644,N_7244,N_7367);
and U7645 (N_7645,N_7410,N_7162);
xor U7646 (N_7646,N_7027,N_7359);
nand U7647 (N_7647,N_7227,N_7473);
and U7648 (N_7648,N_7447,N_7187);
and U7649 (N_7649,N_7422,N_7479);
nor U7650 (N_7650,N_7079,N_7224);
nand U7651 (N_7651,N_7472,N_7111);
nand U7652 (N_7652,N_7018,N_7383);
nor U7653 (N_7653,N_7290,N_7388);
nand U7654 (N_7654,N_7141,N_7372);
or U7655 (N_7655,N_7328,N_7446);
nand U7656 (N_7656,N_7361,N_7331);
nor U7657 (N_7657,N_7483,N_7270);
or U7658 (N_7658,N_7403,N_7303);
or U7659 (N_7659,N_7278,N_7379);
xnor U7660 (N_7660,N_7434,N_7474);
nand U7661 (N_7661,N_7069,N_7476);
or U7662 (N_7662,N_7486,N_7437);
xor U7663 (N_7663,N_7319,N_7045);
and U7664 (N_7664,N_7332,N_7020);
nor U7665 (N_7665,N_7288,N_7204);
nand U7666 (N_7666,N_7399,N_7428);
nand U7667 (N_7667,N_7180,N_7435);
and U7668 (N_7668,N_7339,N_7404);
xor U7669 (N_7669,N_7234,N_7487);
and U7670 (N_7670,N_7211,N_7133);
or U7671 (N_7671,N_7485,N_7430);
nor U7672 (N_7672,N_7392,N_7450);
nor U7673 (N_7673,N_7236,N_7245);
nor U7674 (N_7674,N_7261,N_7123);
nor U7675 (N_7675,N_7181,N_7117);
and U7676 (N_7676,N_7030,N_7377);
nor U7677 (N_7677,N_7070,N_7107);
nand U7678 (N_7678,N_7257,N_7341);
and U7679 (N_7679,N_7009,N_7296);
nand U7680 (N_7680,N_7477,N_7040);
and U7681 (N_7681,N_7130,N_7412);
and U7682 (N_7682,N_7042,N_7413);
and U7683 (N_7683,N_7321,N_7044);
nor U7684 (N_7684,N_7212,N_7307);
or U7685 (N_7685,N_7346,N_7373);
or U7686 (N_7686,N_7469,N_7480);
and U7687 (N_7687,N_7397,N_7120);
or U7688 (N_7688,N_7190,N_7077);
or U7689 (N_7689,N_7252,N_7438);
and U7690 (N_7690,N_7342,N_7062);
or U7691 (N_7691,N_7182,N_7084);
or U7692 (N_7692,N_7344,N_7254);
nor U7693 (N_7693,N_7431,N_7118);
nor U7694 (N_7694,N_7432,N_7497);
xor U7695 (N_7695,N_7402,N_7049);
or U7696 (N_7696,N_7013,N_7396);
and U7697 (N_7697,N_7135,N_7223);
and U7698 (N_7698,N_7186,N_7439);
or U7699 (N_7699,N_7058,N_7196);
and U7700 (N_7700,N_7276,N_7418);
nand U7701 (N_7701,N_7443,N_7240);
and U7702 (N_7702,N_7317,N_7226);
or U7703 (N_7703,N_7154,N_7097);
nor U7704 (N_7704,N_7014,N_7115);
or U7705 (N_7705,N_7179,N_7038);
nor U7706 (N_7706,N_7499,N_7424);
or U7707 (N_7707,N_7258,N_7121);
xnor U7708 (N_7708,N_7064,N_7417);
and U7709 (N_7709,N_7371,N_7368);
or U7710 (N_7710,N_7110,N_7184);
and U7711 (N_7711,N_7421,N_7262);
xnor U7712 (N_7712,N_7140,N_7488);
nor U7713 (N_7713,N_7337,N_7168);
nor U7714 (N_7714,N_7429,N_7381);
xnor U7715 (N_7715,N_7033,N_7041);
xor U7716 (N_7716,N_7493,N_7026);
nand U7717 (N_7717,N_7185,N_7323);
nand U7718 (N_7718,N_7449,N_7148);
or U7719 (N_7719,N_7085,N_7459);
and U7720 (N_7720,N_7308,N_7167);
nor U7721 (N_7721,N_7011,N_7081);
nor U7722 (N_7722,N_7259,N_7175);
xnor U7723 (N_7723,N_7183,N_7202);
xor U7724 (N_7724,N_7461,N_7394);
nand U7725 (N_7725,N_7409,N_7363);
or U7726 (N_7726,N_7155,N_7151);
or U7727 (N_7727,N_7059,N_7061);
and U7728 (N_7728,N_7340,N_7237);
xor U7729 (N_7729,N_7285,N_7351);
xor U7730 (N_7730,N_7297,N_7445);
and U7731 (N_7731,N_7222,N_7213);
nand U7732 (N_7732,N_7228,N_7495);
nor U7733 (N_7733,N_7076,N_7375);
xor U7734 (N_7734,N_7178,N_7452);
xor U7735 (N_7735,N_7002,N_7071);
or U7736 (N_7736,N_7153,N_7494);
nand U7737 (N_7737,N_7478,N_7074);
or U7738 (N_7738,N_7005,N_7048);
xnor U7739 (N_7739,N_7277,N_7051);
and U7740 (N_7740,N_7075,N_7322);
nand U7741 (N_7741,N_7463,N_7335);
nand U7742 (N_7742,N_7306,N_7268);
or U7743 (N_7743,N_7132,N_7126);
xor U7744 (N_7744,N_7143,N_7127);
and U7745 (N_7745,N_7147,N_7218);
and U7746 (N_7746,N_7489,N_7454);
nand U7747 (N_7747,N_7400,N_7103);
xor U7748 (N_7748,N_7295,N_7360);
nor U7749 (N_7749,N_7164,N_7299);
nor U7750 (N_7750,N_7367,N_7365);
xor U7751 (N_7751,N_7490,N_7035);
nand U7752 (N_7752,N_7069,N_7156);
or U7753 (N_7753,N_7099,N_7325);
nand U7754 (N_7754,N_7237,N_7306);
nor U7755 (N_7755,N_7308,N_7080);
xor U7756 (N_7756,N_7438,N_7221);
xnor U7757 (N_7757,N_7219,N_7327);
xor U7758 (N_7758,N_7119,N_7365);
nand U7759 (N_7759,N_7210,N_7013);
and U7760 (N_7760,N_7263,N_7315);
nand U7761 (N_7761,N_7348,N_7013);
and U7762 (N_7762,N_7473,N_7295);
nor U7763 (N_7763,N_7381,N_7051);
or U7764 (N_7764,N_7097,N_7085);
nor U7765 (N_7765,N_7365,N_7487);
and U7766 (N_7766,N_7015,N_7093);
xnor U7767 (N_7767,N_7479,N_7224);
xnor U7768 (N_7768,N_7495,N_7088);
or U7769 (N_7769,N_7413,N_7416);
nor U7770 (N_7770,N_7061,N_7192);
xnor U7771 (N_7771,N_7498,N_7237);
nor U7772 (N_7772,N_7133,N_7339);
xnor U7773 (N_7773,N_7043,N_7492);
xnor U7774 (N_7774,N_7226,N_7334);
nand U7775 (N_7775,N_7403,N_7497);
nand U7776 (N_7776,N_7037,N_7165);
and U7777 (N_7777,N_7044,N_7397);
xor U7778 (N_7778,N_7224,N_7160);
xor U7779 (N_7779,N_7191,N_7390);
and U7780 (N_7780,N_7023,N_7408);
nand U7781 (N_7781,N_7004,N_7088);
nand U7782 (N_7782,N_7264,N_7417);
or U7783 (N_7783,N_7387,N_7047);
and U7784 (N_7784,N_7447,N_7114);
nand U7785 (N_7785,N_7244,N_7172);
and U7786 (N_7786,N_7162,N_7233);
nand U7787 (N_7787,N_7368,N_7149);
or U7788 (N_7788,N_7438,N_7249);
nor U7789 (N_7789,N_7423,N_7222);
and U7790 (N_7790,N_7240,N_7208);
nand U7791 (N_7791,N_7088,N_7333);
nor U7792 (N_7792,N_7317,N_7098);
and U7793 (N_7793,N_7275,N_7052);
or U7794 (N_7794,N_7143,N_7355);
nor U7795 (N_7795,N_7318,N_7198);
or U7796 (N_7796,N_7117,N_7006);
or U7797 (N_7797,N_7370,N_7303);
xor U7798 (N_7798,N_7156,N_7408);
nor U7799 (N_7799,N_7122,N_7164);
and U7800 (N_7800,N_7032,N_7423);
xnor U7801 (N_7801,N_7372,N_7235);
xor U7802 (N_7802,N_7321,N_7156);
xnor U7803 (N_7803,N_7250,N_7199);
or U7804 (N_7804,N_7070,N_7430);
nand U7805 (N_7805,N_7085,N_7082);
nor U7806 (N_7806,N_7368,N_7448);
and U7807 (N_7807,N_7183,N_7187);
nand U7808 (N_7808,N_7323,N_7407);
nor U7809 (N_7809,N_7019,N_7294);
and U7810 (N_7810,N_7323,N_7495);
or U7811 (N_7811,N_7018,N_7425);
xnor U7812 (N_7812,N_7359,N_7256);
or U7813 (N_7813,N_7185,N_7070);
nor U7814 (N_7814,N_7126,N_7338);
xnor U7815 (N_7815,N_7405,N_7211);
nor U7816 (N_7816,N_7306,N_7119);
nor U7817 (N_7817,N_7497,N_7233);
nor U7818 (N_7818,N_7367,N_7034);
xnor U7819 (N_7819,N_7194,N_7017);
or U7820 (N_7820,N_7278,N_7367);
nor U7821 (N_7821,N_7057,N_7291);
and U7822 (N_7822,N_7430,N_7439);
xnor U7823 (N_7823,N_7271,N_7066);
nor U7824 (N_7824,N_7494,N_7172);
nor U7825 (N_7825,N_7077,N_7364);
or U7826 (N_7826,N_7415,N_7428);
or U7827 (N_7827,N_7475,N_7236);
and U7828 (N_7828,N_7050,N_7492);
or U7829 (N_7829,N_7461,N_7245);
nand U7830 (N_7830,N_7343,N_7426);
xor U7831 (N_7831,N_7340,N_7022);
nand U7832 (N_7832,N_7331,N_7157);
and U7833 (N_7833,N_7463,N_7252);
nand U7834 (N_7834,N_7061,N_7158);
nand U7835 (N_7835,N_7278,N_7432);
and U7836 (N_7836,N_7201,N_7449);
nor U7837 (N_7837,N_7065,N_7202);
nor U7838 (N_7838,N_7172,N_7132);
or U7839 (N_7839,N_7330,N_7073);
nand U7840 (N_7840,N_7435,N_7467);
xor U7841 (N_7841,N_7487,N_7432);
or U7842 (N_7842,N_7185,N_7261);
xor U7843 (N_7843,N_7470,N_7250);
or U7844 (N_7844,N_7423,N_7449);
nand U7845 (N_7845,N_7393,N_7348);
nand U7846 (N_7846,N_7248,N_7256);
or U7847 (N_7847,N_7067,N_7082);
xnor U7848 (N_7848,N_7267,N_7135);
nor U7849 (N_7849,N_7093,N_7316);
and U7850 (N_7850,N_7492,N_7253);
and U7851 (N_7851,N_7440,N_7137);
nor U7852 (N_7852,N_7487,N_7328);
nand U7853 (N_7853,N_7362,N_7366);
xnor U7854 (N_7854,N_7222,N_7009);
and U7855 (N_7855,N_7269,N_7011);
or U7856 (N_7856,N_7130,N_7489);
or U7857 (N_7857,N_7099,N_7399);
and U7858 (N_7858,N_7029,N_7243);
xor U7859 (N_7859,N_7148,N_7208);
nand U7860 (N_7860,N_7448,N_7457);
nand U7861 (N_7861,N_7105,N_7030);
and U7862 (N_7862,N_7001,N_7339);
xnor U7863 (N_7863,N_7342,N_7122);
xor U7864 (N_7864,N_7364,N_7098);
and U7865 (N_7865,N_7076,N_7121);
and U7866 (N_7866,N_7301,N_7165);
nor U7867 (N_7867,N_7123,N_7381);
nand U7868 (N_7868,N_7094,N_7214);
nand U7869 (N_7869,N_7350,N_7082);
nand U7870 (N_7870,N_7297,N_7395);
xnor U7871 (N_7871,N_7076,N_7408);
nand U7872 (N_7872,N_7410,N_7367);
xnor U7873 (N_7873,N_7356,N_7068);
xor U7874 (N_7874,N_7136,N_7288);
nand U7875 (N_7875,N_7362,N_7411);
nand U7876 (N_7876,N_7050,N_7037);
nor U7877 (N_7877,N_7272,N_7421);
or U7878 (N_7878,N_7132,N_7151);
xnor U7879 (N_7879,N_7078,N_7112);
xor U7880 (N_7880,N_7009,N_7312);
nand U7881 (N_7881,N_7499,N_7458);
or U7882 (N_7882,N_7420,N_7476);
nor U7883 (N_7883,N_7087,N_7388);
nand U7884 (N_7884,N_7429,N_7152);
or U7885 (N_7885,N_7237,N_7149);
xnor U7886 (N_7886,N_7295,N_7031);
nor U7887 (N_7887,N_7139,N_7112);
nor U7888 (N_7888,N_7070,N_7193);
nand U7889 (N_7889,N_7340,N_7287);
or U7890 (N_7890,N_7393,N_7284);
xor U7891 (N_7891,N_7300,N_7307);
nand U7892 (N_7892,N_7087,N_7094);
and U7893 (N_7893,N_7127,N_7332);
nand U7894 (N_7894,N_7272,N_7169);
nor U7895 (N_7895,N_7445,N_7450);
xnor U7896 (N_7896,N_7150,N_7315);
or U7897 (N_7897,N_7159,N_7313);
and U7898 (N_7898,N_7011,N_7326);
or U7899 (N_7899,N_7186,N_7215);
nand U7900 (N_7900,N_7255,N_7326);
and U7901 (N_7901,N_7166,N_7266);
and U7902 (N_7902,N_7323,N_7260);
xnor U7903 (N_7903,N_7119,N_7493);
nor U7904 (N_7904,N_7083,N_7338);
and U7905 (N_7905,N_7491,N_7212);
and U7906 (N_7906,N_7234,N_7002);
or U7907 (N_7907,N_7349,N_7388);
nor U7908 (N_7908,N_7270,N_7119);
nor U7909 (N_7909,N_7201,N_7391);
nand U7910 (N_7910,N_7364,N_7452);
or U7911 (N_7911,N_7225,N_7048);
xnor U7912 (N_7912,N_7327,N_7353);
nor U7913 (N_7913,N_7001,N_7060);
xnor U7914 (N_7914,N_7433,N_7251);
xor U7915 (N_7915,N_7300,N_7246);
and U7916 (N_7916,N_7400,N_7242);
or U7917 (N_7917,N_7067,N_7098);
or U7918 (N_7918,N_7242,N_7127);
and U7919 (N_7919,N_7184,N_7030);
and U7920 (N_7920,N_7015,N_7247);
and U7921 (N_7921,N_7486,N_7445);
nor U7922 (N_7922,N_7363,N_7379);
and U7923 (N_7923,N_7140,N_7376);
nor U7924 (N_7924,N_7228,N_7178);
xor U7925 (N_7925,N_7329,N_7019);
xnor U7926 (N_7926,N_7045,N_7483);
nor U7927 (N_7927,N_7304,N_7107);
and U7928 (N_7928,N_7283,N_7331);
and U7929 (N_7929,N_7323,N_7339);
or U7930 (N_7930,N_7120,N_7430);
or U7931 (N_7931,N_7386,N_7038);
xor U7932 (N_7932,N_7037,N_7478);
or U7933 (N_7933,N_7223,N_7499);
or U7934 (N_7934,N_7061,N_7225);
nor U7935 (N_7935,N_7364,N_7465);
or U7936 (N_7936,N_7181,N_7304);
nor U7937 (N_7937,N_7140,N_7195);
or U7938 (N_7938,N_7184,N_7210);
nand U7939 (N_7939,N_7105,N_7043);
or U7940 (N_7940,N_7441,N_7045);
xnor U7941 (N_7941,N_7060,N_7117);
nand U7942 (N_7942,N_7178,N_7125);
nand U7943 (N_7943,N_7035,N_7099);
or U7944 (N_7944,N_7441,N_7160);
nor U7945 (N_7945,N_7019,N_7431);
nor U7946 (N_7946,N_7424,N_7151);
nand U7947 (N_7947,N_7473,N_7240);
nor U7948 (N_7948,N_7045,N_7134);
xor U7949 (N_7949,N_7450,N_7470);
xor U7950 (N_7950,N_7485,N_7103);
nand U7951 (N_7951,N_7014,N_7235);
nor U7952 (N_7952,N_7387,N_7492);
or U7953 (N_7953,N_7497,N_7201);
nand U7954 (N_7954,N_7485,N_7197);
nand U7955 (N_7955,N_7202,N_7493);
or U7956 (N_7956,N_7107,N_7403);
and U7957 (N_7957,N_7169,N_7153);
and U7958 (N_7958,N_7236,N_7383);
and U7959 (N_7959,N_7373,N_7196);
nand U7960 (N_7960,N_7445,N_7448);
nor U7961 (N_7961,N_7371,N_7438);
xnor U7962 (N_7962,N_7385,N_7031);
or U7963 (N_7963,N_7088,N_7470);
and U7964 (N_7964,N_7451,N_7499);
xor U7965 (N_7965,N_7234,N_7434);
xor U7966 (N_7966,N_7376,N_7279);
or U7967 (N_7967,N_7170,N_7193);
nand U7968 (N_7968,N_7477,N_7412);
and U7969 (N_7969,N_7120,N_7240);
nand U7970 (N_7970,N_7181,N_7127);
xnor U7971 (N_7971,N_7359,N_7469);
and U7972 (N_7972,N_7461,N_7031);
nor U7973 (N_7973,N_7314,N_7046);
nand U7974 (N_7974,N_7409,N_7330);
or U7975 (N_7975,N_7292,N_7172);
nor U7976 (N_7976,N_7077,N_7275);
nor U7977 (N_7977,N_7417,N_7143);
nor U7978 (N_7978,N_7019,N_7432);
nand U7979 (N_7979,N_7349,N_7258);
xnor U7980 (N_7980,N_7404,N_7457);
or U7981 (N_7981,N_7118,N_7204);
nand U7982 (N_7982,N_7345,N_7016);
xor U7983 (N_7983,N_7357,N_7456);
or U7984 (N_7984,N_7085,N_7181);
nor U7985 (N_7985,N_7348,N_7278);
nand U7986 (N_7986,N_7358,N_7388);
nand U7987 (N_7987,N_7168,N_7040);
nand U7988 (N_7988,N_7360,N_7147);
or U7989 (N_7989,N_7073,N_7082);
xor U7990 (N_7990,N_7025,N_7407);
xor U7991 (N_7991,N_7245,N_7484);
nor U7992 (N_7992,N_7176,N_7060);
and U7993 (N_7993,N_7394,N_7256);
or U7994 (N_7994,N_7337,N_7319);
nand U7995 (N_7995,N_7460,N_7136);
or U7996 (N_7996,N_7054,N_7476);
nor U7997 (N_7997,N_7309,N_7098);
nand U7998 (N_7998,N_7452,N_7492);
nor U7999 (N_7999,N_7481,N_7164);
or U8000 (N_8000,N_7779,N_7891);
nor U8001 (N_8001,N_7778,N_7500);
and U8002 (N_8002,N_7707,N_7659);
nor U8003 (N_8003,N_7772,N_7857);
and U8004 (N_8004,N_7591,N_7911);
nand U8005 (N_8005,N_7641,N_7550);
xnor U8006 (N_8006,N_7664,N_7933);
xnor U8007 (N_8007,N_7810,N_7975);
nor U8008 (N_8008,N_7681,N_7558);
nand U8009 (N_8009,N_7946,N_7639);
nand U8010 (N_8010,N_7851,N_7807);
and U8011 (N_8011,N_7642,N_7669);
nor U8012 (N_8012,N_7740,N_7897);
and U8013 (N_8013,N_7949,N_7632);
nor U8014 (N_8014,N_7756,N_7717);
or U8015 (N_8015,N_7845,N_7593);
or U8016 (N_8016,N_7997,N_7678);
nor U8017 (N_8017,N_7568,N_7829);
or U8018 (N_8018,N_7917,N_7978);
nand U8019 (N_8019,N_7588,N_7923);
and U8020 (N_8020,N_7753,N_7804);
or U8021 (N_8021,N_7977,N_7723);
nand U8022 (N_8022,N_7823,N_7687);
xor U8023 (N_8023,N_7899,N_7648);
xor U8024 (N_8024,N_7542,N_7688);
or U8025 (N_8025,N_7657,N_7529);
or U8026 (N_8026,N_7791,N_7602);
and U8027 (N_8027,N_7822,N_7575);
xor U8028 (N_8028,N_7530,N_7511);
and U8029 (N_8029,N_7821,N_7840);
nand U8030 (N_8030,N_7661,N_7879);
nor U8031 (N_8031,N_7920,N_7535);
xor U8032 (N_8032,N_7759,N_7514);
and U8033 (N_8033,N_7979,N_7704);
and U8034 (N_8034,N_7878,N_7670);
nand U8035 (N_8035,N_7900,N_7745);
xor U8036 (N_8036,N_7819,N_7839);
or U8037 (N_8037,N_7865,N_7658);
xor U8038 (N_8038,N_7972,N_7769);
nand U8039 (N_8039,N_7718,N_7518);
or U8040 (N_8040,N_7677,N_7733);
and U8041 (N_8041,N_7995,N_7962);
or U8042 (N_8042,N_7501,N_7502);
xnor U8043 (N_8043,N_7864,N_7884);
nand U8044 (N_8044,N_7746,N_7951);
nor U8045 (N_8045,N_7767,N_7721);
or U8046 (N_8046,N_7872,N_7633);
or U8047 (N_8047,N_7686,N_7950);
nor U8048 (N_8048,N_7729,N_7757);
xor U8049 (N_8049,N_7883,N_7607);
nand U8050 (N_8050,N_7656,N_7699);
nor U8051 (N_8051,N_7915,N_7574);
and U8052 (N_8052,N_7627,N_7800);
and U8053 (N_8053,N_7705,N_7999);
nor U8054 (N_8054,N_7521,N_7713);
xor U8055 (N_8055,N_7635,N_7604);
xnor U8056 (N_8056,N_7566,N_7939);
or U8057 (N_8057,N_7562,N_7787);
and U8058 (N_8058,N_7832,N_7945);
xnor U8059 (N_8059,N_7506,N_7918);
nand U8060 (N_8060,N_7833,N_7731);
or U8061 (N_8061,N_7974,N_7934);
nand U8062 (N_8062,N_7820,N_7595);
or U8063 (N_8063,N_7689,N_7662);
or U8064 (N_8064,N_7871,N_7725);
nor U8065 (N_8065,N_7583,N_7838);
xor U8066 (N_8066,N_7780,N_7634);
and U8067 (N_8067,N_7960,N_7785);
nor U8068 (N_8068,N_7598,N_7924);
nor U8069 (N_8069,N_7674,N_7853);
xnor U8070 (N_8070,N_7700,N_7647);
xnor U8071 (N_8071,N_7957,N_7777);
and U8072 (N_8072,N_7904,N_7844);
nor U8073 (N_8073,N_7580,N_7628);
xor U8074 (N_8074,N_7711,N_7947);
or U8075 (N_8075,N_7675,N_7524);
nand U8076 (N_8076,N_7512,N_7630);
or U8077 (N_8077,N_7750,N_7741);
nand U8078 (N_8078,N_7836,N_7567);
nor U8079 (N_8079,N_7783,N_7697);
and U8080 (N_8080,N_7561,N_7594);
nor U8081 (N_8081,N_7654,N_7991);
nand U8082 (N_8082,N_7646,N_7549);
or U8083 (N_8083,N_7541,N_7818);
or U8084 (N_8084,N_7993,N_7855);
xnor U8085 (N_8085,N_7766,N_7551);
nand U8086 (N_8086,N_7761,N_7560);
and U8087 (N_8087,N_7868,N_7533);
or U8088 (N_8088,N_7968,N_7963);
or U8089 (N_8089,N_7902,N_7895);
nor U8090 (N_8090,N_7816,N_7784);
xnor U8091 (N_8091,N_7969,N_7651);
xor U8092 (N_8092,N_7732,N_7532);
xnor U8093 (N_8093,N_7861,N_7616);
nand U8094 (N_8094,N_7742,N_7712);
nor U8095 (N_8095,N_7536,N_7623);
xor U8096 (N_8096,N_7672,N_7764);
xnor U8097 (N_8097,N_7796,N_7912);
xor U8098 (N_8098,N_7929,N_7914);
nor U8099 (N_8099,N_7528,N_7813);
and U8100 (N_8100,N_7749,N_7652);
nor U8101 (N_8101,N_7621,N_7507);
xnor U8102 (N_8102,N_7852,N_7587);
nand U8103 (N_8103,N_7916,N_7660);
or U8104 (N_8104,N_7637,N_7600);
nand U8105 (N_8105,N_7626,N_7624);
and U8106 (N_8106,N_7534,N_7565);
or U8107 (N_8107,N_7638,N_7788);
nor U8108 (N_8108,N_7692,N_7928);
and U8109 (N_8109,N_7906,N_7811);
or U8110 (N_8110,N_7727,N_7965);
and U8111 (N_8111,N_7622,N_7792);
nand U8112 (N_8112,N_7998,N_7927);
nand U8113 (N_8113,N_7570,N_7983);
nor U8114 (N_8114,N_7510,N_7763);
or U8115 (N_8115,N_7954,N_7752);
nor U8116 (N_8116,N_7955,N_7668);
xnor U8117 (N_8117,N_7538,N_7655);
nor U8118 (N_8118,N_7556,N_7937);
nor U8119 (N_8119,N_7971,N_7798);
or U8120 (N_8120,N_7619,N_7990);
xor U8121 (N_8121,N_7599,N_7751);
nor U8122 (N_8122,N_7826,N_7696);
or U8123 (N_8123,N_7931,N_7776);
nor U8124 (N_8124,N_7958,N_7544);
xor U8125 (N_8125,N_7980,N_7548);
or U8126 (N_8126,N_7747,N_7932);
nor U8127 (N_8127,N_7846,N_7671);
nand U8128 (N_8128,N_7610,N_7708);
and U8129 (N_8129,N_7824,N_7873);
nor U8130 (N_8130,N_7618,N_7590);
nand U8131 (N_8131,N_7869,N_7984);
xnor U8132 (N_8132,N_7612,N_7629);
or U8133 (N_8133,N_7601,N_7578);
or U8134 (N_8134,N_7774,N_7701);
nand U8135 (N_8135,N_7649,N_7910);
nand U8136 (N_8136,N_7909,N_7519);
nand U8137 (N_8137,N_7793,N_7941);
and U8138 (N_8138,N_7715,N_7513);
nand U8139 (N_8139,N_7503,N_7554);
nand U8140 (N_8140,N_7809,N_7867);
or U8141 (N_8141,N_7617,N_7653);
nand U8142 (N_8142,N_7765,N_7706);
nor U8143 (N_8143,N_7908,N_7794);
xor U8144 (N_8144,N_7702,N_7806);
or U8145 (N_8145,N_7921,N_7959);
nor U8146 (N_8146,N_7515,N_7889);
or U8147 (N_8147,N_7812,N_7814);
nand U8148 (N_8148,N_7537,N_7684);
or U8149 (N_8149,N_7572,N_7760);
and U8150 (N_8150,N_7893,N_7735);
and U8151 (N_8151,N_7584,N_7966);
nand U8152 (N_8152,N_7625,N_7683);
xor U8153 (N_8153,N_7986,N_7837);
and U8154 (N_8154,N_7830,N_7640);
nand U8155 (N_8155,N_7650,N_7539);
and U8156 (N_8156,N_7898,N_7797);
xnor U8157 (N_8157,N_7948,N_7860);
xnor U8158 (N_8158,N_7736,N_7738);
nor U8159 (N_8159,N_7509,N_7645);
xor U8160 (N_8160,N_7863,N_7782);
and U8161 (N_8161,N_7586,N_7976);
nand U8162 (N_8162,N_7803,N_7720);
nand U8163 (N_8163,N_7665,N_7527);
xor U8164 (N_8164,N_7882,N_7722);
nor U8165 (N_8165,N_7885,N_7926);
xnor U8166 (N_8166,N_7636,N_7589);
and U8167 (N_8167,N_7847,N_7953);
nor U8168 (N_8168,N_7922,N_7956);
or U8169 (N_8169,N_7952,N_7981);
and U8170 (N_8170,N_7944,N_7862);
and U8171 (N_8171,N_7547,N_7710);
and U8172 (N_8172,N_7543,N_7730);
or U8173 (N_8173,N_7992,N_7724);
and U8174 (N_8174,N_7808,N_7771);
xor U8175 (N_8175,N_7691,N_7552);
and U8176 (N_8176,N_7935,N_7890);
or U8177 (N_8177,N_7775,N_7802);
or U8178 (N_8178,N_7907,N_7781);
nor U8179 (N_8179,N_7754,N_7611);
nor U8180 (N_8180,N_7795,N_7605);
nor U8181 (N_8181,N_7834,N_7758);
nand U8182 (N_8182,N_7881,N_7545);
nand U8183 (N_8183,N_7614,N_7508);
and U8184 (N_8184,N_7925,N_7987);
or U8185 (N_8185,N_7936,N_7714);
and U8186 (N_8186,N_7526,N_7842);
nand U8187 (N_8187,N_7576,N_7734);
nand U8188 (N_8188,N_7825,N_7563);
or U8189 (N_8189,N_7880,N_7643);
nor U8190 (N_8190,N_7970,N_7703);
xnor U8191 (N_8191,N_7673,N_7553);
and U8192 (N_8192,N_7849,N_7856);
xnor U8193 (N_8193,N_7737,N_7597);
nand U8194 (N_8194,N_7698,N_7919);
and U8195 (N_8195,N_7517,N_7892);
or U8196 (N_8196,N_7557,N_7743);
nor U8197 (N_8197,N_7613,N_7996);
and U8198 (N_8198,N_7546,N_7581);
or U8199 (N_8199,N_7690,N_7680);
nand U8200 (N_8200,N_7985,N_7559);
xnor U8201 (N_8201,N_7505,N_7815);
nor U8202 (N_8202,N_7644,N_7603);
and U8203 (N_8203,N_7913,N_7942);
xor U8204 (N_8204,N_7967,N_7859);
nand U8205 (N_8205,N_7801,N_7666);
xor U8206 (N_8206,N_7522,N_7989);
xor U8207 (N_8207,N_7685,N_7994);
and U8208 (N_8208,N_7964,N_7905);
and U8209 (N_8209,N_7585,N_7679);
or U8210 (N_8210,N_7982,N_7877);
or U8211 (N_8211,N_7827,N_7573);
nand U8212 (N_8212,N_7555,N_7676);
nand U8213 (N_8213,N_7748,N_7516);
and U8214 (N_8214,N_7841,N_7564);
or U8215 (N_8215,N_7768,N_7773);
and U8216 (N_8216,N_7854,N_7799);
nor U8217 (N_8217,N_7888,N_7726);
nor U8218 (N_8218,N_7961,N_7835);
and U8219 (N_8219,N_7943,N_7858);
nand U8220 (N_8220,N_7886,N_7786);
xnor U8221 (N_8221,N_7938,N_7523);
or U8222 (N_8222,N_7988,N_7631);
nand U8223 (N_8223,N_7728,N_7831);
and U8224 (N_8224,N_7805,N_7504);
or U8225 (N_8225,N_7716,N_7828);
and U8226 (N_8226,N_7744,N_7577);
xor U8227 (N_8227,N_7894,N_7596);
or U8228 (N_8228,N_7770,N_7667);
xor U8229 (N_8229,N_7848,N_7615);
xor U8230 (N_8230,N_7663,N_7875);
nand U8231 (N_8231,N_7739,N_7609);
xnor U8232 (N_8232,N_7693,N_7896);
nor U8233 (N_8233,N_7709,N_7540);
nor U8234 (N_8234,N_7592,N_7682);
or U8235 (N_8235,N_7850,N_7843);
or U8236 (N_8236,N_7694,N_7525);
and U8237 (N_8237,N_7930,N_7579);
or U8238 (N_8238,N_7695,N_7789);
or U8239 (N_8239,N_7903,N_7876);
nor U8240 (N_8240,N_7817,N_7973);
or U8241 (N_8241,N_7620,N_7870);
nand U8242 (N_8242,N_7866,N_7606);
nand U8243 (N_8243,N_7874,N_7520);
nand U8244 (N_8244,N_7571,N_7608);
nand U8245 (N_8245,N_7790,N_7719);
xor U8246 (N_8246,N_7887,N_7582);
xnor U8247 (N_8247,N_7531,N_7755);
nand U8248 (N_8248,N_7940,N_7762);
nand U8249 (N_8249,N_7901,N_7569);
nand U8250 (N_8250,N_7562,N_7726);
xnor U8251 (N_8251,N_7962,N_7940);
nor U8252 (N_8252,N_7882,N_7719);
or U8253 (N_8253,N_7924,N_7793);
nor U8254 (N_8254,N_7615,N_7576);
xor U8255 (N_8255,N_7866,N_7640);
or U8256 (N_8256,N_7862,N_7821);
nand U8257 (N_8257,N_7576,N_7604);
xor U8258 (N_8258,N_7938,N_7599);
xor U8259 (N_8259,N_7518,N_7724);
and U8260 (N_8260,N_7720,N_7840);
xor U8261 (N_8261,N_7812,N_7887);
nor U8262 (N_8262,N_7555,N_7696);
and U8263 (N_8263,N_7879,N_7854);
nor U8264 (N_8264,N_7616,N_7829);
xor U8265 (N_8265,N_7909,N_7617);
xnor U8266 (N_8266,N_7741,N_7749);
xor U8267 (N_8267,N_7629,N_7702);
nor U8268 (N_8268,N_7927,N_7593);
xor U8269 (N_8269,N_7966,N_7920);
or U8270 (N_8270,N_7587,N_7983);
and U8271 (N_8271,N_7659,N_7857);
xnor U8272 (N_8272,N_7964,N_7755);
nor U8273 (N_8273,N_7675,N_7682);
and U8274 (N_8274,N_7786,N_7723);
xor U8275 (N_8275,N_7552,N_7870);
and U8276 (N_8276,N_7554,N_7506);
nor U8277 (N_8277,N_7773,N_7745);
xnor U8278 (N_8278,N_7559,N_7936);
or U8279 (N_8279,N_7503,N_7659);
and U8280 (N_8280,N_7656,N_7697);
and U8281 (N_8281,N_7502,N_7693);
and U8282 (N_8282,N_7870,N_7740);
or U8283 (N_8283,N_7604,N_7941);
nor U8284 (N_8284,N_7541,N_7544);
and U8285 (N_8285,N_7528,N_7579);
or U8286 (N_8286,N_7567,N_7882);
nor U8287 (N_8287,N_7611,N_7678);
nor U8288 (N_8288,N_7693,N_7855);
nand U8289 (N_8289,N_7772,N_7766);
xnor U8290 (N_8290,N_7716,N_7801);
and U8291 (N_8291,N_7764,N_7937);
xnor U8292 (N_8292,N_7708,N_7562);
nand U8293 (N_8293,N_7581,N_7952);
nand U8294 (N_8294,N_7607,N_7976);
and U8295 (N_8295,N_7938,N_7715);
and U8296 (N_8296,N_7908,N_7641);
nand U8297 (N_8297,N_7948,N_7811);
or U8298 (N_8298,N_7706,N_7723);
nand U8299 (N_8299,N_7892,N_7672);
or U8300 (N_8300,N_7531,N_7967);
or U8301 (N_8301,N_7615,N_7724);
nand U8302 (N_8302,N_7573,N_7672);
xor U8303 (N_8303,N_7536,N_7680);
xnor U8304 (N_8304,N_7679,N_7966);
or U8305 (N_8305,N_7540,N_7847);
nor U8306 (N_8306,N_7688,N_7808);
or U8307 (N_8307,N_7505,N_7785);
nor U8308 (N_8308,N_7904,N_7697);
nand U8309 (N_8309,N_7781,N_7955);
xnor U8310 (N_8310,N_7697,N_7820);
xnor U8311 (N_8311,N_7682,N_7576);
nand U8312 (N_8312,N_7804,N_7513);
and U8313 (N_8313,N_7699,N_7966);
nor U8314 (N_8314,N_7724,N_7760);
nor U8315 (N_8315,N_7871,N_7777);
xnor U8316 (N_8316,N_7787,N_7601);
and U8317 (N_8317,N_7786,N_7908);
nor U8318 (N_8318,N_7866,N_7832);
nand U8319 (N_8319,N_7620,N_7766);
nor U8320 (N_8320,N_7725,N_7678);
nor U8321 (N_8321,N_7724,N_7623);
xor U8322 (N_8322,N_7817,N_7771);
xor U8323 (N_8323,N_7914,N_7785);
and U8324 (N_8324,N_7566,N_7840);
xnor U8325 (N_8325,N_7674,N_7644);
xor U8326 (N_8326,N_7509,N_7532);
and U8327 (N_8327,N_7836,N_7573);
or U8328 (N_8328,N_7793,N_7536);
or U8329 (N_8329,N_7810,N_7878);
and U8330 (N_8330,N_7617,N_7546);
and U8331 (N_8331,N_7908,N_7851);
or U8332 (N_8332,N_7926,N_7887);
or U8333 (N_8333,N_7923,N_7874);
nor U8334 (N_8334,N_7771,N_7691);
or U8335 (N_8335,N_7988,N_7923);
nor U8336 (N_8336,N_7985,N_7806);
nor U8337 (N_8337,N_7658,N_7746);
or U8338 (N_8338,N_7915,N_7963);
or U8339 (N_8339,N_7998,N_7629);
and U8340 (N_8340,N_7503,N_7708);
and U8341 (N_8341,N_7715,N_7935);
and U8342 (N_8342,N_7598,N_7845);
nor U8343 (N_8343,N_7855,N_7515);
and U8344 (N_8344,N_7751,N_7958);
nor U8345 (N_8345,N_7567,N_7533);
nand U8346 (N_8346,N_7952,N_7889);
nor U8347 (N_8347,N_7586,N_7969);
or U8348 (N_8348,N_7638,N_7564);
xor U8349 (N_8349,N_7885,N_7526);
nand U8350 (N_8350,N_7997,N_7766);
or U8351 (N_8351,N_7532,N_7650);
or U8352 (N_8352,N_7721,N_7888);
nand U8353 (N_8353,N_7956,N_7643);
or U8354 (N_8354,N_7647,N_7583);
and U8355 (N_8355,N_7543,N_7725);
nand U8356 (N_8356,N_7595,N_7840);
nand U8357 (N_8357,N_7726,N_7623);
and U8358 (N_8358,N_7882,N_7850);
xnor U8359 (N_8359,N_7728,N_7720);
nor U8360 (N_8360,N_7747,N_7678);
nor U8361 (N_8361,N_7775,N_7619);
nor U8362 (N_8362,N_7516,N_7725);
nor U8363 (N_8363,N_7784,N_7869);
nand U8364 (N_8364,N_7891,N_7802);
nor U8365 (N_8365,N_7646,N_7800);
or U8366 (N_8366,N_7882,N_7762);
xnor U8367 (N_8367,N_7741,N_7644);
xor U8368 (N_8368,N_7800,N_7643);
nor U8369 (N_8369,N_7941,N_7694);
nand U8370 (N_8370,N_7959,N_7885);
xnor U8371 (N_8371,N_7618,N_7777);
nand U8372 (N_8372,N_7652,N_7525);
or U8373 (N_8373,N_7764,N_7881);
xor U8374 (N_8374,N_7897,N_7658);
nand U8375 (N_8375,N_7907,N_7776);
and U8376 (N_8376,N_7746,N_7825);
and U8377 (N_8377,N_7926,N_7844);
nand U8378 (N_8378,N_7814,N_7587);
or U8379 (N_8379,N_7512,N_7687);
or U8380 (N_8380,N_7828,N_7987);
xnor U8381 (N_8381,N_7984,N_7800);
xnor U8382 (N_8382,N_7705,N_7889);
nor U8383 (N_8383,N_7995,N_7514);
or U8384 (N_8384,N_7662,N_7614);
and U8385 (N_8385,N_7531,N_7725);
and U8386 (N_8386,N_7780,N_7920);
and U8387 (N_8387,N_7685,N_7649);
or U8388 (N_8388,N_7897,N_7685);
nand U8389 (N_8389,N_7795,N_7596);
nand U8390 (N_8390,N_7682,N_7665);
nand U8391 (N_8391,N_7659,N_7957);
or U8392 (N_8392,N_7861,N_7988);
nand U8393 (N_8393,N_7633,N_7505);
nor U8394 (N_8394,N_7614,N_7827);
xnor U8395 (N_8395,N_7524,N_7626);
nand U8396 (N_8396,N_7567,N_7773);
or U8397 (N_8397,N_7509,N_7603);
or U8398 (N_8398,N_7985,N_7890);
and U8399 (N_8399,N_7902,N_7713);
xor U8400 (N_8400,N_7628,N_7712);
or U8401 (N_8401,N_7730,N_7906);
and U8402 (N_8402,N_7703,N_7732);
and U8403 (N_8403,N_7747,N_7695);
nand U8404 (N_8404,N_7698,N_7956);
xnor U8405 (N_8405,N_7544,N_7753);
nor U8406 (N_8406,N_7709,N_7830);
and U8407 (N_8407,N_7875,N_7552);
nor U8408 (N_8408,N_7932,N_7816);
nor U8409 (N_8409,N_7946,N_7867);
and U8410 (N_8410,N_7730,N_7894);
or U8411 (N_8411,N_7677,N_7529);
nor U8412 (N_8412,N_7944,N_7632);
nand U8413 (N_8413,N_7670,N_7611);
xor U8414 (N_8414,N_7828,N_7999);
nand U8415 (N_8415,N_7996,N_7768);
nor U8416 (N_8416,N_7788,N_7712);
xnor U8417 (N_8417,N_7960,N_7790);
or U8418 (N_8418,N_7798,N_7910);
and U8419 (N_8419,N_7981,N_7639);
nor U8420 (N_8420,N_7797,N_7901);
nor U8421 (N_8421,N_7560,N_7509);
or U8422 (N_8422,N_7514,N_7754);
nor U8423 (N_8423,N_7557,N_7706);
and U8424 (N_8424,N_7956,N_7973);
nor U8425 (N_8425,N_7826,N_7819);
nand U8426 (N_8426,N_7919,N_7918);
xnor U8427 (N_8427,N_7657,N_7817);
or U8428 (N_8428,N_7553,N_7799);
nand U8429 (N_8429,N_7555,N_7821);
or U8430 (N_8430,N_7501,N_7761);
and U8431 (N_8431,N_7790,N_7548);
nor U8432 (N_8432,N_7905,N_7945);
or U8433 (N_8433,N_7689,N_7969);
nor U8434 (N_8434,N_7774,N_7759);
nand U8435 (N_8435,N_7789,N_7942);
and U8436 (N_8436,N_7610,N_7743);
nor U8437 (N_8437,N_7684,N_7594);
and U8438 (N_8438,N_7558,N_7685);
and U8439 (N_8439,N_7611,N_7842);
or U8440 (N_8440,N_7843,N_7682);
and U8441 (N_8441,N_7851,N_7614);
nand U8442 (N_8442,N_7524,N_7761);
and U8443 (N_8443,N_7772,N_7575);
nand U8444 (N_8444,N_7725,N_7675);
nor U8445 (N_8445,N_7839,N_7759);
nand U8446 (N_8446,N_7987,N_7845);
or U8447 (N_8447,N_7743,N_7762);
xor U8448 (N_8448,N_7543,N_7900);
nand U8449 (N_8449,N_7566,N_7693);
or U8450 (N_8450,N_7816,N_7992);
nand U8451 (N_8451,N_7568,N_7803);
nand U8452 (N_8452,N_7670,N_7696);
nand U8453 (N_8453,N_7784,N_7844);
and U8454 (N_8454,N_7589,N_7990);
nand U8455 (N_8455,N_7791,N_7553);
xor U8456 (N_8456,N_7701,N_7804);
nor U8457 (N_8457,N_7559,N_7960);
nor U8458 (N_8458,N_7907,N_7956);
nor U8459 (N_8459,N_7762,N_7540);
and U8460 (N_8460,N_7937,N_7594);
xor U8461 (N_8461,N_7932,N_7795);
and U8462 (N_8462,N_7703,N_7881);
nor U8463 (N_8463,N_7925,N_7815);
or U8464 (N_8464,N_7598,N_7913);
xnor U8465 (N_8465,N_7591,N_7926);
nand U8466 (N_8466,N_7618,N_7725);
xnor U8467 (N_8467,N_7855,N_7765);
nor U8468 (N_8468,N_7883,N_7554);
or U8469 (N_8469,N_7722,N_7770);
nor U8470 (N_8470,N_7914,N_7821);
nand U8471 (N_8471,N_7546,N_7948);
xnor U8472 (N_8472,N_7767,N_7914);
nor U8473 (N_8473,N_7766,N_7653);
nand U8474 (N_8474,N_7994,N_7523);
nand U8475 (N_8475,N_7646,N_7871);
nor U8476 (N_8476,N_7765,N_7540);
nor U8477 (N_8477,N_7522,N_7891);
nand U8478 (N_8478,N_7820,N_7979);
xnor U8479 (N_8479,N_7608,N_7638);
nor U8480 (N_8480,N_7724,N_7534);
nand U8481 (N_8481,N_7807,N_7958);
xor U8482 (N_8482,N_7524,N_7701);
and U8483 (N_8483,N_7717,N_7724);
nand U8484 (N_8484,N_7622,N_7979);
xor U8485 (N_8485,N_7943,N_7727);
nand U8486 (N_8486,N_7992,N_7970);
nand U8487 (N_8487,N_7950,N_7906);
and U8488 (N_8488,N_7604,N_7719);
and U8489 (N_8489,N_7560,N_7821);
nor U8490 (N_8490,N_7843,N_7897);
or U8491 (N_8491,N_7848,N_7886);
nand U8492 (N_8492,N_7885,N_7533);
and U8493 (N_8493,N_7941,N_7956);
or U8494 (N_8494,N_7515,N_7682);
xor U8495 (N_8495,N_7662,N_7966);
or U8496 (N_8496,N_7668,N_7715);
or U8497 (N_8497,N_7793,N_7535);
and U8498 (N_8498,N_7821,N_7876);
or U8499 (N_8499,N_7682,N_7595);
or U8500 (N_8500,N_8017,N_8347);
nand U8501 (N_8501,N_8218,N_8316);
or U8502 (N_8502,N_8479,N_8093);
nor U8503 (N_8503,N_8443,N_8380);
or U8504 (N_8504,N_8451,N_8005);
and U8505 (N_8505,N_8014,N_8225);
nor U8506 (N_8506,N_8373,N_8107);
xor U8507 (N_8507,N_8294,N_8145);
and U8508 (N_8508,N_8400,N_8047);
nand U8509 (N_8509,N_8421,N_8442);
or U8510 (N_8510,N_8423,N_8362);
xnor U8511 (N_8511,N_8063,N_8169);
nand U8512 (N_8512,N_8385,N_8016);
or U8513 (N_8513,N_8110,N_8072);
or U8514 (N_8514,N_8130,N_8279);
and U8515 (N_8515,N_8139,N_8413);
or U8516 (N_8516,N_8010,N_8492);
nor U8517 (N_8517,N_8303,N_8314);
xor U8518 (N_8518,N_8231,N_8357);
and U8519 (N_8519,N_8418,N_8074);
or U8520 (N_8520,N_8354,N_8160);
or U8521 (N_8521,N_8336,N_8037);
and U8522 (N_8522,N_8235,N_8477);
or U8523 (N_8523,N_8219,N_8481);
or U8524 (N_8524,N_8104,N_8426);
nor U8525 (N_8525,N_8468,N_8482);
nand U8526 (N_8526,N_8226,N_8113);
and U8527 (N_8527,N_8197,N_8004);
nor U8528 (N_8528,N_8064,N_8236);
or U8529 (N_8529,N_8199,N_8419);
and U8530 (N_8530,N_8227,N_8365);
and U8531 (N_8531,N_8048,N_8174);
xnor U8532 (N_8532,N_8080,N_8390);
nor U8533 (N_8533,N_8313,N_8458);
xnor U8534 (N_8534,N_8209,N_8150);
nor U8535 (N_8535,N_8252,N_8499);
nor U8536 (N_8536,N_8353,N_8082);
nand U8537 (N_8537,N_8059,N_8285);
nand U8538 (N_8538,N_8292,N_8310);
nand U8539 (N_8539,N_8340,N_8319);
nor U8540 (N_8540,N_8154,N_8360);
or U8541 (N_8541,N_8432,N_8325);
nand U8542 (N_8542,N_8301,N_8156);
nor U8543 (N_8543,N_8166,N_8454);
or U8544 (N_8544,N_8031,N_8214);
nand U8545 (N_8545,N_8062,N_8051);
nor U8546 (N_8546,N_8484,N_8459);
and U8547 (N_8547,N_8223,N_8403);
nor U8548 (N_8548,N_8321,N_8341);
or U8549 (N_8549,N_8186,N_8024);
xor U8550 (N_8550,N_8015,N_8368);
nor U8551 (N_8551,N_8159,N_8351);
or U8552 (N_8552,N_8053,N_8241);
and U8553 (N_8553,N_8355,N_8034);
nor U8554 (N_8554,N_8431,N_8334);
xor U8555 (N_8555,N_8006,N_8411);
or U8556 (N_8556,N_8297,N_8405);
nand U8557 (N_8557,N_8305,N_8125);
nor U8558 (N_8558,N_8018,N_8455);
xnor U8559 (N_8559,N_8069,N_8149);
nor U8560 (N_8560,N_8138,N_8157);
and U8561 (N_8561,N_8302,N_8307);
or U8562 (N_8562,N_8030,N_8120);
or U8563 (N_8563,N_8194,N_8094);
and U8564 (N_8564,N_8488,N_8372);
nor U8565 (N_8565,N_8245,N_8165);
nor U8566 (N_8566,N_8021,N_8466);
or U8567 (N_8567,N_8119,N_8280);
xnor U8568 (N_8568,N_8461,N_8193);
or U8569 (N_8569,N_8060,N_8367);
and U8570 (N_8570,N_8128,N_8212);
and U8571 (N_8571,N_8115,N_8439);
nor U8572 (N_8572,N_8124,N_8498);
or U8573 (N_8573,N_8260,N_8433);
nand U8574 (N_8574,N_8382,N_8295);
xnor U8575 (N_8575,N_8487,N_8050);
xnor U8576 (N_8576,N_8163,N_8425);
nand U8577 (N_8577,N_8134,N_8198);
or U8578 (N_8578,N_8462,N_8167);
and U8579 (N_8579,N_8386,N_8127);
or U8580 (N_8580,N_8438,N_8478);
and U8581 (N_8581,N_8299,N_8108);
nand U8582 (N_8582,N_8079,N_8338);
and U8583 (N_8583,N_8315,N_8333);
or U8584 (N_8584,N_8464,N_8114);
nand U8585 (N_8585,N_8475,N_8417);
and U8586 (N_8586,N_8308,N_8287);
xor U8587 (N_8587,N_8217,N_8269);
nor U8588 (N_8588,N_8249,N_8262);
nor U8589 (N_8589,N_8078,N_8320);
nand U8590 (N_8590,N_8151,N_8181);
nor U8591 (N_8591,N_8486,N_8456);
nand U8592 (N_8592,N_8126,N_8045);
nor U8593 (N_8593,N_8187,N_8137);
xor U8594 (N_8594,N_8268,N_8201);
nand U8595 (N_8595,N_8039,N_8026);
nor U8596 (N_8596,N_8389,N_8027);
nor U8597 (N_8597,N_8440,N_8102);
nand U8598 (N_8598,N_8324,N_8189);
and U8599 (N_8599,N_8258,N_8391);
nand U8600 (N_8600,N_8452,N_8396);
or U8601 (N_8601,N_8270,N_8012);
xnor U8602 (N_8602,N_8422,N_8264);
or U8603 (N_8603,N_8066,N_8098);
and U8604 (N_8604,N_8430,N_8318);
xnor U8605 (N_8605,N_8011,N_8434);
nor U8606 (N_8606,N_8331,N_8061);
xnor U8607 (N_8607,N_8447,N_8207);
nand U8608 (N_8608,N_8146,N_8106);
xnor U8609 (N_8609,N_8091,N_8083);
xor U8610 (N_8610,N_8490,N_8099);
nor U8611 (N_8611,N_8042,N_8469);
xnor U8612 (N_8612,N_8428,N_8095);
nor U8613 (N_8613,N_8435,N_8029);
or U8614 (N_8614,N_8398,N_8195);
or U8615 (N_8615,N_8075,N_8446);
or U8616 (N_8616,N_8046,N_8058);
xor U8617 (N_8617,N_8474,N_8101);
and U8618 (N_8618,N_8261,N_8376);
nand U8619 (N_8619,N_8276,N_8494);
nand U8620 (N_8620,N_8179,N_8040);
nor U8621 (N_8621,N_8228,N_8483);
nor U8622 (N_8622,N_8142,N_8077);
nor U8623 (N_8623,N_8412,N_8274);
xor U8624 (N_8624,N_8265,N_8123);
nor U8625 (N_8625,N_8144,N_8222);
nor U8626 (N_8626,N_8416,N_8089);
nand U8627 (N_8627,N_8251,N_8164);
or U8628 (N_8628,N_8073,N_8346);
nor U8629 (N_8629,N_8344,N_8387);
nand U8630 (N_8630,N_8076,N_8087);
or U8631 (N_8631,N_8259,N_8323);
nor U8632 (N_8632,N_8208,N_8190);
nand U8633 (N_8633,N_8381,N_8103);
nand U8634 (N_8634,N_8427,N_8086);
nand U8635 (N_8635,N_8022,N_8003);
nor U8636 (N_8636,N_8122,N_8304);
and U8637 (N_8637,N_8441,N_8306);
and U8638 (N_8638,N_8178,N_8415);
nand U8639 (N_8639,N_8445,N_8001);
or U8640 (N_8640,N_8211,N_8298);
nand U8641 (N_8641,N_8350,N_8049);
nor U8642 (N_8642,N_8096,N_8052);
and U8643 (N_8643,N_8343,N_8491);
nor U8644 (N_8644,N_8028,N_8172);
nand U8645 (N_8645,N_8448,N_8131);
and U8646 (N_8646,N_8271,N_8256);
or U8647 (N_8647,N_8352,N_8369);
nor U8648 (N_8648,N_8023,N_8255);
or U8649 (N_8649,N_8007,N_8129);
and U8650 (N_8650,N_8329,N_8202);
nand U8651 (N_8651,N_8132,N_8224);
xnor U8652 (N_8652,N_8035,N_8311);
nand U8653 (N_8653,N_8230,N_8170);
and U8654 (N_8654,N_8493,N_8221);
and U8655 (N_8655,N_8084,N_8229);
nand U8656 (N_8656,N_8210,N_8277);
nand U8657 (N_8657,N_8288,N_8008);
xnor U8658 (N_8658,N_8100,N_8188);
and U8659 (N_8659,N_8240,N_8032);
or U8660 (N_8660,N_8092,N_8238);
nor U8661 (N_8661,N_8196,N_8476);
or U8662 (N_8662,N_8286,N_8359);
nor U8663 (N_8663,N_8410,N_8135);
and U8664 (N_8664,N_8436,N_8081);
xnor U8665 (N_8665,N_8266,N_8097);
xor U8666 (N_8666,N_8000,N_8065);
xnor U8667 (N_8667,N_8384,N_8056);
nor U8668 (N_8668,N_8054,N_8192);
and U8669 (N_8669,N_8275,N_8019);
xor U8670 (N_8670,N_8383,N_8471);
nand U8671 (N_8671,N_8257,N_8473);
and U8672 (N_8672,N_8183,N_8282);
nor U8673 (N_8673,N_8267,N_8239);
nand U8674 (N_8674,N_8155,N_8407);
nor U8675 (N_8675,N_8068,N_8133);
or U8676 (N_8676,N_8044,N_8116);
or U8677 (N_8677,N_8401,N_8013);
and U8678 (N_8678,N_8363,N_8136);
and U8679 (N_8679,N_8215,N_8370);
and U8680 (N_8680,N_8033,N_8450);
and U8681 (N_8681,N_8467,N_8495);
nand U8682 (N_8682,N_8345,N_8220);
or U8683 (N_8683,N_8420,N_8278);
nand U8684 (N_8684,N_8472,N_8109);
and U8685 (N_8685,N_8337,N_8379);
and U8686 (N_8686,N_8168,N_8088);
and U8687 (N_8687,N_8457,N_8200);
or U8688 (N_8688,N_8090,N_8254);
nand U8689 (N_8689,N_8429,N_8025);
nor U8690 (N_8690,N_8247,N_8496);
nand U8691 (N_8691,N_8465,N_8444);
nand U8692 (N_8692,N_8205,N_8289);
nand U8693 (N_8693,N_8140,N_8147);
and U8694 (N_8694,N_8161,N_8424);
or U8695 (N_8695,N_8206,N_8349);
nor U8696 (N_8696,N_8284,N_8180);
nor U8697 (N_8697,N_8148,N_8393);
xor U8698 (N_8698,N_8002,N_8191);
nor U8699 (N_8699,N_8463,N_8406);
or U8700 (N_8700,N_8071,N_8300);
or U8701 (N_8701,N_8041,N_8397);
nand U8702 (N_8702,N_8453,N_8118);
or U8703 (N_8703,N_8246,N_8317);
or U8704 (N_8704,N_8158,N_8296);
nand U8705 (N_8705,N_8105,N_8204);
and U8706 (N_8706,N_8348,N_8009);
nor U8707 (N_8707,N_8489,N_8171);
or U8708 (N_8708,N_8460,N_8408);
xor U8709 (N_8709,N_8480,N_8244);
xor U8710 (N_8710,N_8162,N_8470);
nor U8711 (N_8711,N_8392,N_8233);
nand U8712 (N_8712,N_8366,N_8388);
nand U8713 (N_8713,N_8273,N_8356);
nor U8714 (N_8714,N_8243,N_8020);
nor U8715 (N_8715,N_8332,N_8112);
and U8716 (N_8716,N_8043,N_8409);
nand U8717 (N_8717,N_8399,N_8248);
nor U8718 (N_8718,N_8377,N_8326);
and U8719 (N_8719,N_8358,N_8152);
nand U8720 (N_8720,N_8404,N_8177);
or U8721 (N_8721,N_8290,N_8036);
xor U8722 (N_8722,N_8361,N_8485);
xnor U8723 (N_8723,N_8395,N_8176);
and U8724 (N_8724,N_8414,N_8253);
nand U8725 (N_8725,N_8272,N_8281);
nor U8726 (N_8726,N_8242,N_8234);
nor U8727 (N_8727,N_8497,N_8213);
xnor U8728 (N_8728,N_8143,N_8291);
and U8729 (N_8729,N_8250,N_8309);
nand U8730 (N_8730,N_8070,N_8216);
or U8731 (N_8731,N_8339,N_8182);
xor U8732 (N_8732,N_8237,N_8312);
and U8733 (N_8733,N_8085,N_8111);
and U8734 (N_8734,N_8184,N_8371);
and U8735 (N_8735,N_8394,N_8117);
nand U8736 (N_8736,N_8038,N_8330);
nor U8737 (N_8737,N_8402,N_8232);
nand U8738 (N_8738,N_8283,N_8327);
or U8739 (N_8739,N_8374,N_8437);
nor U8740 (N_8740,N_8364,N_8449);
or U8741 (N_8741,N_8057,N_8378);
nand U8742 (N_8742,N_8203,N_8342);
and U8743 (N_8743,N_8322,N_8335);
and U8744 (N_8744,N_8067,N_8055);
nand U8745 (N_8745,N_8141,N_8175);
nand U8746 (N_8746,N_8375,N_8328);
nand U8747 (N_8747,N_8293,N_8185);
xnor U8748 (N_8748,N_8263,N_8173);
or U8749 (N_8749,N_8153,N_8121);
and U8750 (N_8750,N_8095,N_8485);
nor U8751 (N_8751,N_8373,N_8109);
xor U8752 (N_8752,N_8050,N_8241);
xnor U8753 (N_8753,N_8302,N_8010);
nand U8754 (N_8754,N_8116,N_8415);
xor U8755 (N_8755,N_8434,N_8450);
and U8756 (N_8756,N_8006,N_8366);
nand U8757 (N_8757,N_8182,N_8021);
nand U8758 (N_8758,N_8362,N_8354);
and U8759 (N_8759,N_8359,N_8143);
or U8760 (N_8760,N_8195,N_8054);
nand U8761 (N_8761,N_8098,N_8325);
nand U8762 (N_8762,N_8353,N_8426);
and U8763 (N_8763,N_8197,N_8457);
or U8764 (N_8764,N_8017,N_8087);
and U8765 (N_8765,N_8124,N_8000);
or U8766 (N_8766,N_8123,N_8414);
nor U8767 (N_8767,N_8495,N_8356);
nor U8768 (N_8768,N_8281,N_8386);
and U8769 (N_8769,N_8123,N_8344);
xnor U8770 (N_8770,N_8012,N_8110);
or U8771 (N_8771,N_8288,N_8351);
xor U8772 (N_8772,N_8337,N_8390);
nand U8773 (N_8773,N_8135,N_8429);
nor U8774 (N_8774,N_8084,N_8275);
and U8775 (N_8775,N_8327,N_8209);
or U8776 (N_8776,N_8272,N_8208);
nand U8777 (N_8777,N_8245,N_8026);
and U8778 (N_8778,N_8241,N_8489);
xnor U8779 (N_8779,N_8033,N_8179);
nand U8780 (N_8780,N_8367,N_8442);
nand U8781 (N_8781,N_8318,N_8445);
nand U8782 (N_8782,N_8049,N_8448);
or U8783 (N_8783,N_8326,N_8095);
or U8784 (N_8784,N_8499,N_8114);
nor U8785 (N_8785,N_8122,N_8021);
or U8786 (N_8786,N_8267,N_8118);
and U8787 (N_8787,N_8188,N_8189);
and U8788 (N_8788,N_8441,N_8034);
nor U8789 (N_8789,N_8368,N_8420);
and U8790 (N_8790,N_8361,N_8200);
xnor U8791 (N_8791,N_8078,N_8440);
nand U8792 (N_8792,N_8222,N_8241);
or U8793 (N_8793,N_8017,N_8301);
or U8794 (N_8794,N_8094,N_8408);
xnor U8795 (N_8795,N_8087,N_8234);
and U8796 (N_8796,N_8093,N_8018);
nor U8797 (N_8797,N_8226,N_8026);
or U8798 (N_8798,N_8111,N_8370);
or U8799 (N_8799,N_8174,N_8387);
and U8800 (N_8800,N_8135,N_8444);
or U8801 (N_8801,N_8109,N_8264);
nand U8802 (N_8802,N_8364,N_8026);
nand U8803 (N_8803,N_8198,N_8218);
or U8804 (N_8804,N_8264,N_8483);
or U8805 (N_8805,N_8043,N_8071);
nand U8806 (N_8806,N_8394,N_8372);
nand U8807 (N_8807,N_8012,N_8337);
or U8808 (N_8808,N_8275,N_8059);
and U8809 (N_8809,N_8241,N_8483);
or U8810 (N_8810,N_8318,N_8195);
and U8811 (N_8811,N_8025,N_8451);
or U8812 (N_8812,N_8392,N_8118);
nor U8813 (N_8813,N_8107,N_8415);
nand U8814 (N_8814,N_8111,N_8278);
nand U8815 (N_8815,N_8152,N_8483);
nand U8816 (N_8816,N_8314,N_8353);
or U8817 (N_8817,N_8358,N_8254);
nor U8818 (N_8818,N_8029,N_8442);
nor U8819 (N_8819,N_8238,N_8374);
or U8820 (N_8820,N_8497,N_8225);
or U8821 (N_8821,N_8119,N_8327);
nor U8822 (N_8822,N_8144,N_8102);
and U8823 (N_8823,N_8172,N_8035);
xnor U8824 (N_8824,N_8478,N_8298);
or U8825 (N_8825,N_8228,N_8110);
and U8826 (N_8826,N_8086,N_8276);
and U8827 (N_8827,N_8400,N_8491);
nor U8828 (N_8828,N_8096,N_8351);
or U8829 (N_8829,N_8437,N_8439);
or U8830 (N_8830,N_8192,N_8235);
nor U8831 (N_8831,N_8257,N_8322);
nand U8832 (N_8832,N_8391,N_8381);
nor U8833 (N_8833,N_8455,N_8098);
xor U8834 (N_8834,N_8155,N_8053);
and U8835 (N_8835,N_8293,N_8115);
nand U8836 (N_8836,N_8185,N_8254);
xor U8837 (N_8837,N_8050,N_8243);
xor U8838 (N_8838,N_8414,N_8366);
nand U8839 (N_8839,N_8487,N_8346);
and U8840 (N_8840,N_8448,N_8288);
and U8841 (N_8841,N_8255,N_8399);
nand U8842 (N_8842,N_8093,N_8355);
nand U8843 (N_8843,N_8435,N_8272);
or U8844 (N_8844,N_8406,N_8457);
or U8845 (N_8845,N_8468,N_8154);
and U8846 (N_8846,N_8228,N_8417);
or U8847 (N_8847,N_8067,N_8274);
or U8848 (N_8848,N_8264,N_8148);
or U8849 (N_8849,N_8069,N_8087);
nor U8850 (N_8850,N_8112,N_8432);
and U8851 (N_8851,N_8220,N_8141);
and U8852 (N_8852,N_8086,N_8195);
and U8853 (N_8853,N_8001,N_8088);
and U8854 (N_8854,N_8454,N_8311);
nand U8855 (N_8855,N_8109,N_8492);
or U8856 (N_8856,N_8143,N_8002);
nand U8857 (N_8857,N_8415,N_8031);
xor U8858 (N_8858,N_8151,N_8007);
xor U8859 (N_8859,N_8185,N_8152);
xor U8860 (N_8860,N_8252,N_8375);
xor U8861 (N_8861,N_8301,N_8280);
nor U8862 (N_8862,N_8342,N_8150);
and U8863 (N_8863,N_8322,N_8344);
or U8864 (N_8864,N_8276,N_8332);
or U8865 (N_8865,N_8242,N_8250);
xnor U8866 (N_8866,N_8388,N_8201);
nor U8867 (N_8867,N_8037,N_8033);
and U8868 (N_8868,N_8010,N_8320);
nand U8869 (N_8869,N_8354,N_8486);
and U8870 (N_8870,N_8198,N_8061);
nor U8871 (N_8871,N_8062,N_8095);
or U8872 (N_8872,N_8473,N_8023);
nand U8873 (N_8873,N_8492,N_8142);
or U8874 (N_8874,N_8362,N_8474);
and U8875 (N_8875,N_8089,N_8430);
xnor U8876 (N_8876,N_8012,N_8457);
nand U8877 (N_8877,N_8132,N_8077);
xnor U8878 (N_8878,N_8352,N_8312);
or U8879 (N_8879,N_8137,N_8135);
and U8880 (N_8880,N_8057,N_8373);
or U8881 (N_8881,N_8382,N_8047);
nand U8882 (N_8882,N_8069,N_8433);
nand U8883 (N_8883,N_8467,N_8130);
nor U8884 (N_8884,N_8062,N_8262);
and U8885 (N_8885,N_8284,N_8255);
nand U8886 (N_8886,N_8167,N_8094);
or U8887 (N_8887,N_8096,N_8048);
xnor U8888 (N_8888,N_8109,N_8145);
nand U8889 (N_8889,N_8322,N_8408);
nor U8890 (N_8890,N_8327,N_8163);
nand U8891 (N_8891,N_8003,N_8238);
nand U8892 (N_8892,N_8249,N_8190);
and U8893 (N_8893,N_8292,N_8457);
and U8894 (N_8894,N_8099,N_8315);
xor U8895 (N_8895,N_8309,N_8346);
and U8896 (N_8896,N_8320,N_8292);
or U8897 (N_8897,N_8066,N_8413);
nor U8898 (N_8898,N_8316,N_8214);
and U8899 (N_8899,N_8134,N_8210);
xnor U8900 (N_8900,N_8152,N_8298);
or U8901 (N_8901,N_8146,N_8029);
nand U8902 (N_8902,N_8077,N_8242);
nor U8903 (N_8903,N_8369,N_8154);
nand U8904 (N_8904,N_8120,N_8224);
or U8905 (N_8905,N_8407,N_8122);
and U8906 (N_8906,N_8012,N_8240);
nand U8907 (N_8907,N_8344,N_8240);
nor U8908 (N_8908,N_8147,N_8030);
and U8909 (N_8909,N_8306,N_8404);
nand U8910 (N_8910,N_8423,N_8307);
nor U8911 (N_8911,N_8299,N_8301);
xor U8912 (N_8912,N_8351,N_8327);
nand U8913 (N_8913,N_8148,N_8155);
nand U8914 (N_8914,N_8170,N_8071);
nand U8915 (N_8915,N_8069,N_8155);
or U8916 (N_8916,N_8473,N_8235);
and U8917 (N_8917,N_8243,N_8130);
nand U8918 (N_8918,N_8198,N_8157);
and U8919 (N_8919,N_8194,N_8228);
or U8920 (N_8920,N_8014,N_8255);
nand U8921 (N_8921,N_8273,N_8066);
and U8922 (N_8922,N_8333,N_8043);
or U8923 (N_8923,N_8194,N_8251);
nor U8924 (N_8924,N_8006,N_8048);
nor U8925 (N_8925,N_8473,N_8223);
or U8926 (N_8926,N_8483,N_8319);
nand U8927 (N_8927,N_8319,N_8241);
nand U8928 (N_8928,N_8433,N_8155);
xor U8929 (N_8929,N_8377,N_8330);
xnor U8930 (N_8930,N_8430,N_8450);
xor U8931 (N_8931,N_8445,N_8320);
nor U8932 (N_8932,N_8340,N_8454);
and U8933 (N_8933,N_8193,N_8233);
xor U8934 (N_8934,N_8071,N_8493);
and U8935 (N_8935,N_8350,N_8214);
xnor U8936 (N_8936,N_8284,N_8437);
xnor U8937 (N_8937,N_8038,N_8233);
nand U8938 (N_8938,N_8091,N_8002);
and U8939 (N_8939,N_8029,N_8306);
xnor U8940 (N_8940,N_8353,N_8342);
or U8941 (N_8941,N_8252,N_8171);
xor U8942 (N_8942,N_8433,N_8025);
and U8943 (N_8943,N_8287,N_8403);
nand U8944 (N_8944,N_8108,N_8214);
nor U8945 (N_8945,N_8393,N_8363);
xnor U8946 (N_8946,N_8301,N_8352);
nand U8947 (N_8947,N_8102,N_8175);
nand U8948 (N_8948,N_8201,N_8219);
or U8949 (N_8949,N_8452,N_8353);
nor U8950 (N_8950,N_8246,N_8356);
xnor U8951 (N_8951,N_8044,N_8134);
nand U8952 (N_8952,N_8153,N_8183);
and U8953 (N_8953,N_8391,N_8395);
nand U8954 (N_8954,N_8246,N_8490);
and U8955 (N_8955,N_8107,N_8334);
nand U8956 (N_8956,N_8135,N_8321);
nand U8957 (N_8957,N_8005,N_8386);
or U8958 (N_8958,N_8013,N_8107);
nor U8959 (N_8959,N_8454,N_8133);
xnor U8960 (N_8960,N_8439,N_8042);
nand U8961 (N_8961,N_8227,N_8443);
and U8962 (N_8962,N_8300,N_8106);
xor U8963 (N_8963,N_8148,N_8086);
nand U8964 (N_8964,N_8228,N_8411);
or U8965 (N_8965,N_8072,N_8070);
nand U8966 (N_8966,N_8087,N_8114);
and U8967 (N_8967,N_8032,N_8036);
nand U8968 (N_8968,N_8392,N_8141);
and U8969 (N_8969,N_8344,N_8021);
nor U8970 (N_8970,N_8201,N_8063);
xor U8971 (N_8971,N_8362,N_8200);
and U8972 (N_8972,N_8063,N_8214);
xor U8973 (N_8973,N_8193,N_8395);
xnor U8974 (N_8974,N_8051,N_8386);
xor U8975 (N_8975,N_8198,N_8395);
nor U8976 (N_8976,N_8462,N_8420);
nand U8977 (N_8977,N_8463,N_8028);
or U8978 (N_8978,N_8382,N_8254);
or U8979 (N_8979,N_8468,N_8374);
nand U8980 (N_8980,N_8071,N_8144);
nand U8981 (N_8981,N_8194,N_8264);
nor U8982 (N_8982,N_8055,N_8347);
xor U8983 (N_8983,N_8067,N_8007);
and U8984 (N_8984,N_8051,N_8274);
xor U8985 (N_8985,N_8195,N_8155);
nand U8986 (N_8986,N_8011,N_8466);
nor U8987 (N_8987,N_8058,N_8435);
nand U8988 (N_8988,N_8385,N_8139);
or U8989 (N_8989,N_8272,N_8094);
or U8990 (N_8990,N_8053,N_8273);
or U8991 (N_8991,N_8362,N_8482);
xor U8992 (N_8992,N_8394,N_8217);
xor U8993 (N_8993,N_8330,N_8404);
nor U8994 (N_8994,N_8134,N_8416);
or U8995 (N_8995,N_8449,N_8219);
xor U8996 (N_8996,N_8269,N_8349);
nor U8997 (N_8997,N_8099,N_8198);
and U8998 (N_8998,N_8128,N_8095);
nand U8999 (N_8999,N_8071,N_8160);
or U9000 (N_9000,N_8708,N_8858);
xor U9001 (N_9001,N_8726,N_8873);
nand U9002 (N_9002,N_8599,N_8997);
nor U9003 (N_9003,N_8821,N_8638);
or U9004 (N_9004,N_8665,N_8981);
or U9005 (N_9005,N_8856,N_8768);
nor U9006 (N_9006,N_8794,N_8795);
or U9007 (N_9007,N_8644,N_8790);
xor U9008 (N_9008,N_8612,N_8639);
nor U9009 (N_9009,N_8525,N_8719);
nor U9010 (N_9010,N_8829,N_8597);
nand U9011 (N_9011,N_8540,N_8667);
or U9012 (N_9012,N_8986,N_8811);
nand U9013 (N_9013,N_8890,N_8658);
nor U9014 (N_9014,N_8534,N_8961);
xor U9015 (N_9015,N_8637,N_8578);
and U9016 (N_9016,N_8931,N_8527);
xor U9017 (N_9017,N_8993,N_8572);
or U9018 (N_9018,N_8879,N_8753);
xnor U9019 (N_9019,N_8636,N_8867);
nand U9020 (N_9020,N_8985,N_8747);
xor U9021 (N_9021,N_8505,N_8625);
and U9022 (N_9022,N_8860,N_8514);
and U9023 (N_9023,N_8691,N_8940);
or U9024 (N_9024,N_8610,N_8656);
or U9025 (N_9025,N_8617,N_8769);
and U9026 (N_9026,N_8774,N_8882);
nor U9027 (N_9027,N_8998,N_8586);
nand U9028 (N_9028,N_8960,N_8651);
or U9029 (N_9029,N_8508,N_8573);
or U9030 (N_9030,N_8903,N_8511);
xor U9031 (N_9031,N_8634,N_8593);
or U9032 (N_9032,N_8605,N_8977);
nand U9033 (N_9033,N_8800,N_8789);
and U9034 (N_9034,N_8904,N_8681);
and U9035 (N_9035,N_8854,N_8934);
and U9036 (N_9036,N_8584,N_8976);
or U9037 (N_9037,N_8746,N_8884);
nor U9038 (N_9038,N_8711,N_8836);
nor U9039 (N_9039,N_8996,N_8580);
or U9040 (N_9040,N_8878,N_8504);
or U9041 (N_9041,N_8616,N_8751);
nor U9042 (N_9042,N_8863,N_8921);
nor U9043 (N_9043,N_8798,N_8547);
nor U9044 (N_9044,N_8980,N_8883);
nand U9045 (N_9045,N_8892,N_8978);
nand U9046 (N_9046,N_8835,N_8861);
nand U9047 (N_9047,N_8692,N_8728);
xnor U9048 (N_9048,N_8518,N_8660);
nand U9049 (N_9049,N_8603,N_8994);
or U9050 (N_9050,N_8913,N_8569);
nand U9051 (N_9051,N_8696,N_8783);
and U9052 (N_9052,N_8983,N_8995);
and U9053 (N_9053,N_8515,N_8770);
and U9054 (N_9054,N_8955,N_8833);
or U9055 (N_9055,N_8530,N_8552);
or U9056 (N_9056,N_8912,N_8686);
nand U9057 (N_9057,N_8548,N_8677);
or U9058 (N_9058,N_8652,N_8812);
xnor U9059 (N_9059,N_8763,N_8744);
nand U9060 (N_9060,N_8909,N_8704);
nand U9061 (N_9061,N_8896,N_8988);
xor U9062 (N_9062,N_8564,N_8533);
and U9063 (N_9063,N_8732,N_8780);
nor U9064 (N_9064,N_8643,N_8982);
or U9065 (N_9065,N_8698,N_8952);
or U9066 (N_9066,N_8999,N_8671);
xor U9067 (N_9067,N_8754,N_8619);
nand U9068 (N_9068,N_8694,N_8685);
xor U9069 (N_9069,N_8925,N_8648);
or U9070 (N_9070,N_8885,N_8672);
and U9071 (N_9071,N_8590,N_8874);
and U9072 (N_9072,N_8852,N_8693);
and U9073 (N_9073,N_8864,N_8814);
xnor U9074 (N_9074,N_8663,N_8826);
or U9075 (N_9075,N_8822,N_8908);
or U9076 (N_9076,N_8970,N_8801);
and U9077 (N_9077,N_8958,N_8992);
nor U9078 (N_9078,N_8521,N_8537);
and U9079 (N_9079,N_8777,N_8741);
xor U9080 (N_9080,N_8778,N_8897);
xor U9081 (N_9081,N_8804,N_8549);
nand U9082 (N_9082,N_8797,N_8556);
xor U9083 (N_9083,N_8635,N_8779);
or U9084 (N_9084,N_8786,N_8933);
xor U9085 (N_9085,N_8510,N_8872);
nand U9086 (N_9086,N_8680,N_8771);
nand U9087 (N_9087,N_8881,N_8784);
nand U9088 (N_9088,N_8932,N_8529);
or U9089 (N_9089,N_8966,N_8501);
or U9090 (N_9090,N_8760,N_8850);
or U9091 (N_9091,N_8902,N_8875);
and U9092 (N_9092,N_8948,N_8526);
or U9093 (N_9093,N_8827,N_8936);
or U9094 (N_9094,N_8690,N_8738);
xor U9095 (N_9095,N_8653,N_8733);
or U9096 (N_9096,N_8718,N_8642);
nor U9097 (N_9097,N_8848,N_8722);
or U9098 (N_9098,N_8766,N_8791);
xnor U9099 (N_9099,N_8944,N_8736);
nor U9100 (N_9100,N_8570,N_8755);
or U9101 (N_9101,N_8927,N_8624);
or U9102 (N_9102,N_8602,N_8938);
nor U9103 (N_9103,N_8654,N_8868);
nor U9104 (N_9104,N_8673,N_8893);
xnor U9105 (N_9105,N_8614,N_8689);
nand U9106 (N_9106,N_8825,N_8926);
and U9107 (N_9107,N_8946,N_8803);
or U9108 (N_9108,N_8675,N_8554);
or U9109 (N_9109,N_8661,N_8739);
and U9110 (N_9110,N_8703,N_8945);
or U9111 (N_9111,N_8532,N_8506);
nor U9112 (N_9112,N_8720,N_8713);
nand U9113 (N_9113,N_8965,N_8608);
nand U9114 (N_9114,N_8969,N_8664);
nand U9115 (N_9115,N_8849,N_8792);
nand U9116 (N_9116,N_8531,N_8716);
xnor U9117 (N_9117,N_8715,N_8595);
nand U9118 (N_9118,N_8757,N_8939);
nor U9119 (N_9119,N_8840,N_8895);
nand U9120 (N_9120,N_8851,N_8891);
nor U9121 (N_9121,N_8923,N_8846);
xor U9122 (N_9122,N_8581,N_8582);
xor U9123 (N_9123,N_8717,N_8973);
or U9124 (N_9124,N_8793,N_8576);
or U9125 (N_9125,N_8523,N_8679);
or U9126 (N_9126,N_8628,N_8669);
nor U9127 (N_9127,N_8745,N_8700);
or U9128 (N_9128,N_8963,N_8536);
or U9129 (N_9129,N_8916,N_8742);
xor U9130 (N_9130,N_8561,N_8641);
or U9131 (N_9131,N_8767,N_8839);
nor U9132 (N_9132,N_8919,N_8706);
or U9133 (N_9133,N_8756,N_8806);
nand U9134 (N_9134,N_8630,N_8830);
nor U9135 (N_9135,N_8964,N_8761);
nor U9136 (N_9136,N_8743,N_8551);
nand U9137 (N_9137,N_8606,N_8979);
or U9138 (N_9138,N_8705,N_8615);
or U9139 (N_9139,N_8538,N_8905);
nand U9140 (N_9140,N_8942,N_8750);
nor U9141 (N_9141,N_8772,N_8828);
xor U9142 (N_9142,N_8562,N_8972);
xor U9143 (N_9143,N_8947,N_8631);
or U9144 (N_9144,N_8735,N_8968);
nor U9145 (N_9145,N_8618,N_8596);
nand U9146 (N_9146,N_8729,N_8898);
xnor U9147 (N_9147,N_8876,N_8967);
or U9148 (N_9148,N_8853,N_8585);
and U9149 (N_9149,N_8598,N_8918);
or U9150 (N_9150,N_8799,N_8601);
nand U9151 (N_9151,N_8666,N_8781);
and U9152 (N_9152,N_8862,N_8687);
or U9153 (N_9153,N_8500,N_8502);
or U9154 (N_9154,N_8808,N_8727);
or U9155 (N_9155,N_8869,N_8503);
xnor U9156 (N_9156,N_8683,N_8871);
or U9157 (N_9157,N_8699,N_8640);
and U9158 (N_9158,N_8566,N_8843);
nor U9159 (N_9159,N_8920,N_8563);
or U9160 (N_9160,N_8788,N_8632);
nor U9161 (N_9161,N_8842,N_8915);
or U9162 (N_9162,N_8962,N_8818);
nand U9163 (N_9163,N_8650,N_8857);
or U9164 (N_9164,N_8588,N_8838);
nand U9165 (N_9165,N_8901,N_8560);
and U9166 (N_9166,N_8817,N_8620);
nor U9167 (N_9167,N_8987,N_8668);
nand U9168 (N_9168,N_8600,N_8712);
nand U9169 (N_9169,N_8541,N_8545);
xnor U9170 (N_9170,N_8579,N_8626);
nor U9171 (N_9171,N_8816,N_8522);
nor U9172 (N_9172,N_8906,N_8859);
and U9173 (N_9173,N_8929,N_8607);
xor U9174 (N_9174,N_8832,N_8855);
nand U9175 (N_9175,N_8678,N_8880);
and U9176 (N_9176,N_8975,N_8734);
or U9177 (N_9177,N_8701,N_8943);
and U9178 (N_9178,N_8785,N_8847);
and U9179 (N_9179,N_8834,N_8592);
or U9180 (N_9180,N_8819,N_8937);
nor U9181 (N_9181,N_8950,N_8910);
nor U9182 (N_9182,N_8528,N_8949);
nand U9183 (N_9183,N_8688,N_8609);
xnor U9184 (N_9184,N_8810,N_8623);
and U9185 (N_9185,N_8555,N_8796);
and U9186 (N_9186,N_8991,N_8737);
and U9187 (N_9187,N_8762,N_8622);
nor U9188 (N_9188,N_8647,N_8577);
nand U9189 (N_9189,N_8587,N_8574);
and U9190 (N_9190,N_8765,N_8759);
nor U9191 (N_9191,N_8613,N_8509);
or U9192 (N_9192,N_8928,N_8544);
or U9193 (N_9193,N_8894,N_8621);
xnor U9194 (N_9194,N_8655,N_8845);
or U9195 (N_9195,N_8870,N_8513);
or U9196 (N_9196,N_8813,N_8589);
xnor U9197 (N_9197,N_8917,N_8568);
nor U9198 (N_9198,N_8707,N_8752);
and U9199 (N_9199,N_8594,N_8725);
nor U9200 (N_9200,N_8709,N_8591);
or U9201 (N_9201,N_8740,N_8542);
and U9202 (N_9202,N_8990,N_8764);
and U9203 (N_9203,N_8837,N_8721);
nor U9204 (N_9204,N_8697,N_8831);
or U9205 (N_9205,N_8886,N_8900);
or U9206 (N_9206,N_8866,N_8517);
nand U9207 (N_9207,N_8558,N_8731);
or U9208 (N_9208,N_8604,N_8682);
and U9209 (N_9209,N_8662,N_8553);
xnor U9210 (N_9210,N_8714,N_8805);
xor U9211 (N_9211,N_8935,N_8889);
nor U9212 (N_9212,N_8914,N_8749);
nand U9213 (N_9213,N_8841,N_8565);
and U9214 (N_9214,N_8877,N_8670);
nand U9215 (N_9215,N_8758,N_8657);
and U9216 (N_9216,N_8611,N_8550);
xor U9217 (N_9217,N_8730,N_8695);
nor U9218 (N_9218,N_8512,N_8649);
xor U9219 (N_9219,N_8684,N_8802);
and U9220 (N_9220,N_8543,N_8951);
or U9221 (N_9221,N_8507,N_8748);
or U9222 (N_9222,N_8710,N_8559);
nand U9223 (N_9223,N_8844,N_8820);
xnor U9224 (N_9224,N_8899,N_8773);
or U9225 (N_9225,N_8583,N_8984);
and U9226 (N_9226,N_8887,N_8953);
nor U9227 (N_9227,N_8807,N_8930);
and U9228 (N_9228,N_8782,N_8775);
or U9229 (N_9229,N_8546,N_8865);
nor U9230 (N_9230,N_8645,N_8888);
or U9231 (N_9231,N_8776,N_8974);
xor U9232 (N_9232,N_8702,N_8646);
xnor U9233 (N_9233,N_8520,N_8557);
nor U9234 (N_9234,N_8956,N_8907);
or U9235 (N_9235,N_8823,N_8959);
nor U9236 (N_9236,N_8575,N_8824);
nand U9237 (N_9237,N_8659,N_8922);
nor U9238 (N_9238,N_8676,N_8629);
nand U9239 (N_9239,N_8535,N_8787);
and U9240 (N_9240,N_8539,N_8627);
or U9241 (N_9241,N_8519,N_8723);
xor U9242 (N_9242,N_8524,N_8571);
and U9243 (N_9243,N_8674,N_8724);
nand U9244 (N_9244,N_8815,N_8941);
or U9245 (N_9245,N_8633,N_8989);
or U9246 (N_9246,N_8911,N_8957);
nand U9247 (N_9247,N_8954,N_8971);
nand U9248 (N_9248,N_8809,N_8924);
and U9249 (N_9249,N_8516,N_8567);
nor U9250 (N_9250,N_8714,N_8539);
xnor U9251 (N_9251,N_8889,N_8726);
nor U9252 (N_9252,N_8511,N_8741);
nand U9253 (N_9253,N_8975,N_8959);
nand U9254 (N_9254,N_8510,N_8774);
nand U9255 (N_9255,N_8635,N_8905);
and U9256 (N_9256,N_8930,N_8591);
xnor U9257 (N_9257,N_8701,N_8791);
nand U9258 (N_9258,N_8912,N_8931);
xnor U9259 (N_9259,N_8901,N_8644);
xor U9260 (N_9260,N_8669,N_8651);
xnor U9261 (N_9261,N_8531,N_8940);
and U9262 (N_9262,N_8538,N_8570);
or U9263 (N_9263,N_8916,N_8943);
or U9264 (N_9264,N_8780,N_8614);
or U9265 (N_9265,N_8614,N_8817);
nand U9266 (N_9266,N_8978,N_8692);
and U9267 (N_9267,N_8874,N_8533);
or U9268 (N_9268,N_8936,N_8733);
xor U9269 (N_9269,N_8718,N_8907);
nand U9270 (N_9270,N_8579,N_8938);
or U9271 (N_9271,N_8873,N_8681);
xor U9272 (N_9272,N_8599,N_8662);
nand U9273 (N_9273,N_8851,N_8603);
or U9274 (N_9274,N_8710,N_8735);
or U9275 (N_9275,N_8981,N_8747);
nor U9276 (N_9276,N_8627,N_8978);
nand U9277 (N_9277,N_8787,N_8640);
nor U9278 (N_9278,N_8980,N_8648);
nand U9279 (N_9279,N_8596,N_8712);
and U9280 (N_9280,N_8512,N_8564);
nand U9281 (N_9281,N_8858,N_8849);
nand U9282 (N_9282,N_8609,N_8866);
nand U9283 (N_9283,N_8644,N_8600);
nor U9284 (N_9284,N_8515,N_8592);
and U9285 (N_9285,N_8990,N_8638);
or U9286 (N_9286,N_8871,N_8998);
nand U9287 (N_9287,N_8603,N_8589);
xor U9288 (N_9288,N_8775,N_8904);
nand U9289 (N_9289,N_8587,N_8521);
nand U9290 (N_9290,N_8692,N_8992);
and U9291 (N_9291,N_8730,N_8842);
or U9292 (N_9292,N_8956,N_8770);
nand U9293 (N_9293,N_8623,N_8893);
and U9294 (N_9294,N_8647,N_8576);
nor U9295 (N_9295,N_8916,N_8763);
nor U9296 (N_9296,N_8980,N_8718);
nor U9297 (N_9297,N_8919,N_8806);
or U9298 (N_9298,N_8751,N_8725);
nor U9299 (N_9299,N_8592,N_8528);
nand U9300 (N_9300,N_8778,N_8851);
xor U9301 (N_9301,N_8734,N_8877);
xor U9302 (N_9302,N_8965,N_8760);
nand U9303 (N_9303,N_8617,N_8788);
xnor U9304 (N_9304,N_8844,N_8704);
or U9305 (N_9305,N_8625,N_8984);
and U9306 (N_9306,N_8527,N_8778);
and U9307 (N_9307,N_8859,N_8516);
nor U9308 (N_9308,N_8886,N_8805);
and U9309 (N_9309,N_8640,N_8945);
or U9310 (N_9310,N_8898,N_8668);
and U9311 (N_9311,N_8650,N_8736);
xnor U9312 (N_9312,N_8823,N_8982);
nor U9313 (N_9313,N_8635,N_8990);
and U9314 (N_9314,N_8990,N_8675);
nand U9315 (N_9315,N_8529,N_8745);
or U9316 (N_9316,N_8630,N_8736);
nor U9317 (N_9317,N_8745,N_8886);
nor U9318 (N_9318,N_8626,N_8765);
nand U9319 (N_9319,N_8781,N_8563);
nand U9320 (N_9320,N_8593,N_8787);
xnor U9321 (N_9321,N_8793,N_8783);
or U9322 (N_9322,N_8907,N_8805);
nor U9323 (N_9323,N_8952,N_8609);
xnor U9324 (N_9324,N_8631,N_8629);
nor U9325 (N_9325,N_8811,N_8850);
nand U9326 (N_9326,N_8923,N_8803);
and U9327 (N_9327,N_8658,N_8757);
and U9328 (N_9328,N_8892,N_8854);
and U9329 (N_9329,N_8890,N_8514);
xnor U9330 (N_9330,N_8987,N_8741);
and U9331 (N_9331,N_8655,N_8540);
and U9332 (N_9332,N_8787,N_8745);
xnor U9333 (N_9333,N_8655,N_8501);
nand U9334 (N_9334,N_8896,N_8957);
or U9335 (N_9335,N_8953,N_8770);
nor U9336 (N_9336,N_8620,N_8673);
or U9337 (N_9337,N_8734,N_8567);
nand U9338 (N_9338,N_8697,N_8790);
or U9339 (N_9339,N_8728,N_8881);
nor U9340 (N_9340,N_8795,N_8812);
nand U9341 (N_9341,N_8997,N_8996);
nor U9342 (N_9342,N_8565,N_8582);
nor U9343 (N_9343,N_8799,N_8699);
and U9344 (N_9344,N_8975,N_8788);
xor U9345 (N_9345,N_8976,N_8847);
and U9346 (N_9346,N_8975,N_8726);
nor U9347 (N_9347,N_8698,N_8576);
nand U9348 (N_9348,N_8781,N_8952);
or U9349 (N_9349,N_8862,N_8514);
and U9350 (N_9350,N_8706,N_8689);
and U9351 (N_9351,N_8557,N_8652);
and U9352 (N_9352,N_8875,N_8663);
nand U9353 (N_9353,N_8930,N_8943);
nand U9354 (N_9354,N_8589,N_8742);
or U9355 (N_9355,N_8688,N_8676);
nor U9356 (N_9356,N_8571,N_8888);
nor U9357 (N_9357,N_8506,N_8835);
and U9358 (N_9358,N_8902,N_8883);
and U9359 (N_9359,N_8770,N_8797);
xor U9360 (N_9360,N_8833,N_8689);
xor U9361 (N_9361,N_8706,N_8835);
and U9362 (N_9362,N_8854,N_8613);
nor U9363 (N_9363,N_8728,N_8694);
xor U9364 (N_9364,N_8548,N_8719);
or U9365 (N_9365,N_8995,N_8818);
and U9366 (N_9366,N_8761,N_8996);
xnor U9367 (N_9367,N_8620,N_8505);
nand U9368 (N_9368,N_8712,N_8874);
and U9369 (N_9369,N_8990,N_8837);
nand U9370 (N_9370,N_8838,N_8615);
or U9371 (N_9371,N_8919,N_8784);
xnor U9372 (N_9372,N_8519,N_8838);
or U9373 (N_9373,N_8712,N_8954);
nor U9374 (N_9374,N_8796,N_8966);
and U9375 (N_9375,N_8536,N_8549);
nand U9376 (N_9376,N_8839,N_8671);
nand U9377 (N_9377,N_8515,N_8826);
nand U9378 (N_9378,N_8522,N_8671);
or U9379 (N_9379,N_8615,N_8825);
nor U9380 (N_9380,N_8620,N_8744);
nor U9381 (N_9381,N_8723,N_8604);
or U9382 (N_9382,N_8634,N_8566);
or U9383 (N_9383,N_8672,N_8503);
or U9384 (N_9384,N_8847,N_8784);
xor U9385 (N_9385,N_8609,N_8555);
nor U9386 (N_9386,N_8849,N_8778);
xnor U9387 (N_9387,N_8904,N_8999);
or U9388 (N_9388,N_8900,N_8996);
or U9389 (N_9389,N_8854,N_8858);
or U9390 (N_9390,N_8563,N_8561);
nor U9391 (N_9391,N_8700,N_8755);
xor U9392 (N_9392,N_8713,N_8975);
and U9393 (N_9393,N_8508,N_8565);
or U9394 (N_9394,N_8956,N_8889);
nor U9395 (N_9395,N_8609,N_8637);
xor U9396 (N_9396,N_8584,N_8776);
nor U9397 (N_9397,N_8767,N_8506);
nor U9398 (N_9398,N_8579,N_8655);
nor U9399 (N_9399,N_8881,N_8564);
xnor U9400 (N_9400,N_8927,N_8955);
xnor U9401 (N_9401,N_8587,N_8909);
nor U9402 (N_9402,N_8623,N_8874);
xor U9403 (N_9403,N_8768,N_8780);
nor U9404 (N_9404,N_8933,N_8603);
xnor U9405 (N_9405,N_8519,N_8966);
and U9406 (N_9406,N_8670,N_8765);
and U9407 (N_9407,N_8609,N_8913);
and U9408 (N_9408,N_8599,N_8858);
nor U9409 (N_9409,N_8925,N_8935);
nand U9410 (N_9410,N_8566,N_8625);
or U9411 (N_9411,N_8632,N_8686);
xor U9412 (N_9412,N_8612,N_8538);
or U9413 (N_9413,N_8798,N_8823);
and U9414 (N_9414,N_8711,N_8681);
nor U9415 (N_9415,N_8901,N_8671);
nor U9416 (N_9416,N_8615,N_8827);
nor U9417 (N_9417,N_8697,N_8868);
xor U9418 (N_9418,N_8979,N_8657);
nand U9419 (N_9419,N_8911,N_8734);
nand U9420 (N_9420,N_8977,N_8595);
nor U9421 (N_9421,N_8657,N_8745);
nand U9422 (N_9422,N_8773,N_8683);
nand U9423 (N_9423,N_8524,N_8691);
and U9424 (N_9424,N_8993,N_8733);
or U9425 (N_9425,N_8900,N_8532);
nand U9426 (N_9426,N_8711,N_8700);
nor U9427 (N_9427,N_8800,N_8675);
or U9428 (N_9428,N_8880,N_8784);
nand U9429 (N_9429,N_8704,N_8808);
or U9430 (N_9430,N_8587,N_8550);
and U9431 (N_9431,N_8911,N_8660);
nand U9432 (N_9432,N_8686,N_8522);
nor U9433 (N_9433,N_8598,N_8957);
nor U9434 (N_9434,N_8582,N_8596);
xnor U9435 (N_9435,N_8992,N_8676);
or U9436 (N_9436,N_8558,N_8965);
nor U9437 (N_9437,N_8598,N_8783);
nor U9438 (N_9438,N_8638,N_8908);
and U9439 (N_9439,N_8950,N_8587);
or U9440 (N_9440,N_8716,N_8735);
nor U9441 (N_9441,N_8695,N_8591);
nand U9442 (N_9442,N_8630,N_8986);
and U9443 (N_9443,N_8669,N_8782);
xnor U9444 (N_9444,N_8666,N_8651);
or U9445 (N_9445,N_8623,N_8581);
or U9446 (N_9446,N_8882,N_8775);
or U9447 (N_9447,N_8723,N_8731);
and U9448 (N_9448,N_8983,N_8790);
nand U9449 (N_9449,N_8513,N_8774);
nor U9450 (N_9450,N_8869,N_8997);
and U9451 (N_9451,N_8560,N_8777);
nor U9452 (N_9452,N_8849,N_8703);
nand U9453 (N_9453,N_8517,N_8670);
and U9454 (N_9454,N_8863,N_8678);
nand U9455 (N_9455,N_8754,N_8569);
nor U9456 (N_9456,N_8905,N_8739);
xnor U9457 (N_9457,N_8877,N_8975);
xor U9458 (N_9458,N_8763,N_8680);
nor U9459 (N_9459,N_8881,N_8703);
nand U9460 (N_9460,N_8920,N_8867);
or U9461 (N_9461,N_8784,N_8855);
nand U9462 (N_9462,N_8989,N_8870);
nor U9463 (N_9463,N_8566,N_8860);
or U9464 (N_9464,N_8872,N_8542);
or U9465 (N_9465,N_8787,N_8791);
or U9466 (N_9466,N_8793,N_8546);
nor U9467 (N_9467,N_8998,N_8985);
and U9468 (N_9468,N_8739,N_8625);
nand U9469 (N_9469,N_8999,N_8669);
or U9470 (N_9470,N_8932,N_8684);
xor U9471 (N_9471,N_8696,N_8942);
or U9472 (N_9472,N_8915,N_8640);
nand U9473 (N_9473,N_8776,N_8932);
nor U9474 (N_9474,N_8974,N_8658);
xnor U9475 (N_9475,N_8573,N_8951);
xor U9476 (N_9476,N_8958,N_8918);
or U9477 (N_9477,N_8725,N_8656);
nand U9478 (N_9478,N_8558,N_8980);
nand U9479 (N_9479,N_8691,N_8853);
or U9480 (N_9480,N_8629,N_8906);
and U9481 (N_9481,N_8503,N_8581);
and U9482 (N_9482,N_8665,N_8798);
xnor U9483 (N_9483,N_8754,N_8732);
xnor U9484 (N_9484,N_8795,N_8858);
xor U9485 (N_9485,N_8681,N_8961);
and U9486 (N_9486,N_8852,N_8995);
and U9487 (N_9487,N_8523,N_8693);
nand U9488 (N_9488,N_8762,N_8922);
or U9489 (N_9489,N_8867,N_8824);
nand U9490 (N_9490,N_8844,N_8527);
xor U9491 (N_9491,N_8694,N_8595);
or U9492 (N_9492,N_8511,N_8959);
xnor U9493 (N_9493,N_8517,N_8530);
xor U9494 (N_9494,N_8900,N_8788);
nand U9495 (N_9495,N_8915,N_8703);
or U9496 (N_9496,N_8838,N_8521);
xnor U9497 (N_9497,N_8990,N_8845);
xor U9498 (N_9498,N_8708,N_8548);
xnor U9499 (N_9499,N_8963,N_8712);
xor U9500 (N_9500,N_9132,N_9163);
xor U9501 (N_9501,N_9431,N_9112);
and U9502 (N_9502,N_9092,N_9340);
or U9503 (N_9503,N_9426,N_9359);
nand U9504 (N_9504,N_9331,N_9411);
xor U9505 (N_9505,N_9399,N_9377);
and U9506 (N_9506,N_9020,N_9376);
xor U9507 (N_9507,N_9014,N_9486);
and U9508 (N_9508,N_9094,N_9382);
and U9509 (N_9509,N_9462,N_9019);
and U9510 (N_9510,N_9236,N_9117);
xnor U9511 (N_9511,N_9494,N_9338);
xor U9512 (N_9512,N_9362,N_9196);
nand U9513 (N_9513,N_9490,N_9296);
xnor U9514 (N_9514,N_9123,N_9394);
nor U9515 (N_9515,N_9071,N_9146);
or U9516 (N_9516,N_9316,N_9120);
and U9517 (N_9517,N_9397,N_9499);
and U9518 (N_9518,N_9349,N_9450);
nor U9519 (N_9519,N_9385,N_9217);
nand U9520 (N_9520,N_9157,N_9484);
or U9521 (N_9521,N_9429,N_9233);
xor U9522 (N_9522,N_9179,N_9198);
nor U9523 (N_9523,N_9269,N_9048);
or U9524 (N_9524,N_9015,N_9281);
nand U9525 (N_9525,N_9025,N_9416);
nor U9526 (N_9526,N_9354,N_9300);
xnor U9527 (N_9527,N_9045,N_9479);
or U9528 (N_9528,N_9036,N_9312);
nand U9529 (N_9529,N_9148,N_9278);
and U9530 (N_9530,N_9439,N_9118);
or U9531 (N_9531,N_9289,N_9465);
and U9532 (N_9532,N_9031,N_9044);
nand U9533 (N_9533,N_9337,N_9032);
nor U9534 (N_9534,N_9352,N_9070);
nor U9535 (N_9535,N_9063,N_9068);
or U9536 (N_9536,N_9309,N_9151);
or U9537 (N_9537,N_9261,N_9154);
xnor U9538 (N_9538,N_9201,N_9024);
or U9539 (N_9539,N_9401,N_9268);
or U9540 (N_9540,N_9298,N_9249);
or U9541 (N_9541,N_9164,N_9466);
xnor U9542 (N_9542,N_9073,N_9083);
nor U9543 (N_9543,N_9041,N_9229);
xor U9544 (N_9544,N_9413,N_9442);
xnor U9545 (N_9545,N_9027,N_9095);
xnor U9546 (N_9546,N_9271,N_9226);
nor U9547 (N_9547,N_9344,N_9001);
nor U9548 (N_9548,N_9364,N_9257);
xor U9549 (N_9549,N_9402,N_9414);
xnor U9550 (N_9550,N_9434,N_9131);
nor U9551 (N_9551,N_9320,N_9000);
nand U9552 (N_9552,N_9188,N_9369);
xnor U9553 (N_9553,N_9483,N_9141);
nor U9554 (N_9554,N_9457,N_9476);
and U9555 (N_9555,N_9144,N_9389);
or U9556 (N_9556,N_9202,N_9080);
nor U9557 (N_9557,N_9234,N_9177);
nand U9558 (N_9558,N_9206,N_9053);
or U9559 (N_9559,N_9308,N_9358);
xor U9560 (N_9560,N_9203,N_9323);
and U9561 (N_9561,N_9314,N_9055);
nor U9562 (N_9562,N_9356,N_9400);
and U9563 (N_9563,N_9345,N_9247);
nand U9564 (N_9564,N_9475,N_9241);
nand U9565 (N_9565,N_9446,N_9158);
or U9566 (N_9566,N_9299,N_9138);
nor U9567 (N_9567,N_9142,N_9496);
nand U9568 (N_9568,N_9473,N_9087);
xor U9569 (N_9569,N_9108,N_9210);
or U9570 (N_9570,N_9265,N_9365);
nor U9571 (N_9571,N_9432,N_9113);
and U9572 (N_9572,N_9424,N_9435);
and U9573 (N_9573,N_9197,N_9322);
nand U9574 (N_9574,N_9443,N_9495);
or U9575 (N_9575,N_9363,N_9464);
and U9576 (N_9576,N_9445,N_9018);
or U9577 (N_9577,N_9379,N_9405);
xor U9578 (N_9578,N_9448,N_9291);
nor U9579 (N_9579,N_9449,N_9168);
nand U9580 (N_9580,N_9319,N_9033);
nor U9581 (N_9581,N_9213,N_9129);
and U9582 (N_9582,N_9122,N_9391);
nand U9583 (N_9583,N_9304,N_9311);
nor U9584 (N_9584,N_9343,N_9245);
or U9585 (N_9585,N_9485,N_9351);
nor U9586 (N_9586,N_9286,N_9487);
nand U9587 (N_9587,N_9103,N_9250);
nand U9588 (N_9588,N_9488,N_9075);
xor U9589 (N_9589,N_9016,N_9292);
and U9590 (N_9590,N_9355,N_9270);
nor U9591 (N_9591,N_9180,N_9136);
or U9592 (N_9592,N_9366,N_9101);
nand U9593 (N_9593,N_9433,N_9470);
xor U9594 (N_9594,N_9253,N_9403);
xnor U9595 (N_9595,N_9115,N_9461);
nand U9596 (N_9596,N_9452,N_9127);
xor U9597 (N_9597,N_9339,N_9190);
nand U9598 (N_9598,N_9360,N_9105);
or U9599 (N_9599,N_9267,N_9310);
and U9600 (N_9600,N_9116,N_9329);
and U9601 (N_9601,N_9460,N_9248);
nor U9602 (N_9602,N_9463,N_9378);
nand U9603 (N_9603,N_9037,N_9240);
and U9604 (N_9604,N_9350,N_9189);
xnor U9605 (N_9605,N_9128,N_9121);
nor U9606 (N_9606,N_9474,N_9317);
nor U9607 (N_9607,N_9017,N_9006);
xnor U9608 (N_9608,N_9491,N_9126);
xnor U9609 (N_9609,N_9227,N_9022);
xnor U9610 (N_9610,N_9221,N_9009);
xnor U9611 (N_9611,N_9147,N_9178);
or U9612 (N_9612,N_9357,N_9183);
nand U9613 (N_9613,N_9028,N_9187);
nor U9614 (N_9614,N_9035,N_9417);
or U9615 (N_9615,N_9273,N_9302);
xor U9616 (N_9616,N_9393,N_9155);
xnor U9617 (N_9617,N_9353,N_9341);
or U9618 (N_9618,N_9199,N_9419);
nor U9619 (N_9619,N_9029,N_9346);
nor U9620 (N_9620,N_9230,N_9471);
or U9621 (N_9621,N_9256,N_9325);
nand U9622 (N_9622,N_9161,N_9301);
nor U9623 (N_9623,N_9328,N_9214);
nand U9624 (N_9624,N_9079,N_9266);
nand U9625 (N_9625,N_9372,N_9060);
xor U9626 (N_9626,N_9477,N_9192);
and U9627 (N_9627,N_9374,N_9407);
xor U9628 (N_9628,N_9420,N_9380);
nand U9629 (N_9629,N_9447,N_9093);
or U9630 (N_9630,N_9481,N_9396);
nand U9631 (N_9631,N_9072,N_9049);
or U9632 (N_9632,N_9056,N_9412);
nand U9633 (N_9633,N_9171,N_9246);
xor U9634 (N_9634,N_9336,N_9386);
and U9635 (N_9635,N_9225,N_9150);
or U9636 (N_9636,N_9427,N_9091);
nand U9637 (N_9637,N_9318,N_9347);
nand U9638 (N_9638,N_9294,N_9110);
and U9639 (N_9639,N_9493,N_9334);
or U9640 (N_9640,N_9276,N_9454);
and U9641 (N_9641,N_9004,N_9425);
and U9642 (N_9642,N_9408,N_9170);
or U9643 (N_9643,N_9050,N_9260);
and U9644 (N_9644,N_9280,N_9455);
or U9645 (N_9645,N_9390,N_9472);
nand U9646 (N_9646,N_9173,N_9238);
or U9647 (N_9647,N_9172,N_9251);
or U9648 (N_9648,N_9066,N_9102);
xor U9649 (N_9649,N_9235,N_9287);
nand U9650 (N_9650,N_9130,N_9263);
and U9651 (N_9651,N_9096,N_9283);
xor U9652 (N_9652,N_9264,N_9114);
xnor U9653 (N_9653,N_9143,N_9159);
nand U9654 (N_9654,N_9458,N_9051);
xnor U9655 (N_9655,N_9216,N_9133);
nand U9656 (N_9656,N_9451,N_9232);
nor U9657 (N_9657,N_9330,N_9002);
nor U9658 (N_9658,N_9104,N_9005);
nor U9659 (N_9659,N_9277,N_9367);
or U9660 (N_9660,N_9089,N_9212);
or U9661 (N_9661,N_9058,N_9193);
nand U9662 (N_9662,N_9444,N_9368);
and U9663 (N_9663,N_9139,N_9167);
nor U9664 (N_9664,N_9497,N_9086);
nand U9665 (N_9665,N_9284,N_9211);
nor U9666 (N_9666,N_9428,N_9406);
xor U9667 (N_9667,N_9224,N_9181);
and U9668 (N_9668,N_9067,N_9034);
xnor U9669 (N_9669,N_9410,N_9040);
xor U9670 (N_9670,N_9026,N_9162);
or U9671 (N_9671,N_9272,N_9194);
nor U9672 (N_9672,N_9332,N_9057);
or U9673 (N_9673,N_9418,N_9046);
nand U9674 (N_9674,N_9489,N_9438);
or U9675 (N_9675,N_9423,N_9109);
and U9676 (N_9676,N_9415,N_9293);
and U9677 (N_9677,N_9371,N_9469);
nand U9678 (N_9678,N_9315,N_9169);
and U9679 (N_9679,N_9084,N_9321);
xnor U9680 (N_9680,N_9052,N_9011);
and U9681 (N_9681,N_9174,N_9007);
xnor U9682 (N_9682,N_9384,N_9137);
xor U9683 (N_9683,N_9111,N_9059);
nor U9684 (N_9684,N_9498,N_9492);
xnor U9685 (N_9685,N_9279,N_9327);
or U9686 (N_9686,N_9003,N_9303);
or U9687 (N_9687,N_9135,N_9153);
or U9688 (N_9688,N_9456,N_9107);
or U9689 (N_9689,N_9274,N_9218);
xor U9690 (N_9690,N_9326,N_9076);
or U9691 (N_9691,N_9307,N_9088);
and U9692 (N_9692,N_9078,N_9065);
xor U9693 (N_9693,N_9152,N_9195);
xor U9694 (N_9694,N_9054,N_9219);
nor U9695 (N_9695,N_9098,N_9042);
or U9696 (N_9696,N_9013,N_9043);
xor U9697 (N_9697,N_9134,N_9228);
xor U9698 (N_9698,N_9395,N_9008);
nand U9699 (N_9699,N_9124,N_9480);
or U9700 (N_9700,N_9453,N_9254);
or U9701 (N_9701,N_9288,N_9237);
and U9702 (N_9702,N_9215,N_9231);
or U9703 (N_9703,N_9239,N_9436);
or U9704 (N_9704,N_9335,N_9061);
xnor U9705 (N_9705,N_9165,N_9306);
or U9706 (N_9706,N_9404,N_9074);
xor U9707 (N_9707,N_9010,N_9200);
or U9708 (N_9708,N_9145,N_9333);
or U9709 (N_9709,N_9208,N_9220);
and U9710 (N_9710,N_9459,N_9097);
nor U9711 (N_9711,N_9243,N_9186);
or U9712 (N_9712,N_9119,N_9275);
xnor U9713 (N_9713,N_9090,N_9182);
nand U9714 (N_9714,N_9100,N_9285);
and U9715 (N_9715,N_9478,N_9392);
or U9716 (N_9716,N_9383,N_9038);
or U9717 (N_9717,N_9175,N_9324);
xor U9718 (N_9718,N_9258,N_9437);
nor U9719 (N_9719,N_9209,N_9062);
nor U9720 (N_9720,N_9184,N_9106);
or U9721 (N_9721,N_9223,N_9422);
nor U9722 (N_9722,N_9023,N_9149);
or U9723 (N_9723,N_9255,N_9030);
nand U9724 (N_9724,N_9468,N_9125);
nor U9725 (N_9725,N_9305,N_9099);
or U9726 (N_9726,N_9409,N_9262);
and U9727 (N_9727,N_9012,N_9205);
nor U9728 (N_9728,N_9166,N_9361);
nand U9729 (N_9729,N_9160,N_9176);
nand U9730 (N_9730,N_9482,N_9242);
or U9731 (N_9731,N_9039,N_9373);
nand U9732 (N_9732,N_9297,N_9047);
or U9733 (N_9733,N_9021,N_9207);
nor U9734 (N_9734,N_9191,N_9064);
and U9735 (N_9735,N_9441,N_9140);
nand U9736 (N_9736,N_9156,N_9421);
or U9737 (N_9737,N_9381,N_9348);
nand U9738 (N_9738,N_9244,N_9222);
xnor U9739 (N_9739,N_9085,N_9204);
or U9740 (N_9740,N_9375,N_9077);
and U9741 (N_9741,N_9398,N_9387);
or U9742 (N_9742,N_9082,N_9467);
nand U9743 (N_9743,N_9342,N_9430);
xor U9744 (N_9744,N_9282,N_9388);
nand U9745 (N_9745,N_9252,N_9259);
xnor U9746 (N_9746,N_9440,N_9081);
xor U9747 (N_9747,N_9295,N_9290);
or U9748 (N_9748,N_9069,N_9185);
nor U9749 (N_9749,N_9313,N_9370);
nand U9750 (N_9750,N_9064,N_9431);
xor U9751 (N_9751,N_9222,N_9358);
and U9752 (N_9752,N_9284,N_9107);
nor U9753 (N_9753,N_9274,N_9040);
nand U9754 (N_9754,N_9164,N_9232);
nor U9755 (N_9755,N_9434,N_9336);
nand U9756 (N_9756,N_9334,N_9346);
nand U9757 (N_9757,N_9454,N_9128);
nand U9758 (N_9758,N_9261,N_9235);
and U9759 (N_9759,N_9442,N_9158);
xor U9760 (N_9760,N_9117,N_9441);
or U9761 (N_9761,N_9326,N_9459);
nor U9762 (N_9762,N_9170,N_9072);
nor U9763 (N_9763,N_9180,N_9471);
xnor U9764 (N_9764,N_9174,N_9002);
and U9765 (N_9765,N_9407,N_9181);
nand U9766 (N_9766,N_9015,N_9471);
nor U9767 (N_9767,N_9478,N_9257);
nand U9768 (N_9768,N_9402,N_9178);
and U9769 (N_9769,N_9088,N_9093);
and U9770 (N_9770,N_9355,N_9266);
nor U9771 (N_9771,N_9386,N_9008);
nand U9772 (N_9772,N_9135,N_9333);
nand U9773 (N_9773,N_9364,N_9087);
and U9774 (N_9774,N_9177,N_9253);
and U9775 (N_9775,N_9046,N_9348);
and U9776 (N_9776,N_9305,N_9358);
and U9777 (N_9777,N_9205,N_9140);
nor U9778 (N_9778,N_9262,N_9303);
and U9779 (N_9779,N_9094,N_9248);
or U9780 (N_9780,N_9459,N_9194);
or U9781 (N_9781,N_9481,N_9450);
and U9782 (N_9782,N_9167,N_9160);
nand U9783 (N_9783,N_9284,N_9396);
or U9784 (N_9784,N_9405,N_9155);
xnor U9785 (N_9785,N_9401,N_9340);
and U9786 (N_9786,N_9344,N_9006);
nor U9787 (N_9787,N_9007,N_9357);
nor U9788 (N_9788,N_9428,N_9015);
nand U9789 (N_9789,N_9217,N_9076);
nor U9790 (N_9790,N_9332,N_9327);
and U9791 (N_9791,N_9416,N_9234);
and U9792 (N_9792,N_9328,N_9277);
nor U9793 (N_9793,N_9010,N_9017);
or U9794 (N_9794,N_9447,N_9133);
xor U9795 (N_9795,N_9062,N_9248);
nand U9796 (N_9796,N_9031,N_9147);
or U9797 (N_9797,N_9410,N_9416);
and U9798 (N_9798,N_9435,N_9191);
nand U9799 (N_9799,N_9138,N_9033);
or U9800 (N_9800,N_9415,N_9140);
nor U9801 (N_9801,N_9338,N_9136);
nand U9802 (N_9802,N_9425,N_9009);
xnor U9803 (N_9803,N_9115,N_9064);
or U9804 (N_9804,N_9104,N_9484);
or U9805 (N_9805,N_9270,N_9328);
xnor U9806 (N_9806,N_9298,N_9239);
nand U9807 (N_9807,N_9315,N_9106);
nor U9808 (N_9808,N_9362,N_9162);
nor U9809 (N_9809,N_9382,N_9368);
xor U9810 (N_9810,N_9080,N_9491);
and U9811 (N_9811,N_9412,N_9062);
or U9812 (N_9812,N_9136,N_9044);
nor U9813 (N_9813,N_9407,N_9247);
xor U9814 (N_9814,N_9046,N_9298);
xnor U9815 (N_9815,N_9271,N_9343);
or U9816 (N_9816,N_9060,N_9006);
and U9817 (N_9817,N_9485,N_9210);
and U9818 (N_9818,N_9158,N_9034);
xnor U9819 (N_9819,N_9027,N_9061);
nand U9820 (N_9820,N_9372,N_9024);
or U9821 (N_9821,N_9218,N_9436);
or U9822 (N_9822,N_9230,N_9042);
nor U9823 (N_9823,N_9026,N_9492);
and U9824 (N_9824,N_9168,N_9273);
and U9825 (N_9825,N_9260,N_9483);
and U9826 (N_9826,N_9255,N_9435);
nand U9827 (N_9827,N_9448,N_9151);
and U9828 (N_9828,N_9459,N_9427);
xnor U9829 (N_9829,N_9424,N_9491);
nand U9830 (N_9830,N_9013,N_9268);
or U9831 (N_9831,N_9440,N_9251);
and U9832 (N_9832,N_9358,N_9389);
or U9833 (N_9833,N_9138,N_9335);
or U9834 (N_9834,N_9322,N_9132);
xor U9835 (N_9835,N_9055,N_9381);
xor U9836 (N_9836,N_9059,N_9004);
nor U9837 (N_9837,N_9355,N_9250);
or U9838 (N_9838,N_9403,N_9150);
and U9839 (N_9839,N_9476,N_9168);
and U9840 (N_9840,N_9473,N_9165);
nor U9841 (N_9841,N_9240,N_9178);
nor U9842 (N_9842,N_9082,N_9088);
nand U9843 (N_9843,N_9414,N_9175);
xnor U9844 (N_9844,N_9048,N_9162);
and U9845 (N_9845,N_9078,N_9211);
nor U9846 (N_9846,N_9360,N_9410);
xor U9847 (N_9847,N_9497,N_9251);
nor U9848 (N_9848,N_9445,N_9343);
nand U9849 (N_9849,N_9188,N_9235);
and U9850 (N_9850,N_9495,N_9416);
nor U9851 (N_9851,N_9400,N_9172);
nand U9852 (N_9852,N_9461,N_9209);
nand U9853 (N_9853,N_9089,N_9081);
nand U9854 (N_9854,N_9212,N_9004);
nand U9855 (N_9855,N_9267,N_9422);
and U9856 (N_9856,N_9473,N_9325);
and U9857 (N_9857,N_9468,N_9067);
nor U9858 (N_9858,N_9185,N_9253);
and U9859 (N_9859,N_9315,N_9293);
nor U9860 (N_9860,N_9160,N_9131);
and U9861 (N_9861,N_9247,N_9194);
nand U9862 (N_9862,N_9190,N_9257);
xor U9863 (N_9863,N_9143,N_9103);
or U9864 (N_9864,N_9223,N_9275);
nand U9865 (N_9865,N_9280,N_9197);
nand U9866 (N_9866,N_9386,N_9043);
nand U9867 (N_9867,N_9255,N_9323);
or U9868 (N_9868,N_9092,N_9044);
and U9869 (N_9869,N_9193,N_9097);
and U9870 (N_9870,N_9294,N_9192);
nor U9871 (N_9871,N_9386,N_9213);
nor U9872 (N_9872,N_9294,N_9410);
or U9873 (N_9873,N_9275,N_9045);
and U9874 (N_9874,N_9384,N_9124);
or U9875 (N_9875,N_9244,N_9446);
or U9876 (N_9876,N_9150,N_9114);
or U9877 (N_9877,N_9170,N_9079);
xnor U9878 (N_9878,N_9042,N_9282);
xnor U9879 (N_9879,N_9217,N_9153);
nand U9880 (N_9880,N_9432,N_9255);
and U9881 (N_9881,N_9351,N_9006);
and U9882 (N_9882,N_9000,N_9134);
nand U9883 (N_9883,N_9113,N_9339);
nand U9884 (N_9884,N_9009,N_9155);
nand U9885 (N_9885,N_9400,N_9348);
and U9886 (N_9886,N_9499,N_9450);
nor U9887 (N_9887,N_9270,N_9442);
nand U9888 (N_9888,N_9025,N_9468);
nor U9889 (N_9889,N_9309,N_9094);
or U9890 (N_9890,N_9080,N_9085);
or U9891 (N_9891,N_9011,N_9077);
and U9892 (N_9892,N_9123,N_9431);
nor U9893 (N_9893,N_9462,N_9191);
nand U9894 (N_9894,N_9382,N_9274);
xor U9895 (N_9895,N_9417,N_9145);
xnor U9896 (N_9896,N_9443,N_9145);
and U9897 (N_9897,N_9196,N_9215);
or U9898 (N_9898,N_9280,N_9160);
and U9899 (N_9899,N_9110,N_9045);
and U9900 (N_9900,N_9403,N_9297);
nor U9901 (N_9901,N_9057,N_9231);
or U9902 (N_9902,N_9137,N_9340);
nand U9903 (N_9903,N_9082,N_9418);
nand U9904 (N_9904,N_9278,N_9084);
nand U9905 (N_9905,N_9377,N_9313);
and U9906 (N_9906,N_9363,N_9074);
or U9907 (N_9907,N_9148,N_9399);
xor U9908 (N_9908,N_9416,N_9365);
or U9909 (N_9909,N_9451,N_9497);
xnor U9910 (N_9910,N_9339,N_9033);
xor U9911 (N_9911,N_9267,N_9480);
xor U9912 (N_9912,N_9004,N_9342);
and U9913 (N_9913,N_9120,N_9382);
nand U9914 (N_9914,N_9266,N_9444);
and U9915 (N_9915,N_9487,N_9146);
and U9916 (N_9916,N_9106,N_9444);
nor U9917 (N_9917,N_9494,N_9132);
xnor U9918 (N_9918,N_9124,N_9125);
nor U9919 (N_9919,N_9043,N_9319);
xor U9920 (N_9920,N_9437,N_9431);
nor U9921 (N_9921,N_9146,N_9112);
nand U9922 (N_9922,N_9475,N_9272);
nor U9923 (N_9923,N_9239,N_9265);
or U9924 (N_9924,N_9178,N_9059);
nand U9925 (N_9925,N_9001,N_9249);
or U9926 (N_9926,N_9254,N_9304);
nor U9927 (N_9927,N_9049,N_9444);
and U9928 (N_9928,N_9178,N_9310);
xnor U9929 (N_9929,N_9102,N_9294);
xor U9930 (N_9930,N_9463,N_9171);
nor U9931 (N_9931,N_9211,N_9278);
nand U9932 (N_9932,N_9224,N_9345);
xnor U9933 (N_9933,N_9398,N_9079);
xor U9934 (N_9934,N_9307,N_9380);
and U9935 (N_9935,N_9164,N_9435);
or U9936 (N_9936,N_9007,N_9420);
or U9937 (N_9937,N_9150,N_9365);
xor U9938 (N_9938,N_9393,N_9269);
or U9939 (N_9939,N_9073,N_9462);
xnor U9940 (N_9940,N_9032,N_9295);
nand U9941 (N_9941,N_9390,N_9138);
xnor U9942 (N_9942,N_9278,N_9029);
nor U9943 (N_9943,N_9033,N_9129);
xor U9944 (N_9944,N_9231,N_9039);
or U9945 (N_9945,N_9097,N_9370);
nor U9946 (N_9946,N_9294,N_9323);
or U9947 (N_9947,N_9297,N_9387);
xnor U9948 (N_9948,N_9180,N_9262);
xnor U9949 (N_9949,N_9288,N_9488);
nor U9950 (N_9950,N_9223,N_9064);
or U9951 (N_9951,N_9357,N_9271);
nand U9952 (N_9952,N_9111,N_9264);
nor U9953 (N_9953,N_9305,N_9335);
xnor U9954 (N_9954,N_9494,N_9304);
nand U9955 (N_9955,N_9248,N_9334);
and U9956 (N_9956,N_9404,N_9131);
nor U9957 (N_9957,N_9116,N_9187);
nand U9958 (N_9958,N_9450,N_9030);
nor U9959 (N_9959,N_9140,N_9204);
or U9960 (N_9960,N_9015,N_9084);
nand U9961 (N_9961,N_9395,N_9429);
nor U9962 (N_9962,N_9063,N_9186);
or U9963 (N_9963,N_9102,N_9126);
or U9964 (N_9964,N_9382,N_9044);
and U9965 (N_9965,N_9213,N_9269);
xnor U9966 (N_9966,N_9320,N_9016);
xnor U9967 (N_9967,N_9084,N_9257);
and U9968 (N_9968,N_9150,N_9066);
and U9969 (N_9969,N_9217,N_9161);
or U9970 (N_9970,N_9294,N_9107);
or U9971 (N_9971,N_9257,N_9208);
and U9972 (N_9972,N_9281,N_9265);
and U9973 (N_9973,N_9202,N_9151);
and U9974 (N_9974,N_9236,N_9470);
or U9975 (N_9975,N_9176,N_9235);
nand U9976 (N_9976,N_9030,N_9045);
nor U9977 (N_9977,N_9465,N_9340);
nand U9978 (N_9978,N_9270,N_9218);
and U9979 (N_9979,N_9052,N_9215);
nand U9980 (N_9980,N_9025,N_9268);
and U9981 (N_9981,N_9064,N_9287);
nand U9982 (N_9982,N_9180,N_9474);
nor U9983 (N_9983,N_9466,N_9014);
nand U9984 (N_9984,N_9278,N_9169);
and U9985 (N_9985,N_9448,N_9382);
or U9986 (N_9986,N_9373,N_9152);
and U9987 (N_9987,N_9009,N_9344);
and U9988 (N_9988,N_9116,N_9444);
nand U9989 (N_9989,N_9345,N_9145);
nand U9990 (N_9990,N_9008,N_9381);
and U9991 (N_9991,N_9484,N_9359);
xnor U9992 (N_9992,N_9056,N_9133);
xor U9993 (N_9993,N_9088,N_9298);
and U9994 (N_9994,N_9094,N_9097);
and U9995 (N_9995,N_9420,N_9157);
nor U9996 (N_9996,N_9120,N_9101);
nor U9997 (N_9997,N_9209,N_9305);
nor U9998 (N_9998,N_9057,N_9045);
or U9999 (N_9999,N_9446,N_9245);
and UO_0 (O_0,N_9822,N_9760);
nand UO_1 (O_1,N_9647,N_9722);
xor UO_2 (O_2,N_9993,N_9530);
nand UO_3 (O_3,N_9969,N_9548);
xor UO_4 (O_4,N_9711,N_9723);
and UO_5 (O_5,N_9585,N_9895);
and UO_6 (O_6,N_9902,N_9538);
nor UO_7 (O_7,N_9938,N_9770);
and UO_8 (O_8,N_9677,N_9640);
and UO_9 (O_9,N_9662,N_9783);
nand UO_10 (O_10,N_9545,N_9680);
nand UO_11 (O_11,N_9625,N_9910);
nand UO_12 (O_12,N_9686,N_9540);
xnor UO_13 (O_13,N_9911,N_9520);
xnor UO_14 (O_14,N_9663,N_9652);
nor UO_15 (O_15,N_9637,N_9606);
and UO_16 (O_16,N_9959,N_9758);
or UO_17 (O_17,N_9805,N_9963);
nor UO_18 (O_18,N_9617,N_9668);
or UO_19 (O_19,N_9628,N_9961);
or UO_20 (O_20,N_9999,N_9856);
nand UO_21 (O_21,N_9750,N_9932);
nand UO_22 (O_22,N_9656,N_9528);
nand UO_23 (O_23,N_9554,N_9735);
nor UO_24 (O_24,N_9622,N_9743);
or UO_25 (O_25,N_9714,N_9840);
xnor UO_26 (O_26,N_9900,N_9982);
or UO_27 (O_27,N_9874,N_9777);
or UO_28 (O_28,N_9854,N_9966);
nand UO_29 (O_29,N_9605,N_9789);
or UO_30 (O_30,N_9919,N_9522);
nor UO_31 (O_31,N_9697,N_9563);
xnor UO_32 (O_32,N_9987,N_9672);
and UO_33 (O_33,N_9573,N_9521);
xnor UO_34 (O_34,N_9817,N_9692);
nor UO_35 (O_35,N_9514,N_9810);
and UO_36 (O_36,N_9803,N_9772);
nand UO_37 (O_37,N_9517,N_9892);
xnor UO_38 (O_38,N_9526,N_9825);
nor UO_39 (O_39,N_9983,N_9655);
xnor UO_40 (O_40,N_9535,N_9508);
or UO_41 (O_41,N_9844,N_9748);
nor UO_42 (O_42,N_9918,N_9587);
nand UO_43 (O_43,N_9733,N_9609);
and UO_44 (O_44,N_9747,N_9721);
and UO_45 (O_45,N_9509,N_9518);
nand UO_46 (O_46,N_9867,N_9980);
or UO_47 (O_47,N_9669,N_9962);
xor UO_48 (O_48,N_9763,N_9568);
or UO_49 (O_49,N_9594,N_9581);
or UO_50 (O_50,N_9600,N_9820);
nand UO_51 (O_51,N_9674,N_9519);
nand UO_52 (O_52,N_9981,N_9688);
nand UO_53 (O_53,N_9607,N_9591);
or UO_54 (O_54,N_9884,N_9572);
nand UO_55 (O_55,N_9727,N_9561);
xnor UO_56 (O_56,N_9970,N_9537);
or UO_57 (O_57,N_9761,N_9940);
or UO_58 (O_58,N_9984,N_9831);
nor UO_59 (O_59,N_9604,N_9658);
and UO_60 (O_60,N_9951,N_9565);
or UO_61 (O_61,N_9539,N_9724);
xnor UO_62 (O_62,N_9541,N_9815);
nand UO_63 (O_63,N_9944,N_9971);
or UO_64 (O_64,N_9745,N_9795);
nor UO_65 (O_65,N_9929,N_9931);
xor UO_66 (O_66,N_9593,N_9927);
nor UO_67 (O_67,N_9757,N_9713);
nor UO_68 (O_68,N_9569,N_9602);
nand UO_69 (O_69,N_9644,N_9878);
nand UO_70 (O_70,N_9730,N_9752);
nor UO_71 (O_71,N_9690,N_9923);
xnor UO_72 (O_72,N_9975,N_9619);
xor UO_73 (O_73,N_9995,N_9952);
or UO_74 (O_74,N_9731,N_9801);
nand UO_75 (O_75,N_9855,N_9564);
nor UO_76 (O_76,N_9865,N_9876);
and UO_77 (O_77,N_9994,N_9653);
and UO_78 (O_78,N_9556,N_9779);
nand UO_79 (O_79,N_9813,N_9542);
xor UO_80 (O_80,N_9888,N_9659);
or UO_81 (O_81,N_9504,N_9797);
nand UO_82 (O_82,N_9755,N_9916);
nand UO_83 (O_83,N_9873,N_9764);
and UO_84 (O_84,N_9558,N_9703);
xnor UO_85 (O_85,N_9861,N_9943);
nand UO_86 (O_86,N_9776,N_9798);
xnor UO_87 (O_87,N_9645,N_9551);
xnor UO_88 (O_88,N_9712,N_9978);
or UO_89 (O_89,N_9749,N_9853);
xnor UO_90 (O_90,N_9829,N_9579);
nand UO_91 (O_91,N_9899,N_9904);
nand UO_92 (O_92,N_9958,N_9986);
nor UO_93 (O_93,N_9784,N_9802);
nand UO_94 (O_94,N_9661,N_9863);
nand UO_95 (O_95,N_9678,N_9588);
xnor UO_96 (O_96,N_9950,N_9774);
or UO_97 (O_97,N_9555,N_9570);
and UO_98 (O_98,N_9917,N_9821);
and UO_99 (O_99,N_9634,N_9681);
xnor UO_100 (O_100,N_9704,N_9553);
xnor UO_101 (O_101,N_9960,N_9837);
nor UO_102 (O_102,N_9636,N_9737);
or UO_103 (O_103,N_9529,N_9510);
nand UO_104 (O_104,N_9543,N_9567);
nand UO_105 (O_105,N_9756,N_9527);
nor UO_106 (O_106,N_9997,N_9560);
and UO_107 (O_107,N_9500,N_9939);
or UO_108 (O_108,N_9624,N_9501);
or UO_109 (O_109,N_9574,N_9566);
or UO_110 (O_110,N_9794,N_9885);
and UO_111 (O_111,N_9557,N_9869);
xnor UO_112 (O_112,N_9592,N_9699);
nor UO_113 (O_113,N_9954,N_9946);
and UO_114 (O_114,N_9616,N_9985);
xor UO_115 (O_115,N_9872,N_9965);
or UO_116 (O_116,N_9934,N_9691);
nand UO_117 (O_117,N_9546,N_9875);
nand UO_118 (O_118,N_9597,N_9702);
nand UO_119 (O_119,N_9897,N_9889);
xor UO_120 (O_120,N_9671,N_9838);
nor UO_121 (O_121,N_9552,N_9968);
and UO_122 (O_122,N_9576,N_9785);
or UO_123 (O_123,N_9870,N_9908);
and UO_124 (O_124,N_9513,N_9786);
nand UO_125 (O_125,N_9660,N_9685);
nor UO_126 (O_126,N_9738,N_9626);
nor UO_127 (O_127,N_9544,N_9860);
or UO_128 (O_128,N_9614,N_9759);
and UO_129 (O_129,N_9926,N_9957);
nor UO_130 (O_130,N_9868,N_9808);
xor UO_131 (O_131,N_9766,N_9534);
xor UO_132 (O_132,N_9502,N_9532);
and UO_133 (O_133,N_9835,N_9913);
xnor UO_134 (O_134,N_9695,N_9967);
nand UO_135 (O_135,N_9611,N_9608);
nor UO_136 (O_136,N_9953,N_9709);
or UO_137 (O_137,N_9700,N_9780);
nor UO_138 (O_138,N_9618,N_9603);
xor UO_139 (O_139,N_9828,N_9819);
nor UO_140 (O_140,N_9804,N_9696);
nand UO_141 (O_141,N_9834,N_9862);
nand UO_142 (O_142,N_9955,N_9682);
or UO_143 (O_143,N_9881,N_9920);
nand UO_144 (O_144,N_9880,N_9753);
nand UO_145 (O_145,N_9523,N_9621);
and UO_146 (O_146,N_9687,N_9942);
or UO_147 (O_147,N_9654,N_9858);
or UO_148 (O_148,N_9717,N_9836);
nand UO_149 (O_149,N_9891,N_9924);
and UO_150 (O_150,N_9977,N_9974);
and UO_151 (O_151,N_9689,N_9765);
or UO_152 (O_152,N_9547,N_9638);
nor UO_153 (O_153,N_9914,N_9988);
nand UO_154 (O_154,N_9941,N_9947);
and UO_155 (O_155,N_9912,N_9814);
and UO_156 (O_156,N_9790,N_9679);
xor UO_157 (O_157,N_9612,N_9506);
or UO_158 (O_158,N_9898,N_9922);
xnor UO_159 (O_159,N_9976,N_9744);
or UO_160 (O_160,N_9751,N_9676);
and UO_161 (O_161,N_9507,N_9586);
nor UO_162 (O_162,N_9726,N_9590);
nor UO_163 (O_163,N_9596,N_9824);
or UO_164 (O_164,N_9627,N_9851);
xor UO_165 (O_165,N_9716,N_9890);
or UO_166 (O_166,N_9599,N_9812);
or UO_167 (O_167,N_9613,N_9710);
or UO_168 (O_168,N_9793,N_9531);
and UO_169 (O_169,N_9937,N_9809);
nor UO_170 (O_170,N_9571,N_9754);
or UO_171 (O_171,N_9578,N_9732);
nand UO_172 (O_172,N_9882,N_9610);
nor UO_173 (O_173,N_9577,N_9893);
or UO_174 (O_174,N_9623,N_9620);
xor UO_175 (O_175,N_9683,N_9788);
or UO_176 (O_176,N_9833,N_9848);
nand UO_177 (O_177,N_9762,N_9511);
nand UO_178 (O_178,N_9734,N_9816);
nand UO_179 (O_179,N_9649,N_9907);
nor UO_180 (O_180,N_9807,N_9707);
xor UO_181 (O_181,N_9549,N_9849);
xnor UO_182 (O_182,N_9742,N_9639);
xnor UO_183 (O_183,N_9675,N_9575);
nand UO_184 (O_184,N_9857,N_9580);
and UO_185 (O_185,N_9740,N_9693);
xnor UO_186 (O_186,N_9964,N_9706);
and UO_187 (O_187,N_9665,N_9818);
and UO_188 (O_188,N_9925,N_9845);
xor UO_189 (O_189,N_9670,N_9792);
nor UO_190 (O_190,N_9928,N_9642);
xnor UO_191 (O_191,N_9843,N_9823);
and UO_192 (O_192,N_9641,N_9650);
or UO_193 (O_193,N_9991,N_9533);
or UO_194 (O_194,N_9505,N_9989);
and UO_195 (O_195,N_9524,N_9635);
nor UO_196 (O_196,N_9515,N_9583);
or UO_197 (O_197,N_9503,N_9992);
nor UO_198 (O_198,N_9562,N_9615);
or UO_199 (O_199,N_9701,N_9990);
or UO_200 (O_200,N_9827,N_9694);
or UO_201 (O_201,N_9787,N_9718);
or UO_202 (O_202,N_9973,N_9972);
and UO_203 (O_203,N_9516,N_9896);
xnor UO_204 (O_204,N_9633,N_9811);
nand UO_205 (O_205,N_9598,N_9741);
nor UO_206 (O_206,N_9877,N_9806);
nand UO_207 (O_207,N_9768,N_9630);
nor UO_208 (O_208,N_9646,N_9852);
or UO_209 (O_209,N_9536,N_9842);
nor UO_210 (O_210,N_9945,N_9719);
or UO_211 (O_211,N_9906,N_9512);
xor UO_212 (O_212,N_9956,N_9582);
or UO_213 (O_213,N_9998,N_9739);
nand UO_214 (O_214,N_9631,N_9996);
or UO_215 (O_215,N_9930,N_9728);
and UO_216 (O_216,N_9841,N_9915);
xor UO_217 (O_217,N_9847,N_9705);
and UO_218 (O_218,N_9894,N_9859);
xnor UO_219 (O_219,N_9736,N_9715);
nor UO_220 (O_220,N_9657,N_9781);
xor UO_221 (O_221,N_9832,N_9883);
and UO_222 (O_222,N_9800,N_9864);
nand UO_223 (O_223,N_9589,N_9673);
nand UO_224 (O_224,N_9866,N_9632);
and UO_225 (O_225,N_9903,N_9651);
xnor UO_226 (O_226,N_9648,N_9886);
nand UO_227 (O_227,N_9595,N_9601);
xor UO_228 (O_228,N_9850,N_9826);
nor UO_229 (O_229,N_9871,N_9773);
or UO_230 (O_230,N_9775,N_9729);
nor UO_231 (O_231,N_9909,N_9791);
and UO_232 (O_232,N_9879,N_9935);
nor UO_233 (O_233,N_9664,N_9666);
or UO_234 (O_234,N_9901,N_9771);
nor UO_235 (O_235,N_9629,N_9746);
or UO_236 (O_236,N_9936,N_9559);
and UO_237 (O_237,N_9830,N_9667);
nand UO_238 (O_238,N_9698,N_9905);
or UO_239 (O_239,N_9839,N_9782);
or UO_240 (O_240,N_9767,N_9684);
nor UO_241 (O_241,N_9550,N_9846);
nor UO_242 (O_242,N_9725,N_9778);
or UO_243 (O_243,N_9799,N_9921);
nand UO_244 (O_244,N_9949,N_9979);
or UO_245 (O_245,N_9720,N_9643);
nor UO_246 (O_246,N_9796,N_9708);
nand UO_247 (O_247,N_9584,N_9933);
or UO_248 (O_248,N_9525,N_9948);
or UO_249 (O_249,N_9769,N_9887);
nand UO_250 (O_250,N_9662,N_9860);
and UO_251 (O_251,N_9767,N_9766);
nand UO_252 (O_252,N_9924,N_9680);
nor UO_253 (O_253,N_9922,N_9956);
nand UO_254 (O_254,N_9793,N_9873);
xor UO_255 (O_255,N_9858,N_9584);
nand UO_256 (O_256,N_9899,N_9961);
xnor UO_257 (O_257,N_9766,N_9725);
nand UO_258 (O_258,N_9587,N_9559);
and UO_259 (O_259,N_9917,N_9866);
nand UO_260 (O_260,N_9920,N_9764);
xnor UO_261 (O_261,N_9814,N_9785);
nor UO_262 (O_262,N_9900,N_9581);
nor UO_263 (O_263,N_9506,N_9562);
xor UO_264 (O_264,N_9747,N_9728);
xor UO_265 (O_265,N_9615,N_9847);
and UO_266 (O_266,N_9602,N_9889);
or UO_267 (O_267,N_9699,N_9944);
nor UO_268 (O_268,N_9957,N_9879);
and UO_269 (O_269,N_9553,N_9560);
and UO_270 (O_270,N_9962,N_9829);
nand UO_271 (O_271,N_9913,N_9702);
nor UO_272 (O_272,N_9927,N_9531);
and UO_273 (O_273,N_9665,N_9561);
or UO_274 (O_274,N_9633,N_9711);
and UO_275 (O_275,N_9933,N_9872);
and UO_276 (O_276,N_9946,N_9577);
or UO_277 (O_277,N_9894,N_9934);
or UO_278 (O_278,N_9552,N_9560);
or UO_279 (O_279,N_9723,N_9797);
and UO_280 (O_280,N_9806,N_9503);
or UO_281 (O_281,N_9574,N_9585);
nor UO_282 (O_282,N_9609,N_9675);
or UO_283 (O_283,N_9652,N_9917);
and UO_284 (O_284,N_9692,N_9629);
nor UO_285 (O_285,N_9606,N_9851);
and UO_286 (O_286,N_9871,N_9673);
nand UO_287 (O_287,N_9976,N_9942);
nand UO_288 (O_288,N_9662,N_9909);
nor UO_289 (O_289,N_9958,N_9910);
or UO_290 (O_290,N_9733,N_9680);
xnor UO_291 (O_291,N_9759,N_9572);
and UO_292 (O_292,N_9900,N_9856);
xnor UO_293 (O_293,N_9759,N_9722);
nand UO_294 (O_294,N_9784,N_9924);
and UO_295 (O_295,N_9897,N_9806);
xnor UO_296 (O_296,N_9945,N_9904);
and UO_297 (O_297,N_9547,N_9569);
or UO_298 (O_298,N_9957,N_9795);
nand UO_299 (O_299,N_9721,N_9935);
nor UO_300 (O_300,N_9841,N_9753);
xnor UO_301 (O_301,N_9750,N_9992);
nand UO_302 (O_302,N_9584,N_9770);
or UO_303 (O_303,N_9800,N_9868);
and UO_304 (O_304,N_9697,N_9595);
nor UO_305 (O_305,N_9796,N_9563);
xor UO_306 (O_306,N_9568,N_9644);
nor UO_307 (O_307,N_9529,N_9959);
nand UO_308 (O_308,N_9954,N_9623);
nor UO_309 (O_309,N_9509,N_9571);
nand UO_310 (O_310,N_9663,N_9617);
or UO_311 (O_311,N_9794,N_9633);
xnor UO_312 (O_312,N_9523,N_9561);
nor UO_313 (O_313,N_9879,N_9936);
nand UO_314 (O_314,N_9942,N_9876);
and UO_315 (O_315,N_9858,N_9994);
and UO_316 (O_316,N_9641,N_9702);
nor UO_317 (O_317,N_9701,N_9872);
or UO_318 (O_318,N_9616,N_9820);
nand UO_319 (O_319,N_9528,N_9601);
xor UO_320 (O_320,N_9907,N_9935);
and UO_321 (O_321,N_9754,N_9884);
or UO_322 (O_322,N_9589,N_9520);
xor UO_323 (O_323,N_9815,N_9532);
nand UO_324 (O_324,N_9615,N_9824);
and UO_325 (O_325,N_9727,N_9511);
and UO_326 (O_326,N_9791,N_9929);
nor UO_327 (O_327,N_9795,N_9661);
or UO_328 (O_328,N_9621,N_9930);
nor UO_329 (O_329,N_9793,N_9838);
nand UO_330 (O_330,N_9914,N_9576);
xor UO_331 (O_331,N_9655,N_9939);
nand UO_332 (O_332,N_9679,N_9581);
nor UO_333 (O_333,N_9601,N_9585);
nand UO_334 (O_334,N_9961,N_9643);
nor UO_335 (O_335,N_9976,N_9574);
or UO_336 (O_336,N_9908,N_9984);
xnor UO_337 (O_337,N_9994,N_9698);
or UO_338 (O_338,N_9781,N_9590);
nor UO_339 (O_339,N_9900,N_9801);
and UO_340 (O_340,N_9677,N_9594);
nand UO_341 (O_341,N_9945,N_9757);
and UO_342 (O_342,N_9988,N_9742);
nand UO_343 (O_343,N_9550,N_9763);
nor UO_344 (O_344,N_9895,N_9975);
xor UO_345 (O_345,N_9931,N_9581);
and UO_346 (O_346,N_9748,N_9636);
nor UO_347 (O_347,N_9645,N_9611);
or UO_348 (O_348,N_9520,N_9878);
or UO_349 (O_349,N_9710,N_9514);
xor UO_350 (O_350,N_9598,N_9550);
and UO_351 (O_351,N_9938,N_9953);
and UO_352 (O_352,N_9714,N_9574);
xnor UO_353 (O_353,N_9744,N_9987);
nand UO_354 (O_354,N_9932,N_9858);
nand UO_355 (O_355,N_9917,N_9646);
nor UO_356 (O_356,N_9961,N_9959);
and UO_357 (O_357,N_9505,N_9849);
nor UO_358 (O_358,N_9867,N_9744);
nor UO_359 (O_359,N_9649,N_9988);
nand UO_360 (O_360,N_9549,N_9766);
or UO_361 (O_361,N_9584,N_9518);
nand UO_362 (O_362,N_9949,N_9811);
and UO_363 (O_363,N_9747,N_9891);
and UO_364 (O_364,N_9529,N_9773);
nand UO_365 (O_365,N_9749,N_9886);
nand UO_366 (O_366,N_9912,N_9826);
xnor UO_367 (O_367,N_9796,N_9986);
and UO_368 (O_368,N_9510,N_9715);
or UO_369 (O_369,N_9865,N_9857);
nor UO_370 (O_370,N_9515,N_9789);
xnor UO_371 (O_371,N_9720,N_9927);
and UO_372 (O_372,N_9507,N_9733);
nand UO_373 (O_373,N_9763,N_9686);
or UO_374 (O_374,N_9738,N_9535);
xnor UO_375 (O_375,N_9601,N_9582);
nand UO_376 (O_376,N_9709,N_9672);
or UO_377 (O_377,N_9680,N_9691);
nor UO_378 (O_378,N_9939,N_9683);
or UO_379 (O_379,N_9802,N_9958);
nand UO_380 (O_380,N_9565,N_9637);
and UO_381 (O_381,N_9971,N_9861);
xnor UO_382 (O_382,N_9607,N_9715);
xor UO_383 (O_383,N_9908,N_9816);
or UO_384 (O_384,N_9755,N_9752);
nand UO_385 (O_385,N_9851,N_9784);
nand UO_386 (O_386,N_9505,N_9724);
nor UO_387 (O_387,N_9945,N_9986);
nand UO_388 (O_388,N_9990,N_9860);
nor UO_389 (O_389,N_9824,N_9774);
nor UO_390 (O_390,N_9629,N_9611);
and UO_391 (O_391,N_9729,N_9821);
and UO_392 (O_392,N_9835,N_9794);
nor UO_393 (O_393,N_9816,N_9569);
and UO_394 (O_394,N_9844,N_9963);
xnor UO_395 (O_395,N_9862,N_9674);
nor UO_396 (O_396,N_9869,N_9991);
or UO_397 (O_397,N_9623,N_9900);
xnor UO_398 (O_398,N_9709,N_9905);
or UO_399 (O_399,N_9580,N_9539);
xor UO_400 (O_400,N_9901,N_9850);
nor UO_401 (O_401,N_9547,N_9650);
xnor UO_402 (O_402,N_9585,N_9920);
nor UO_403 (O_403,N_9730,N_9861);
nor UO_404 (O_404,N_9946,N_9803);
or UO_405 (O_405,N_9770,N_9824);
nor UO_406 (O_406,N_9746,N_9522);
and UO_407 (O_407,N_9637,N_9863);
or UO_408 (O_408,N_9866,N_9537);
nor UO_409 (O_409,N_9872,N_9912);
nor UO_410 (O_410,N_9990,N_9921);
xor UO_411 (O_411,N_9873,N_9771);
xor UO_412 (O_412,N_9782,N_9525);
xor UO_413 (O_413,N_9537,N_9627);
or UO_414 (O_414,N_9671,N_9728);
xor UO_415 (O_415,N_9818,N_9901);
nand UO_416 (O_416,N_9960,N_9540);
nor UO_417 (O_417,N_9953,N_9550);
and UO_418 (O_418,N_9697,N_9648);
and UO_419 (O_419,N_9695,N_9638);
or UO_420 (O_420,N_9911,N_9737);
nand UO_421 (O_421,N_9923,N_9999);
nand UO_422 (O_422,N_9993,N_9565);
or UO_423 (O_423,N_9767,N_9926);
or UO_424 (O_424,N_9765,N_9888);
nor UO_425 (O_425,N_9556,N_9928);
xnor UO_426 (O_426,N_9567,N_9841);
nor UO_427 (O_427,N_9628,N_9566);
or UO_428 (O_428,N_9510,N_9587);
nand UO_429 (O_429,N_9688,N_9892);
or UO_430 (O_430,N_9659,N_9807);
xnor UO_431 (O_431,N_9656,N_9610);
and UO_432 (O_432,N_9719,N_9988);
and UO_433 (O_433,N_9863,N_9969);
or UO_434 (O_434,N_9990,N_9797);
xnor UO_435 (O_435,N_9817,N_9695);
nor UO_436 (O_436,N_9968,N_9759);
nand UO_437 (O_437,N_9604,N_9594);
nor UO_438 (O_438,N_9559,N_9922);
or UO_439 (O_439,N_9737,N_9669);
nand UO_440 (O_440,N_9899,N_9974);
xnor UO_441 (O_441,N_9942,N_9908);
and UO_442 (O_442,N_9867,N_9933);
nand UO_443 (O_443,N_9976,N_9949);
nand UO_444 (O_444,N_9898,N_9596);
nor UO_445 (O_445,N_9611,N_9711);
nor UO_446 (O_446,N_9719,N_9994);
nor UO_447 (O_447,N_9800,N_9940);
and UO_448 (O_448,N_9868,N_9939);
nor UO_449 (O_449,N_9689,N_9740);
or UO_450 (O_450,N_9891,N_9854);
nor UO_451 (O_451,N_9693,N_9569);
or UO_452 (O_452,N_9980,N_9960);
xnor UO_453 (O_453,N_9651,N_9582);
and UO_454 (O_454,N_9812,N_9581);
xor UO_455 (O_455,N_9867,N_9690);
nand UO_456 (O_456,N_9614,N_9879);
nor UO_457 (O_457,N_9718,N_9781);
xnor UO_458 (O_458,N_9665,N_9957);
and UO_459 (O_459,N_9707,N_9522);
and UO_460 (O_460,N_9618,N_9680);
and UO_461 (O_461,N_9931,N_9563);
or UO_462 (O_462,N_9530,N_9812);
xnor UO_463 (O_463,N_9627,N_9692);
and UO_464 (O_464,N_9879,N_9990);
or UO_465 (O_465,N_9961,N_9515);
xnor UO_466 (O_466,N_9724,N_9681);
nor UO_467 (O_467,N_9565,N_9560);
xnor UO_468 (O_468,N_9851,N_9986);
nand UO_469 (O_469,N_9591,N_9555);
and UO_470 (O_470,N_9881,N_9772);
xor UO_471 (O_471,N_9580,N_9660);
xor UO_472 (O_472,N_9993,N_9648);
xor UO_473 (O_473,N_9948,N_9694);
and UO_474 (O_474,N_9859,N_9759);
nand UO_475 (O_475,N_9590,N_9770);
xor UO_476 (O_476,N_9896,N_9777);
nand UO_477 (O_477,N_9660,N_9511);
nand UO_478 (O_478,N_9682,N_9883);
nand UO_479 (O_479,N_9920,N_9620);
nor UO_480 (O_480,N_9677,N_9727);
nor UO_481 (O_481,N_9889,N_9922);
xor UO_482 (O_482,N_9981,N_9553);
nor UO_483 (O_483,N_9731,N_9626);
nand UO_484 (O_484,N_9746,N_9942);
nand UO_485 (O_485,N_9845,N_9948);
or UO_486 (O_486,N_9865,N_9740);
nor UO_487 (O_487,N_9808,N_9513);
nor UO_488 (O_488,N_9715,N_9762);
or UO_489 (O_489,N_9618,N_9694);
nand UO_490 (O_490,N_9606,N_9632);
xnor UO_491 (O_491,N_9588,N_9630);
or UO_492 (O_492,N_9743,N_9776);
nor UO_493 (O_493,N_9834,N_9761);
and UO_494 (O_494,N_9786,N_9936);
and UO_495 (O_495,N_9769,N_9523);
and UO_496 (O_496,N_9733,N_9833);
nand UO_497 (O_497,N_9720,N_9917);
xor UO_498 (O_498,N_9900,N_9985);
nand UO_499 (O_499,N_9553,N_9684);
and UO_500 (O_500,N_9510,N_9872);
nor UO_501 (O_501,N_9658,N_9695);
and UO_502 (O_502,N_9791,N_9953);
xor UO_503 (O_503,N_9561,N_9541);
nand UO_504 (O_504,N_9697,N_9510);
nor UO_505 (O_505,N_9889,N_9784);
or UO_506 (O_506,N_9537,N_9581);
and UO_507 (O_507,N_9972,N_9705);
nand UO_508 (O_508,N_9662,N_9586);
nand UO_509 (O_509,N_9980,N_9966);
nand UO_510 (O_510,N_9688,N_9725);
nor UO_511 (O_511,N_9796,N_9890);
nand UO_512 (O_512,N_9765,N_9585);
and UO_513 (O_513,N_9502,N_9857);
xor UO_514 (O_514,N_9698,N_9696);
and UO_515 (O_515,N_9699,N_9629);
nor UO_516 (O_516,N_9848,N_9901);
and UO_517 (O_517,N_9905,N_9815);
xor UO_518 (O_518,N_9815,N_9789);
nand UO_519 (O_519,N_9641,N_9646);
xor UO_520 (O_520,N_9633,N_9660);
or UO_521 (O_521,N_9502,N_9910);
nand UO_522 (O_522,N_9633,N_9568);
nand UO_523 (O_523,N_9533,N_9929);
nor UO_524 (O_524,N_9611,N_9730);
nor UO_525 (O_525,N_9666,N_9597);
nor UO_526 (O_526,N_9645,N_9623);
nor UO_527 (O_527,N_9569,N_9838);
or UO_528 (O_528,N_9939,N_9562);
nor UO_529 (O_529,N_9579,N_9572);
nor UO_530 (O_530,N_9894,N_9649);
or UO_531 (O_531,N_9831,N_9785);
nand UO_532 (O_532,N_9991,N_9544);
nor UO_533 (O_533,N_9508,N_9570);
nand UO_534 (O_534,N_9890,N_9952);
and UO_535 (O_535,N_9917,N_9563);
or UO_536 (O_536,N_9675,N_9612);
or UO_537 (O_537,N_9819,N_9718);
xor UO_538 (O_538,N_9757,N_9835);
nand UO_539 (O_539,N_9869,N_9523);
xnor UO_540 (O_540,N_9817,N_9592);
xor UO_541 (O_541,N_9557,N_9625);
nor UO_542 (O_542,N_9599,N_9523);
nand UO_543 (O_543,N_9955,N_9750);
or UO_544 (O_544,N_9734,N_9946);
and UO_545 (O_545,N_9686,N_9918);
or UO_546 (O_546,N_9852,N_9691);
nor UO_547 (O_547,N_9788,N_9516);
or UO_548 (O_548,N_9960,N_9686);
and UO_549 (O_549,N_9989,N_9941);
and UO_550 (O_550,N_9532,N_9554);
nand UO_551 (O_551,N_9803,N_9774);
and UO_552 (O_552,N_9644,N_9506);
nand UO_553 (O_553,N_9894,N_9588);
xnor UO_554 (O_554,N_9773,N_9878);
and UO_555 (O_555,N_9973,N_9649);
xnor UO_556 (O_556,N_9689,N_9652);
nor UO_557 (O_557,N_9693,N_9975);
nor UO_558 (O_558,N_9577,N_9655);
or UO_559 (O_559,N_9970,N_9580);
nand UO_560 (O_560,N_9823,N_9870);
xor UO_561 (O_561,N_9710,N_9868);
nand UO_562 (O_562,N_9866,N_9673);
nor UO_563 (O_563,N_9967,N_9713);
xor UO_564 (O_564,N_9518,N_9990);
and UO_565 (O_565,N_9930,N_9707);
nand UO_566 (O_566,N_9800,N_9554);
xnor UO_567 (O_567,N_9948,N_9633);
nor UO_568 (O_568,N_9768,N_9587);
nor UO_569 (O_569,N_9849,N_9791);
nor UO_570 (O_570,N_9712,N_9523);
nor UO_571 (O_571,N_9892,N_9985);
nor UO_572 (O_572,N_9854,N_9894);
or UO_573 (O_573,N_9782,N_9764);
and UO_574 (O_574,N_9723,N_9570);
or UO_575 (O_575,N_9819,N_9549);
and UO_576 (O_576,N_9736,N_9650);
and UO_577 (O_577,N_9958,N_9753);
and UO_578 (O_578,N_9674,N_9506);
or UO_579 (O_579,N_9590,N_9549);
nand UO_580 (O_580,N_9847,N_9614);
nand UO_581 (O_581,N_9916,N_9860);
or UO_582 (O_582,N_9919,N_9811);
nor UO_583 (O_583,N_9903,N_9762);
or UO_584 (O_584,N_9535,N_9672);
or UO_585 (O_585,N_9853,N_9542);
and UO_586 (O_586,N_9796,N_9524);
nand UO_587 (O_587,N_9909,N_9562);
and UO_588 (O_588,N_9999,N_9588);
and UO_589 (O_589,N_9602,N_9769);
xor UO_590 (O_590,N_9709,N_9560);
or UO_591 (O_591,N_9832,N_9737);
nand UO_592 (O_592,N_9577,N_9801);
nand UO_593 (O_593,N_9876,N_9925);
and UO_594 (O_594,N_9591,N_9993);
and UO_595 (O_595,N_9713,N_9901);
nand UO_596 (O_596,N_9650,N_9762);
or UO_597 (O_597,N_9726,N_9915);
xnor UO_598 (O_598,N_9718,N_9527);
or UO_599 (O_599,N_9815,N_9749);
nand UO_600 (O_600,N_9772,N_9509);
xor UO_601 (O_601,N_9769,N_9550);
or UO_602 (O_602,N_9511,N_9662);
nor UO_603 (O_603,N_9785,N_9588);
xor UO_604 (O_604,N_9846,N_9519);
or UO_605 (O_605,N_9734,N_9680);
nand UO_606 (O_606,N_9596,N_9880);
nor UO_607 (O_607,N_9933,N_9540);
nand UO_608 (O_608,N_9650,N_9959);
or UO_609 (O_609,N_9590,N_9769);
or UO_610 (O_610,N_9837,N_9904);
or UO_611 (O_611,N_9873,N_9600);
nand UO_612 (O_612,N_9710,N_9607);
nand UO_613 (O_613,N_9735,N_9641);
and UO_614 (O_614,N_9604,N_9606);
nand UO_615 (O_615,N_9941,N_9601);
nand UO_616 (O_616,N_9608,N_9576);
xnor UO_617 (O_617,N_9839,N_9606);
xnor UO_618 (O_618,N_9608,N_9520);
nand UO_619 (O_619,N_9801,N_9505);
nand UO_620 (O_620,N_9939,N_9661);
xnor UO_621 (O_621,N_9785,N_9506);
nor UO_622 (O_622,N_9962,N_9898);
and UO_623 (O_623,N_9768,N_9697);
nand UO_624 (O_624,N_9925,N_9866);
xor UO_625 (O_625,N_9558,N_9606);
nor UO_626 (O_626,N_9707,N_9954);
nand UO_627 (O_627,N_9834,N_9650);
nor UO_628 (O_628,N_9968,N_9683);
and UO_629 (O_629,N_9611,N_9767);
and UO_630 (O_630,N_9964,N_9537);
xor UO_631 (O_631,N_9622,N_9562);
nand UO_632 (O_632,N_9719,N_9750);
or UO_633 (O_633,N_9594,N_9772);
xnor UO_634 (O_634,N_9839,N_9757);
nand UO_635 (O_635,N_9837,N_9970);
nor UO_636 (O_636,N_9662,N_9524);
nor UO_637 (O_637,N_9693,N_9932);
nand UO_638 (O_638,N_9890,N_9879);
nand UO_639 (O_639,N_9916,N_9800);
and UO_640 (O_640,N_9812,N_9694);
or UO_641 (O_641,N_9814,N_9777);
and UO_642 (O_642,N_9757,N_9654);
xnor UO_643 (O_643,N_9585,N_9609);
nor UO_644 (O_644,N_9665,N_9732);
and UO_645 (O_645,N_9835,N_9993);
and UO_646 (O_646,N_9859,N_9593);
or UO_647 (O_647,N_9615,N_9623);
xnor UO_648 (O_648,N_9845,N_9680);
xnor UO_649 (O_649,N_9562,N_9977);
and UO_650 (O_650,N_9991,N_9877);
xnor UO_651 (O_651,N_9728,N_9863);
xnor UO_652 (O_652,N_9705,N_9949);
nor UO_653 (O_653,N_9946,N_9603);
nor UO_654 (O_654,N_9934,N_9989);
or UO_655 (O_655,N_9853,N_9860);
nor UO_656 (O_656,N_9963,N_9754);
xnor UO_657 (O_657,N_9534,N_9899);
and UO_658 (O_658,N_9635,N_9889);
and UO_659 (O_659,N_9666,N_9541);
or UO_660 (O_660,N_9599,N_9866);
xor UO_661 (O_661,N_9972,N_9887);
nor UO_662 (O_662,N_9549,N_9516);
or UO_663 (O_663,N_9838,N_9896);
xnor UO_664 (O_664,N_9805,N_9915);
xnor UO_665 (O_665,N_9690,N_9751);
xnor UO_666 (O_666,N_9695,N_9840);
nor UO_667 (O_667,N_9910,N_9569);
or UO_668 (O_668,N_9519,N_9959);
xor UO_669 (O_669,N_9820,N_9611);
or UO_670 (O_670,N_9851,N_9580);
nand UO_671 (O_671,N_9967,N_9626);
or UO_672 (O_672,N_9525,N_9715);
or UO_673 (O_673,N_9731,N_9839);
xnor UO_674 (O_674,N_9885,N_9578);
xor UO_675 (O_675,N_9963,N_9707);
xor UO_676 (O_676,N_9900,N_9835);
and UO_677 (O_677,N_9655,N_9828);
nor UO_678 (O_678,N_9991,N_9740);
nor UO_679 (O_679,N_9926,N_9533);
or UO_680 (O_680,N_9997,N_9660);
nor UO_681 (O_681,N_9851,N_9683);
xnor UO_682 (O_682,N_9969,N_9881);
nand UO_683 (O_683,N_9813,N_9559);
nor UO_684 (O_684,N_9874,N_9597);
nand UO_685 (O_685,N_9593,N_9766);
nor UO_686 (O_686,N_9746,N_9985);
or UO_687 (O_687,N_9744,N_9835);
xor UO_688 (O_688,N_9646,N_9857);
or UO_689 (O_689,N_9813,N_9867);
xnor UO_690 (O_690,N_9777,N_9970);
and UO_691 (O_691,N_9715,N_9708);
and UO_692 (O_692,N_9522,N_9753);
and UO_693 (O_693,N_9738,N_9879);
nor UO_694 (O_694,N_9766,N_9734);
xor UO_695 (O_695,N_9502,N_9861);
nand UO_696 (O_696,N_9743,N_9961);
and UO_697 (O_697,N_9917,N_9521);
and UO_698 (O_698,N_9546,N_9801);
nand UO_699 (O_699,N_9513,N_9989);
and UO_700 (O_700,N_9906,N_9654);
nor UO_701 (O_701,N_9694,N_9624);
and UO_702 (O_702,N_9666,N_9841);
and UO_703 (O_703,N_9552,N_9599);
and UO_704 (O_704,N_9597,N_9730);
nand UO_705 (O_705,N_9565,N_9866);
and UO_706 (O_706,N_9618,N_9590);
nand UO_707 (O_707,N_9938,N_9972);
or UO_708 (O_708,N_9650,N_9895);
nand UO_709 (O_709,N_9985,N_9545);
xor UO_710 (O_710,N_9578,N_9862);
nand UO_711 (O_711,N_9619,N_9755);
nand UO_712 (O_712,N_9780,N_9584);
xor UO_713 (O_713,N_9879,N_9661);
nor UO_714 (O_714,N_9762,N_9936);
or UO_715 (O_715,N_9695,N_9782);
and UO_716 (O_716,N_9681,N_9984);
xor UO_717 (O_717,N_9990,N_9925);
or UO_718 (O_718,N_9710,N_9546);
nand UO_719 (O_719,N_9620,N_9519);
nor UO_720 (O_720,N_9591,N_9619);
nand UO_721 (O_721,N_9983,N_9869);
nand UO_722 (O_722,N_9857,N_9639);
xor UO_723 (O_723,N_9763,N_9724);
and UO_724 (O_724,N_9870,N_9969);
nand UO_725 (O_725,N_9904,N_9738);
nand UO_726 (O_726,N_9505,N_9542);
nand UO_727 (O_727,N_9509,N_9858);
or UO_728 (O_728,N_9637,N_9935);
xnor UO_729 (O_729,N_9836,N_9574);
xor UO_730 (O_730,N_9597,N_9924);
or UO_731 (O_731,N_9800,N_9789);
xor UO_732 (O_732,N_9864,N_9618);
and UO_733 (O_733,N_9864,N_9944);
or UO_734 (O_734,N_9854,N_9705);
xor UO_735 (O_735,N_9625,N_9809);
or UO_736 (O_736,N_9839,N_9790);
xnor UO_737 (O_737,N_9745,N_9896);
nor UO_738 (O_738,N_9616,N_9996);
and UO_739 (O_739,N_9776,N_9532);
and UO_740 (O_740,N_9572,N_9768);
nand UO_741 (O_741,N_9744,N_9917);
xor UO_742 (O_742,N_9956,N_9554);
nor UO_743 (O_743,N_9691,N_9948);
nand UO_744 (O_744,N_9533,N_9517);
nand UO_745 (O_745,N_9645,N_9829);
or UO_746 (O_746,N_9770,N_9705);
or UO_747 (O_747,N_9764,N_9592);
nor UO_748 (O_748,N_9999,N_9788);
xor UO_749 (O_749,N_9805,N_9833);
and UO_750 (O_750,N_9841,N_9842);
or UO_751 (O_751,N_9895,N_9958);
nand UO_752 (O_752,N_9839,N_9829);
or UO_753 (O_753,N_9619,N_9898);
xnor UO_754 (O_754,N_9780,N_9662);
nor UO_755 (O_755,N_9581,N_9752);
and UO_756 (O_756,N_9868,N_9615);
xnor UO_757 (O_757,N_9653,N_9556);
and UO_758 (O_758,N_9754,N_9938);
and UO_759 (O_759,N_9924,N_9968);
and UO_760 (O_760,N_9759,N_9606);
nor UO_761 (O_761,N_9564,N_9890);
nor UO_762 (O_762,N_9551,N_9697);
or UO_763 (O_763,N_9695,N_9607);
or UO_764 (O_764,N_9586,N_9613);
xnor UO_765 (O_765,N_9831,N_9815);
nor UO_766 (O_766,N_9554,N_9689);
or UO_767 (O_767,N_9866,N_9933);
nor UO_768 (O_768,N_9549,N_9511);
nor UO_769 (O_769,N_9791,N_9868);
xnor UO_770 (O_770,N_9531,N_9526);
xnor UO_771 (O_771,N_9670,N_9731);
xnor UO_772 (O_772,N_9625,N_9529);
nor UO_773 (O_773,N_9894,N_9904);
nand UO_774 (O_774,N_9845,N_9895);
xnor UO_775 (O_775,N_9705,N_9666);
xnor UO_776 (O_776,N_9550,N_9966);
xor UO_777 (O_777,N_9809,N_9684);
nor UO_778 (O_778,N_9732,N_9575);
or UO_779 (O_779,N_9626,N_9629);
xor UO_780 (O_780,N_9915,N_9942);
or UO_781 (O_781,N_9551,N_9932);
or UO_782 (O_782,N_9820,N_9772);
and UO_783 (O_783,N_9919,N_9793);
or UO_784 (O_784,N_9894,N_9687);
and UO_785 (O_785,N_9979,N_9610);
or UO_786 (O_786,N_9917,N_9714);
nand UO_787 (O_787,N_9828,N_9981);
or UO_788 (O_788,N_9700,N_9602);
nor UO_789 (O_789,N_9788,N_9770);
or UO_790 (O_790,N_9739,N_9615);
or UO_791 (O_791,N_9521,N_9616);
xor UO_792 (O_792,N_9784,N_9779);
nand UO_793 (O_793,N_9569,N_9839);
nand UO_794 (O_794,N_9941,N_9886);
nor UO_795 (O_795,N_9504,N_9853);
or UO_796 (O_796,N_9899,N_9733);
or UO_797 (O_797,N_9652,N_9691);
nor UO_798 (O_798,N_9667,N_9984);
xor UO_799 (O_799,N_9913,N_9829);
nand UO_800 (O_800,N_9951,N_9632);
xnor UO_801 (O_801,N_9763,N_9752);
and UO_802 (O_802,N_9991,N_9592);
or UO_803 (O_803,N_9822,N_9808);
nor UO_804 (O_804,N_9923,N_9868);
and UO_805 (O_805,N_9743,N_9778);
nand UO_806 (O_806,N_9546,N_9615);
or UO_807 (O_807,N_9889,N_9972);
xnor UO_808 (O_808,N_9664,N_9774);
nor UO_809 (O_809,N_9624,N_9884);
or UO_810 (O_810,N_9679,N_9552);
xor UO_811 (O_811,N_9952,N_9504);
nor UO_812 (O_812,N_9605,N_9963);
and UO_813 (O_813,N_9849,N_9646);
or UO_814 (O_814,N_9870,N_9631);
xnor UO_815 (O_815,N_9844,N_9973);
xnor UO_816 (O_816,N_9569,N_9772);
nand UO_817 (O_817,N_9560,N_9636);
and UO_818 (O_818,N_9527,N_9763);
xnor UO_819 (O_819,N_9927,N_9994);
nand UO_820 (O_820,N_9726,N_9575);
xor UO_821 (O_821,N_9868,N_9670);
and UO_822 (O_822,N_9597,N_9989);
xnor UO_823 (O_823,N_9752,N_9641);
nor UO_824 (O_824,N_9635,N_9899);
nand UO_825 (O_825,N_9706,N_9922);
nand UO_826 (O_826,N_9896,N_9766);
xnor UO_827 (O_827,N_9988,N_9755);
or UO_828 (O_828,N_9829,N_9574);
nand UO_829 (O_829,N_9581,N_9710);
nor UO_830 (O_830,N_9945,N_9962);
nand UO_831 (O_831,N_9747,N_9505);
nor UO_832 (O_832,N_9706,N_9544);
nand UO_833 (O_833,N_9912,N_9577);
or UO_834 (O_834,N_9590,N_9699);
xor UO_835 (O_835,N_9958,N_9761);
or UO_836 (O_836,N_9717,N_9532);
or UO_837 (O_837,N_9978,N_9965);
or UO_838 (O_838,N_9690,N_9765);
xor UO_839 (O_839,N_9674,N_9704);
or UO_840 (O_840,N_9920,N_9696);
and UO_841 (O_841,N_9538,N_9947);
or UO_842 (O_842,N_9625,N_9915);
xor UO_843 (O_843,N_9786,N_9689);
or UO_844 (O_844,N_9925,N_9576);
nand UO_845 (O_845,N_9936,N_9979);
xnor UO_846 (O_846,N_9816,N_9603);
nor UO_847 (O_847,N_9865,N_9994);
xor UO_848 (O_848,N_9882,N_9968);
and UO_849 (O_849,N_9843,N_9911);
or UO_850 (O_850,N_9517,N_9776);
xor UO_851 (O_851,N_9742,N_9926);
and UO_852 (O_852,N_9639,N_9762);
nor UO_853 (O_853,N_9830,N_9522);
or UO_854 (O_854,N_9699,N_9563);
or UO_855 (O_855,N_9994,N_9694);
or UO_856 (O_856,N_9943,N_9636);
and UO_857 (O_857,N_9509,N_9826);
xnor UO_858 (O_858,N_9563,N_9883);
xor UO_859 (O_859,N_9962,N_9774);
and UO_860 (O_860,N_9630,N_9812);
or UO_861 (O_861,N_9526,N_9680);
nand UO_862 (O_862,N_9893,N_9631);
xnor UO_863 (O_863,N_9721,N_9531);
nand UO_864 (O_864,N_9623,N_9730);
nor UO_865 (O_865,N_9502,N_9840);
nand UO_866 (O_866,N_9528,N_9706);
or UO_867 (O_867,N_9658,N_9971);
nor UO_868 (O_868,N_9694,N_9510);
or UO_869 (O_869,N_9952,N_9862);
or UO_870 (O_870,N_9888,N_9678);
xnor UO_871 (O_871,N_9799,N_9760);
xnor UO_872 (O_872,N_9697,N_9660);
or UO_873 (O_873,N_9718,N_9594);
and UO_874 (O_874,N_9880,N_9623);
xor UO_875 (O_875,N_9987,N_9783);
xnor UO_876 (O_876,N_9873,N_9965);
nor UO_877 (O_877,N_9638,N_9862);
or UO_878 (O_878,N_9809,N_9632);
or UO_879 (O_879,N_9634,N_9932);
xnor UO_880 (O_880,N_9709,N_9539);
xnor UO_881 (O_881,N_9946,N_9607);
or UO_882 (O_882,N_9646,N_9618);
and UO_883 (O_883,N_9884,N_9961);
nor UO_884 (O_884,N_9941,N_9698);
nand UO_885 (O_885,N_9533,N_9718);
nand UO_886 (O_886,N_9726,N_9913);
xor UO_887 (O_887,N_9865,N_9917);
or UO_888 (O_888,N_9864,N_9966);
nand UO_889 (O_889,N_9682,N_9972);
nand UO_890 (O_890,N_9580,N_9552);
and UO_891 (O_891,N_9978,N_9829);
and UO_892 (O_892,N_9576,N_9657);
xnor UO_893 (O_893,N_9556,N_9910);
nand UO_894 (O_894,N_9789,N_9555);
xor UO_895 (O_895,N_9601,N_9824);
nor UO_896 (O_896,N_9830,N_9845);
and UO_897 (O_897,N_9654,N_9794);
nand UO_898 (O_898,N_9827,N_9877);
nor UO_899 (O_899,N_9583,N_9762);
and UO_900 (O_900,N_9551,N_9992);
xor UO_901 (O_901,N_9833,N_9973);
nand UO_902 (O_902,N_9809,N_9713);
nor UO_903 (O_903,N_9532,N_9668);
nand UO_904 (O_904,N_9785,N_9636);
nand UO_905 (O_905,N_9890,N_9574);
or UO_906 (O_906,N_9813,N_9539);
xnor UO_907 (O_907,N_9703,N_9791);
or UO_908 (O_908,N_9855,N_9740);
nand UO_909 (O_909,N_9851,N_9556);
and UO_910 (O_910,N_9865,N_9529);
or UO_911 (O_911,N_9624,N_9828);
nand UO_912 (O_912,N_9973,N_9814);
nand UO_913 (O_913,N_9897,N_9681);
and UO_914 (O_914,N_9757,N_9707);
xor UO_915 (O_915,N_9564,N_9587);
xnor UO_916 (O_916,N_9786,N_9846);
xnor UO_917 (O_917,N_9539,N_9521);
and UO_918 (O_918,N_9965,N_9609);
and UO_919 (O_919,N_9864,N_9580);
or UO_920 (O_920,N_9809,N_9683);
xor UO_921 (O_921,N_9539,N_9950);
nor UO_922 (O_922,N_9598,N_9830);
nor UO_923 (O_923,N_9863,N_9660);
and UO_924 (O_924,N_9622,N_9565);
and UO_925 (O_925,N_9958,N_9737);
nand UO_926 (O_926,N_9770,N_9603);
nor UO_927 (O_927,N_9963,N_9730);
or UO_928 (O_928,N_9754,N_9854);
or UO_929 (O_929,N_9585,N_9683);
or UO_930 (O_930,N_9671,N_9513);
and UO_931 (O_931,N_9882,N_9513);
or UO_932 (O_932,N_9981,N_9652);
nand UO_933 (O_933,N_9793,N_9533);
xnor UO_934 (O_934,N_9940,N_9938);
and UO_935 (O_935,N_9579,N_9543);
and UO_936 (O_936,N_9797,N_9934);
and UO_937 (O_937,N_9814,N_9552);
and UO_938 (O_938,N_9768,N_9843);
and UO_939 (O_939,N_9565,N_9799);
xnor UO_940 (O_940,N_9734,N_9765);
nor UO_941 (O_941,N_9924,N_9616);
or UO_942 (O_942,N_9624,N_9656);
and UO_943 (O_943,N_9845,N_9573);
xor UO_944 (O_944,N_9579,N_9763);
nor UO_945 (O_945,N_9866,N_9525);
or UO_946 (O_946,N_9637,N_9584);
xor UO_947 (O_947,N_9621,N_9761);
and UO_948 (O_948,N_9969,N_9629);
or UO_949 (O_949,N_9578,N_9707);
xnor UO_950 (O_950,N_9796,N_9508);
or UO_951 (O_951,N_9939,N_9989);
and UO_952 (O_952,N_9623,N_9823);
nor UO_953 (O_953,N_9609,N_9554);
nand UO_954 (O_954,N_9599,N_9638);
xnor UO_955 (O_955,N_9540,N_9977);
xor UO_956 (O_956,N_9772,N_9732);
nand UO_957 (O_957,N_9806,N_9934);
xnor UO_958 (O_958,N_9807,N_9536);
xor UO_959 (O_959,N_9960,N_9738);
or UO_960 (O_960,N_9712,N_9839);
xnor UO_961 (O_961,N_9874,N_9610);
xor UO_962 (O_962,N_9935,N_9727);
and UO_963 (O_963,N_9615,N_9756);
or UO_964 (O_964,N_9893,N_9747);
nor UO_965 (O_965,N_9708,N_9648);
nor UO_966 (O_966,N_9673,N_9693);
or UO_967 (O_967,N_9620,N_9954);
nor UO_968 (O_968,N_9636,N_9837);
xor UO_969 (O_969,N_9980,N_9584);
nor UO_970 (O_970,N_9618,N_9832);
nor UO_971 (O_971,N_9887,N_9832);
nand UO_972 (O_972,N_9540,N_9641);
and UO_973 (O_973,N_9600,N_9770);
nand UO_974 (O_974,N_9885,N_9925);
xnor UO_975 (O_975,N_9821,N_9534);
or UO_976 (O_976,N_9773,N_9937);
and UO_977 (O_977,N_9699,N_9824);
and UO_978 (O_978,N_9661,N_9687);
nand UO_979 (O_979,N_9607,N_9684);
or UO_980 (O_980,N_9718,N_9602);
or UO_981 (O_981,N_9847,N_9796);
xnor UO_982 (O_982,N_9989,N_9573);
xnor UO_983 (O_983,N_9985,N_9949);
nand UO_984 (O_984,N_9608,N_9716);
and UO_985 (O_985,N_9636,N_9706);
xnor UO_986 (O_986,N_9941,N_9818);
nor UO_987 (O_987,N_9768,N_9979);
and UO_988 (O_988,N_9608,N_9788);
xor UO_989 (O_989,N_9643,N_9973);
nor UO_990 (O_990,N_9724,N_9811);
xor UO_991 (O_991,N_9511,N_9646);
and UO_992 (O_992,N_9875,N_9854);
or UO_993 (O_993,N_9598,N_9841);
xor UO_994 (O_994,N_9615,N_9801);
or UO_995 (O_995,N_9564,N_9783);
or UO_996 (O_996,N_9967,N_9730);
nand UO_997 (O_997,N_9743,N_9966);
and UO_998 (O_998,N_9940,N_9841);
xnor UO_999 (O_999,N_9510,N_9757);
nor UO_1000 (O_1000,N_9518,N_9793);
nand UO_1001 (O_1001,N_9892,N_9752);
xnor UO_1002 (O_1002,N_9861,N_9646);
and UO_1003 (O_1003,N_9786,N_9913);
nand UO_1004 (O_1004,N_9779,N_9641);
xor UO_1005 (O_1005,N_9865,N_9815);
xnor UO_1006 (O_1006,N_9682,N_9813);
nand UO_1007 (O_1007,N_9754,N_9613);
xor UO_1008 (O_1008,N_9693,N_9562);
nor UO_1009 (O_1009,N_9950,N_9939);
xnor UO_1010 (O_1010,N_9883,N_9810);
xnor UO_1011 (O_1011,N_9696,N_9879);
nand UO_1012 (O_1012,N_9807,N_9612);
xor UO_1013 (O_1013,N_9713,N_9665);
nand UO_1014 (O_1014,N_9708,N_9789);
nor UO_1015 (O_1015,N_9526,N_9713);
and UO_1016 (O_1016,N_9906,N_9874);
xnor UO_1017 (O_1017,N_9776,N_9978);
nor UO_1018 (O_1018,N_9684,N_9975);
or UO_1019 (O_1019,N_9504,N_9906);
nand UO_1020 (O_1020,N_9675,N_9932);
nand UO_1021 (O_1021,N_9774,N_9657);
or UO_1022 (O_1022,N_9770,N_9724);
nor UO_1023 (O_1023,N_9883,N_9671);
xor UO_1024 (O_1024,N_9919,N_9752);
nand UO_1025 (O_1025,N_9718,N_9854);
nand UO_1026 (O_1026,N_9626,N_9841);
or UO_1027 (O_1027,N_9822,N_9964);
xnor UO_1028 (O_1028,N_9850,N_9946);
xnor UO_1029 (O_1029,N_9907,N_9741);
and UO_1030 (O_1030,N_9872,N_9843);
nor UO_1031 (O_1031,N_9863,N_9753);
nand UO_1032 (O_1032,N_9809,N_9817);
xnor UO_1033 (O_1033,N_9790,N_9659);
and UO_1034 (O_1034,N_9812,N_9718);
and UO_1035 (O_1035,N_9921,N_9566);
and UO_1036 (O_1036,N_9676,N_9899);
xor UO_1037 (O_1037,N_9700,N_9644);
nor UO_1038 (O_1038,N_9587,N_9591);
nand UO_1039 (O_1039,N_9679,N_9555);
and UO_1040 (O_1040,N_9758,N_9698);
and UO_1041 (O_1041,N_9637,N_9973);
xnor UO_1042 (O_1042,N_9754,N_9733);
nand UO_1043 (O_1043,N_9782,N_9888);
or UO_1044 (O_1044,N_9877,N_9932);
nand UO_1045 (O_1045,N_9644,N_9754);
xor UO_1046 (O_1046,N_9767,N_9994);
or UO_1047 (O_1047,N_9678,N_9675);
nand UO_1048 (O_1048,N_9920,N_9748);
nand UO_1049 (O_1049,N_9878,N_9944);
or UO_1050 (O_1050,N_9797,N_9592);
or UO_1051 (O_1051,N_9992,N_9792);
nand UO_1052 (O_1052,N_9606,N_9981);
or UO_1053 (O_1053,N_9672,N_9974);
nand UO_1054 (O_1054,N_9925,N_9950);
nor UO_1055 (O_1055,N_9720,N_9622);
or UO_1056 (O_1056,N_9754,N_9922);
and UO_1057 (O_1057,N_9922,N_9763);
nand UO_1058 (O_1058,N_9657,N_9700);
and UO_1059 (O_1059,N_9745,N_9994);
or UO_1060 (O_1060,N_9879,N_9512);
nand UO_1061 (O_1061,N_9549,N_9730);
xor UO_1062 (O_1062,N_9947,N_9551);
and UO_1063 (O_1063,N_9549,N_9978);
nor UO_1064 (O_1064,N_9867,N_9962);
and UO_1065 (O_1065,N_9696,N_9637);
or UO_1066 (O_1066,N_9699,N_9810);
xnor UO_1067 (O_1067,N_9692,N_9732);
nor UO_1068 (O_1068,N_9880,N_9738);
xnor UO_1069 (O_1069,N_9609,N_9980);
nand UO_1070 (O_1070,N_9504,N_9815);
nand UO_1071 (O_1071,N_9690,N_9825);
xor UO_1072 (O_1072,N_9635,N_9963);
xor UO_1073 (O_1073,N_9809,N_9969);
nor UO_1074 (O_1074,N_9755,N_9784);
nor UO_1075 (O_1075,N_9773,N_9846);
xor UO_1076 (O_1076,N_9587,N_9611);
and UO_1077 (O_1077,N_9781,N_9999);
nor UO_1078 (O_1078,N_9898,N_9537);
and UO_1079 (O_1079,N_9782,N_9940);
xnor UO_1080 (O_1080,N_9546,N_9642);
nor UO_1081 (O_1081,N_9548,N_9617);
and UO_1082 (O_1082,N_9862,N_9720);
nand UO_1083 (O_1083,N_9984,N_9807);
nand UO_1084 (O_1084,N_9780,N_9594);
and UO_1085 (O_1085,N_9865,N_9770);
or UO_1086 (O_1086,N_9593,N_9718);
nor UO_1087 (O_1087,N_9812,N_9945);
and UO_1088 (O_1088,N_9781,N_9808);
nand UO_1089 (O_1089,N_9691,N_9870);
xor UO_1090 (O_1090,N_9637,N_9596);
xor UO_1091 (O_1091,N_9987,N_9789);
or UO_1092 (O_1092,N_9766,N_9856);
nor UO_1093 (O_1093,N_9976,N_9531);
and UO_1094 (O_1094,N_9518,N_9570);
nor UO_1095 (O_1095,N_9892,N_9730);
and UO_1096 (O_1096,N_9729,N_9647);
or UO_1097 (O_1097,N_9508,N_9626);
xnor UO_1098 (O_1098,N_9608,N_9929);
xor UO_1099 (O_1099,N_9766,N_9605);
xor UO_1100 (O_1100,N_9729,N_9677);
nor UO_1101 (O_1101,N_9736,N_9832);
xnor UO_1102 (O_1102,N_9736,N_9870);
or UO_1103 (O_1103,N_9690,N_9991);
or UO_1104 (O_1104,N_9959,N_9600);
xnor UO_1105 (O_1105,N_9788,N_9824);
nand UO_1106 (O_1106,N_9723,N_9922);
nand UO_1107 (O_1107,N_9899,N_9856);
nor UO_1108 (O_1108,N_9656,N_9831);
nor UO_1109 (O_1109,N_9936,N_9646);
nor UO_1110 (O_1110,N_9565,N_9831);
nor UO_1111 (O_1111,N_9990,N_9894);
nor UO_1112 (O_1112,N_9568,N_9550);
nand UO_1113 (O_1113,N_9961,N_9842);
and UO_1114 (O_1114,N_9957,N_9659);
nor UO_1115 (O_1115,N_9842,N_9558);
nor UO_1116 (O_1116,N_9861,N_9617);
xor UO_1117 (O_1117,N_9665,N_9568);
nor UO_1118 (O_1118,N_9531,N_9629);
nand UO_1119 (O_1119,N_9630,N_9658);
or UO_1120 (O_1120,N_9825,N_9523);
nor UO_1121 (O_1121,N_9605,N_9839);
and UO_1122 (O_1122,N_9709,N_9755);
nor UO_1123 (O_1123,N_9749,N_9851);
xor UO_1124 (O_1124,N_9649,N_9573);
xnor UO_1125 (O_1125,N_9868,N_9653);
nor UO_1126 (O_1126,N_9584,N_9790);
nand UO_1127 (O_1127,N_9555,N_9557);
or UO_1128 (O_1128,N_9996,N_9682);
nand UO_1129 (O_1129,N_9874,N_9612);
xor UO_1130 (O_1130,N_9837,N_9649);
xnor UO_1131 (O_1131,N_9672,N_9528);
nand UO_1132 (O_1132,N_9869,N_9848);
and UO_1133 (O_1133,N_9965,N_9618);
nand UO_1134 (O_1134,N_9880,N_9865);
or UO_1135 (O_1135,N_9812,N_9738);
or UO_1136 (O_1136,N_9740,N_9661);
and UO_1137 (O_1137,N_9686,N_9985);
nor UO_1138 (O_1138,N_9818,N_9981);
nand UO_1139 (O_1139,N_9742,N_9857);
nor UO_1140 (O_1140,N_9645,N_9582);
xor UO_1141 (O_1141,N_9881,N_9746);
nor UO_1142 (O_1142,N_9548,N_9864);
or UO_1143 (O_1143,N_9735,N_9520);
and UO_1144 (O_1144,N_9614,N_9907);
nand UO_1145 (O_1145,N_9832,N_9802);
nand UO_1146 (O_1146,N_9991,N_9723);
nand UO_1147 (O_1147,N_9816,N_9842);
nand UO_1148 (O_1148,N_9713,N_9982);
nor UO_1149 (O_1149,N_9713,N_9947);
or UO_1150 (O_1150,N_9613,N_9908);
or UO_1151 (O_1151,N_9811,N_9909);
nand UO_1152 (O_1152,N_9664,N_9852);
xnor UO_1153 (O_1153,N_9912,N_9925);
or UO_1154 (O_1154,N_9613,N_9723);
xnor UO_1155 (O_1155,N_9701,N_9857);
and UO_1156 (O_1156,N_9889,N_9620);
or UO_1157 (O_1157,N_9600,N_9822);
nor UO_1158 (O_1158,N_9650,N_9786);
or UO_1159 (O_1159,N_9757,N_9996);
xnor UO_1160 (O_1160,N_9891,N_9905);
and UO_1161 (O_1161,N_9865,N_9874);
and UO_1162 (O_1162,N_9906,N_9711);
nor UO_1163 (O_1163,N_9580,N_9900);
nand UO_1164 (O_1164,N_9524,N_9922);
xor UO_1165 (O_1165,N_9930,N_9967);
and UO_1166 (O_1166,N_9610,N_9559);
xor UO_1167 (O_1167,N_9934,N_9725);
or UO_1168 (O_1168,N_9721,N_9507);
xor UO_1169 (O_1169,N_9603,N_9645);
and UO_1170 (O_1170,N_9729,N_9540);
xnor UO_1171 (O_1171,N_9920,N_9622);
xor UO_1172 (O_1172,N_9515,N_9952);
or UO_1173 (O_1173,N_9965,N_9693);
nand UO_1174 (O_1174,N_9533,N_9565);
xor UO_1175 (O_1175,N_9825,N_9504);
nand UO_1176 (O_1176,N_9609,N_9687);
nand UO_1177 (O_1177,N_9931,N_9823);
xnor UO_1178 (O_1178,N_9892,N_9563);
nand UO_1179 (O_1179,N_9634,N_9604);
nor UO_1180 (O_1180,N_9563,N_9615);
nand UO_1181 (O_1181,N_9634,N_9941);
nor UO_1182 (O_1182,N_9880,N_9693);
nand UO_1183 (O_1183,N_9871,N_9710);
nand UO_1184 (O_1184,N_9925,N_9910);
and UO_1185 (O_1185,N_9749,N_9601);
nor UO_1186 (O_1186,N_9997,N_9597);
xor UO_1187 (O_1187,N_9948,N_9584);
nor UO_1188 (O_1188,N_9756,N_9676);
and UO_1189 (O_1189,N_9761,N_9980);
nand UO_1190 (O_1190,N_9844,N_9831);
and UO_1191 (O_1191,N_9691,N_9727);
nor UO_1192 (O_1192,N_9645,N_9983);
nand UO_1193 (O_1193,N_9639,N_9992);
or UO_1194 (O_1194,N_9588,N_9806);
xor UO_1195 (O_1195,N_9661,N_9852);
xnor UO_1196 (O_1196,N_9576,N_9689);
and UO_1197 (O_1197,N_9517,N_9973);
nand UO_1198 (O_1198,N_9637,N_9933);
and UO_1199 (O_1199,N_9660,N_9950);
and UO_1200 (O_1200,N_9767,N_9789);
nor UO_1201 (O_1201,N_9703,N_9737);
xor UO_1202 (O_1202,N_9508,N_9595);
nor UO_1203 (O_1203,N_9542,N_9506);
nor UO_1204 (O_1204,N_9563,N_9888);
xnor UO_1205 (O_1205,N_9645,N_9970);
nor UO_1206 (O_1206,N_9764,N_9565);
nand UO_1207 (O_1207,N_9817,N_9783);
nor UO_1208 (O_1208,N_9580,N_9574);
nand UO_1209 (O_1209,N_9575,N_9591);
or UO_1210 (O_1210,N_9653,N_9821);
or UO_1211 (O_1211,N_9586,N_9598);
or UO_1212 (O_1212,N_9642,N_9523);
nor UO_1213 (O_1213,N_9609,N_9647);
and UO_1214 (O_1214,N_9955,N_9679);
nor UO_1215 (O_1215,N_9522,N_9556);
nand UO_1216 (O_1216,N_9628,N_9873);
nor UO_1217 (O_1217,N_9556,N_9609);
nor UO_1218 (O_1218,N_9578,N_9831);
or UO_1219 (O_1219,N_9572,N_9733);
xnor UO_1220 (O_1220,N_9954,N_9576);
xor UO_1221 (O_1221,N_9836,N_9619);
or UO_1222 (O_1222,N_9894,N_9769);
and UO_1223 (O_1223,N_9914,N_9541);
or UO_1224 (O_1224,N_9907,N_9538);
nor UO_1225 (O_1225,N_9509,N_9746);
xnor UO_1226 (O_1226,N_9659,N_9917);
xor UO_1227 (O_1227,N_9851,N_9810);
or UO_1228 (O_1228,N_9792,N_9926);
or UO_1229 (O_1229,N_9925,N_9522);
or UO_1230 (O_1230,N_9915,N_9842);
nor UO_1231 (O_1231,N_9525,N_9707);
or UO_1232 (O_1232,N_9719,N_9794);
and UO_1233 (O_1233,N_9801,N_9929);
xor UO_1234 (O_1234,N_9713,N_9850);
and UO_1235 (O_1235,N_9763,N_9990);
xnor UO_1236 (O_1236,N_9738,N_9811);
nand UO_1237 (O_1237,N_9563,N_9932);
or UO_1238 (O_1238,N_9693,N_9820);
and UO_1239 (O_1239,N_9902,N_9923);
and UO_1240 (O_1240,N_9968,N_9930);
and UO_1241 (O_1241,N_9594,N_9566);
and UO_1242 (O_1242,N_9506,N_9679);
xnor UO_1243 (O_1243,N_9919,N_9597);
nor UO_1244 (O_1244,N_9660,N_9995);
or UO_1245 (O_1245,N_9807,N_9637);
or UO_1246 (O_1246,N_9820,N_9536);
nor UO_1247 (O_1247,N_9896,N_9682);
and UO_1248 (O_1248,N_9609,N_9869);
and UO_1249 (O_1249,N_9869,N_9982);
and UO_1250 (O_1250,N_9522,N_9745);
nor UO_1251 (O_1251,N_9818,N_9848);
nand UO_1252 (O_1252,N_9861,N_9811);
nor UO_1253 (O_1253,N_9767,N_9571);
nand UO_1254 (O_1254,N_9765,N_9716);
or UO_1255 (O_1255,N_9765,N_9662);
nand UO_1256 (O_1256,N_9962,N_9555);
nor UO_1257 (O_1257,N_9865,N_9615);
or UO_1258 (O_1258,N_9774,N_9567);
xor UO_1259 (O_1259,N_9561,N_9833);
nand UO_1260 (O_1260,N_9945,N_9741);
xnor UO_1261 (O_1261,N_9882,N_9947);
xor UO_1262 (O_1262,N_9714,N_9895);
or UO_1263 (O_1263,N_9659,N_9934);
nor UO_1264 (O_1264,N_9549,N_9811);
or UO_1265 (O_1265,N_9517,N_9596);
and UO_1266 (O_1266,N_9928,N_9888);
or UO_1267 (O_1267,N_9950,N_9514);
xor UO_1268 (O_1268,N_9992,N_9515);
nand UO_1269 (O_1269,N_9551,N_9512);
nor UO_1270 (O_1270,N_9940,N_9538);
or UO_1271 (O_1271,N_9558,N_9756);
xor UO_1272 (O_1272,N_9711,N_9518);
and UO_1273 (O_1273,N_9951,N_9784);
xor UO_1274 (O_1274,N_9876,N_9551);
or UO_1275 (O_1275,N_9997,N_9831);
or UO_1276 (O_1276,N_9542,N_9501);
nor UO_1277 (O_1277,N_9982,N_9961);
and UO_1278 (O_1278,N_9919,N_9502);
and UO_1279 (O_1279,N_9640,N_9766);
or UO_1280 (O_1280,N_9919,N_9519);
and UO_1281 (O_1281,N_9622,N_9673);
nand UO_1282 (O_1282,N_9717,N_9556);
nand UO_1283 (O_1283,N_9959,N_9752);
xnor UO_1284 (O_1284,N_9914,N_9900);
and UO_1285 (O_1285,N_9853,N_9990);
and UO_1286 (O_1286,N_9620,N_9553);
nor UO_1287 (O_1287,N_9899,N_9790);
and UO_1288 (O_1288,N_9579,N_9870);
or UO_1289 (O_1289,N_9858,N_9577);
nor UO_1290 (O_1290,N_9650,N_9885);
nor UO_1291 (O_1291,N_9664,N_9613);
xor UO_1292 (O_1292,N_9773,N_9507);
and UO_1293 (O_1293,N_9932,N_9701);
and UO_1294 (O_1294,N_9899,N_9834);
nor UO_1295 (O_1295,N_9614,N_9642);
nor UO_1296 (O_1296,N_9923,N_9955);
nand UO_1297 (O_1297,N_9699,N_9514);
or UO_1298 (O_1298,N_9834,N_9811);
nand UO_1299 (O_1299,N_9667,N_9856);
nor UO_1300 (O_1300,N_9834,N_9861);
and UO_1301 (O_1301,N_9531,N_9599);
and UO_1302 (O_1302,N_9956,N_9648);
nand UO_1303 (O_1303,N_9705,N_9641);
and UO_1304 (O_1304,N_9916,N_9826);
nor UO_1305 (O_1305,N_9721,N_9847);
nor UO_1306 (O_1306,N_9698,N_9640);
nand UO_1307 (O_1307,N_9524,N_9715);
nor UO_1308 (O_1308,N_9938,N_9694);
xnor UO_1309 (O_1309,N_9722,N_9527);
or UO_1310 (O_1310,N_9977,N_9620);
xnor UO_1311 (O_1311,N_9907,N_9610);
xor UO_1312 (O_1312,N_9947,N_9982);
and UO_1313 (O_1313,N_9764,N_9654);
nor UO_1314 (O_1314,N_9779,N_9841);
and UO_1315 (O_1315,N_9679,N_9830);
or UO_1316 (O_1316,N_9920,N_9946);
nor UO_1317 (O_1317,N_9625,N_9857);
nor UO_1318 (O_1318,N_9647,N_9760);
xnor UO_1319 (O_1319,N_9767,N_9915);
and UO_1320 (O_1320,N_9791,N_9939);
xor UO_1321 (O_1321,N_9912,N_9980);
or UO_1322 (O_1322,N_9836,N_9952);
and UO_1323 (O_1323,N_9591,N_9825);
nand UO_1324 (O_1324,N_9666,N_9714);
or UO_1325 (O_1325,N_9505,N_9563);
or UO_1326 (O_1326,N_9784,N_9686);
nor UO_1327 (O_1327,N_9857,N_9829);
and UO_1328 (O_1328,N_9535,N_9879);
xor UO_1329 (O_1329,N_9676,N_9867);
and UO_1330 (O_1330,N_9928,N_9707);
and UO_1331 (O_1331,N_9656,N_9625);
nand UO_1332 (O_1332,N_9532,N_9604);
nor UO_1333 (O_1333,N_9722,N_9649);
and UO_1334 (O_1334,N_9949,N_9827);
and UO_1335 (O_1335,N_9870,N_9718);
xor UO_1336 (O_1336,N_9526,N_9811);
or UO_1337 (O_1337,N_9726,N_9779);
and UO_1338 (O_1338,N_9944,N_9682);
nor UO_1339 (O_1339,N_9700,N_9840);
or UO_1340 (O_1340,N_9612,N_9837);
or UO_1341 (O_1341,N_9839,N_9631);
or UO_1342 (O_1342,N_9584,N_9815);
nor UO_1343 (O_1343,N_9929,N_9910);
nand UO_1344 (O_1344,N_9536,N_9771);
xnor UO_1345 (O_1345,N_9518,N_9827);
xnor UO_1346 (O_1346,N_9828,N_9581);
or UO_1347 (O_1347,N_9740,N_9804);
xnor UO_1348 (O_1348,N_9607,N_9786);
nor UO_1349 (O_1349,N_9882,N_9972);
nand UO_1350 (O_1350,N_9977,N_9754);
or UO_1351 (O_1351,N_9641,N_9826);
or UO_1352 (O_1352,N_9947,N_9925);
xor UO_1353 (O_1353,N_9873,N_9701);
and UO_1354 (O_1354,N_9927,N_9878);
xor UO_1355 (O_1355,N_9858,N_9715);
and UO_1356 (O_1356,N_9886,N_9667);
nand UO_1357 (O_1357,N_9856,N_9718);
xnor UO_1358 (O_1358,N_9841,N_9614);
xor UO_1359 (O_1359,N_9892,N_9738);
and UO_1360 (O_1360,N_9847,N_9722);
xor UO_1361 (O_1361,N_9606,N_9679);
or UO_1362 (O_1362,N_9592,N_9962);
or UO_1363 (O_1363,N_9897,N_9940);
nand UO_1364 (O_1364,N_9709,N_9913);
nor UO_1365 (O_1365,N_9547,N_9542);
nor UO_1366 (O_1366,N_9592,N_9518);
nand UO_1367 (O_1367,N_9677,N_9865);
xnor UO_1368 (O_1368,N_9590,N_9546);
and UO_1369 (O_1369,N_9536,N_9978);
and UO_1370 (O_1370,N_9760,N_9982);
nand UO_1371 (O_1371,N_9548,N_9634);
xnor UO_1372 (O_1372,N_9543,N_9704);
or UO_1373 (O_1373,N_9843,N_9776);
and UO_1374 (O_1374,N_9703,N_9640);
nand UO_1375 (O_1375,N_9614,N_9675);
nor UO_1376 (O_1376,N_9690,N_9852);
xnor UO_1377 (O_1377,N_9584,N_9821);
or UO_1378 (O_1378,N_9530,N_9691);
nor UO_1379 (O_1379,N_9851,N_9988);
nand UO_1380 (O_1380,N_9988,N_9787);
nand UO_1381 (O_1381,N_9535,N_9831);
and UO_1382 (O_1382,N_9764,N_9578);
xnor UO_1383 (O_1383,N_9662,N_9544);
and UO_1384 (O_1384,N_9706,N_9750);
or UO_1385 (O_1385,N_9604,N_9622);
and UO_1386 (O_1386,N_9806,N_9524);
or UO_1387 (O_1387,N_9767,N_9883);
or UO_1388 (O_1388,N_9520,N_9562);
or UO_1389 (O_1389,N_9691,N_9914);
or UO_1390 (O_1390,N_9969,N_9667);
nand UO_1391 (O_1391,N_9648,N_9939);
nand UO_1392 (O_1392,N_9844,N_9823);
nand UO_1393 (O_1393,N_9515,N_9836);
nand UO_1394 (O_1394,N_9979,N_9507);
and UO_1395 (O_1395,N_9744,N_9695);
or UO_1396 (O_1396,N_9511,N_9941);
and UO_1397 (O_1397,N_9504,N_9675);
xnor UO_1398 (O_1398,N_9591,N_9894);
xor UO_1399 (O_1399,N_9761,N_9784);
or UO_1400 (O_1400,N_9832,N_9809);
nor UO_1401 (O_1401,N_9540,N_9940);
or UO_1402 (O_1402,N_9938,N_9535);
or UO_1403 (O_1403,N_9843,N_9877);
xnor UO_1404 (O_1404,N_9914,N_9581);
nor UO_1405 (O_1405,N_9727,N_9579);
nand UO_1406 (O_1406,N_9807,N_9973);
or UO_1407 (O_1407,N_9520,N_9982);
nand UO_1408 (O_1408,N_9752,N_9926);
nor UO_1409 (O_1409,N_9799,N_9910);
and UO_1410 (O_1410,N_9948,N_9524);
nor UO_1411 (O_1411,N_9845,N_9518);
nand UO_1412 (O_1412,N_9651,N_9933);
nor UO_1413 (O_1413,N_9992,N_9953);
or UO_1414 (O_1414,N_9557,N_9617);
nor UO_1415 (O_1415,N_9712,N_9813);
nand UO_1416 (O_1416,N_9855,N_9745);
or UO_1417 (O_1417,N_9594,N_9542);
or UO_1418 (O_1418,N_9916,N_9908);
nor UO_1419 (O_1419,N_9965,N_9827);
xor UO_1420 (O_1420,N_9730,N_9907);
nand UO_1421 (O_1421,N_9901,N_9745);
xor UO_1422 (O_1422,N_9611,N_9533);
or UO_1423 (O_1423,N_9746,N_9926);
nor UO_1424 (O_1424,N_9732,N_9868);
nand UO_1425 (O_1425,N_9717,N_9956);
and UO_1426 (O_1426,N_9735,N_9811);
nand UO_1427 (O_1427,N_9552,N_9559);
nor UO_1428 (O_1428,N_9634,N_9891);
or UO_1429 (O_1429,N_9763,N_9578);
nor UO_1430 (O_1430,N_9504,N_9839);
nand UO_1431 (O_1431,N_9691,N_9790);
and UO_1432 (O_1432,N_9872,N_9795);
nor UO_1433 (O_1433,N_9500,N_9744);
nand UO_1434 (O_1434,N_9905,N_9658);
nand UO_1435 (O_1435,N_9699,N_9532);
nor UO_1436 (O_1436,N_9527,N_9706);
or UO_1437 (O_1437,N_9673,N_9686);
xnor UO_1438 (O_1438,N_9647,N_9858);
xnor UO_1439 (O_1439,N_9787,N_9528);
or UO_1440 (O_1440,N_9699,N_9708);
nor UO_1441 (O_1441,N_9790,N_9667);
or UO_1442 (O_1442,N_9892,N_9862);
and UO_1443 (O_1443,N_9802,N_9539);
xor UO_1444 (O_1444,N_9911,N_9531);
nor UO_1445 (O_1445,N_9856,N_9628);
xor UO_1446 (O_1446,N_9577,N_9684);
and UO_1447 (O_1447,N_9865,N_9709);
xor UO_1448 (O_1448,N_9524,N_9800);
or UO_1449 (O_1449,N_9575,N_9956);
nand UO_1450 (O_1450,N_9624,N_9542);
or UO_1451 (O_1451,N_9711,N_9969);
nand UO_1452 (O_1452,N_9581,N_9533);
or UO_1453 (O_1453,N_9511,N_9529);
or UO_1454 (O_1454,N_9667,N_9953);
or UO_1455 (O_1455,N_9990,N_9998);
or UO_1456 (O_1456,N_9727,N_9702);
nor UO_1457 (O_1457,N_9911,N_9809);
nor UO_1458 (O_1458,N_9845,N_9846);
xnor UO_1459 (O_1459,N_9680,N_9518);
xor UO_1460 (O_1460,N_9537,N_9797);
and UO_1461 (O_1461,N_9709,N_9625);
nand UO_1462 (O_1462,N_9826,N_9862);
xor UO_1463 (O_1463,N_9550,N_9587);
or UO_1464 (O_1464,N_9827,N_9664);
xnor UO_1465 (O_1465,N_9595,N_9745);
nor UO_1466 (O_1466,N_9524,N_9992);
and UO_1467 (O_1467,N_9601,N_9835);
nor UO_1468 (O_1468,N_9682,N_9722);
nor UO_1469 (O_1469,N_9758,N_9857);
xnor UO_1470 (O_1470,N_9613,N_9881);
nor UO_1471 (O_1471,N_9967,N_9618);
or UO_1472 (O_1472,N_9662,N_9526);
nor UO_1473 (O_1473,N_9917,N_9716);
or UO_1474 (O_1474,N_9799,N_9964);
or UO_1475 (O_1475,N_9562,N_9925);
or UO_1476 (O_1476,N_9756,N_9865);
xnor UO_1477 (O_1477,N_9638,N_9836);
xnor UO_1478 (O_1478,N_9552,N_9777);
nor UO_1479 (O_1479,N_9716,N_9837);
nor UO_1480 (O_1480,N_9828,N_9872);
and UO_1481 (O_1481,N_9958,N_9658);
nor UO_1482 (O_1482,N_9732,N_9883);
nand UO_1483 (O_1483,N_9789,N_9861);
or UO_1484 (O_1484,N_9907,N_9721);
nand UO_1485 (O_1485,N_9731,N_9921);
nor UO_1486 (O_1486,N_9726,N_9708);
and UO_1487 (O_1487,N_9771,N_9973);
or UO_1488 (O_1488,N_9787,N_9743);
or UO_1489 (O_1489,N_9615,N_9889);
xnor UO_1490 (O_1490,N_9535,N_9841);
or UO_1491 (O_1491,N_9899,N_9583);
or UO_1492 (O_1492,N_9984,N_9792);
xnor UO_1493 (O_1493,N_9602,N_9890);
or UO_1494 (O_1494,N_9698,N_9975);
or UO_1495 (O_1495,N_9753,N_9659);
xnor UO_1496 (O_1496,N_9783,N_9914);
and UO_1497 (O_1497,N_9514,N_9549);
and UO_1498 (O_1498,N_9973,N_9658);
nand UO_1499 (O_1499,N_9942,N_9629);
endmodule