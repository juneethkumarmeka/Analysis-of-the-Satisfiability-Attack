module basic_1500_15000_2000_15_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_82,In_884);
nand U1 (N_1,In_162,In_890);
xor U2 (N_2,In_669,In_245);
or U3 (N_3,In_205,In_1048);
nor U4 (N_4,In_1003,In_883);
nand U5 (N_5,In_399,In_249);
and U6 (N_6,In_1401,In_308);
and U7 (N_7,In_144,In_1483);
or U8 (N_8,In_630,In_27);
nand U9 (N_9,In_58,In_659);
or U10 (N_10,In_812,In_637);
xnor U11 (N_11,In_1001,In_747);
xor U12 (N_12,In_843,In_209);
nand U13 (N_13,In_1245,In_1239);
or U14 (N_14,In_83,In_1074);
and U15 (N_15,In_688,In_1312);
nand U16 (N_16,In_993,In_514);
or U17 (N_17,In_1167,In_856);
nand U18 (N_18,In_732,In_877);
xnor U19 (N_19,In_849,In_605);
or U20 (N_20,In_1413,In_227);
xor U21 (N_21,In_210,In_7);
nor U22 (N_22,In_1147,In_445);
or U23 (N_23,In_655,In_789);
or U24 (N_24,In_1259,In_534);
nand U25 (N_25,In_93,In_1263);
and U26 (N_26,In_486,In_173);
or U27 (N_27,In_1327,In_982);
xor U28 (N_28,In_979,In_721);
nand U29 (N_29,In_692,In_527);
xnor U30 (N_30,In_525,In_932);
xnor U31 (N_31,In_1301,In_1258);
xor U32 (N_32,In_412,In_97);
nor U33 (N_33,In_99,In_914);
nand U34 (N_34,In_78,In_295);
and U35 (N_35,In_766,In_1212);
nand U36 (N_36,In_171,In_679);
nor U37 (N_37,In_850,In_744);
and U38 (N_38,In_1362,In_1075);
or U39 (N_39,In_323,In_45);
xnor U40 (N_40,In_670,In_892);
nand U41 (N_41,In_651,In_1410);
or U42 (N_42,In_95,In_204);
nor U43 (N_43,In_56,In_14);
xnor U44 (N_44,In_453,In_1382);
xor U45 (N_45,In_950,In_522);
xnor U46 (N_46,In_1468,In_600);
and U47 (N_47,In_864,In_1027);
and U48 (N_48,In_328,In_132);
and U49 (N_49,In_1170,In_919);
or U50 (N_50,In_1324,In_963);
nor U51 (N_51,In_889,In_1023);
nand U52 (N_52,In_1024,In_943);
nor U53 (N_53,In_1415,In_594);
or U54 (N_54,In_134,In_322);
and U55 (N_55,In_573,In_625);
or U56 (N_56,In_777,In_108);
nand U57 (N_57,In_248,In_549);
nand U58 (N_58,In_438,In_1015);
and U59 (N_59,In_832,In_432);
and U60 (N_60,In_974,In_555);
xnor U61 (N_61,In_332,In_1206);
or U62 (N_62,In_1252,In_846);
xnor U63 (N_63,In_1179,In_735);
or U64 (N_64,In_192,In_619);
or U65 (N_65,In_513,In_265);
and U66 (N_66,In_775,In_269);
and U67 (N_67,In_301,In_1274);
or U68 (N_68,In_1223,In_660);
nand U69 (N_69,In_1095,In_1232);
xor U70 (N_70,In_1225,In_949);
nor U71 (N_71,In_1266,In_1041);
nand U72 (N_72,In_303,In_163);
nor U73 (N_73,In_575,In_583);
xnor U74 (N_74,In_211,In_1283);
nand U75 (N_75,In_1000,In_218);
nor U76 (N_76,In_1113,In_553);
nor U77 (N_77,In_327,In_566);
xnor U78 (N_78,In_639,In_1273);
and U79 (N_79,In_13,In_723);
xor U80 (N_80,In_1143,In_570);
and U81 (N_81,In_120,In_1172);
or U82 (N_82,In_256,In_1151);
nand U83 (N_83,In_1036,In_1211);
xor U84 (N_84,In_543,In_1062);
or U85 (N_85,In_1103,In_447);
and U86 (N_86,In_800,In_425);
nor U87 (N_87,In_598,In_1496);
nor U88 (N_88,In_469,In_1220);
xor U89 (N_89,In_546,In_562);
and U90 (N_90,In_48,In_776);
xnor U91 (N_91,In_745,In_764);
nand U92 (N_92,In_729,In_741);
and U93 (N_93,In_417,In_661);
nor U94 (N_94,In_400,In_719);
nand U95 (N_95,In_101,In_885);
or U96 (N_96,In_1008,In_935);
or U97 (N_97,In_1017,In_253);
nand U98 (N_98,In_1213,In_1304);
or U99 (N_99,In_1313,In_881);
nor U100 (N_100,In_581,In_39);
or U101 (N_101,In_678,In_848);
nand U102 (N_102,In_451,In_589);
or U103 (N_103,In_1426,In_467);
nand U104 (N_104,In_1291,In_809);
and U105 (N_105,In_1254,In_1489);
nand U106 (N_106,In_448,In_16);
or U107 (N_107,In_636,In_668);
nor U108 (N_108,In_740,In_972);
xor U109 (N_109,In_717,In_1116);
or U110 (N_110,In_393,In_175);
xor U111 (N_111,In_1108,In_1309);
xnor U112 (N_112,In_333,In_786);
and U113 (N_113,In_1169,In_395);
or U114 (N_114,In_371,In_457);
and U115 (N_115,In_1215,In_1011);
and U116 (N_116,In_704,In_81);
nand U117 (N_117,In_1390,In_827);
and U118 (N_118,In_808,In_1499);
or U119 (N_119,In_79,In_1141);
xor U120 (N_120,In_533,In_738);
xnor U121 (N_121,In_861,In_1288);
nor U122 (N_122,In_749,In_646);
and U123 (N_123,In_456,In_307);
xnor U124 (N_124,In_813,In_362);
xor U125 (N_125,In_202,In_606);
or U126 (N_126,In_554,In_1352);
and U127 (N_127,In_998,In_1233);
or U128 (N_128,In_627,In_897);
nand U129 (N_129,In_1201,In_604);
nand U130 (N_130,In_862,In_858);
or U131 (N_131,In_112,In_422);
nand U132 (N_132,In_531,In_185);
and U133 (N_133,In_965,In_302);
xor U134 (N_134,In_1078,In_894);
xor U135 (N_135,In_1334,In_12);
nand U136 (N_136,In_1257,In_869);
nor U137 (N_137,In_722,In_177);
or U138 (N_138,In_561,In_1424);
and U139 (N_139,In_454,In_762);
and U140 (N_140,In_1367,In_226);
xor U141 (N_141,In_318,In_128);
xor U142 (N_142,In_916,In_10);
nand U143 (N_143,In_169,In_1185);
xnor U144 (N_144,In_53,In_1490);
nor U145 (N_145,In_542,In_321);
nand U146 (N_146,In_1429,In_953);
nor U147 (N_147,In_460,In_1081);
or U148 (N_148,In_608,In_491);
nor U149 (N_149,In_1430,In_420);
xor U150 (N_150,In_948,In_336);
and U151 (N_151,In_164,In_1261);
nor U152 (N_152,In_1280,In_1482);
or U153 (N_153,In_330,In_603);
or U154 (N_154,In_551,In_1308);
or U155 (N_155,In_266,In_1355);
and U156 (N_156,In_1067,In_33);
and U157 (N_157,In_443,In_1047);
xor U158 (N_158,In_1091,In_1403);
and U159 (N_159,In_18,In_751);
and U160 (N_160,In_1210,In_1423);
xor U161 (N_161,In_1256,In_1150);
and U162 (N_162,In_1454,In_122);
xor U163 (N_163,In_556,In_76);
nor U164 (N_164,In_1442,In_1061);
and U165 (N_165,In_633,In_615);
xor U166 (N_166,In_37,In_703);
xor U167 (N_167,In_587,In_923);
nor U168 (N_168,In_1123,In_1006);
nand U169 (N_169,In_465,In_1432);
nor U170 (N_170,In_300,In_440);
and U171 (N_171,In_288,In_136);
or U172 (N_172,In_271,In_524);
nor U173 (N_173,In_274,In_797);
and U174 (N_174,In_487,In_1384);
nor U175 (N_175,In_1359,In_1350);
nand U176 (N_176,In_1237,In_1181);
nor U177 (N_177,In_535,In_857);
nor U178 (N_178,In_641,In_154);
or U179 (N_179,In_23,In_331);
nor U180 (N_180,In_1255,In_584);
and U181 (N_181,In_1441,In_879);
nand U182 (N_182,In_1456,In_1360);
and U183 (N_183,In_805,In_273);
nand U184 (N_184,In_1431,In_756);
or U185 (N_185,In_268,In_787);
xor U186 (N_186,In_284,In_1194);
nor U187 (N_187,In_252,In_282);
and U188 (N_188,In_126,In_100);
nand U189 (N_189,In_544,In_552);
and U190 (N_190,In_874,In_1231);
or U191 (N_191,In_1109,In_1495);
and U192 (N_192,In_1180,In_232);
and U193 (N_193,In_221,In_985);
nand U194 (N_194,In_1411,In_1425);
xnor U195 (N_195,In_1096,In_355);
nand U196 (N_196,In_1,In_1476);
xor U197 (N_197,In_803,In_726);
and U198 (N_198,In_1380,In_642);
xnor U199 (N_199,In_1406,In_842);
xor U200 (N_200,In_389,In_822);
and U201 (N_201,In_876,In_1397);
or U202 (N_202,In_290,In_1251);
nor U203 (N_203,In_1458,In_1228);
xnor U204 (N_204,In_1337,In_314);
nand U205 (N_205,In_701,In_286);
or U206 (N_206,In_1464,In_579);
or U207 (N_207,In_85,In_153);
nor U208 (N_208,In_541,In_41);
nand U209 (N_209,In_1402,In_357);
nand U210 (N_210,In_1347,In_1230);
or U211 (N_211,In_1162,In_815);
and U212 (N_212,In_699,In_381);
or U213 (N_213,In_94,In_1404);
and U214 (N_214,In_1176,In_1160);
nor U215 (N_215,In_313,In_230);
xnor U216 (N_216,In_277,In_1089);
nand U217 (N_217,In_161,In_143);
or U218 (N_218,In_29,In_64);
nand U219 (N_219,In_1277,In_398);
nor U220 (N_220,In_1282,In_1012);
nand U221 (N_221,In_1018,In_621);
xor U222 (N_222,In_997,In_996);
or U223 (N_223,In_306,In_969);
and U224 (N_224,In_930,In_1193);
nor U225 (N_225,In_538,In_903);
or U226 (N_226,In_667,In_358);
and U227 (N_227,In_151,In_200);
nand U228 (N_228,In_1467,In_1022);
nand U229 (N_229,In_1224,In_505);
and U230 (N_230,In_394,In_127);
xor U231 (N_231,In_473,In_700);
nor U232 (N_232,In_966,In_289);
nand U233 (N_233,In_1217,In_560);
nand U234 (N_234,In_1372,In_17);
nand U235 (N_235,In_962,In_1065);
nand U236 (N_236,In_69,In_459);
nor U237 (N_237,In_900,In_1445);
nor U238 (N_238,In_572,In_337);
nor U239 (N_239,In_616,In_937);
nor U240 (N_240,In_196,In_20);
and U241 (N_241,In_86,In_326);
xor U242 (N_242,In_658,In_1272);
nor U243 (N_243,In_801,In_353);
nand U244 (N_244,In_939,In_582);
xor U245 (N_245,In_298,In_1448);
nand U246 (N_246,In_1434,In_779);
nor U247 (N_247,In_868,In_504);
and U248 (N_248,In_114,In_882);
nand U249 (N_249,In_638,In_1242);
and U250 (N_250,In_1058,In_278);
xor U251 (N_251,In_565,In_1294);
nand U252 (N_252,In_1025,In_1443);
or U253 (N_253,In_1122,In_372);
nand U254 (N_254,In_329,In_437);
nor U255 (N_255,In_155,In_66);
nand U256 (N_256,In_1192,In_261);
and U257 (N_257,In_622,In_1057);
xor U258 (N_258,In_1357,In_375);
nor U259 (N_259,In_413,In_70);
or U260 (N_260,In_1407,In_835);
and U261 (N_261,In_429,In_891);
xor U262 (N_262,In_135,In_1064);
nor U263 (N_263,In_989,In_590);
nand U264 (N_264,In_1378,In_568);
and U265 (N_265,In_71,In_599);
and U266 (N_266,In_474,In_1115);
or U267 (N_267,In_1440,In_1159);
nand U268 (N_268,In_1154,In_926);
nor U269 (N_269,In_63,In_1447);
nor U270 (N_270,In_404,In_267);
nand U271 (N_271,In_961,In_392);
or U272 (N_272,In_219,In_1034);
or U273 (N_273,In_578,In_1336);
or U274 (N_274,In_246,In_1140);
nand U275 (N_275,In_1052,In_516);
xnor U276 (N_276,In_1284,In_770);
xor U277 (N_277,In_475,In_536);
and U278 (N_278,In_1131,In_145);
or U279 (N_279,In_1374,In_917);
or U280 (N_280,In_526,In_152);
nand U281 (N_281,In_1264,In_880);
xor U282 (N_282,In_825,In_833);
or U283 (N_283,In_1385,In_349);
xor U284 (N_284,In_377,In_571);
and U285 (N_285,In_411,In_506);
or U286 (N_286,In_1016,In_893);
nor U287 (N_287,In_148,In_481);
nor U288 (N_288,In_1085,In_1102);
nand U289 (N_289,In_1144,In_1219);
or U290 (N_290,In_38,In_1369);
nor U291 (N_291,In_558,In_981);
nor U292 (N_292,In_887,In_1148);
nand U293 (N_293,In_793,In_1325);
xor U294 (N_294,In_710,In_416);
or U295 (N_295,In_778,In_913);
xor U296 (N_296,In_1361,In_947);
or U297 (N_297,In_1437,In_229);
nor U298 (N_298,In_195,In_925);
nand U299 (N_299,In_896,In_244);
nand U300 (N_300,In_1182,In_1416);
xnor U301 (N_301,In_1241,In_40);
nand U302 (N_302,In_21,In_987);
nor U303 (N_303,In_414,In_240);
nand U304 (N_304,In_147,In_1340);
nand U305 (N_305,In_1296,In_761);
nand U306 (N_306,In_360,In_67);
nor U307 (N_307,In_264,In_1040);
or U308 (N_308,In_73,In_1435);
or U309 (N_309,In_1297,In_1346);
and U310 (N_310,In_520,In_1107);
nand U311 (N_311,In_1267,In_847);
nor U312 (N_312,In_720,In_225);
xnor U313 (N_313,In_190,In_1135);
or U314 (N_314,In_715,In_597);
xor U315 (N_315,In_74,In_458);
xnor U316 (N_316,In_1342,In_396);
nor U317 (N_317,In_208,In_1472);
and U318 (N_318,In_1487,In_55);
xnor U319 (N_319,In_956,In_992);
or U320 (N_320,In_1279,In_693);
xor U321 (N_321,In_449,In_632);
or U322 (N_322,In_1449,In_257);
and U323 (N_323,In_673,In_921);
nand U324 (N_324,In_283,In_611);
xnor U325 (N_325,In_180,In_662);
or U326 (N_326,In_576,In_117);
nor U327 (N_327,In_410,In_61);
and U328 (N_328,In_348,In_1226);
and U329 (N_329,In_315,In_1097);
and U330 (N_330,In_51,In_166);
or U331 (N_331,In_287,In_905);
nand U332 (N_332,In_401,In_1293);
nor U333 (N_333,In_291,In_484);
or U334 (N_334,In_821,In_121);
nor U335 (N_335,In_757,In_933);
or U336 (N_336,In_772,In_109);
xnor U337 (N_337,In_1079,In_1243);
or U338 (N_338,In_577,In_1009);
nand U339 (N_339,In_1262,In_958);
xnor U340 (N_340,In_1265,In_1019);
or U341 (N_341,In_471,In_1285);
nor U342 (N_342,In_1491,In_816);
xor U343 (N_343,In_77,In_694);
and U344 (N_344,In_1335,In_1238);
nor U345 (N_345,In_702,In_782);
and U346 (N_346,In_1298,In_87);
and U347 (N_347,In_1268,In_111);
or U348 (N_348,In_494,In_380);
nor U349 (N_349,In_72,In_901);
and U350 (N_350,In_30,In_1494);
xor U351 (N_351,In_507,In_837);
nor U352 (N_352,In_384,In_928);
nand U353 (N_353,In_1111,In_1059);
and U354 (N_354,In_493,In_1186);
and U355 (N_355,In_243,In_957);
xor U356 (N_356,In_36,In_968);
or U357 (N_357,In_1486,In_512);
nor U358 (N_358,In_1492,In_1035);
and U359 (N_359,In_807,In_653);
xor U360 (N_360,In_3,In_983);
nand U361 (N_361,In_497,In_319);
and U362 (N_362,In_676,In_378);
nand U363 (N_363,In_304,In_1168);
nand U364 (N_364,In_643,In_174);
xnor U365 (N_365,In_140,In_442);
nor U366 (N_366,In_1187,In_366);
xor U367 (N_367,In_430,In_1094);
nand U368 (N_368,In_1086,In_1249);
or U369 (N_369,In_924,In_888);
nand U370 (N_370,In_994,In_387);
nor U371 (N_371,In_1375,In_1465);
nand U372 (N_372,In_47,In_233);
xnor U373 (N_373,In_1260,In_737);
xnor U374 (N_374,In_1196,In_150);
xor U375 (N_375,In_485,In_385);
and U376 (N_376,In_718,In_539);
nor U377 (N_377,In_755,In_1339);
and U378 (N_378,In_344,In_1177);
xnor U379 (N_379,In_472,In_379);
nor U380 (N_380,In_1234,In_1333);
or U381 (N_381,In_102,In_648);
and U382 (N_382,In_292,In_91);
and U383 (N_383,In_316,In_463);
or U384 (N_384,In_1142,In_68);
nand U385 (N_385,In_1152,In_1127);
xor U386 (N_386,In_60,In_1156);
xor U387 (N_387,In_811,In_1010);
or U388 (N_388,In_1099,In_503);
xor U389 (N_389,In_285,In_629);
xnor U390 (N_390,In_920,In_1269);
and U391 (N_391,In_1171,In_325);
and U392 (N_392,In_1105,In_1341);
and U393 (N_393,In_191,In_783);
or U394 (N_394,In_1110,In_895);
nand U395 (N_395,In_1137,In_674);
and U396 (N_396,In_1028,In_1412);
xor U397 (N_397,In_946,In_428);
xor U398 (N_398,In_1202,In_508);
and U399 (N_399,In_1038,In_197);
xor U400 (N_400,In_716,In_1414);
or U401 (N_401,In_836,In_1207);
xnor U402 (N_402,In_839,In_1497);
xor U403 (N_403,In_343,In_382);
and U404 (N_404,In_272,In_1120);
xor U405 (N_405,In_435,In_517);
xnor U406 (N_406,In_1066,In_1145);
and U407 (N_407,In_376,In_647);
nand U408 (N_408,In_1005,In_125);
nor U409 (N_409,In_580,In_1043);
nand U410 (N_410,In_1275,In_1104);
xnor U411 (N_411,In_515,In_652);
nor U412 (N_412,In_626,In_780);
nor U413 (N_413,In_1363,In_234);
nand U414 (N_414,In_402,In_370);
xnor U415 (N_415,In_359,In_774);
or U416 (N_416,In_142,In_1399);
nand U417 (N_417,In_1190,In_1118);
nand U418 (N_418,In_1128,In_408);
or U419 (N_419,In_557,In_532);
or U420 (N_420,In_1364,In_1029);
nor U421 (N_421,In_80,In_686);
xor U422 (N_422,In_275,In_339);
or U423 (N_423,In_671,In_1485);
nor U424 (N_424,In_1271,In_1316);
and U425 (N_425,In_730,In_1370);
and U426 (N_426,In_806,In_1033);
nand U427 (N_427,In_609,In_1049);
nor U428 (N_428,In_324,In_1130);
or U429 (N_429,In_773,In_624);
and U430 (N_430,In_564,In_46);
and U431 (N_431,In_1218,In_19);
and U432 (N_432,In_1319,In_1462);
and U433 (N_433,In_886,In_1227);
xnor U434 (N_434,In_52,In_912);
nand U435 (N_435,In_1209,In_1157);
xor U436 (N_436,In_262,In_518);
nor U437 (N_437,In_824,In_75);
nor U438 (N_438,In_354,In_592);
and U439 (N_439,In_238,In_1306);
xor U440 (N_440,In_476,In_1365);
nor U441 (N_441,In_159,In_254);
and U442 (N_442,In_975,In_1221);
or U443 (N_443,In_365,In_116);
and U444 (N_444,In_904,In_338);
xor U445 (N_445,In_421,In_707);
and U446 (N_446,In_672,In_407);
nand U447 (N_447,In_1292,In_1229);
xnor U448 (N_448,In_1068,In_96);
or U449 (N_449,In_320,In_1463);
xnor U450 (N_450,In_1175,In_1393);
or U451 (N_451,In_1101,In_1453);
or U452 (N_452,In_6,In_1344);
nor U453 (N_453,In_510,In_1338);
or U454 (N_454,In_1433,In_317);
xor U455 (N_455,In_1060,In_203);
xnor U456 (N_456,In_834,In_1373);
nand U457 (N_457,In_1484,In_118);
or U458 (N_458,In_352,In_231);
xor U459 (N_459,In_1371,In_1470);
xnor U460 (N_460,In_452,In_388);
nand U461 (N_461,In_260,In_1072);
xor U462 (N_462,In_199,In_569);
nor U463 (N_463,In_767,In_1459);
nor U464 (N_464,In_25,In_567);
nand U465 (N_465,In_409,In_613);
nor U466 (N_466,In_259,In_754);
and U467 (N_467,In_426,In_258);
or U468 (N_468,In_753,In_540);
nand U469 (N_469,In_1084,In_820);
xnor U470 (N_470,In_733,In_24);
nand U471 (N_471,In_875,In_680);
and U472 (N_472,In_1153,In_689);
nand U473 (N_473,In_724,In_439);
or U474 (N_474,In_1368,In_511);
nand U475 (N_475,In_129,In_841);
nand U476 (N_476,In_201,In_383);
and U477 (N_477,In_1106,In_529);
nor U478 (N_478,In_665,In_1134);
nand U479 (N_479,In_1199,In_363);
and U480 (N_480,In_984,In_1455);
nor U481 (N_481,In_663,In_586);
xnor U482 (N_482,In_844,In_691);
nor U483 (N_483,In_635,In_139);
and U484 (N_484,In_1165,In_237);
and U485 (N_485,In_1329,In_1400);
xnor U486 (N_486,In_446,In_851);
nor U487 (N_487,In_480,In_477);
or U488 (N_488,In_623,In_1139);
nor U489 (N_489,In_908,In_910);
nand U490 (N_490,In_785,In_911);
nor U491 (N_491,In_938,In_1093);
nor U492 (N_492,In_1444,In_976);
and U493 (N_493,In_312,In_714);
and U494 (N_494,In_138,In_769);
and U495 (N_495,In_1244,In_305);
and U496 (N_496,In_1323,In_944);
nand U497 (N_497,In_479,In_1138);
xor U498 (N_498,In_464,In_1421);
and U499 (N_499,In_470,In_1287);
nor U500 (N_500,In_951,In_1450);
or U501 (N_501,In_973,In_645);
nor U502 (N_502,In_490,In_43);
xor U503 (N_503,In_1114,In_977);
xnor U504 (N_504,In_902,In_872);
and U505 (N_505,In_1351,In_1124);
and U506 (N_506,In_342,In_478);
and U507 (N_507,In_796,In_1133);
nand U508 (N_508,In_133,In_1032);
or U509 (N_509,In_959,In_1418);
nor U510 (N_510,In_734,In_1331);
nor U511 (N_511,In_489,In_854);
xor U512 (N_512,In_1366,In_675);
xnor U513 (N_513,In_364,In_1055);
nor U514 (N_514,In_1044,In_792);
nand U515 (N_515,In_44,In_242);
nor U516 (N_516,In_1200,In_42);
or U517 (N_517,In_373,In_2);
nand U518 (N_518,In_853,In_748);
nor U519 (N_519,In_397,In_1408);
nor U520 (N_520,In_1387,In_548);
xnor U521 (N_521,In_1117,In_165);
or U522 (N_522,In_1250,In_1222);
nand U523 (N_523,In_696,In_631);
xor U524 (N_524,In_1488,In_340);
xor U525 (N_525,In_537,In_967);
nand U526 (N_526,In_1419,In_818);
and U527 (N_527,In_1457,In_1322);
xnor U528 (N_528,In_9,In_115);
and U529 (N_529,In_1112,In_870);
and U530 (N_530,In_945,In_433);
and U531 (N_531,In_1161,In_1381);
nand U532 (N_532,In_293,In_0);
and U533 (N_533,In_954,In_1163);
nand U534 (N_534,In_251,In_547);
nand U535 (N_535,In_212,In_137);
xor U536 (N_536,In_934,In_1051);
nor U537 (N_537,In_1475,In_759);
nor U538 (N_538,In_1173,In_4);
and U539 (N_539,In_865,In_1303);
nand U540 (N_540,In_999,In_1042);
xnor U541 (N_541,In_28,In_57);
and U542 (N_542,In_499,In_742);
nor U543 (N_543,In_170,In_831);
xor U544 (N_544,In_711,In_654);
and U545 (N_545,In_906,In_666);
and U546 (N_546,In_1278,In_113);
and U547 (N_547,In_1466,In_995);
nand U548 (N_548,In_198,In_610);
nor U549 (N_549,In_1083,In_829);
or U550 (N_550,In_620,In_1166);
nor U551 (N_551,In_172,In_15);
or U552 (N_552,In_496,In_1348);
xnor U553 (N_553,In_1203,In_419);
and U554 (N_554,In_105,In_618);
and U555 (N_555,In_223,In_104);
nand U556 (N_556,In_591,In_819);
nor U557 (N_557,In_794,In_1191);
or U558 (N_558,In_585,In_183);
and U559 (N_559,In_1080,In_107);
and U560 (N_560,In_84,In_878);
xnor U561 (N_561,In_840,In_1092);
xnor U562 (N_562,In_574,In_682);
or U563 (N_563,In_1205,In_461);
nor U564 (N_564,In_369,In_178);
xor U565 (N_565,In_179,In_1014);
nor U566 (N_566,In_215,In_1427);
or U567 (N_567,In_131,In_1417);
and U568 (N_568,In_607,In_690);
nor U569 (N_569,In_495,In_50);
nand U570 (N_570,In_1343,In_1132);
and U571 (N_571,In_1039,In_1149);
or U572 (N_572,In_1332,In_588);
and U573 (N_573,In_32,In_1326);
nand U574 (N_574,In_873,In_498);
nand U575 (N_575,In_771,In_1436);
nor U576 (N_576,In_1345,In_1452);
and U577 (N_577,In_1031,In_563);
or U578 (N_578,In_34,In_1349);
and U579 (N_579,In_1070,In_250);
nand U580 (N_580,In_863,In_1146);
or U581 (N_581,In_970,In_991);
nand U582 (N_582,In_1471,In_1054);
or U583 (N_583,In_1314,In_1077);
nor U584 (N_584,In_852,In_441);
nand U585 (N_585,In_1469,In_311);
xnor U586 (N_586,In_1063,In_758);
or U587 (N_587,In_1395,In_224);
nand U588 (N_588,In_750,In_860);
and U589 (N_589,In_482,In_54);
or U590 (N_590,In_1037,In_123);
xnor U591 (N_591,In_186,In_664);
nand U592 (N_592,In_739,In_1354);
or U593 (N_593,In_182,In_502);
nor U594 (N_594,In_255,In_1216);
nor U595 (N_595,In_299,In_802);
nand U596 (N_596,In_1356,In_1396);
and U597 (N_597,In_978,In_390);
and U598 (N_598,In_768,In_931);
nor U599 (N_599,In_89,In_156);
and U600 (N_600,In_450,In_521);
and U601 (N_601,In_1358,In_697);
nor U602 (N_602,In_1236,In_898);
nor U603 (N_603,In_434,In_791);
or U604 (N_604,In_915,In_110);
or U605 (N_605,In_640,In_980);
and U606 (N_606,In_119,In_228);
nor U607 (N_607,In_1253,In_644);
nor U608 (N_608,In_1480,In_1214);
nand U609 (N_609,In_712,In_5);
or U610 (N_610,In_59,In_1087);
nor U611 (N_611,In_500,In_649);
nor U612 (N_612,In_222,In_194);
nor U613 (N_613,In_922,In_1178);
or U614 (N_614,In_657,In_1088);
xor U615 (N_615,In_1204,In_415);
nand U616 (N_616,In_971,In_988);
xnor U617 (N_617,In_1376,In_1289);
nor U618 (N_618,In_188,In_1300);
xnor U619 (N_619,In_294,In_367);
and U620 (N_620,In_1481,In_1197);
or U621 (N_621,In_1136,In_614);
and U622 (N_622,In_149,In_1428);
nor U623 (N_623,In_523,In_828);
xor U624 (N_624,In_1405,In_1391);
xor U625 (N_625,In_1321,In_810);
or U626 (N_626,In_1090,In_727);
and U627 (N_627,In_11,In_909);
xor U628 (N_628,In_270,In_26);
or U629 (N_629,In_35,In_940);
or U630 (N_630,In_207,In_942);
and U631 (N_631,In_677,In_1281);
nor U632 (N_632,In_62,In_705);
or U633 (N_633,In_168,In_466);
and U634 (N_634,In_374,In_709);
and U635 (N_635,In_418,In_859);
or U636 (N_636,In_423,In_1121);
and U637 (N_637,In_368,In_628);
nand U638 (N_638,In_1353,In_386);
nor U639 (N_639,In_927,In_296);
and U640 (N_640,In_1479,In_1305);
nor U641 (N_641,In_1460,In_804);
xor U642 (N_642,In_867,In_1439);
xnor U643 (N_643,In_167,In_1020);
xnor U644 (N_644,In_1286,In_1310);
nand U645 (N_645,In_350,In_405);
nand U646 (N_646,In_687,In_601);
xor U647 (N_647,In_1446,In_280);
nand U648 (N_648,In_130,In_826);
and U649 (N_649,In_236,In_685);
or U650 (N_650,In_929,In_1299);
nor U651 (N_651,In_1155,In_1474);
and U652 (N_652,In_1004,In_334);
or U653 (N_653,In_617,In_431);
or U654 (N_654,In_941,In_936);
and U655 (N_655,In_88,In_1389);
nand U656 (N_656,In_1183,In_1302);
xor U657 (N_657,In_684,In_346);
nand U658 (N_658,In_1125,In_1071);
nand U659 (N_659,In_595,In_276);
or U660 (N_660,In_1420,In_1493);
xnor U661 (N_661,In_1409,In_1328);
nand U662 (N_662,In_746,In_955);
or U663 (N_663,In_1053,In_335);
and U664 (N_664,In_1198,In_263);
xnor U665 (N_665,In_683,In_141);
xnor U666 (N_666,In_455,In_798);
or U667 (N_667,In_103,In_281);
and U668 (N_668,In_65,In_1126);
xnor U669 (N_669,In_550,In_90);
and U670 (N_670,In_1045,In_899);
and U671 (N_671,In_1438,In_743);
xor U672 (N_672,In_49,In_1311);
and U673 (N_673,In_1129,In_347);
nor U674 (N_674,In_1477,In_1007);
nand U675 (N_675,In_1498,In_176);
and U676 (N_676,In_1247,In_187);
xor U677 (N_677,In_1386,In_1394);
or U678 (N_678,In_279,In_184);
xnor U679 (N_679,In_1235,In_612);
nand U680 (N_680,In_361,In_1002);
nor U681 (N_681,In_650,In_1164);
nor U682 (N_682,In_310,In_845);
or U683 (N_683,In_681,In_1195);
and U684 (N_684,In_31,In_698);
xnor U685 (N_685,In_725,In_765);
and U686 (N_686,In_157,In_708);
and U687 (N_687,In_781,In_1295);
and U688 (N_688,In_1082,In_1030);
xnor U689 (N_689,In_602,In_92);
nor U690 (N_690,In_436,In_1388);
xor U691 (N_691,In_1451,In_345);
nand U692 (N_692,In_241,In_695);
and U693 (N_693,In_214,In_1246);
or U694 (N_694,In_341,In_468);
nand U695 (N_695,In_952,In_814);
nor U696 (N_696,In_960,In_1473);
and U697 (N_697,In_656,In_1069);
xnor U698 (N_698,In_713,In_530);
nor U699 (N_699,In_817,In_160);
or U700 (N_700,In_731,In_1189);
and U701 (N_701,In_1046,In_1076);
and U702 (N_702,In_855,In_1398);
nor U703 (N_703,In_1158,In_752);
nand U704 (N_704,In_22,In_1422);
or U705 (N_705,In_1276,In_509);
nor U706 (N_706,In_1026,In_356);
and U707 (N_707,In_8,In_444);
nand U708 (N_708,In_106,In_124);
nor U709 (N_709,In_545,In_297);
or U710 (N_710,In_760,In_990);
and U711 (N_711,In_189,In_1073);
nor U712 (N_712,In_1379,In_1383);
and U713 (N_713,In_1478,In_1315);
or U714 (N_714,In_838,In_1307);
xor U715 (N_715,In_634,In_763);
nand U716 (N_716,In_1270,In_596);
nor U717 (N_717,In_247,In_217);
xor U718 (N_718,In_1208,In_528);
and U719 (N_719,In_1317,In_1240);
nor U720 (N_720,In_406,In_220);
nor U721 (N_721,In_181,In_1184);
or U722 (N_722,In_213,In_351);
nor U723 (N_723,In_1377,In_799);
xor U724 (N_724,In_1330,In_559);
nor U725 (N_725,In_1174,In_309);
xor U726 (N_726,In_427,In_1290);
xor U727 (N_727,In_728,In_1098);
or U728 (N_728,In_918,In_462);
xnor U729 (N_729,In_146,In_492);
nand U730 (N_730,In_216,In_736);
and U731 (N_731,In_795,In_1013);
or U732 (N_732,In_403,In_1392);
nand U733 (N_733,In_788,In_866);
or U734 (N_734,In_424,In_1248);
nand U735 (N_735,In_1461,In_158);
nand U736 (N_736,In_193,In_1100);
or U737 (N_737,In_823,In_964);
nor U738 (N_738,In_1021,In_488);
or U739 (N_739,In_1320,In_784);
nand U740 (N_740,In_206,In_391);
nand U741 (N_741,In_1188,In_1119);
nand U742 (N_742,In_235,In_907);
and U743 (N_743,In_1050,In_790);
or U744 (N_744,In_871,In_830);
nand U745 (N_745,In_239,In_519);
nor U746 (N_746,In_1056,In_593);
or U747 (N_747,In_1318,In_483);
nor U748 (N_748,In_501,In_98);
nand U749 (N_749,In_706,In_986);
xnor U750 (N_750,In_230,In_1116);
and U751 (N_751,In_804,In_1326);
nor U752 (N_752,In_562,In_1373);
or U753 (N_753,In_1080,In_1002);
xor U754 (N_754,In_723,In_1182);
and U755 (N_755,In_240,In_491);
nor U756 (N_756,In_584,In_219);
nor U757 (N_757,In_1057,In_1086);
and U758 (N_758,In_1433,In_146);
nor U759 (N_759,In_1123,In_1049);
and U760 (N_760,In_441,In_563);
and U761 (N_761,In_736,In_352);
nand U762 (N_762,In_396,In_783);
nor U763 (N_763,In_806,In_634);
and U764 (N_764,In_1247,In_0);
or U765 (N_765,In_112,In_1070);
nand U766 (N_766,In_1146,In_110);
and U767 (N_767,In_950,In_457);
nor U768 (N_768,In_1395,In_577);
or U769 (N_769,In_135,In_1353);
nand U770 (N_770,In_1358,In_709);
or U771 (N_771,In_383,In_279);
nor U772 (N_772,In_812,In_508);
and U773 (N_773,In_835,In_1422);
or U774 (N_774,In_385,In_894);
xnor U775 (N_775,In_334,In_1090);
or U776 (N_776,In_599,In_1007);
or U777 (N_777,In_1005,In_615);
nor U778 (N_778,In_331,In_1290);
nand U779 (N_779,In_1183,In_1008);
or U780 (N_780,In_673,In_775);
or U781 (N_781,In_1433,In_209);
and U782 (N_782,In_924,In_738);
xor U783 (N_783,In_1354,In_984);
and U784 (N_784,In_1490,In_54);
xnor U785 (N_785,In_353,In_607);
or U786 (N_786,In_479,In_6);
nor U787 (N_787,In_528,In_25);
nand U788 (N_788,In_534,In_324);
nor U789 (N_789,In_894,In_366);
and U790 (N_790,In_390,In_504);
or U791 (N_791,In_6,In_1419);
or U792 (N_792,In_1128,In_705);
or U793 (N_793,In_1024,In_964);
nor U794 (N_794,In_319,In_489);
or U795 (N_795,In_255,In_1416);
nor U796 (N_796,In_1071,In_1277);
or U797 (N_797,In_882,In_827);
and U798 (N_798,In_468,In_498);
nand U799 (N_799,In_86,In_349);
or U800 (N_800,In_468,In_892);
nand U801 (N_801,In_187,In_1058);
or U802 (N_802,In_586,In_153);
nor U803 (N_803,In_87,In_105);
xnor U804 (N_804,In_1480,In_375);
and U805 (N_805,In_515,In_131);
xor U806 (N_806,In_58,In_1389);
xnor U807 (N_807,In_1388,In_526);
and U808 (N_808,In_1171,In_1335);
nand U809 (N_809,In_98,In_490);
nand U810 (N_810,In_88,In_432);
nor U811 (N_811,In_280,In_1066);
or U812 (N_812,In_1334,In_1460);
nor U813 (N_813,In_431,In_1025);
and U814 (N_814,In_682,In_1120);
and U815 (N_815,In_872,In_151);
and U816 (N_816,In_1394,In_186);
nor U817 (N_817,In_621,In_1390);
or U818 (N_818,In_241,In_1387);
or U819 (N_819,In_625,In_1250);
nand U820 (N_820,In_316,In_265);
xor U821 (N_821,In_184,In_914);
nand U822 (N_822,In_1277,In_224);
xnor U823 (N_823,In_418,In_1331);
or U824 (N_824,In_1091,In_1432);
nand U825 (N_825,In_806,In_1279);
nor U826 (N_826,In_1154,In_1005);
nand U827 (N_827,In_1146,In_575);
and U828 (N_828,In_756,In_72);
xor U829 (N_829,In_56,In_114);
nand U830 (N_830,In_953,In_845);
and U831 (N_831,In_1218,In_46);
or U832 (N_832,In_713,In_56);
nand U833 (N_833,In_1310,In_1038);
nand U834 (N_834,In_618,In_695);
xor U835 (N_835,In_751,In_118);
nor U836 (N_836,In_1478,In_865);
nor U837 (N_837,In_1294,In_684);
and U838 (N_838,In_1070,In_800);
nand U839 (N_839,In_1449,In_1441);
xor U840 (N_840,In_655,In_1182);
nor U841 (N_841,In_1234,In_1398);
nor U842 (N_842,In_670,In_1407);
xnor U843 (N_843,In_1236,In_885);
xnor U844 (N_844,In_522,In_144);
nor U845 (N_845,In_222,In_1123);
or U846 (N_846,In_61,In_1164);
nor U847 (N_847,In_681,In_1038);
nor U848 (N_848,In_175,In_1455);
xnor U849 (N_849,In_1126,In_31);
or U850 (N_850,In_1333,In_759);
xnor U851 (N_851,In_436,In_539);
nand U852 (N_852,In_93,In_888);
xor U853 (N_853,In_1295,In_923);
and U854 (N_854,In_1318,In_1116);
or U855 (N_855,In_265,In_744);
xnor U856 (N_856,In_74,In_299);
xnor U857 (N_857,In_1346,In_407);
xor U858 (N_858,In_1308,In_1349);
nor U859 (N_859,In_335,In_767);
and U860 (N_860,In_535,In_650);
nor U861 (N_861,In_762,In_1095);
or U862 (N_862,In_212,In_653);
or U863 (N_863,In_946,In_1225);
or U864 (N_864,In_1005,In_684);
and U865 (N_865,In_83,In_551);
xor U866 (N_866,In_62,In_260);
or U867 (N_867,In_1311,In_909);
nand U868 (N_868,In_1234,In_239);
nor U869 (N_869,In_978,In_663);
and U870 (N_870,In_306,In_566);
nand U871 (N_871,In_1067,In_537);
or U872 (N_872,In_1340,In_416);
and U873 (N_873,In_198,In_1089);
nor U874 (N_874,In_1371,In_484);
nor U875 (N_875,In_1379,In_584);
or U876 (N_876,In_524,In_134);
nand U877 (N_877,In_789,In_8);
and U878 (N_878,In_1078,In_1464);
nor U879 (N_879,In_201,In_138);
and U880 (N_880,In_1485,In_1487);
or U881 (N_881,In_1215,In_982);
nand U882 (N_882,In_1437,In_1332);
nand U883 (N_883,In_859,In_363);
nor U884 (N_884,In_516,In_609);
and U885 (N_885,In_739,In_585);
or U886 (N_886,In_208,In_1388);
nor U887 (N_887,In_1463,In_275);
nor U888 (N_888,In_1069,In_176);
or U889 (N_889,In_297,In_4);
or U890 (N_890,In_1142,In_74);
and U891 (N_891,In_209,In_583);
nor U892 (N_892,In_719,In_131);
or U893 (N_893,In_72,In_503);
nor U894 (N_894,In_342,In_305);
nand U895 (N_895,In_1005,In_1072);
or U896 (N_896,In_17,In_1096);
or U897 (N_897,In_853,In_1345);
and U898 (N_898,In_831,In_1117);
nand U899 (N_899,In_943,In_307);
or U900 (N_900,In_1334,In_247);
nand U901 (N_901,In_660,In_570);
nor U902 (N_902,In_223,In_1370);
xnor U903 (N_903,In_378,In_1345);
or U904 (N_904,In_287,In_1364);
xor U905 (N_905,In_1033,In_170);
and U906 (N_906,In_1150,In_419);
and U907 (N_907,In_704,In_523);
or U908 (N_908,In_1231,In_890);
nor U909 (N_909,In_1195,In_773);
nor U910 (N_910,In_1069,In_608);
xnor U911 (N_911,In_1164,In_260);
nor U912 (N_912,In_218,In_1010);
nor U913 (N_913,In_737,In_851);
or U914 (N_914,In_709,In_365);
and U915 (N_915,In_656,In_1286);
nand U916 (N_916,In_599,In_1246);
and U917 (N_917,In_53,In_1056);
and U918 (N_918,In_56,In_936);
nor U919 (N_919,In_1028,In_509);
nor U920 (N_920,In_995,In_1029);
xnor U921 (N_921,In_1168,In_1044);
or U922 (N_922,In_428,In_1499);
and U923 (N_923,In_40,In_935);
or U924 (N_924,In_95,In_55);
nand U925 (N_925,In_1384,In_242);
nand U926 (N_926,In_1055,In_499);
and U927 (N_927,In_851,In_866);
nand U928 (N_928,In_427,In_233);
or U929 (N_929,In_626,In_1307);
and U930 (N_930,In_931,In_1280);
or U931 (N_931,In_1243,In_231);
and U932 (N_932,In_557,In_370);
nand U933 (N_933,In_1004,In_985);
and U934 (N_934,In_619,In_1078);
nand U935 (N_935,In_689,In_233);
nand U936 (N_936,In_472,In_540);
or U937 (N_937,In_1321,In_421);
nor U938 (N_938,In_279,In_485);
or U939 (N_939,In_757,In_1253);
or U940 (N_940,In_439,In_942);
or U941 (N_941,In_884,In_982);
or U942 (N_942,In_677,In_44);
or U943 (N_943,In_838,In_1116);
xnor U944 (N_944,In_461,In_247);
nor U945 (N_945,In_382,In_278);
nand U946 (N_946,In_208,In_703);
xor U947 (N_947,In_211,In_859);
nand U948 (N_948,In_669,In_77);
or U949 (N_949,In_866,In_571);
nor U950 (N_950,In_1462,In_192);
nor U951 (N_951,In_797,In_374);
nor U952 (N_952,In_907,In_1270);
and U953 (N_953,In_85,In_474);
nand U954 (N_954,In_626,In_9);
nand U955 (N_955,In_711,In_238);
nor U956 (N_956,In_493,In_1187);
and U957 (N_957,In_314,In_1148);
nand U958 (N_958,In_68,In_143);
nor U959 (N_959,In_337,In_48);
nand U960 (N_960,In_442,In_1252);
and U961 (N_961,In_319,In_1369);
xor U962 (N_962,In_570,In_1364);
and U963 (N_963,In_473,In_1007);
xor U964 (N_964,In_350,In_1213);
nand U965 (N_965,In_7,In_477);
and U966 (N_966,In_375,In_949);
nand U967 (N_967,In_345,In_262);
nor U968 (N_968,In_97,In_730);
and U969 (N_969,In_391,In_172);
and U970 (N_970,In_1443,In_1017);
nor U971 (N_971,In_42,In_996);
nand U972 (N_972,In_1327,In_1161);
xor U973 (N_973,In_475,In_735);
nor U974 (N_974,In_660,In_1053);
and U975 (N_975,In_575,In_523);
nand U976 (N_976,In_1344,In_619);
nand U977 (N_977,In_1115,In_1141);
or U978 (N_978,In_529,In_750);
nand U979 (N_979,In_487,In_1076);
xor U980 (N_980,In_1069,In_735);
nor U981 (N_981,In_350,In_1365);
and U982 (N_982,In_1081,In_278);
xor U983 (N_983,In_1075,In_620);
nand U984 (N_984,In_1280,In_981);
nor U985 (N_985,In_107,In_1051);
nand U986 (N_986,In_885,In_1036);
xor U987 (N_987,In_639,In_672);
and U988 (N_988,In_1222,In_285);
nand U989 (N_989,In_703,In_280);
xnor U990 (N_990,In_1034,In_1140);
and U991 (N_991,In_45,In_561);
nor U992 (N_992,In_1013,In_1480);
and U993 (N_993,In_1263,In_1441);
nor U994 (N_994,In_314,In_279);
nor U995 (N_995,In_1075,In_435);
and U996 (N_996,In_193,In_647);
and U997 (N_997,In_794,In_1435);
and U998 (N_998,In_1348,In_696);
nor U999 (N_999,In_387,In_585);
and U1000 (N_1000,N_266,N_313);
xor U1001 (N_1001,N_850,N_440);
or U1002 (N_1002,N_265,N_445);
and U1003 (N_1003,N_388,N_281);
xor U1004 (N_1004,N_561,N_237);
and U1005 (N_1005,N_157,N_24);
xor U1006 (N_1006,N_420,N_697);
and U1007 (N_1007,N_733,N_162);
and U1008 (N_1008,N_206,N_377);
xnor U1009 (N_1009,N_438,N_400);
and U1010 (N_1010,N_36,N_169);
xnor U1011 (N_1011,N_855,N_120);
and U1012 (N_1012,N_607,N_17);
and U1013 (N_1013,N_702,N_522);
or U1014 (N_1014,N_890,N_614);
xor U1015 (N_1015,N_884,N_27);
nor U1016 (N_1016,N_182,N_340);
and U1017 (N_1017,N_798,N_109);
nand U1018 (N_1018,N_19,N_306);
and U1019 (N_1019,N_970,N_544);
and U1020 (N_1020,N_200,N_848);
nand U1021 (N_1021,N_465,N_564);
nand U1022 (N_1022,N_512,N_367);
xnor U1023 (N_1023,N_565,N_920);
nand U1024 (N_1024,N_339,N_108);
and U1025 (N_1025,N_251,N_156);
nand U1026 (N_1026,N_241,N_669);
nor U1027 (N_1027,N_292,N_310);
nand U1028 (N_1028,N_750,N_551);
xnor U1029 (N_1029,N_977,N_463);
xnor U1030 (N_1030,N_272,N_989);
and U1031 (N_1031,N_662,N_815);
nand U1032 (N_1032,N_436,N_449);
nor U1033 (N_1033,N_26,N_100);
and U1034 (N_1034,N_70,N_466);
xor U1035 (N_1035,N_208,N_913);
nand U1036 (N_1036,N_394,N_350);
nor U1037 (N_1037,N_950,N_974);
or U1038 (N_1038,N_124,N_742);
nand U1039 (N_1039,N_902,N_164);
nand U1040 (N_1040,N_82,N_282);
xor U1041 (N_1041,N_193,N_961);
nor U1042 (N_1042,N_195,N_378);
nand U1043 (N_1043,N_907,N_773);
nand U1044 (N_1044,N_389,N_938);
nand U1045 (N_1045,N_321,N_98);
nor U1046 (N_1046,N_633,N_588);
xnor U1047 (N_1047,N_179,N_579);
or U1048 (N_1048,N_910,N_152);
or U1049 (N_1049,N_427,N_705);
xnor U1050 (N_1050,N_572,N_991);
nor U1051 (N_1051,N_868,N_460);
nand U1052 (N_1052,N_520,N_804);
xor U1053 (N_1053,N_117,N_694);
nand U1054 (N_1054,N_771,N_239);
and U1055 (N_1055,N_777,N_791);
or U1056 (N_1056,N_379,N_918);
xnor U1057 (N_1057,N_550,N_63);
xnor U1058 (N_1058,N_895,N_186);
nor U1059 (N_1059,N_140,N_879);
and U1060 (N_1060,N_28,N_844);
or U1061 (N_1061,N_46,N_188);
or U1062 (N_1062,N_255,N_976);
and U1063 (N_1063,N_91,N_232);
and U1064 (N_1064,N_178,N_358);
nor U1065 (N_1065,N_660,N_13);
or U1066 (N_1066,N_691,N_990);
nand U1067 (N_1067,N_885,N_993);
nor U1068 (N_1068,N_782,N_801);
nand U1069 (N_1069,N_995,N_318);
xnor U1070 (N_1070,N_270,N_31);
nand U1071 (N_1071,N_403,N_645);
xnor U1072 (N_1072,N_227,N_606);
and U1073 (N_1073,N_137,N_897);
or U1074 (N_1074,N_754,N_617);
and U1075 (N_1075,N_308,N_37);
nor U1076 (N_1076,N_395,N_861);
and U1077 (N_1077,N_570,N_542);
or U1078 (N_1078,N_558,N_821);
nor U1079 (N_1079,N_635,N_627);
or U1080 (N_1080,N_61,N_332);
nand U1081 (N_1081,N_877,N_757);
nor U1082 (N_1082,N_826,N_829);
and U1083 (N_1083,N_881,N_221);
xnor U1084 (N_1084,N_835,N_327);
nand U1085 (N_1085,N_153,N_53);
nor U1086 (N_1086,N_215,N_293);
or U1087 (N_1087,N_923,N_426);
xor U1088 (N_1088,N_904,N_811);
nand U1089 (N_1089,N_537,N_611);
or U1090 (N_1090,N_368,N_830);
and U1091 (N_1091,N_837,N_706);
nand U1092 (N_1092,N_207,N_498);
nor U1093 (N_1093,N_184,N_62);
xnor U1094 (N_1094,N_887,N_381);
nand U1095 (N_1095,N_354,N_613);
or U1096 (N_1096,N_925,N_50);
and U1097 (N_1097,N_390,N_841);
nand U1098 (N_1098,N_119,N_9);
nand U1099 (N_1099,N_183,N_736);
nor U1100 (N_1100,N_129,N_434);
xor U1101 (N_1101,N_851,N_446);
xnor U1102 (N_1102,N_527,N_4);
nand U1103 (N_1103,N_344,N_245);
xor U1104 (N_1104,N_431,N_181);
or U1105 (N_1105,N_235,N_787);
nor U1106 (N_1106,N_934,N_889);
or U1107 (N_1107,N_765,N_911);
and U1108 (N_1108,N_796,N_16);
or U1109 (N_1109,N_853,N_719);
xor U1110 (N_1110,N_328,N_842);
nand U1111 (N_1111,N_761,N_2);
xnor U1112 (N_1112,N_286,N_59);
xnor U1113 (N_1113,N_22,N_205);
xnor U1114 (N_1114,N_203,N_809);
or U1115 (N_1115,N_198,N_102);
nor U1116 (N_1116,N_975,N_644);
or U1117 (N_1117,N_875,N_894);
or U1118 (N_1118,N_172,N_979);
nor U1119 (N_1119,N_778,N_472);
or U1120 (N_1120,N_985,N_593);
nor U1121 (N_1121,N_30,N_210);
and U1122 (N_1122,N_836,N_219);
nor U1123 (N_1123,N_248,N_847);
or U1124 (N_1124,N_309,N_770);
and U1125 (N_1125,N_684,N_277);
or U1126 (N_1126,N_74,N_196);
nor U1127 (N_1127,N_418,N_479);
or U1128 (N_1128,N_271,N_682);
xnor U1129 (N_1129,N_679,N_280);
or U1130 (N_1130,N_173,N_238);
nor U1131 (N_1131,N_538,N_903);
or U1132 (N_1132,N_408,N_322);
or U1133 (N_1133,N_988,N_176);
xor U1134 (N_1134,N_663,N_111);
and U1135 (N_1135,N_526,N_118);
nor U1136 (N_1136,N_678,N_780);
and U1137 (N_1137,N_387,N_450);
nor U1138 (N_1138,N_715,N_941);
nor U1139 (N_1139,N_489,N_501);
or U1140 (N_1140,N_139,N_680);
and U1141 (N_1141,N_797,N_529);
or U1142 (N_1142,N_171,N_949);
xnor U1143 (N_1143,N_89,N_159);
or U1144 (N_1144,N_452,N_738);
and U1145 (N_1145,N_566,N_269);
or U1146 (N_1146,N_352,N_581);
xor U1147 (N_1147,N_838,N_739);
or U1148 (N_1148,N_447,N_957);
nor U1149 (N_1149,N_900,N_155);
and U1150 (N_1150,N_189,N_643);
nand U1151 (N_1151,N_143,N_901);
nor U1152 (N_1152,N_960,N_756);
and U1153 (N_1153,N_363,N_414);
nor U1154 (N_1154,N_568,N_375);
and U1155 (N_1155,N_559,N_672);
and U1156 (N_1156,N_486,N_421);
nor U1157 (N_1157,N_982,N_752);
xnor U1158 (N_1158,N_928,N_681);
and U1159 (N_1159,N_927,N_469);
nand U1160 (N_1160,N_213,N_315);
and U1161 (N_1161,N_790,N_312);
nand U1162 (N_1162,N_25,N_576);
nand U1163 (N_1163,N_299,N_583);
and U1164 (N_1164,N_734,N_393);
nand U1165 (N_1165,N_290,N_29);
or U1166 (N_1166,N_912,N_823);
and U1167 (N_1167,N_492,N_260);
nand U1168 (N_1168,N_698,N_197);
and U1169 (N_1169,N_940,N_513);
xor U1170 (N_1170,N_168,N_759);
nor U1171 (N_1171,N_355,N_464);
nor U1172 (N_1172,N_35,N_864);
nor U1173 (N_1173,N_236,N_657);
or U1174 (N_1174,N_185,N_824);
or U1175 (N_1175,N_926,N_401);
and U1176 (N_1176,N_969,N_749);
xor U1177 (N_1177,N_630,N_582);
nor U1178 (N_1178,N_710,N_998);
and U1179 (N_1179,N_839,N_86);
and U1180 (N_1180,N_362,N_936);
and U1181 (N_1181,N_14,N_685);
or U1182 (N_1182,N_714,N_64);
or U1183 (N_1183,N_433,N_649);
nand U1184 (N_1184,N_603,N_632);
nand U1185 (N_1185,N_495,N_812);
nand U1186 (N_1186,N_488,N_626);
and U1187 (N_1187,N_654,N_474);
nand U1188 (N_1188,N_870,N_202);
nor U1189 (N_1189,N_744,N_814);
xor U1190 (N_1190,N_786,N_921);
nand U1191 (N_1191,N_231,N_43);
or U1192 (N_1192,N_783,N_718);
nor U1193 (N_1193,N_240,N_964);
nor U1194 (N_1194,N_667,N_924);
nor U1195 (N_1195,N_1,N_799);
nor U1196 (N_1196,N_351,N_605);
nor U1197 (N_1197,N_298,N_955);
or U1198 (N_1198,N_822,N_406);
and U1199 (N_1199,N_932,N_741);
nand U1200 (N_1200,N_141,N_775);
nand U1201 (N_1201,N_737,N_211);
nor U1202 (N_1202,N_437,N_647);
nand U1203 (N_1203,N_573,N_547);
or U1204 (N_1204,N_45,N_999);
or U1205 (N_1205,N_865,N_873);
nand U1206 (N_1206,N_106,N_914);
nor U1207 (N_1207,N_301,N_404);
or U1208 (N_1208,N_937,N_968);
and U1209 (N_1209,N_3,N_813);
xor U1210 (N_1210,N_48,N_589);
or U1211 (N_1211,N_233,N_220);
nor U1212 (N_1212,N_166,N_5);
nand U1213 (N_1213,N_112,N_668);
nor U1214 (N_1214,N_768,N_349);
nor U1215 (N_1215,N_341,N_661);
nor U1216 (N_1216,N_674,N_66);
nand U1217 (N_1217,N_478,N_508);
xor U1218 (N_1218,N_410,N_229);
nand U1219 (N_1219,N_631,N_323);
or U1220 (N_1220,N_507,N_735);
nor U1221 (N_1221,N_333,N_781);
nor U1222 (N_1222,N_8,N_874);
nor U1223 (N_1223,N_345,N_133);
nand U1224 (N_1224,N_546,N_963);
nor U1225 (N_1225,N_10,N_732);
nor U1226 (N_1226,N_85,N_296);
nand U1227 (N_1227,N_514,N_125);
or U1228 (N_1228,N_800,N_67);
or U1229 (N_1229,N_994,N_658);
nand U1230 (N_1230,N_32,N_721);
or U1231 (N_1231,N_348,N_533);
xnor U1232 (N_1232,N_521,N_655);
nand U1233 (N_1233,N_114,N_575);
and U1234 (N_1234,N_857,N_121);
or U1235 (N_1235,N_97,N_33);
nor U1236 (N_1236,N_257,N_451);
and U1237 (N_1237,N_675,N_729);
or U1238 (N_1238,N_412,N_476);
or U1239 (N_1239,N_524,N_56);
or U1240 (N_1240,N_223,N_893);
nand U1241 (N_1241,N_872,N_840);
nand U1242 (N_1242,N_453,N_996);
xnor U1243 (N_1243,N_316,N_723);
or U1244 (N_1244,N_543,N_399);
or U1245 (N_1245,N_984,N_898);
nand U1246 (N_1246,N_148,N_651);
and U1247 (N_1247,N_78,N_247);
nand U1248 (N_1248,N_578,N_549);
and U1249 (N_1249,N_218,N_856);
and U1250 (N_1250,N_413,N_99);
or U1251 (N_1251,N_65,N_134);
xor U1252 (N_1252,N_769,N_625);
and U1253 (N_1253,N_105,N_860);
and U1254 (N_1254,N_515,N_665);
nand U1255 (N_1255,N_353,N_191);
nand U1256 (N_1256,N_49,N_131);
nand U1257 (N_1257,N_428,N_242);
xnor U1258 (N_1258,N_642,N_429);
xor U1259 (N_1259,N_256,N_361);
and U1260 (N_1260,N_51,N_448);
nand U1261 (N_1261,N_320,N_136);
and U1262 (N_1262,N_335,N_487);
nand U1263 (N_1263,N_300,N_326);
xor U1264 (N_1264,N_187,N_371);
or U1265 (N_1265,N_845,N_808);
nand U1266 (N_1266,N_194,N_90);
nand U1267 (N_1267,N_424,N_594);
or U1268 (N_1268,N_454,N_832);
nor U1269 (N_1269,N_528,N_986);
xor U1270 (N_1270,N_192,N_38);
nor U1271 (N_1271,N_494,N_916);
nor U1272 (N_1272,N_405,N_283);
or U1273 (N_1273,N_666,N_959);
or U1274 (N_1274,N_273,N_289);
or U1275 (N_1275,N_711,N_810);
or U1276 (N_1276,N_422,N_288);
nor U1277 (N_1277,N_122,N_442);
nand U1278 (N_1278,N_596,N_652);
and U1279 (N_1279,N_638,N_621);
and U1280 (N_1280,N_212,N_577);
and U1281 (N_1281,N_688,N_262);
xnor U1282 (N_1282,N_276,N_6);
or U1283 (N_1283,N_356,N_693);
nand U1284 (N_1284,N_336,N_939);
and U1285 (N_1285,N_539,N_158);
and U1286 (N_1286,N_556,N_639);
nor U1287 (N_1287,N_407,N_699);
or U1288 (N_1288,N_915,N_641);
nor U1289 (N_1289,N_149,N_965);
nand U1290 (N_1290,N_720,N_724);
nand U1291 (N_1291,N_967,N_461);
nand U1292 (N_1292,N_180,N_480);
nand U1293 (N_1293,N_966,N_73);
and U1294 (N_1294,N_252,N_497);
or U1295 (N_1295,N_767,N_34);
and U1296 (N_1296,N_789,N_945);
or U1297 (N_1297,N_689,N_250);
and U1298 (N_1298,N_52,N_331);
nor U1299 (N_1299,N_519,N_0);
nor U1300 (N_1300,N_792,N_946);
nand U1301 (N_1301,N_415,N_818);
nor U1302 (N_1302,N_444,N_858);
xnor U1303 (N_1303,N_468,N_712);
nor U1304 (N_1304,N_859,N_372);
xnor U1305 (N_1305,N_511,N_295);
or U1306 (N_1306,N_287,N_337);
or U1307 (N_1307,N_816,N_84);
nor U1308 (N_1308,N_228,N_294);
and U1309 (N_1309,N_615,N_243);
nor U1310 (N_1310,N_888,N_398);
nand U1311 (N_1311,N_828,N_703);
and U1312 (N_1312,N_716,N_972);
or U1313 (N_1313,N_640,N_555);
and U1314 (N_1314,N_766,N_366);
nand U1315 (N_1315,N_762,N_81);
nand U1316 (N_1316,N_929,N_500);
nand U1317 (N_1317,N_676,N_755);
or U1318 (N_1318,N_75,N_740);
nor U1319 (N_1319,N_284,N_935);
nand U1320 (N_1320,N_96,N_677);
and U1321 (N_1321,N_785,N_704);
nor U1322 (N_1322,N_443,N_883);
or U1323 (N_1323,N_541,N_268);
xor U1324 (N_1324,N_933,N_425);
nand U1325 (N_1325,N_833,N_113);
xnor U1326 (N_1326,N_653,N_943);
nor U1327 (N_1327,N_40,N_899);
and U1328 (N_1328,N_160,N_60);
nor U1329 (N_1329,N_584,N_458);
xnor U1330 (N_1330,N_628,N_346);
nor U1331 (N_1331,N_76,N_216);
nand U1332 (N_1332,N_731,N_609);
nand U1333 (N_1333,N_509,N_760);
nor U1334 (N_1334,N_909,N_462);
and U1335 (N_1335,N_285,N_825);
nand U1336 (N_1336,N_382,N_138);
nor U1337 (N_1337,N_263,N_499);
xnor U1338 (N_1338,N_93,N_88);
xnor U1339 (N_1339,N_562,N_545);
nor U1340 (N_1340,N_128,N_886);
or U1341 (N_1341,N_330,N_535);
xnor U1342 (N_1342,N_673,N_973);
nand U1343 (N_1343,N_254,N_696);
xor U1344 (N_1344,N_360,N_147);
or U1345 (N_1345,N_142,N_68);
nand U1346 (N_1346,N_167,N_12);
xor U1347 (N_1347,N_634,N_214);
xor U1348 (N_1348,N_905,N_163);
xor U1349 (N_1349,N_278,N_717);
nand U1350 (N_1350,N_144,N_636);
nand U1351 (N_1351,N_803,N_230);
or U1352 (N_1352,N_774,N_574);
nor U1353 (N_1353,N_587,N_264);
xnor U1354 (N_1354,N_779,N_484);
nor U1355 (N_1355,N_103,N_843);
xnor U1356 (N_1356,N_386,N_80);
xnor U1357 (N_1357,N_342,N_601);
and U1358 (N_1358,N_600,N_906);
or U1359 (N_1359,N_314,N_931);
or U1360 (N_1360,N_987,N_58);
xor U1361 (N_1361,N_225,N_18);
nor U1362 (N_1362,N_126,N_204);
nand U1363 (N_1363,N_146,N_145);
and U1364 (N_1364,N_954,N_701);
or U1365 (N_1365,N_548,N_21);
and U1366 (N_1366,N_980,N_629);
nor U1367 (N_1367,N_127,N_599);
nand U1368 (N_1368,N_540,N_908);
xor U1369 (N_1369,N_457,N_523);
or U1370 (N_1370,N_592,N_170);
xor U1371 (N_1371,N_319,N_485);
and U1372 (N_1372,N_534,N_477);
nand U1373 (N_1373,N_880,N_585);
xnor U1374 (N_1374,N_569,N_567);
and U1375 (N_1375,N_92,N_258);
nor U1376 (N_1376,N_831,N_608);
and U1377 (N_1377,N_116,N_686);
or U1378 (N_1378,N_597,N_303);
or U1379 (N_1379,N_123,N_307);
and U1380 (N_1380,N_467,N_338);
or U1381 (N_1381,N_659,N_151);
and U1382 (N_1382,N_619,N_610);
and U1383 (N_1383,N_878,N_552);
or U1384 (N_1384,N_23,N_304);
and U1385 (N_1385,N_275,N_867);
nor U1386 (N_1386,N_317,N_199);
xnor U1387 (N_1387,N_951,N_805);
and U1388 (N_1388,N_764,N_94);
and U1389 (N_1389,N_150,N_11);
xor U1390 (N_1390,N_505,N_590);
nand U1391 (N_1391,N_776,N_598);
xor U1392 (N_1392,N_795,N_637);
nor U1393 (N_1393,N_802,N_201);
xnor U1394 (N_1394,N_224,N_591);
xnor U1395 (N_1395,N_325,N_646);
xor U1396 (N_1396,N_869,N_42);
nand U1397 (N_1397,N_305,N_919);
nand U1398 (N_1398,N_671,N_396);
nor U1399 (N_1399,N_7,N_948);
nand U1400 (N_1400,N_69,N_846);
nor U1401 (N_1401,N_525,N_553);
and U1402 (N_1402,N_435,N_624);
nand U1403 (N_1403,N_324,N_560);
nand U1404 (N_1404,N_730,N_922);
and U1405 (N_1405,N_725,N_419);
or U1406 (N_1406,N_690,N_311);
and U1407 (N_1407,N_77,N_374);
nor U1408 (N_1408,N_110,N_246);
nor U1409 (N_1409,N_482,N_602);
nand U1410 (N_1410,N_47,N_820);
nor U1411 (N_1411,N_506,N_863);
and U1412 (N_1412,N_57,N_683);
or U1413 (N_1413,N_370,N_15);
or U1414 (N_1414,N_473,N_347);
xnor U1415 (N_1415,N_135,N_174);
xor U1416 (N_1416,N_397,N_384);
or U1417 (N_1417,N_177,N_978);
or U1418 (N_1418,N_481,N_334);
xor U1419 (N_1419,N_751,N_101);
and U1420 (N_1420,N_748,N_417);
or U1421 (N_1421,N_648,N_896);
and U1422 (N_1422,N_794,N_536);
xor U1423 (N_1423,N_154,N_373);
or U1424 (N_1424,N_962,N_743);
and U1425 (N_1425,N_83,N_259);
xor U1426 (N_1426,N_249,N_297);
xnor U1427 (N_1427,N_217,N_475);
and U1428 (N_1428,N_244,N_554);
or U1429 (N_1429,N_892,N_917);
or U1430 (N_1430,N_380,N_209);
nand U1431 (N_1431,N_793,N_483);
nand U1432 (N_1432,N_595,N_496);
or U1433 (N_1433,N_71,N_502);
xor U1434 (N_1434,N_518,N_226);
nand U1435 (N_1435,N_871,N_981);
xnor U1436 (N_1436,N_107,N_747);
nor U1437 (N_1437,N_490,N_854);
or U1438 (N_1438,N_95,N_728);
or U1439 (N_1439,N_175,N_456);
xor U1440 (N_1440,N_997,N_618);
and U1441 (N_1441,N_876,N_439);
nor U1442 (N_1442,N_707,N_953);
or U1443 (N_1443,N_132,N_491);
nor U1444 (N_1444,N_416,N_343);
and U1445 (N_1445,N_758,N_557);
nand U1446 (N_1446,N_623,N_687);
nand U1447 (N_1447,N_261,N_862);
or U1448 (N_1448,N_274,N_411);
nand U1449 (N_1449,N_20,N_402);
xnor U1450 (N_1450,N_942,N_722);
nor U1451 (N_1451,N_849,N_992);
and U1452 (N_1452,N_531,N_39);
and U1453 (N_1453,N_763,N_455);
nand U1454 (N_1454,N_891,N_604);
xor U1455 (N_1455,N_656,N_291);
nand U1456 (N_1456,N_385,N_616);
and U1457 (N_1457,N_586,N_392);
or U1458 (N_1458,N_504,N_563);
or U1459 (N_1459,N_620,N_234);
or U1460 (N_1460,N_708,N_470);
or U1461 (N_1461,N_930,N_516);
nor U1462 (N_1462,N_834,N_79);
and U1463 (N_1463,N_882,N_357);
nor U1464 (N_1464,N_819,N_788);
nand U1465 (N_1465,N_532,N_530);
xnor U1466 (N_1466,N_650,N_726);
and U1467 (N_1467,N_329,N_971);
and U1468 (N_1468,N_772,N_115);
nor U1469 (N_1469,N_44,N_41);
or U1470 (N_1470,N_423,N_302);
nor U1471 (N_1471,N_517,N_359);
and U1472 (N_1472,N_852,N_510);
nand U1473 (N_1473,N_709,N_104);
nand U1474 (N_1474,N_753,N_365);
xnor U1475 (N_1475,N_866,N_827);
xor U1476 (N_1476,N_459,N_253);
nor U1477 (N_1477,N_713,N_432);
nor U1478 (N_1478,N_222,N_692);
nor U1479 (N_1479,N_441,N_807);
or U1480 (N_1480,N_958,N_503);
nand U1481 (N_1481,N_72,N_409);
or U1482 (N_1482,N_87,N_54);
and U1483 (N_1483,N_383,N_430);
xnor U1484 (N_1484,N_55,N_983);
and U1485 (N_1485,N_817,N_279);
nor U1486 (N_1486,N_745,N_944);
or U1487 (N_1487,N_190,N_727);
nand U1488 (N_1488,N_471,N_391);
or U1489 (N_1489,N_952,N_622);
xor U1490 (N_1490,N_267,N_806);
xnor U1491 (N_1491,N_580,N_670);
and U1492 (N_1492,N_376,N_784);
and U1493 (N_1493,N_364,N_664);
and U1494 (N_1494,N_493,N_695);
nor U1495 (N_1495,N_161,N_369);
nor U1496 (N_1496,N_746,N_956);
or U1497 (N_1497,N_947,N_571);
nand U1498 (N_1498,N_165,N_130);
nand U1499 (N_1499,N_700,N_612);
xnor U1500 (N_1500,N_378,N_390);
xnor U1501 (N_1501,N_225,N_979);
and U1502 (N_1502,N_964,N_579);
nor U1503 (N_1503,N_155,N_88);
and U1504 (N_1504,N_679,N_400);
and U1505 (N_1505,N_317,N_440);
nand U1506 (N_1506,N_743,N_905);
and U1507 (N_1507,N_596,N_13);
nor U1508 (N_1508,N_656,N_961);
or U1509 (N_1509,N_835,N_73);
xor U1510 (N_1510,N_845,N_910);
nor U1511 (N_1511,N_606,N_955);
xor U1512 (N_1512,N_614,N_843);
xor U1513 (N_1513,N_873,N_465);
and U1514 (N_1514,N_975,N_518);
nand U1515 (N_1515,N_609,N_580);
xnor U1516 (N_1516,N_528,N_773);
and U1517 (N_1517,N_49,N_780);
nor U1518 (N_1518,N_669,N_747);
nor U1519 (N_1519,N_430,N_272);
xnor U1520 (N_1520,N_905,N_260);
xnor U1521 (N_1521,N_824,N_986);
or U1522 (N_1522,N_327,N_584);
or U1523 (N_1523,N_71,N_956);
and U1524 (N_1524,N_363,N_271);
xnor U1525 (N_1525,N_221,N_773);
nand U1526 (N_1526,N_954,N_722);
or U1527 (N_1527,N_732,N_911);
nand U1528 (N_1528,N_380,N_475);
nand U1529 (N_1529,N_818,N_85);
xnor U1530 (N_1530,N_181,N_987);
and U1531 (N_1531,N_54,N_653);
nor U1532 (N_1532,N_396,N_479);
nor U1533 (N_1533,N_273,N_641);
nor U1534 (N_1534,N_441,N_976);
nand U1535 (N_1535,N_428,N_278);
nor U1536 (N_1536,N_909,N_993);
nand U1537 (N_1537,N_361,N_105);
nand U1538 (N_1538,N_303,N_715);
and U1539 (N_1539,N_155,N_185);
nand U1540 (N_1540,N_644,N_773);
nand U1541 (N_1541,N_992,N_499);
nor U1542 (N_1542,N_433,N_2);
and U1543 (N_1543,N_642,N_240);
nand U1544 (N_1544,N_280,N_859);
and U1545 (N_1545,N_111,N_654);
xor U1546 (N_1546,N_651,N_307);
xor U1547 (N_1547,N_100,N_459);
nand U1548 (N_1548,N_173,N_593);
xnor U1549 (N_1549,N_536,N_651);
and U1550 (N_1550,N_350,N_567);
and U1551 (N_1551,N_314,N_865);
nand U1552 (N_1552,N_404,N_167);
nor U1553 (N_1553,N_775,N_424);
or U1554 (N_1554,N_37,N_393);
nand U1555 (N_1555,N_971,N_867);
or U1556 (N_1556,N_136,N_374);
xor U1557 (N_1557,N_201,N_221);
or U1558 (N_1558,N_582,N_426);
nand U1559 (N_1559,N_27,N_907);
nand U1560 (N_1560,N_248,N_912);
nor U1561 (N_1561,N_174,N_192);
xnor U1562 (N_1562,N_8,N_313);
and U1563 (N_1563,N_72,N_510);
nand U1564 (N_1564,N_750,N_173);
nand U1565 (N_1565,N_683,N_551);
and U1566 (N_1566,N_36,N_225);
nand U1567 (N_1567,N_293,N_391);
nand U1568 (N_1568,N_803,N_43);
nand U1569 (N_1569,N_858,N_658);
nor U1570 (N_1570,N_279,N_12);
nand U1571 (N_1571,N_142,N_72);
xnor U1572 (N_1572,N_709,N_845);
or U1573 (N_1573,N_885,N_727);
xor U1574 (N_1574,N_88,N_607);
xnor U1575 (N_1575,N_14,N_700);
nand U1576 (N_1576,N_824,N_401);
nand U1577 (N_1577,N_442,N_310);
and U1578 (N_1578,N_401,N_835);
and U1579 (N_1579,N_997,N_12);
and U1580 (N_1580,N_12,N_744);
nor U1581 (N_1581,N_443,N_589);
nand U1582 (N_1582,N_654,N_791);
nand U1583 (N_1583,N_588,N_246);
or U1584 (N_1584,N_176,N_560);
or U1585 (N_1585,N_539,N_333);
or U1586 (N_1586,N_562,N_300);
and U1587 (N_1587,N_511,N_542);
and U1588 (N_1588,N_282,N_339);
nor U1589 (N_1589,N_468,N_684);
nor U1590 (N_1590,N_20,N_791);
nand U1591 (N_1591,N_667,N_312);
xnor U1592 (N_1592,N_593,N_654);
and U1593 (N_1593,N_296,N_640);
xnor U1594 (N_1594,N_349,N_430);
nand U1595 (N_1595,N_954,N_880);
and U1596 (N_1596,N_903,N_51);
and U1597 (N_1597,N_229,N_654);
nand U1598 (N_1598,N_999,N_676);
nor U1599 (N_1599,N_937,N_759);
or U1600 (N_1600,N_621,N_724);
nor U1601 (N_1601,N_529,N_659);
or U1602 (N_1602,N_574,N_722);
xnor U1603 (N_1603,N_753,N_701);
or U1604 (N_1604,N_511,N_581);
or U1605 (N_1605,N_259,N_596);
or U1606 (N_1606,N_747,N_459);
or U1607 (N_1607,N_76,N_718);
nand U1608 (N_1608,N_251,N_324);
and U1609 (N_1609,N_231,N_936);
nor U1610 (N_1610,N_921,N_108);
nand U1611 (N_1611,N_124,N_558);
nand U1612 (N_1612,N_536,N_802);
and U1613 (N_1613,N_783,N_537);
nor U1614 (N_1614,N_767,N_106);
nor U1615 (N_1615,N_90,N_559);
or U1616 (N_1616,N_111,N_937);
nand U1617 (N_1617,N_407,N_620);
nand U1618 (N_1618,N_546,N_742);
nor U1619 (N_1619,N_666,N_789);
or U1620 (N_1620,N_530,N_149);
or U1621 (N_1621,N_603,N_717);
xnor U1622 (N_1622,N_387,N_356);
nand U1623 (N_1623,N_905,N_133);
nand U1624 (N_1624,N_360,N_291);
and U1625 (N_1625,N_893,N_557);
and U1626 (N_1626,N_812,N_298);
xor U1627 (N_1627,N_540,N_143);
or U1628 (N_1628,N_952,N_775);
or U1629 (N_1629,N_614,N_338);
nand U1630 (N_1630,N_118,N_465);
nand U1631 (N_1631,N_292,N_49);
and U1632 (N_1632,N_893,N_769);
nand U1633 (N_1633,N_687,N_373);
and U1634 (N_1634,N_342,N_885);
and U1635 (N_1635,N_949,N_144);
or U1636 (N_1636,N_416,N_604);
nand U1637 (N_1637,N_403,N_641);
nand U1638 (N_1638,N_776,N_286);
nor U1639 (N_1639,N_34,N_137);
or U1640 (N_1640,N_498,N_475);
or U1641 (N_1641,N_621,N_237);
nand U1642 (N_1642,N_605,N_663);
or U1643 (N_1643,N_271,N_471);
and U1644 (N_1644,N_776,N_880);
or U1645 (N_1645,N_819,N_232);
nand U1646 (N_1646,N_51,N_956);
xnor U1647 (N_1647,N_460,N_832);
and U1648 (N_1648,N_982,N_172);
xnor U1649 (N_1649,N_910,N_660);
nor U1650 (N_1650,N_440,N_664);
xor U1651 (N_1651,N_345,N_829);
and U1652 (N_1652,N_696,N_919);
nor U1653 (N_1653,N_885,N_661);
or U1654 (N_1654,N_273,N_386);
and U1655 (N_1655,N_421,N_422);
nand U1656 (N_1656,N_30,N_845);
or U1657 (N_1657,N_931,N_617);
xnor U1658 (N_1658,N_81,N_380);
nand U1659 (N_1659,N_486,N_785);
and U1660 (N_1660,N_86,N_185);
nand U1661 (N_1661,N_601,N_612);
nand U1662 (N_1662,N_99,N_467);
and U1663 (N_1663,N_229,N_237);
xnor U1664 (N_1664,N_279,N_302);
or U1665 (N_1665,N_522,N_994);
xnor U1666 (N_1666,N_973,N_850);
xor U1667 (N_1667,N_643,N_561);
nor U1668 (N_1668,N_126,N_906);
nor U1669 (N_1669,N_58,N_377);
nand U1670 (N_1670,N_67,N_512);
and U1671 (N_1671,N_42,N_119);
xor U1672 (N_1672,N_470,N_87);
and U1673 (N_1673,N_486,N_257);
nor U1674 (N_1674,N_56,N_6);
and U1675 (N_1675,N_336,N_635);
or U1676 (N_1676,N_104,N_744);
xor U1677 (N_1677,N_245,N_968);
or U1678 (N_1678,N_169,N_950);
or U1679 (N_1679,N_184,N_678);
nand U1680 (N_1680,N_601,N_311);
and U1681 (N_1681,N_123,N_36);
and U1682 (N_1682,N_403,N_618);
nor U1683 (N_1683,N_77,N_861);
or U1684 (N_1684,N_308,N_497);
nand U1685 (N_1685,N_192,N_882);
xor U1686 (N_1686,N_159,N_478);
xor U1687 (N_1687,N_115,N_701);
or U1688 (N_1688,N_604,N_338);
and U1689 (N_1689,N_408,N_912);
nor U1690 (N_1690,N_220,N_553);
xnor U1691 (N_1691,N_546,N_610);
and U1692 (N_1692,N_990,N_685);
nor U1693 (N_1693,N_333,N_766);
nor U1694 (N_1694,N_477,N_427);
or U1695 (N_1695,N_524,N_503);
xor U1696 (N_1696,N_571,N_478);
and U1697 (N_1697,N_329,N_27);
and U1698 (N_1698,N_100,N_113);
nor U1699 (N_1699,N_272,N_113);
nand U1700 (N_1700,N_773,N_384);
nand U1701 (N_1701,N_511,N_985);
nand U1702 (N_1702,N_4,N_194);
nor U1703 (N_1703,N_450,N_74);
nor U1704 (N_1704,N_194,N_5);
and U1705 (N_1705,N_117,N_732);
nor U1706 (N_1706,N_143,N_4);
nor U1707 (N_1707,N_264,N_806);
nand U1708 (N_1708,N_602,N_780);
xor U1709 (N_1709,N_860,N_848);
nand U1710 (N_1710,N_307,N_953);
nand U1711 (N_1711,N_748,N_173);
or U1712 (N_1712,N_946,N_874);
nor U1713 (N_1713,N_187,N_648);
nand U1714 (N_1714,N_479,N_467);
or U1715 (N_1715,N_911,N_162);
and U1716 (N_1716,N_364,N_927);
xor U1717 (N_1717,N_239,N_572);
or U1718 (N_1718,N_118,N_732);
and U1719 (N_1719,N_321,N_189);
and U1720 (N_1720,N_542,N_380);
or U1721 (N_1721,N_441,N_897);
xnor U1722 (N_1722,N_870,N_344);
or U1723 (N_1723,N_34,N_612);
and U1724 (N_1724,N_328,N_388);
xor U1725 (N_1725,N_593,N_553);
xor U1726 (N_1726,N_636,N_452);
or U1727 (N_1727,N_202,N_860);
nand U1728 (N_1728,N_356,N_88);
or U1729 (N_1729,N_231,N_990);
xor U1730 (N_1730,N_296,N_239);
or U1731 (N_1731,N_845,N_561);
or U1732 (N_1732,N_250,N_516);
nor U1733 (N_1733,N_669,N_697);
nand U1734 (N_1734,N_215,N_898);
or U1735 (N_1735,N_713,N_286);
xnor U1736 (N_1736,N_635,N_925);
and U1737 (N_1737,N_819,N_538);
nand U1738 (N_1738,N_267,N_125);
or U1739 (N_1739,N_98,N_745);
nor U1740 (N_1740,N_422,N_550);
nor U1741 (N_1741,N_767,N_117);
or U1742 (N_1742,N_553,N_743);
or U1743 (N_1743,N_871,N_579);
and U1744 (N_1744,N_315,N_170);
xor U1745 (N_1745,N_95,N_786);
nand U1746 (N_1746,N_311,N_223);
and U1747 (N_1747,N_603,N_528);
or U1748 (N_1748,N_762,N_394);
nand U1749 (N_1749,N_175,N_510);
nand U1750 (N_1750,N_608,N_614);
and U1751 (N_1751,N_665,N_781);
nand U1752 (N_1752,N_452,N_286);
and U1753 (N_1753,N_110,N_482);
nor U1754 (N_1754,N_428,N_196);
nand U1755 (N_1755,N_203,N_844);
xor U1756 (N_1756,N_289,N_189);
nor U1757 (N_1757,N_158,N_247);
and U1758 (N_1758,N_937,N_35);
nand U1759 (N_1759,N_912,N_255);
xnor U1760 (N_1760,N_818,N_943);
xnor U1761 (N_1761,N_873,N_503);
or U1762 (N_1762,N_268,N_83);
and U1763 (N_1763,N_715,N_792);
and U1764 (N_1764,N_961,N_11);
or U1765 (N_1765,N_262,N_248);
xnor U1766 (N_1766,N_650,N_100);
and U1767 (N_1767,N_382,N_746);
or U1768 (N_1768,N_937,N_129);
nand U1769 (N_1769,N_98,N_843);
and U1770 (N_1770,N_435,N_738);
nor U1771 (N_1771,N_730,N_468);
nor U1772 (N_1772,N_423,N_219);
nand U1773 (N_1773,N_168,N_669);
or U1774 (N_1774,N_4,N_516);
nor U1775 (N_1775,N_332,N_581);
xnor U1776 (N_1776,N_138,N_372);
nor U1777 (N_1777,N_294,N_317);
or U1778 (N_1778,N_934,N_981);
nor U1779 (N_1779,N_855,N_21);
and U1780 (N_1780,N_34,N_798);
xnor U1781 (N_1781,N_158,N_241);
nand U1782 (N_1782,N_218,N_782);
nand U1783 (N_1783,N_442,N_286);
or U1784 (N_1784,N_220,N_202);
nand U1785 (N_1785,N_209,N_824);
xnor U1786 (N_1786,N_129,N_512);
nand U1787 (N_1787,N_415,N_757);
or U1788 (N_1788,N_772,N_172);
xnor U1789 (N_1789,N_439,N_94);
and U1790 (N_1790,N_352,N_178);
and U1791 (N_1791,N_863,N_611);
or U1792 (N_1792,N_624,N_820);
nand U1793 (N_1793,N_68,N_975);
or U1794 (N_1794,N_158,N_145);
nand U1795 (N_1795,N_604,N_947);
xor U1796 (N_1796,N_147,N_848);
nand U1797 (N_1797,N_544,N_365);
nor U1798 (N_1798,N_621,N_446);
xor U1799 (N_1799,N_295,N_64);
xor U1800 (N_1800,N_603,N_385);
or U1801 (N_1801,N_890,N_47);
nand U1802 (N_1802,N_283,N_903);
and U1803 (N_1803,N_786,N_624);
and U1804 (N_1804,N_933,N_811);
or U1805 (N_1805,N_788,N_367);
or U1806 (N_1806,N_481,N_423);
and U1807 (N_1807,N_133,N_491);
nor U1808 (N_1808,N_138,N_410);
nand U1809 (N_1809,N_548,N_260);
nand U1810 (N_1810,N_417,N_134);
nand U1811 (N_1811,N_255,N_286);
xnor U1812 (N_1812,N_655,N_875);
xor U1813 (N_1813,N_148,N_142);
nand U1814 (N_1814,N_903,N_591);
nor U1815 (N_1815,N_592,N_686);
nand U1816 (N_1816,N_347,N_350);
xor U1817 (N_1817,N_372,N_479);
nor U1818 (N_1818,N_548,N_972);
nor U1819 (N_1819,N_379,N_391);
xnor U1820 (N_1820,N_403,N_948);
xor U1821 (N_1821,N_170,N_953);
or U1822 (N_1822,N_267,N_881);
nor U1823 (N_1823,N_263,N_620);
nand U1824 (N_1824,N_156,N_271);
nand U1825 (N_1825,N_41,N_132);
nor U1826 (N_1826,N_245,N_709);
nand U1827 (N_1827,N_118,N_454);
nand U1828 (N_1828,N_438,N_820);
and U1829 (N_1829,N_333,N_227);
nand U1830 (N_1830,N_661,N_134);
nor U1831 (N_1831,N_267,N_874);
or U1832 (N_1832,N_892,N_893);
nor U1833 (N_1833,N_945,N_519);
xnor U1834 (N_1834,N_960,N_22);
xor U1835 (N_1835,N_404,N_398);
xnor U1836 (N_1836,N_840,N_5);
nand U1837 (N_1837,N_279,N_682);
nor U1838 (N_1838,N_824,N_585);
nand U1839 (N_1839,N_489,N_666);
nand U1840 (N_1840,N_671,N_136);
nand U1841 (N_1841,N_347,N_333);
xnor U1842 (N_1842,N_217,N_1);
nand U1843 (N_1843,N_679,N_234);
and U1844 (N_1844,N_389,N_219);
or U1845 (N_1845,N_519,N_11);
and U1846 (N_1846,N_102,N_284);
xor U1847 (N_1847,N_568,N_180);
or U1848 (N_1848,N_116,N_710);
nor U1849 (N_1849,N_922,N_374);
and U1850 (N_1850,N_124,N_105);
and U1851 (N_1851,N_161,N_724);
nor U1852 (N_1852,N_530,N_933);
nor U1853 (N_1853,N_664,N_10);
xnor U1854 (N_1854,N_233,N_143);
nor U1855 (N_1855,N_240,N_400);
or U1856 (N_1856,N_797,N_580);
and U1857 (N_1857,N_943,N_226);
nand U1858 (N_1858,N_661,N_249);
or U1859 (N_1859,N_549,N_884);
and U1860 (N_1860,N_133,N_752);
and U1861 (N_1861,N_184,N_137);
nor U1862 (N_1862,N_482,N_512);
or U1863 (N_1863,N_761,N_496);
nand U1864 (N_1864,N_570,N_947);
and U1865 (N_1865,N_965,N_407);
or U1866 (N_1866,N_837,N_669);
nor U1867 (N_1867,N_733,N_719);
nor U1868 (N_1868,N_622,N_981);
nor U1869 (N_1869,N_82,N_376);
and U1870 (N_1870,N_18,N_959);
nor U1871 (N_1871,N_947,N_164);
or U1872 (N_1872,N_748,N_469);
nand U1873 (N_1873,N_497,N_833);
nand U1874 (N_1874,N_749,N_224);
and U1875 (N_1875,N_303,N_213);
xor U1876 (N_1876,N_852,N_278);
xnor U1877 (N_1877,N_197,N_996);
or U1878 (N_1878,N_921,N_735);
xor U1879 (N_1879,N_850,N_687);
xor U1880 (N_1880,N_615,N_385);
nor U1881 (N_1881,N_460,N_810);
nor U1882 (N_1882,N_375,N_485);
or U1883 (N_1883,N_522,N_806);
nor U1884 (N_1884,N_558,N_78);
xnor U1885 (N_1885,N_475,N_290);
and U1886 (N_1886,N_280,N_177);
and U1887 (N_1887,N_40,N_509);
nor U1888 (N_1888,N_127,N_777);
xnor U1889 (N_1889,N_210,N_457);
or U1890 (N_1890,N_500,N_617);
nand U1891 (N_1891,N_495,N_92);
or U1892 (N_1892,N_168,N_134);
and U1893 (N_1893,N_378,N_730);
nor U1894 (N_1894,N_680,N_112);
and U1895 (N_1895,N_847,N_588);
xnor U1896 (N_1896,N_109,N_917);
or U1897 (N_1897,N_718,N_836);
xor U1898 (N_1898,N_399,N_539);
xnor U1899 (N_1899,N_507,N_371);
and U1900 (N_1900,N_821,N_699);
xor U1901 (N_1901,N_31,N_938);
xnor U1902 (N_1902,N_112,N_442);
or U1903 (N_1903,N_365,N_307);
and U1904 (N_1904,N_577,N_851);
nand U1905 (N_1905,N_180,N_588);
and U1906 (N_1906,N_646,N_450);
or U1907 (N_1907,N_893,N_9);
or U1908 (N_1908,N_483,N_469);
or U1909 (N_1909,N_354,N_307);
xor U1910 (N_1910,N_106,N_682);
nand U1911 (N_1911,N_743,N_394);
nor U1912 (N_1912,N_544,N_424);
and U1913 (N_1913,N_567,N_691);
xor U1914 (N_1914,N_956,N_206);
xnor U1915 (N_1915,N_308,N_981);
or U1916 (N_1916,N_944,N_527);
nor U1917 (N_1917,N_499,N_724);
xor U1918 (N_1918,N_75,N_509);
and U1919 (N_1919,N_805,N_391);
nor U1920 (N_1920,N_442,N_150);
nand U1921 (N_1921,N_542,N_152);
nor U1922 (N_1922,N_11,N_28);
nor U1923 (N_1923,N_394,N_24);
nand U1924 (N_1924,N_755,N_790);
or U1925 (N_1925,N_495,N_464);
or U1926 (N_1926,N_909,N_962);
or U1927 (N_1927,N_382,N_499);
xor U1928 (N_1928,N_921,N_478);
nand U1929 (N_1929,N_239,N_425);
xnor U1930 (N_1930,N_573,N_395);
and U1931 (N_1931,N_173,N_595);
and U1932 (N_1932,N_8,N_468);
and U1933 (N_1933,N_354,N_186);
nand U1934 (N_1934,N_635,N_525);
or U1935 (N_1935,N_20,N_892);
xnor U1936 (N_1936,N_339,N_80);
or U1937 (N_1937,N_508,N_995);
and U1938 (N_1938,N_990,N_281);
nor U1939 (N_1939,N_177,N_564);
nor U1940 (N_1940,N_145,N_960);
or U1941 (N_1941,N_592,N_19);
nand U1942 (N_1942,N_54,N_391);
nor U1943 (N_1943,N_339,N_607);
nand U1944 (N_1944,N_284,N_711);
nand U1945 (N_1945,N_673,N_729);
xor U1946 (N_1946,N_796,N_28);
xor U1947 (N_1947,N_901,N_688);
nand U1948 (N_1948,N_565,N_508);
xnor U1949 (N_1949,N_423,N_789);
nor U1950 (N_1950,N_736,N_894);
xor U1951 (N_1951,N_548,N_475);
and U1952 (N_1952,N_871,N_260);
xnor U1953 (N_1953,N_929,N_878);
or U1954 (N_1954,N_432,N_838);
and U1955 (N_1955,N_487,N_856);
or U1956 (N_1956,N_351,N_655);
or U1957 (N_1957,N_981,N_503);
and U1958 (N_1958,N_780,N_852);
or U1959 (N_1959,N_768,N_727);
nor U1960 (N_1960,N_385,N_192);
xor U1961 (N_1961,N_775,N_198);
nand U1962 (N_1962,N_93,N_135);
nor U1963 (N_1963,N_874,N_766);
xnor U1964 (N_1964,N_119,N_253);
xnor U1965 (N_1965,N_794,N_635);
or U1966 (N_1966,N_785,N_997);
nor U1967 (N_1967,N_979,N_426);
nor U1968 (N_1968,N_93,N_383);
xor U1969 (N_1969,N_766,N_647);
nor U1970 (N_1970,N_20,N_695);
nor U1971 (N_1971,N_641,N_433);
and U1972 (N_1972,N_522,N_18);
and U1973 (N_1973,N_782,N_211);
nor U1974 (N_1974,N_235,N_458);
or U1975 (N_1975,N_239,N_9);
nor U1976 (N_1976,N_394,N_517);
or U1977 (N_1977,N_298,N_418);
nor U1978 (N_1978,N_313,N_556);
and U1979 (N_1979,N_922,N_109);
and U1980 (N_1980,N_796,N_281);
nand U1981 (N_1981,N_425,N_562);
nor U1982 (N_1982,N_336,N_764);
nor U1983 (N_1983,N_207,N_934);
xor U1984 (N_1984,N_100,N_114);
nor U1985 (N_1985,N_557,N_992);
nand U1986 (N_1986,N_253,N_758);
nor U1987 (N_1987,N_904,N_522);
nor U1988 (N_1988,N_993,N_385);
or U1989 (N_1989,N_287,N_303);
or U1990 (N_1990,N_68,N_793);
nand U1991 (N_1991,N_407,N_109);
or U1992 (N_1992,N_840,N_661);
nor U1993 (N_1993,N_236,N_608);
nand U1994 (N_1994,N_765,N_302);
and U1995 (N_1995,N_267,N_724);
nor U1996 (N_1996,N_942,N_514);
nand U1997 (N_1997,N_794,N_735);
or U1998 (N_1998,N_978,N_599);
xnor U1999 (N_1999,N_273,N_497);
and U2000 (N_2000,N_1786,N_1897);
xnor U2001 (N_2001,N_1673,N_1691);
nor U2002 (N_2002,N_1853,N_1543);
nand U2003 (N_2003,N_1357,N_1273);
nand U2004 (N_2004,N_1241,N_1036);
and U2005 (N_2005,N_1911,N_1612);
and U2006 (N_2006,N_1285,N_1568);
nor U2007 (N_2007,N_1584,N_1880);
xnor U2008 (N_2008,N_1839,N_1329);
nor U2009 (N_2009,N_1722,N_1066);
xnor U2010 (N_2010,N_1572,N_1463);
nor U2011 (N_2011,N_1406,N_1184);
xnor U2012 (N_2012,N_1877,N_1057);
xnor U2013 (N_2013,N_1913,N_1434);
nand U2014 (N_2014,N_1305,N_1702);
nand U2015 (N_2015,N_1652,N_1769);
xnor U2016 (N_2016,N_1025,N_1868);
xnor U2017 (N_2017,N_1466,N_1534);
and U2018 (N_2018,N_1738,N_1084);
or U2019 (N_2019,N_1332,N_1481);
or U2020 (N_2020,N_1507,N_1980);
nand U2021 (N_2021,N_1428,N_1016);
xnor U2022 (N_2022,N_1354,N_1969);
xor U2023 (N_2023,N_1894,N_1021);
and U2024 (N_2024,N_1928,N_1429);
nor U2025 (N_2025,N_1808,N_1122);
or U2026 (N_2026,N_1855,N_1148);
and U2027 (N_2027,N_1991,N_1182);
nand U2028 (N_2028,N_1760,N_1884);
xnor U2029 (N_2029,N_1934,N_1843);
nor U2030 (N_2030,N_1658,N_1228);
and U2031 (N_2031,N_1765,N_1633);
nor U2032 (N_2032,N_1154,N_1260);
and U2033 (N_2033,N_1407,N_1856);
and U2034 (N_2034,N_1772,N_1335);
and U2035 (N_2035,N_1915,N_1405);
xor U2036 (N_2036,N_1356,N_1200);
nand U2037 (N_2037,N_1314,N_1779);
or U2038 (N_2038,N_1266,N_1380);
nand U2039 (N_2039,N_1959,N_1918);
nand U2040 (N_2040,N_1456,N_1472);
or U2041 (N_2041,N_1675,N_1008);
nor U2042 (N_2042,N_1791,N_1471);
and U2043 (N_2043,N_1886,N_1920);
nor U2044 (N_2044,N_1660,N_1051);
nand U2045 (N_2045,N_1863,N_1014);
or U2046 (N_2046,N_1866,N_1694);
nand U2047 (N_2047,N_1803,N_1173);
and U2048 (N_2048,N_1500,N_1414);
and U2049 (N_2049,N_1951,N_1004);
nor U2050 (N_2050,N_1515,N_1501);
nand U2051 (N_2051,N_1419,N_1557);
nor U2052 (N_2052,N_1374,N_1056);
xor U2053 (N_2053,N_1152,N_1508);
and U2054 (N_2054,N_1267,N_1194);
nand U2055 (N_2055,N_1069,N_1547);
and U2056 (N_2056,N_1770,N_1806);
xor U2057 (N_2057,N_1616,N_1116);
nand U2058 (N_2058,N_1376,N_1392);
and U2059 (N_2059,N_1007,N_1831);
and U2060 (N_2060,N_1527,N_1889);
nand U2061 (N_2061,N_1771,N_1341);
and U2062 (N_2062,N_1602,N_1207);
or U2063 (N_2063,N_1922,N_1573);
and U2064 (N_2064,N_1859,N_1661);
xor U2065 (N_2065,N_1043,N_1246);
and U2066 (N_2066,N_1972,N_1895);
nor U2067 (N_2067,N_1238,N_1117);
nand U2068 (N_2068,N_1822,N_1902);
or U2069 (N_2069,N_1344,N_1511);
nor U2070 (N_2070,N_1667,N_1337);
nand U2071 (N_2071,N_1411,N_1067);
and U2072 (N_2072,N_1664,N_1430);
nand U2073 (N_2073,N_1119,N_1012);
or U2074 (N_2074,N_1676,N_1597);
xnor U2075 (N_2075,N_1022,N_1706);
or U2076 (N_2076,N_1090,N_1973);
nor U2077 (N_2077,N_1499,N_1916);
or U2078 (N_2078,N_1966,N_1085);
or U2079 (N_2079,N_1377,N_1778);
and U2080 (N_2080,N_1635,N_1999);
or U2081 (N_2081,N_1538,N_1288);
or U2082 (N_2082,N_1340,N_1265);
xnor U2083 (N_2083,N_1402,N_1105);
nand U2084 (N_2084,N_1542,N_1303);
or U2085 (N_2085,N_1869,N_1290);
and U2086 (N_2086,N_1925,N_1565);
or U2087 (N_2087,N_1409,N_1162);
nand U2088 (N_2088,N_1427,N_1514);
xor U2089 (N_2089,N_1359,N_1125);
or U2090 (N_2090,N_1531,N_1593);
nand U2091 (N_2091,N_1133,N_1494);
nor U2092 (N_2092,N_1272,N_1548);
xor U2093 (N_2093,N_1132,N_1968);
and U2094 (N_2094,N_1350,N_1062);
nand U2095 (N_2095,N_1111,N_1741);
or U2096 (N_2096,N_1188,N_1291);
and U2097 (N_2097,N_1214,N_1140);
and U2098 (N_2098,N_1513,N_1537);
nor U2099 (N_2099,N_1686,N_1930);
nor U2100 (N_2100,N_1005,N_1533);
xor U2101 (N_2101,N_1331,N_1330);
or U2102 (N_2102,N_1759,N_1081);
nor U2103 (N_2103,N_1473,N_1395);
nand U2104 (N_2104,N_1300,N_1674);
or U2105 (N_2105,N_1028,N_1035);
nor U2106 (N_2106,N_1165,N_1219);
nand U2107 (N_2107,N_1865,N_1408);
and U2108 (N_2108,N_1361,N_1095);
and U2109 (N_2109,N_1493,N_1669);
nor U2110 (N_2110,N_1996,N_1352);
xnor U2111 (N_2111,N_1933,N_1023);
and U2112 (N_2112,N_1334,N_1243);
or U2113 (N_2113,N_1129,N_1458);
xor U2114 (N_2114,N_1082,N_1432);
nand U2115 (N_2115,N_1417,N_1701);
nand U2116 (N_2116,N_1289,N_1032);
nor U2117 (N_2117,N_1160,N_1202);
or U2118 (N_2118,N_1109,N_1617);
and U2119 (N_2119,N_1452,N_1091);
xor U2120 (N_2120,N_1195,N_1955);
xor U2121 (N_2121,N_1995,N_1447);
and U2122 (N_2122,N_1301,N_1992);
nand U2123 (N_2123,N_1360,N_1242);
or U2124 (N_2124,N_1030,N_1536);
or U2125 (N_2125,N_1775,N_1546);
nand U2126 (N_2126,N_1651,N_1457);
nand U2127 (N_2127,N_1295,N_1298);
and U2128 (N_2128,N_1826,N_1812);
nand U2129 (N_2129,N_1782,N_1224);
nand U2130 (N_2130,N_1994,N_1728);
nor U2131 (N_2131,N_1704,N_1820);
xor U2132 (N_2132,N_1258,N_1807);
nor U2133 (N_2133,N_1550,N_1294);
nor U2134 (N_2134,N_1627,N_1217);
nor U2135 (N_2135,N_1474,N_1156);
nand U2136 (N_2136,N_1710,N_1079);
or U2137 (N_2137,N_1576,N_1271);
or U2138 (N_2138,N_1015,N_1124);
and U2139 (N_2139,N_1167,N_1393);
and U2140 (N_2140,N_1851,N_1997);
and U2141 (N_2141,N_1384,N_1622);
and U2142 (N_2142,N_1656,N_1908);
or U2143 (N_2143,N_1977,N_1465);
and U2144 (N_2144,N_1155,N_1017);
or U2145 (N_2145,N_1440,N_1087);
xor U2146 (N_2146,N_1735,N_1832);
nand U2147 (N_2147,N_1719,N_1445);
nand U2148 (N_2148,N_1179,N_1221);
xor U2149 (N_2149,N_1220,N_1985);
and U2150 (N_2150,N_1990,N_1521);
and U2151 (N_2151,N_1755,N_1787);
or U2152 (N_2152,N_1312,N_1767);
nand U2153 (N_2153,N_1436,N_1919);
nand U2154 (N_2154,N_1906,N_1963);
or U2155 (N_2155,N_1824,N_1752);
or U2156 (N_2156,N_1993,N_1952);
nor U2157 (N_2157,N_1257,N_1403);
nor U2158 (N_2158,N_1668,N_1281);
xor U2159 (N_2159,N_1423,N_1459);
and U2160 (N_2160,N_1496,N_1814);
and U2161 (N_2161,N_1177,N_1147);
or U2162 (N_2162,N_1881,N_1580);
and U2163 (N_2163,N_1603,N_1270);
nor U2164 (N_2164,N_1313,N_1625);
and U2165 (N_2165,N_1921,N_1181);
nand U2166 (N_2166,N_1185,N_1638);
xor U2167 (N_2167,N_1479,N_1401);
and U2168 (N_2168,N_1929,N_1491);
or U2169 (N_2169,N_1108,N_1914);
xnor U2170 (N_2170,N_1011,N_1926);
nand U2171 (N_2171,N_1848,N_1981);
or U2172 (N_2172,N_1239,N_1130);
and U2173 (N_2173,N_1611,N_1591);
nand U2174 (N_2174,N_1757,N_1903);
and U2175 (N_2175,N_1945,N_1149);
or U2176 (N_2176,N_1261,N_1198);
nand U2177 (N_2177,N_1070,N_1852);
or U2178 (N_2178,N_1818,N_1736);
nor U2179 (N_2179,N_1659,N_1366);
nor U2180 (N_2180,N_1323,N_1758);
xnor U2181 (N_2181,N_1749,N_1711);
xnor U2182 (N_2182,N_1747,N_1234);
and U2183 (N_2183,N_1879,N_1415);
nand U2184 (N_2184,N_1449,N_1583);
nand U2185 (N_2185,N_1956,N_1811);
and U2186 (N_2186,N_1932,N_1343);
nor U2187 (N_2187,N_1467,N_1009);
or U2188 (N_2188,N_1448,N_1805);
xnor U2189 (N_2189,N_1634,N_1123);
xnor U2190 (N_2190,N_1336,N_1168);
nor U2191 (N_2191,N_1789,N_1172);
nand U2192 (N_2192,N_1618,N_1784);
xnor U2193 (N_2193,N_1693,N_1316);
nand U2194 (N_2194,N_1699,N_1424);
or U2195 (N_2195,N_1763,N_1950);
nor U2196 (N_2196,N_1682,N_1315);
nor U2197 (N_2197,N_1708,N_1391);
nor U2198 (N_2198,N_1311,N_1225);
or U2199 (N_2199,N_1530,N_1631);
nand U2200 (N_2200,N_1308,N_1358);
and U2201 (N_2201,N_1590,N_1639);
nor U2202 (N_2202,N_1754,N_1072);
xnor U2203 (N_2203,N_1054,N_1827);
or U2204 (N_2204,N_1318,N_1365);
xor U2205 (N_2205,N_1883,N_1485);
xor U2206 (N_2206,N_1324,N_1059);
nor U2207 (N_2207,N_1277,N_1582);
nor U2208 (N_2208,N_1630,N_1042);
or U2209 (N_2209,N_1386,N_1872);
or U2210 (N_2210,N_1558,N_1400);
nand U2211 (N_2211,N_1142,N_1632);
and U2212 (N_2212,N_1662,N_1000);
nor U2213 (N_2213,N_1746,N_1347);
xnor U2214 (N_2214,N_1737,N_1286);
or U2215 (N_2215,N_1138,N_1961);
or U2216 (N_2216,N_1061,N_1716);
or U2217 (N_2217,N_1450,N_1099);
or U2218 (N_2218,N_1655,N_1720);
or U2219 (N_2219,N_1828,N_1846);
nand U2220 (N_2220,N_1605,N_1034);
nor U2221 (N_2221,N_1192,N_1768);
or U2222 (N_2222,N_1068,N_1398);
or U2223 (N_2223,N_1055,N_1954);
or U2224 (N_2224,N_1255,N_1197);
nand U2225 (N_2225,N_1641,N_1263);
nand U2226 (N_2226,N_1064,N_1551);
xor U2227 (N_2227,N_1136,N_1650);
nand U2228 (N_2228,N_1685,N_1975);
or U2229 (N_2229,N_1088,N_1421);
nor U2230 (N_2230,N_1112,N_1413);
nor U2231 (N_2231,N_1753,N_1570);
xnor U2232 (N_2232,N_1029,N_1309);
nand U2233 (N_2233,N_1461,N_1802);
and U2234 (N_2234,N_1924,N_1698);
xor U2235 (N_2235,N_1717,N_1193);
nor U2236 (N_2236,N_1215,N_1180);
nor U2237 (N_2237,N_1328,N_1610);
nor U2238 (N_2238,N_1739,N_1478);
nand U2239 (N_2239,N_1134,N_1891);
xnor U2240 (N_2240,N_1367,N_1205);
and U2241 (N_2241,N_1204,N_1351);
nand U2242 (N_2242,N_1104,N_1060);
xnor U2243 (N_2243,N_1788,N_1037);
and U2244 (N_2244,N_1399,N_1714);
nor U2245 (N_2245,N_1705,N_1212);
nand U2246 (N_2246,N_1126,N_1046);
nor U2247 (N_2247,N_1163,N_1599);
xnor U2248 (N_2248,N_1346,N_1598);
or U2249 (N_2249,N_1890,N_1947);
nand U2250 (N_2250,N_1208,N_1917);
nand U2251 (N_2251,N_1556,N_1766);
and U2252 (N_2252,N_1861,N_1236);
or U2253 (N_2253,N_1744,N_1495);
or U2254 (N_2254,N_1480,N_1909);
or U2255 (N_2255,N_1489,N_1362);
nor U2256 (N_2256,N_1319,N_1077);
xnor U2257 (N_2257,N_1823,N_1483);
nor U2258 (N_2258,N_1844,N_1525);
or U2259 (N_2259,N_1278,N_1885);
and U2260 (N_2260,N_1137,N_1683);
or U2261 (N_2261,N_1539,N_1158);
xor U2262 (N_2262,N_1535,N_1245);
nor U2263 (N_2263,N_1169,N_1426);
or U2264 (N_2264,N_1709,N_1206);
nand U2265 (N_2265,N_1927,N_1707);
or U2266 (N_2266,N_1497,N_1742);
nand U2267 (N_2267,N_1882,N_1027);
xor U2268 (N_2268,N_1703,N_1821);
nor U2269 (N_2269,N_1368,N_1888);
nor U2270 (N_2270,N_1946,N_1971);
nand U2271 (N_2271,N_1781,N_1086);
xnor U2272 (N_2272,N_1488,N_1433);
or U2273 (N_2273,N_1528,N_1498);
or U2274 (N_2274,N_1813,N_1187);
and U2275 (N_2275,N_1503,N_1482);
xor U2276 (N_2276,N_1306,N_1256);
nand U2277 (N_2277,N_1773,N_1732);
nand U2278 (N_2278,N_1250,N_1101);
nor U2279 (N_2279,N_1640,N_1734);
and U2280 (N_2280,N_1559,N_1860);
and U2281 (N_2281,N_1325,N_1190);
nor U2282 (N_2282,N_1191,N_1454);
and U2283 (N_2283,N_1385,N_1578);
xnor U2284 (N_2284,N_1387,N_1743);
or U2285 (N_2285,N_1218,N_1998);
nor U2286 (N_2286,N_1923,N_1562);
nor U2287 (N_2287,N_1199,N_1460);
or U2288 (N_2288,N_1389,N_1983);
nor U2289 (N_2289,N_1887,N_1751);
or U2290 (N_2290,N_1984,N_1608);
and U2291 (N_2291,N_1512,N_1825);
nand U2292 (N_2292,N_1541,N_1135);
nor U2293 (N_2293,N_1912,N_1041);
nor U2294 (N_2294,N_1476,N_1280);
or U2295 (N_2295,N_1937,N_1834);
nand U2296 (N_2296,N_1170,N_1431);
xor U2297 (N_2297,N_1989,N_1150);
nor U2298 (N_2298,N_1438,N_1725);
nand U2299 (N_2299,N_1816,N_1700);
nor U2300 (N_2300,N_1988,N_1183);
nand U2301 (N_2301,N_1339,N_1878);
nor U2302 (N_2302,N_1645,N_1010);
nand U2303 (N_2303,N_1829,N_1692);
xnor U2304 (N_2304,N_1073,N_1626);
or U2305 (N_2305,N_1382,N_1777);
xnor U2306 (N_2306,N_1974,N_1774);
nor U2307 (N_2307,N_1047,N_1412);
nor U2308 (N_2308,N_1441,N_1801);
or U2309 (N_2309,N_1209,N_1321);
nor U2310 (N_2310,N_1904,N_1282);
and U2311 (N_2311,N_1468,N_1678);
xor U2312 (N_2312,N_1127,N_1264);
and U2313 (N_2313,N_1506,N_1577);
nor U2314 (N_2314,N_1240,N_1033);
and U2315 (N_2315,N_1798,N_1874);
nand U2316 (N_2316,N_1592,N_1949);
xnor U2317 (N_2317,N_1785,N_1526);
xnor U2318 (N_2318,N_1681,N_1666);
xor U2319 (N_2319,N_1131,N_1729);
or U2320 (N_2320,N_1231,N_1516);
nor U2321 (N_2321,N_1871,N_1776);
nor U2322 (N_2322,N_1620,N_1048);
xnor U2323 (N_2323,N_1540,N_1435);
or U2324 (N_2324,N_1905,N_1657);
and U2325 (N_2325,N_1796,N_1671);
xnor U2326 (N_2326,N_1201,N_1713);
nor U2327 (N_2327,N_1836,N_1520);
xor U2328 (N_2328,N_1646,N_1939);
xnor U2329 (N_2329,N_1196,N_1561);
nor U2330 (N_2330,N_1484,N_1020);
or U2331 (N_2331,N_1254,N_1670);
xor U2332 (N_2332,N_1092,N_1410);
or U2333 (N_2333,N_1804,N_1372);
nor U2334 (N_2334,N_1970,N_1279);
xor U2335 (N_2335,N_1797,N_1063);
nor U2336 (N_2336,N_1649,N_1726);
nand U2337 (N_2337,N_1875,N_1353);
and U2338 (N_2338,N_1186,N_1519);
or U2339 (N_2339,N_1249,N_1689);
xnor U2340 (N_2340,N_1680,N_1375);
and U2341 (N_2341,N_1900,N_1965);
nand U2342 (N_2342,N_1615,N_1078);
nand U2343 (N_2343,N_1115,N_1274);
nand U2344 (N_2344,N_1120,N_1102);
and U2345 (N_2345,N_1723,N_1227);
nand U2346 (N_2346,N_1672,N_1566);
and U2347 (N_2347,N_1636,N_1600);
xor U2348 (N_2348,N_1838,N_1854);
or U2349 (N_2349,N_1587,N_1850);
xnor U2350 (N_2350,N_1940,N_1013);
nor U2351 (N_2351,N_1830,N_1379);
or U2352 (N_2352,N_1018,N_1810);
and U2353 (N_2353,N_1244,N_1867);
or U2354 (N_2354,N_1297,N_1143);
or U2355 (N_2355,N_1817,N_1727);
nand U2356 (N_2356,N_1750,N_1383);
nand U2357 (N_2357,N_1296,N_1555);
nand U2358 (N_2358,N_1189,N_1761);
xnor U2359 (N_2359,N_1629,N_1342);
or U2360 (N_2360,N_1145,N_1799);
or U2361 (N_2361,N_1322,N_1790);
and U2362 (N_2362,N_1864,N_1841);
and U2363 (N_2363,N_1601,N_1226);
nor U2364 (N_2364,N_1107,N_1718);
or U2365 (N_2365,N_1161,N_1957);
nand U2366 (N_2366,N_1978,N_1840);
xnor U2367 (N_2367,N_1604,N_1545);
and U2368 (N_2368,N_1381,N_1469);
and U2369 (N_2369,N_1229,N_1178);
and U2370 (N_2370,N_1733,N_1024);
and U2371 (N_2371,N_1941,N_1532);
nand U2372 (N_2372,N_1276,N_1210);
and U2373 (N_2373,N_1862,N_1175);
nand U2374 (N_2374,N_1338,N_1058);
or U2375 (N_2375,N_1378,N_1118);
nor U2376 (N_2376,N_1349,N_1006);
nand U2377 (N_2377,N_1490,N_1544);
nand U2378 (N_2378,N_1628,N_1151);
or U2379 (N_2379,N_1783,N_1619);
and U2380 (N_2380,N_1096,N_1232);
nor U2381 (N_2381,N_1019,N_1756);
and U2382 (N_2382,N_1517,N_1222);
or U2383 (N_2383,N_1327,N_1745);
nand U2384 (N_2384,N_1574,N_1644);
and U2385 (N_2385,N_1964,N_1233);
and U2386 (N_2386,N_1462,N_1446);
nand U2387 (N_2387,N_1792,N_1607);
nor U2388 (N_2388,N_1464,N_1213);
xor U2389 (N_2389,N_1893,N_1302);
or U2390 (N_2390,N_1960,N_1040);
and U2391 (N_2391,N_1589,N_1110);
xnor U2392 (N_2392,N_1575,N_1416);
nand U2393 (N_2393,N_1251,N_1800);
and U2394 (N_2394,N_1114,N_1001);
or U2395 (N_2395,N_1748,N_1326);
xnor U2396 (N_2396,N_1363,N_1269);
xor U2397 (N_2397,N_1128,N_1986);
xor U2398 (N_2398,N_1857,N_1690);
nor U2399 (N_2399,N_1938,N_1247);
nor U2400 (N_2400,N_1849,N_1369);
nand U2401 (N_2401,N_1609,N_1696);
or U2402 (N_2402,N_1594,N_1653);
or U2403 (N_2403,N_1262,N_1364);
xnor U2404 (N_2404,N_1404,N_1621);
nand U2405 (N_2405,N_1098,N_1569);
and U2406 (N_2406,N_1453,N_1958);
and U2407 (N_2407,N_1987,N_1420);
or U2408 (N_2408,N_1422,N_1348);
nor U2409 (N_2409,N_1333,N_1809);
nand U2410 (N_2410,N_1388,N_1901);
or U2411 (N_2411,N_1292,N_1795);
nand U2412 (N_2412,N_1371,N_1596);
nand U2413 (N_2413,N_1252,N_1355);
nand U2414 (N_2414,N_1979,N_1505);
nor U2415 (N_2415,N_1654,N_1031);
xnor U2416 (N_2416,N_1815,N_1876);
nor U2417 (N_2417,N_1396,N_1470);
nand U2418 (N_2418,N_1870,N_1284);
and U2419 (N_2419,N_1571,N_1100);
or U2420 (N_2420,N_1648,N_1216);
or U2421 (N_2421,N_1962,N_1093);
xor U2422 (N_2422,N_1071,N_1873);
xor U2423 (N_2423,N_1153,N_1026);
xnor U2424 (N_2424,N_1936,N_1614);
nor U2425 (N_2425,N_1074,N_1982);
and U2426 (N_2426,N_1845,N_1942);
nor U2427 (N_2427,N_1065,N_1475);
xnor U2428 (N_2428,N_1076,N_1268);
nor U2429 (N_2429,N_1439,N_1953);
nor U2430 (N_2430,N_1259,N_1665);
or U2431 (N_2431,N_1451,N_1103);
nor U2432 (N_2432,N_1144,N_1898);
nand U2433 (N_2433,N_1647,N_1299);
nor U2434 (N_2434,N_1684,N_1394);
xnor U2435 (N_2435,N_1842,N_1304);
xor U2436 (N_2436,N_1141,N_1637);
nand U2437 (N_2437,N_1425,N_1522);
nor U2438 (N_2438,N_1724,N_1663);
nor U2439 (N_2439,N_1695,N_1721);
nor U2440 (N_2440,N_1050,N_1345);
nor U2441 (N_2441,N_1039,N_1935);
nor U2442 (N_2442,N_1390,N_1307);
and U2443 (N_2443,N_1171,N_1003);
nor U2444 (N_2444,N_1837,N_1097);
xnor U2445 (N_2445,N_1492,N_1564);
or U2446 (N_2446,N_1677,N_1793);
nand U2447 (N_2447,N_1443,N_1899);
nor U2448 (N_2448,N_1176,N_1283);
xor U2449 (N_2449,N_1948,N_1907);
nor U2450 (N_2450,N_1106,N_1509);
nand U2451 (N_2451,N_1164,N_1455);
nand U2452 (N_2452,N_1211,N_1910);
or U2453 (N_2453,N_1089,N_1524);
and U2454 (N_2454,N_1554,N_1052);
and U2455 (N_2455,N_1643,N_1518);
and U2456 (N_2456,N_1293,N_1080);
and U2457 (N_2457,N_1858,N_1094);
or U2458 (N_2458,N_1679,N_1762);
nand U2459 (N_2459,N_1230,N_1967);
or U2460 (N_2460,N_1563,N_1044);
nand U2461 (N_2461,N_1581,N_1730);
and U2462 (N_2462,N_1253,N_1002);
and U2463 (N_2463,N_1523,N_1976);
and U2464 (N_2464,N_1444,N_1688);
xnor U2465 (N_2465,N_1740,N_1203);
nor U2466 (N_2466,N_1113,N_1248);
or U2467 (N_2467,N_1075,N_1166);
nor U2468 (N_2468,N_1560,N_1320);
and U2469 (N_2469,N_1477,N_1585);
and U2470 (N_2470,N_1606,N_1121);
nand U2471 (N_2471,N_1712,N_1780);
and U2472 (N_2472,N_1045,N_1174);
nand U2473 (N_2473,N_1235,N_1549);
nand U2474 (N_2474,N_1437,N_1624);
nand U2475 (N_2475,N_1139,N_1157);
or U2476 (N_2476,N_1819,N_1896);
and U2477 (N_2477,N_1049,N_1731);
nor U2478 (N_2478,N_1373,N_1159);
nor U2479 (N_2479,N_1038,N_1835);
and U2480 (N_2480,N_1715,N_1586);
and U2481 (N_2481,N_1794,N_1502);
nand U2482 (N_2482,N_1083,N_1579);
and U2483 (N_2483,N_1833,N_1053);
xor U2484 (N_2484,N_1317,N_1504);
and U2485 (N_2485,N_1287,N_1146);
or U2486 (N_2486,N_1944,N_1237);
or U2487 (N_2487,N_1529,N_1931);
xnor U2488 (N_2488,N_1613,N_1418);
and U2489 (N_2489,N_1397,N_1687);
and U2490 (N_2490,N_1487,N_1943);
xor U2491 (N_2491,N_1642,N_1486);
and U2492 (N_2492,N_1552,N_1370);
or U2493 (N_2493,N_1510,N_1764);
or U2494 (N_2494,N_1223,N_1275);
and U2495 (N_2495,N_1588,N_1595);
and U2496 (N_2496,N_1567,N_1847);
or U2497 (N_2497,N_1442,N_1892);
nor U2498 (N_2498,N_1553,N_1310);
xnor U2499 (N_2499,N_1623,N_1697);
nor U2500 (N_2500,N_1570,N_1061);
nor U2501 (N_2501,N_1680,N_1884);
xor U2502 (N_2502,N_1758,N_1363);
xor U2503 (N_2503,N_1529,N_1421);
and U2504 (N_2504,N_1748,N_1619);
or U2505 (N_2505,N_1581,N_1106);
nand U2506 (N_2506,N_1540,N_1615);
nor U2507 (N_2507,N_1478,N_1964);
nand U2508 (N_2508,N_1693,N_1544);
or U2509 (N_2509,N_1111,N_1212);
or U2510 (N_2510,N_1346,N_1656);
nor U2511 (N_2511,N_1986,N_1767);
or U2512 (N_2512,N_1668,N_1639);
nand U2513 (N_2513,N_1613,N_1460);
and U2514 (N_2514,N_1597,N_1134);
or U2515 (N_2515,N_1934,N_1005);
nor U2516 (N_2516,N_1082,N_1387);
xnor U2517 (N_2517,N_1192,N_1462);
nor U2518 (N_2518,N_1038,N_1706);
nor U2519 (N_2519,N_1996,N_1461);
or U2520 (N_2520,N_1152,N_1599);
nand U2521 (N_2521,N_1357,N_1259);
xnor U2522 (N_2522,N_1933,N_1488);
xnor U2523 (N_2523,N_1888,N_1899);
xor U2524 (N_2524,N_1619,N_1499);
and U2525 (N_2525,N_1690,N_1230);
nor U2526 (N_2526,N_1905,N_1065);
or U2527 (N_2527,N_1190,N_1013);
nand U2528 (N_2528,N_1070,N_1158);
and U2529 (N_2529,N_1637,N_1766);
xor U2530 (N_2530,N_1715,N_1983);
nor U2531 (N_2531,N_1319,N_1032);
or U2532 (N_2532,N_1747,N_1555);
and U2533 (N_2533,N_1254,N_1888);
xor U2534 (N_2534,N_1512,N_1647);
nor U2535 (N_2535,N_1880,N_1077);
or U2536 (N_2536,N_1638,N_1346);
nand U2537 (N_2537,N_1923,N_1525);
or U2538 (N_2538,N_1179,N_1160);
or U2539 (N_2539,N_1519,N_1801);
nand U2540 (N_2540,N_1101,N_1696);
and U2541 (N_2541,N_1480,N_1788);
nand U2542 (N_2542,N_1831,N_1175);
nor U2543 (N_2543,N_1539,N_1976);
and U2544 (N_2544,N_1617,N_1418);
nand U2545 (N_2545,N_1141,N_1112);
nand U2546 (N_2546,N_1618,N_1064);
xor U2547 (N_2547,N_1900,N_1705);
xor U2548 (N_2548,N_1231,N_1942);
and U2549 (N_2549,N_1372,N_1243);
or U2550 (N_2550,N_1721,N_1500);
or U2551 (N_2551,N_1560,N_1365);
nand U2552 (N_2552,N_1303,N_1270);
and U2553 (N_2553,N_1530,N_1240);
or U2554 (N_2554,N_1720,N_1432);
or U2555 (N_2555,N_1954,N_1694);
xor U2556 (N_2556,N_1375,N_1834);
nand U2557 (N_2557,N_1691,N_1308);
nor U2558 (N_2558,N_1732,N_1244);
nor U2559 (N_2559,N_1768,N_1450);
and U2560 (N_2560,N_1542,N_1591);
or U2561 (N_2561,N_1074,N_1509);
or U2562 (N_2562,N_1586,N_1029);
nand U2563 (N_2563,N_1526,N_1472);
and U2564 (N_2564,N_1727,N_1844);
nor U2565 (N_2565,N_1589,N_1302);
xor U2566 (N_2566,N_1229,N_1688);
or U2567 (N_2567,N_1841,N_1145);
nand U2568 (N_2568,N_1782,N_1615);
or U2569 (N_2569,N_1295,N_1717);
nand U2570 (N_2570,N_1245,N_1181);
nor U2571 (N_2571,N_1960,N_1072);
and U2572 (N_2572,N_1946,N_1875);
nor U2573 (N_2573,N_1164,N_1024);
and U2574 (N_2574,N_1740,N_1208);
nor U2575 (N_2575,N_1020,N_1243);
nand U2576 (N_2576,N_1747,N_1949);
nor U2577 (N_2577,N_1303,N_1522);
nand U2578 (N_2578,N_1413,N_1545);
and U2579 (N_2579,N_1377,N_1551);
and U2580 (N_2580,N_1231,N_1883);
xor U2581 (N_2581,N_1091,N_1261);
nand U2582 (N_2582,N_1411,N_1596);
or U2583 (N_2583,N_1539,N_1472);
or U2584 (N_2584,N_1981,N_1119);
and U2585 (N_2585,N_1399,N_1999);
xor U2586 (N_2586,N_1245,N_1347);
and U2587 (N_2587,N_1529,N_1522);
or U2588 (N_2588,N_1593,N_1852);
or U2589 (N_2589,N_1030,N_1527);
or U2590 (N_2590,N_1784,N_1503);
and U2591 (N_2591,N_1317,N_1960);
nor U2592 (N_2592,N_1238,N_1125);
xnor U2593 (N_2593,N_1486,N_1076);
and U2594 (N_2594,N_1422,N_1614);
nor U2595 (N_2595,N_1744,N_1601);
nand U2596 (N_2596,N_1298,N_1003);
xnor U2597 (N_2597,N_1399,N_1849);
and U2598 (N_2598,N_1020,N_1199);
nor U2599 (N_2599,N_1375,N_1497);
xnor U2600 (N_2600,N_1938,N_1623);
xnor U2601 (N_2601,N_1239,N_1133);
and U2602 (N_2602,N_1817,N_1939);
or U2603 (N_2603,N_1433,N_1547);
or U2604 (N_2604,N_1528,N_1722);
nand U2605 (N_2605,N_1923,N_1663);
xor U2606 (N_2606,N_1627,N_1892);
nand U2607 (N_2607,N_1786,N_1728);
nand U2608 (N_2608,N_1667,N_1378);
nor U2609 (N_2609,N_1983,N_1112);
nor U2610 (N_2610,N_1970,N_1140);
or U2611 (N_2611,N_1611,N_1224);
xnor U2612 (N_2612,N_1560,N_1029);
and U2613 (N_2613,N_1598,N_1659);
and U2614 (N_2614,N_1492,N_1584);
or U2615 (N_2615,N_1226,N_1943);
or U2616 (N_2616,N_1625,N_1212);
nor U2617 (N_2617,N_1066,N_1161);
xnor U2618 (N_2618,N_1067,N_1096);
and U2619 (N_2619,N_1672,N_1933);
nand U2620 (N_2620,N_1518,N_1867);
and U2621 (N_2621,N_1568,N_1805);
xnor U2622 (N_2622,N_1018,N_1767);
nand U2623 (N_2623,N_1896,N_1138);
nand U2624 (N_2624,N_1423,N_1761);
nor U2625 (N_2625,N_1508,N_1956);
nor U2626 (N_2626,N_1289,N_1208);
and U2627 (N_2627,N_1556,N_1644);
and U2628 (N_2628,N_1077,N_1304);
xor U2629 (N_2629,N_1861,N_1117);
nand U2630 (N_2630,N_1538,N_1345);
xor U2631 (N_2631,N_1103,N_1070);
nand U2632 (N_2632,N_1325,N_1341);
or U2633 (N_2633,N_1475,N_1898);
or U2634 (N_2634,N_1426,N_1635);
or U2635 (N_2635,N_1404,N_1851);
nor U2636 (N_2636,N_1899,N_1862);
nand U2637 (N_2637,N_1787,N_1198);
or U2638 (N_2638,N_1785,N_1207);
nor U2639 (N_2639,N_1477,N_1906);
or U2640 (N_2640,N_1407,N_1678);
and U2641 (N_2641,N_1663,N_1810);
nor U2642 (N_2642,N_1376,N_1996);
nor U2643 (N_2643,N_1576,N_1747);
xnor U2644 (N_2644,N_1375,N_1403);
and U2645 (N_2645,N_1845,N_1022);
and U2646 (N_2646,N_1120,N_1032);
nor U2647 (N_2647,N_1422,N_1162);
or U2648 (N_2648,N_1263,N_1176);
or U2649 (N_2649,N_1389,N_1168);
nand U2650 (N_2650,N_1859,N_1498);
and U2651 (N_2651,N_1898,N_1037);
nand U2652 (N_2652,N_1861,N_1244);
and U2653 (N_2653,N_1324,N_1805);
and U2654 (N_2654,N_1889,N_1950);
and U2655 (N_2655,N_1742,N_1297);
nor U2656 (N_2656,N_1739,N_1261);
xor U2657 (N_2657,N_1317,N_1590);
nor U2658 (N_2658,N_1396,N_1436);
xor U2659 (N_2659,N_1082,N_1095);
or U2660 (N_2660,N_1861,N_1585);
nor U2661 (N_2661,N_1404,N_1516);
nor U2662 (N_2662,N_1381,N_1507);
xor U2663 (N_2663,N_1529,N_1412);
or U2664 (N_2664,N_1358,N_1098);
xor U2665 (N_2665,N_1590,N_1119);
nor U2666 (N_2666,N_1918,N_1913);
and U2667 (N_2667,N_1133,N_1937);
and U2668 (N_2668,N_1536,N_1002);
nor U2669 (N_2669,N_1398,N_1500);
and U2670 (N_2670,N_1254,N_1433);
nand U2671 (N_2671,N_1372,N_1852);
and U2672 (N_2672,N_1954,N_1228);
and U2673 (N_2673,N_1878,N_1841);
or U2674 (N_2674,N_1037,N_1375);
and U2675 (N_2675,N_1413,N_1896);
nor U2676 (N_2676,N_1419,N_1060);
and U2677 (N_2677,N_1770,N_1426);
xnor U2678 (N_2678,N_1977,N_1037);
nand U2679 (N_2679,N_1338,N_1387);
and U2680 (N_2680,N_1527,N_1682);
xor U2681 (N_2681,N_1176,N_1970);
xor U2682 (N_2682,N_1550,N_1251);
nand U2683 (N_2683,N_1225,N_1413);
nand U2684 (N_2684,N_1859,N_1355);
nand U2685 (N_2685,N_1093,N_1881);
or U2686 (N_2686,N_1692,N_1323);
nand U2687 (N_2687,N_1108,N_1464);
nor U2688 (N_2688,N_1225,N_1191);
and U2689 (N_2689,N_1149,N_1079);
and U2690 (N_2690,N_1799,N_1217);
or U2691 (N_2691,N_1918,N_1937);
or U2692 (N_2692,N_1993,N_1245);
nor U2693 (N_2693,N_1600,N_1429);
and U2694 (N_2694,N_1124,N_1698);
nand U2695 (N_2695,N_1043,N_1561);
or U2696 (N_2696,N_1456,N_1158);
and U2697 (N_2697,N_1469,N_1959);
xnor U2698 (N_2698,N_1121,N_1728);
and U2699 (N_2699,N_1867,N_1503);
nor U2700 (N_2700,N_1123,N_1144);
nor U2701 (N_2701,N_1980,N_1074);
nor U2702 (N_2702,N_1819,N_1950);
xor U2703 (N_2703,N_1870,N_1341);
and U2704 (N_2704,N_1619,N_1827);
or U2705 (N_2705,N_1907,N_1734);
and U2706 (N_2706,N_1487,N_1336);
xnor U2707 (N_2707,N_1715,N_1869);
nand U2708 (N_2708,N_1105,N_1736);
and U2709 (N_2709,N_1026,N_1665);
and U2710 (N_2710,N_1436,N_1170);
and U2711 (N_2711,N_1709,N_1743);
xnor U2712 (N_2712,N_1252,N_1694);
nand U2713 (N_2713,N_1322,N_1831);
or U2714 (N_2714,N_1827,N_1561);
xnor U2715 (N_2715,N_1740,N_1687);
nor U2716 (N_2716,N_1701,N_1773);
nor U2717 (N_2717,N_1979,N_1899);
nand U2718 (N_2718,N_1593,N_1400);
nand U2719 (N_2719,N_1616,N_1149);
xnor U2720 (N_2720,N_1585,N_1214);
or U2721 (N_2721,N_1717,N_1012);
nand U2722 (N_2722,N_1998,N_1508);
nor U2723 (N_2723,N_1029,N_1953);
xor U2724 (N_2724,N_1385,N_1918);
or U2725 (N_2725,N_1941,N_1845);
xnor U2726 (N_2726,N_1213,N_1115);
or U2727 (N_2727,N_1278,N_1985);
or U2728 (N_2728,N_1506,N_1526);
nor U2729 (N_2729,N_1518,N_1078);
nand U2730 (N_2730,N_1832,N_1895);
nor U2731 (N_2731,N_1190,N_1877);
and U2732 (N_2732,N_1480,N_1712);
or U2733 (N_2733,N_1787,N_1760);
or U2734 (N_2734,N_1313,N_1202);
nor U2735 (N_2735,N_1322,N_1929);
or U2736 (N_2736,N_1084,N_1552);
nand U2737 (N_2737,N_1184,N_1587);
nor U2738 (N_2738,N_1829,N_1754);
xnor U2739 (N_2739,N_1756,N_1947);
and U2740 (N_2740,N_1457,N_1429);
xnor U2741 (N_2741,N_1715,N_1255);
and U2742 (N_2742,N_1274,N_1773);
nor U2743 (N_2743,N_1241,N_1723);
or U2744 (N_2744,N_1156,N_1286);
and U2745 (N_2745,N_1377,N_1714);
nand U2746 (N_2746,N_1077,N_1938);
and U2747 (N_2747,N_1597,N_1283);
nor U2748 (N_2748,N_1755,N_1660);
xor U2749 (N_2749,N_1059,N_1477);
xnor U2750 (N_2750,N_1768,N_1204);
and U2751 (N_2751,N_1750,N_1713);
nor U2752 (N_2752,N_1166,N_1580);
and U2753 (N_2753,N_1679,N_1970);
nand U2754 (N_2754,N_1618,N_1519);
or U2755 (N_2755,N_1022,N_1177);
and U2756 (N_2756,N_1272,N_1404);
xor U2757 (N_2757,N_1412,N_1830);
nor U2758 (N_2758,N_1670,N_1406);
and U2759 (N_2759,N_1663,N_1417);
nor U2760 (N_2760,N_1114,N_1499);
nand U2761 (N_2761,N_1259,N_1767);
or U2762 (N_2762,N_1117,N_1123);
xor U2763 (N_2763,N_1670,N_1794);
and U2764 (N_2764,N_1331,N_1134);
xnor U2765 (N_2765,N_1000,N_1261);
and U2766 (N_2766,N_1432,N_1050);
xor U2767 (N_2767,N_1362,N_1919);
nor U2768 (N_2768,N_1395,N_1106);
nand U2769 (N_2769,N_1014,N_1191);
nor U2770 (N_2770,N_1908,N_1925);
nor U2771 (N_2771,N_1451,N_1328);
nand U2772 (N_2772,N_1687,N_1336);
xnor U2773 (N_2773,N_1171,N_1769);
nand U2774 (N_2774,N_1440,N_1226);
xor U2775 (N_2775,N_1144,N_1945);
or U2776 (N_2776,N_1017,N_1503);
or U2777 (N_2777,N_1880,N_1243);
xnor U2778 (N_2778,N_1319,N_1540);
xnor U2779 (N_2779,N_1582,N_1390);
or U2780 (N_2780,N_1833,N_1442);
or U2781 (N_2781,N_1399,N_1294);
xnor U2782 (N_2782,N_1055,N_1195);
nand U2783 (N_2783,N_1820,N_1174);
or U2784 (N_2784,N_1401,N_1876);
nand U2785 (N_2785,N_1856,N_1896);
or U2786 (N_2786,N_1755,N_1735);
nor U2787 (N_2787,N_1471,N_1388);
nor U2788 (N_2788,N_1576,N_1040);
and U2789 (N_2789,N_1918,N_1569);
and U2790 (N_2790,N_1387,N_1595);
nor U2791 (N_2791,N_1763,N_1153);
or U2792 (N_2792,N_1549,N_1242);
nand U2793 (N_2793,N_1918,N_1697);
nor U2794 (N_2794,N_1100,N_1188);
nor U2795 (N_2795,N_1916,N_1240);
nor U2796 (N_2796,N_1068,N_1239);
or U2797 (N_2797,N_1483,N_1934);
nor U2798 (N_2798,N_1231,N_1976);
nand U2799 (N_2799,N_1655,N_1233);
nand U2800 (N_2800,N_1949,N_1841);
nand U2801 (N_2801,N_1877,N_1817);
xor U2802 (N_2802,N_1020,N_1202);
xor U2803 (N_2803,N_1144,N_1801);
nor U2804 (N_2804,N_1854,N_1382);
xnor U2805 (N_2805,N_1652,N_1666);
xor U2806 (N_2806,N_1251,N_1432);
xnor U2807 (N_2807,N_1015,N_1866);
or U2808 (N_2808,N_1739,N_1169);
or U2809 (N_2809,N_1864,N_1594);
and U2810 (N_2810,N_1280,N_1870);
xnor U2811 (N_2811,N_1379,N_1736);
nand U2812 (N_2812,N_1519,N_1489);
and U2813 (N_2813,N_1757,N_1582);
or U2814 (N_2814,N_1652,N_1782);
nand U2815 (N_2815,N_1202,N_1464);
and U2816 (N_2816,N_1429,N_1249);
and U2817 (N_2817,N_1248,N_1295);
nor U2818 (N_2818,N_1967,N_1957);
nor U2819 (N_2819,N_1207,N_1265);
nand U2820 (N_2820,N_1170,N_1658);
nand U2821 (N_2821,N_1903,N_1322);
or U2822 (N_2822,N_1451,N_1590);
nor U2823 (N_2823,N_1112,N_1098);
xor U2824 (N_2824,N_1030,N_1566);
nor U2825 (N_2825,N_1764,N_1498);
xnor U2826 (N_2826,N_1170,N_1138);
nand U2827 (N_2827,N_1780,N_1846);
and U2828 (N_2828,N_1365,N_1884);
nand U2829 (N_2829,N_1916,N_1524);
nand U2830 (N_2830,N_1220,N_1862);
xnor U2831 (N_2831,N_1398,N_1618);
nor U2832 (N_2832,N_1502,N_1075);
nand U2833 (N_2833,N_1471,N_1928);
nor U2834 (N_2834,N_1663,N_1106);
or U2835 (N_2835,N_1201,N_1666);
nand U2836 (N_2836,N_1574,N_1974);
or U2837 (N_2837,N_1940,N_1818);
and U2838 (N_2838,N_1513,N_1450);
xor U2839 (N_2839,N_1706,N_1642);
or U2840 (N_2840,N_1778,N_1155);
nand U2841 (N_2841,N_1125,N_1116);
and U2842 (N_2842,N_1467,N_1946);
nand U2843 (N_2843,N_1585,N_1309);
and U2844 (N_2844,N_1179,N_1612);
nor U2845 (N_2845,N_1108,N_1810);
and U2846 (N_2846,N_1904,N_1509);
xnor U2847 (N_2847,N_1870,N_1071);
nand U2848 (N_2848,N_1379,N_1437);
nand U2849 (N_2849,N_1325,N_1241);
nor U2850 (N_2850,N_1421,N_1002);
or U2851 (N_2851,N_1910,N_1007);
nor U2852 (N_2852,N_1254,N_1419);
and U2853 (N_2853,N_1653,N_1113);
nor U2854 (N_2854,N_1849,N_1521);
and U2855 (N_2855,N_1863,N_1492);
nor U2856 (N_2856,N_1826,N_1398);
xor U2857 (N_2857,N_1021,N_1626);
nand U2858 (N_2858,N_1689,N_1270);
nor U2859 (N_2859,N_1333,N_1205);
xnor U2860 (N_2860,N_1328,N_1394);
or U2861 (N_2861,N_1142,N_1010);
or U2862 (N_2862,N_1364,N_1374);
nor U2863 (N_2863,N_1479,N_1651);
xnor U2864 (N_2864,N_1897,N_1859);
or U2865 (N_2865,N_1836,N_1813);
and U2866 (N_2866,N_1943,N_1706);
xor U2867 (N_2867,N_1494,N_1310);
and U2868 (N_2868,N_1076,N_1185);
nand U2869 (N_2869,N_1428,N_1842);
and U2870 (N_2870,N_1444,N_1032);
and U2871 (N_2871,N_1862,N_1833);
or U2872 (N_2872,N_1346,N_1163);
xor U2873 (N_2873,N_1499,N_1065);
nor U2874 (N_2874,N_1949,N_1359);
and U2875 (N_2875,N_1011,N_1514);
and U2876 (N_2876,N_1634,N_1956);
xor U2877 (N_2877,N_1899,N_1972);
nor U2878 (N_2878,N_1580,N_1678);
or U2879 (N_2879,N_1212,N_1258);
or U2880 (N_2880,N_1589,N_1805);
xor U2881 (N_2881,N_1610,N_1059);
or U2882 (N_2882,N_1071,N_1333);
nand U2883 (N_2883,N_1728,N_1861);
or U2884 (N_2884,N_1775,N_1688);
or U2885 (N_2885,N_1810,N_1995);
or U2886 (N_2886,N_1106,N_1239);
and U2887 (N_2887,N_1045,N_1023);
and U2888 (N_2888,N_1389,N_1106);
nor U2889 (N_2889,N_1035,N_1745);
nand U2890 (N_2890,N_1598,N_1366);
or U2891 (N_2891,N_1270,N_1675);
or U2892 (N_2892,N_1805,N_1338);
or U2893 (N_2893,N_1337,N_1025);
nor U2894 (N_2894,N_1991,N_1971);
or U2895 (N_2895,N_1962,N_1018);
nand U2896 (N_2896,N_1851,N_1894);
xnor U2897 (N_2897,N_1199,N_1026);
and U2898 (N_2898,N_1081,N_1293);
xor U2899 (N_2899,N_1559,N_1715);
xor U2900 (N_2900,N_1572,N_1274);
xor U2901 (N_2901,N_1146,N_1144);
nor U2902 (N_2902,N_1066,N_1936);
and U2903 (N_2903,N_1570,N_1544);
xnor U2904 (N_2904,N_1427,N_1455);
nor U2905 (N_2905,N_1339,N_1110);
and U2906 (N_2906,N_1951,N_1073);
nor U2907 (N_2907,N_1287,N_1353);
xor U2908 (N_2908,N_1402,N_1268);
or U2909 (N_2909,N_1921,N_1955);
nor U2910 (N_2910,N_1122,N_1180);
or U2911 (N_2911,N_1284,N_1481);
nor U2912 (N_2912,N_1913,N_1532);
nor U2913 (N_2913,N_1304,N_1544);
and U2914 (N_2914,N_1232,N_1887);
nand U2915 (N_2915,N_1088,N_1222);
and U2916 (N_2916,N_1678,N_1362);
nand U2917 (N_2917,N_1206,N_1236);
or U2918 (N_2918,N_1993,N_1784);
and U2919 (N_2919,N_1686,N_1364);
nor U2920 (N_2920,N_1239,N_1942);
or U2921 (N_2921,N_1488,N_1967);
and U2922 (N_2922,N_1682,N_1998);
nand U2923 (N_2923,N_1269,N_1623);
and U2924 (N_2924,N_1994,N_1134);
nor U2925 (N_2925,N_1329,N_1263);
or U2926 (N_2926,N_1568,N_1033);
nor U2927 (N_2927,N_1537,N_1963);
nor U2928 (N_2928,N_1270,N_1060);
and U2929 (N_2929,N_1164,N_1890);
and U2930 (N_2930,N_1506,N_1510);
nor U2931 (N_2931,N_1482,N_1485);
or U2932 (N_2932,N_1101,N_1919);
or U2933 (N_2933,N_1975,N_1233);
or U2934 (N_2934,N_1718,N_1532);
nand U2935 (N_2935,N_1975,N_1941);
nor U2936 (N_2936,N_1815,N_1524);
nor U2937 (N_2937,N_1227,N_1653);
or U2938 (N_2938,N_1476,N_1739);
or U2939 (N_2939,N_1713,N_1632);
or U2940 (N_2940,N_1586,N_1666);
nand U2941 (N_2941,N_1725,N_1510);
or U2942 (N_2942,N_1713,N_1331);
xnor U2943 (N_2943,N_1110,N_1543);
nor U2944 (N_2944,N_1247,N_1584);
and U2945 (N_2945,N_1226,N_1756);
nor U2946 (N_2946,N_1185,N_1182);
or U2947 (N_2947,N_1508,N_1346);
xnor U2948 (N_2948,N_1711,N_1532);
and U2949 (N_2949,N_1840,N_1000);
nand U2950 (N_2950,N_1154,N_1201);
nor U2951 (N_2951,N_1926,N_1548);
xnor U2952 (N_2952,N_1817,N_1841);
nand U2953 (N_2953,N_1164,N_1500);
and U2954 (N_2954,N_1471,N_1578);
nor U2955 (N_2955,N_1309,N_1871);
nor U2956 (N_2956,N_1152,N_1164);
nor U2957 (N_2957,N_1479,N_1994);
nor U2958 (N_2958,N_1434,N_1219);
or U2959 (N_2959,N_1351,N_1684);
nand U2960 (N_2960,N_1888,N_1924);
and U2961 (N_2961,N_1307,N_1503);
xnor U2962 (N_2962,N_1989,N_1693);
xnor U2963 (N_2963,N_1973,N_1056);
nor U2964 (N_2964,N_1325,N_1050);
xnor U2965 (N_2965,N_1993,N_1222);
nor U2966 (N_2966,N_1839,N_1558);
and U2967 (N_2967,N_1545,N_1877);
xor U2968 (N_2968,N_1094,N_1264);
and U2969 (N_2969,N_1670,N_1261);
nand U2970 (N_2970,N_1778,N_1126);
nor U2971 (N_2971,N_1815,N_1099);
nor U2972 (N_2972,N_1689,N_1525);
nand U2973 (N_2973,N_1259,N_1835);
nor U2974 (N_2974,N_1445,N_1156);
nor U2975 (N_2975,N_1615,N_1183);
and U2976 (N_2976,N_1303,N_1085);
xor U2977 (N_2977,N_1162,N_1728);
and U2978 (N_2978,N_1341,N_1800);
or U2979 (N_2979,N_1681,N_1534);
and U2980 (N_2980,N_1076,N_1431);
xnor U2981 (N_2981,N_1734,N_1395);
nand U2982 (N_2982,N_1928,N_1576);
xnor U2983 (N_2983,N_1606,N_1028);
xor U2984 (N_2984,N_1178,N_1833);
or U2985 (N_2985,N_1814,N_1216);
and U2986 (N_2986,N_1901,N_1790);
nand U2987 (N_2987,N_1943,N_1740);
or U2988 (N_2988,N_1538,N_1141);
and U2989 (N_2989,N_1173,N_1267);
or U2990 (N_2990,N_1261,N_1970);
and U2991 (N_2991,N_1245,N_1890);
nor U2992 (N_2992,N_1826,N_1336);
nor U2993 (N_2993,N_1485,N_1565);
and U2994 (N_2994,N_1394,N_1148);
xnor U2995 (N_2995,N_1925,N_1945);
and U2996 (N_2996,N_1962,N_1246);
xor U2997 (N_2997,N_1658,N_1167);
nor U2998 (N_2998,N_1280,N_1867);
nor U2999 (N_2999,N_1477,N_1727);
xor U3000 (N_3000,N_2352,N_2659);
or U3001 (N_3001,N_2077,N_2584);
or U3002 (N_3002,N_2489,N_2680);
nand U3003 (N_3003,N_2941,N_2065);
and U3004 (N_3004,N_2518,N_2287);
or U3005 (N_3005,N_2530,N_2856);
or U3006 (N_3006,N_2995,N_2138);
nor U3007 (N_3007,N_2321,N_2638);
xnor U3008 (N_3008,N_2246,N_2688);
nand U3009 (N_3009,N_2763,N_2203);
and U3010 (N_3010,N_2987,N_2345);
and U3011 (N_3011,N_2308,N_2340);
nand U3012 (N_3012,N_2473,N_2544);
and U3013 (N_3013,N_2312,N_2209);
or U3014 (N_3014,N_2719,N_2961);
and U3015 (N_3015,N_2061,N_2270);
or U3016 (N_3016,N_2366,N_2132);
xor U3017 (N_3017,N_2798,N_2505);
and U3018 (N_3018,N_2152,N_2539);
nor U3019 (N_3019,N_2383,N_2319);
nor U3020 (N_3020,N_2029,N_2647);
and U3021 (N_3021,N_2067,N_2254);
nor U3022 (N_3022,N_2656,N_2020);
or U3023 (N_3023,N_2674,N_2202);
xor U3024 (N_3024,N_2349,N_2055);
nor U3025 (N_3025,N_2697,N_2780);
nand U3026 (N_3026,N_2163,N_2162);
nand U3027 (N_3027,N_2429,N_2956);
nand U3028 (N_3028,N_2315,N_2768);
xor U3029 (N_3029,N_2420,N_2470);
or U3030 (N_3030,N_2347,N_2227);
nand U3031 (N_3031,N_2616,N_2859);
or U3032 (N_3032,N_2236,N_2015);
xnor U3033 (N_3033,N_2170,N_2298);
xnor U3034 (N_3034,N_2490,N_2915);
nor U3035 (N_3035,N_2813,N_2288);
and U3036 (N_3036,N_2853,N_2501);
or U3037 (N_3037,N_2343,N_2376);
and U3038 (N_3038,N_2750,N_2089);
nor U3039 (N_3039,N_2538,N_2219);
nor U3040 (N_3040,N_2186,N_2592);
and U3041 (N_3041,N_2271,N_2979);
nand U3042 (N_3042,N_2633,N_2892);
xnor U3043 (N_3043,N_2854,N_2278);
nor U3044 (N_3044,N_2223,N_2789);
xor U3045 (N_3045,N_2706,N_2043);
xor U3046 (N_3046,N_2191,N_2310);
xor U3047 (N_3047,N_2985,N_2272);
xnor U3048 (N_3048,N_2147,N_2864);
nand U3049 (N_3049,N_2895,N_2040);
or U3050 (N_3050,N_2556,N_2927);
and U3051 (N_3051,N_2369,N_2066);
nand U3052 (N_3052,N_2078,N_2670);
and U3053 (N_3053,N_2705,N_2788);
and U3054 (N_3054,N_2189,N_2106);
and U3055 (N_3055,N_2962,N_2877);
nand U3056 (N_3056,N_2244,N_2013);
and U3057 (N_3057,N_2045,N_2965);
and U3058 (N_3058,N_2689,N_2296);
and U3059 (N_3059,N_2211,N_2590);
xor U3060 (N_3060,N_2199,N_2739);
nand U3061 (N_3061,N_2918,N_2461);
xnor U3062 (N_3062,N_2615,N_2654);
and U3063 (N_3063,N_2621,N_2221);
nor U3064 (N_3064,N_2041,N_2741);
nor U3065 (N_3065,N_2491,N_2603);
and U3066 (N_3066,N_2746,N_2800);
and U3067 (N_3067,N_2125,N_2431);
nor U3068 (N_3068,N_2586,N_2515);
or U3069 (N_3069,N_2107,N_2377);
and U3070 (N_3070,N_2939,N_2607);
and U3071 (N_3071,N_2392,N_2997);
nand U3072 (N_3072,N_2032,N_2213);
nand U3073 (N_3073,N_2970,N_2000);
nand U3074 (N_3074,N_2806,N_2049);
nor U3075 (N_3075,N_2946,N_2721);
and U3076 (N_3076,N_2968,N_2687);
and U3077 (N_3077,N_2086,N_2472);
and U3078 (N_3078,N_2925,N_2198);
xnor U3079 (N_3079,N_2795,N_2857);
nor U3080 (N_3080,N_2494,N_2649);
nand U3081 (N_3081,N_2467,N_2591);
nand U3082 (N_3082,N_2880,N_2164);
or U3083 (N_3083,N_2963,N_2699);
or U3084 (N_3084,N_2757,N_2333);
and U3085 (N_3085,N_2154,N_2993);
nor U3086 (N_3086,N_2222,N_2532);
xnor U3087 (N_3087,N_2974,N_2861);
xor U3088 (N_3088,N_2560,N_2943);
and U3089 (N_3089,N_2456,N_2942);
nand U3090 (N_3090,N_2522,N_2713);
and U3091 (N_3091,N_2819,N_2835);
nand U3092 (N_3092,N_2769,N_2128);
xor U3093 (N_3093,N_2338,N_2093);
or U3094 (N_3094,N_2930,N_2146);
nor U3095 (N_3095,N_2401,N_2373);
or U3096 (N_3096,N_2513,N_2365);
and U3097 (N_3097,N_2282,N_2975);
xnor U3098 (N_3098,N_2671,N_2395);
nor U3099 (N_3099,N_2869,N_2945);
xor U3100 (N_3100,N_2003,N_2669);
nor U3101 (N_3101,N_2335,N_2393);
and U3102 (N_3102,N_2818,N_2088);
xnor U3103 (N_3103,N_2953,N_2762);
or U3104 (N_3104,N_2541,N_2949);
nor U3105 (N_3105,N_2458,N_2173);
nand U3106 (N_3106,N_2053,N_2973);
nand U3107 (N_3107,N_2115,N_2430);
nor U3108 (N_3108,N_2736,N_2822);
or U3109 (N_3109,N_2913,N_2749);
or U3110 (N_3110,N_2837,N_2150);
nor U3111 (N_3111,N_2573,N_2572);
nand U3112 (N_3112,N_2954,N_2731);
or U3113 (N_3113,N_2039,N_2155);
nor U3114 (N_3114,N_2109,N_2242);
nand U3115 (N_3115,N_2655,N_2339);
xor U3116 (N_3116,N_2113,N_2710);
xnor U3117 (N_3117,N_2047,N_2225);
and U3118 (N_3118,N_2714,N_2433);
and U3119 (N_3119,N_2112,N_2496);
nor U3120 (N_3120,N_2253,N_2667);
nand U3121 (N_3121,N_2156,N_2509);
and U3122 (N_3122,N_2909,N_2297);
nor U3123 (N_3123,N_2836,N_2240);
and U3124 (N_3124,N_2384,N_2305);
nand U3125 (N_3125,N_2397,N_2883);
nor U3126 (N_3126,N_2627,N_2998);
nand U3127 (N_3127,N_2529,N_2448);
and U3128 (N_3128,N_2723,N_2600);
nand U3129 (N_3129,N_2428,N_2964);
nand U3130 (N_3130,N_2829,N_2921);
and U3131 (N_3131,N_2755,N_2525);
or U3132 (N_3132,N_2481,N_2237);
xor U3133 (N_3133,N_2177,N_2465);
xor U3134 (N_3134,N_2809,N_2385);
nand U3135 (N_3135,N_2716,N_2104);
nand U3136 (N_3136,N_2309,N_2738);
xor U3137 (N_3137,N_2359,N_2416);
and U3138 (N_3138,N_2797,N_2380);
and U3139 (N_3139,N_2482,N_2890);
and U3140 (N_3140,N_2404,N_2069);
and U3141 (N_3141,N_2601,N_2062);
nor U3142 (N_3142,N_2438,N_2151);
nand U3143 (N_3143,N_2764,N_2052);
or U3144 (N_3144,N_2702,N_2368);
and U3145 (N_3145,N_2210,N_2316);
or U3146 (N_3146,N_2311,N_2348);
and U3147 (N_3147,N_2457,N_2639);
nor U3148 (N_3148,N_2988,N_2082);
nor U3149 (N_3149,N_2231,N_2855);
nor U3150 (N_3150,N_2666,N_2087);
nor U3151 (N_3151,N_2098,N_2631);
or U3152 (N_3152,N_2827,N_2785);
and U3153 (N_3153,N_2274,N_2678);
xor U3154 (N_3154,N_2512,N_2924);
or U3155 (N_3155,N_2172,N_2766);
nor U3156 (N_3156,N_2537,N_2224);
and U3157 (N_3157,N_2017,N_2907);
or U3158 (N_3158,N_2761,N_2139);
or U3159 (N_3159,N_2387,N_2056);
nand U3160 (N_3160,N_2823,N_2117);
xor U3161 (N_3161,N_2881,N_2035);
and U3162 (N_3162,N_2684,N_2767);
nand U3163 (N_3163,N_2578,N_2418);
nor U3164 (N_3164,N_2743,N_2459);
nor U3165 (N_3165,N_2449,N_2097);
and U3166 (N_3166,N_2928,N_2576);
or U3167 (N_3167,N_2703,N_2846);
nand U3168 (N_3168,N_2228,N_2123);
xnor U3169 (N_3169,N_2059,N_2682);
or U3170 (N_3170,N_2821,N_2011);
nor U3171 (N_3171,N_2405,N_2722);
nor U3172 (N_3172,N_2858,N_2447);
nor U3173 (N_3173,N_2364,N_2103);
nor U3174 (N_3174,N_2137,N_2134);
nor U3175 (N_3175,N_2614,N_2337);
nand U3176 (N_3176,N_2570,N_2632);
nand U3177 (N_3177,N_2101,N_2452);
or U3178 (N_3178,N_2265,N_2552);
and U3179 (N_3179,N_2903,N_2374);
or U3180 (N_3180,N_2812,N_2516);
and U3181 (N_3181,N_2068,N_2840);
nor U3182 (N_3182,N_2398,N_2412);
or U3183 (N_3183,N_2476,N_2732);
xor U3184 (N_3184,N_2197,N_2026);
or U3185 (N_3185,N_2502,N_2808);
or U3186 (N_3186,N_2643,N_2843);
nor U3187 (N_3187,N_2183,N_2712);
nor U3188 (N_3188,N_2867,N_2596);
or U3189 (N_3189,N_2446,N_2024);
or U3190 (N_3190,N_2866,N_2971);
or U3191 (N_3191,N_2126,N_2933);
and U3192 (N_3192,N_2326,N_2926);
xnor U3193 (N_3193,N_2510,N_2526);
xor U3194 (N_3194,N_2775,N_2980);
nand U3195 (N_3195,N_2388,N_2317);
nand U3196 (N_3196,N_2188,N_2878);
nor U3197 (N_3197,N_2568,N_2329);
or U3198 (N_3198,N_2765,N_2451);
and U3199 (N_3199,N_2293,N_2092);
xnor U3200 (N_3200,N_2229,N_2302);
xor U3201 (N_3201,N_2791,N_2874);
nand U3202 (N_3202,N_2929,N_2543);
and U3203 (N_3203,N_2645,N_2200);
and U3204 (N_3204,N_2790,N_2406);
or U3205 (N_3205,N_2624,N_2220);
nor U3206 (N_3206,N_2937,N_2218);
xnor U3207 (N_3207,N_2102,N_2114);
and U3208 (N_3208,N_2175,N_2266);
or U3209 (N_3209,N_2916,N_2834);
nand U3210 (N_3210,N_2331,N_2807);
or U3211 (N_3211,N_2178,N_2038);
nor U3212 (N_3212,N_2625,N_2728);
or U3213 (N_3213,N_2204,N_2908);
xnor U3214 (N_3214,N_2740,N_2653);
nor U3215 (N_3215,N_2528,N_2161);
xor U3216 (N_3216,N_2262,N_2334);
nand U3217 (N_3217,N_2990,N_2579);
nand U3218 (N_3218,N_2439,N_2399);
and U3219 (N_3219,N_2677,N_2517);
xor U3220 (N_3220,N_2497,N_2118);
xnor U3221 (N_3221,N_2711,N_2196);
or U3222 (N_3222,N_2410,N_2546);
nand U3223 (N_3223,N_2460,N_2136);
xnor U3224 (N_3224,N_2727,N_2910);
nand U3225 (N_3225,N_2493,N_2742);
and U3226 (N_3226,N_2879,N_2773);
xnor U3227 (N_3227,N_2286,N_2028);
nand U3228 (N_3228,N_2332,N_2730);
or U3229 (N_3229,N_2301,N_2390);
nand U3230 (N_3230,N_2724,N_2850);
nor U3231 (N_3231,N_2176,N_2935);
or U3232 (N_3232,N_2779,N_2717);
or U3233 (N_3233,N_2900,N_2094);
and U3234 (N_3234,N_2803,N_2726);
nor U3235 (N_3235,N_2683,N_2378);
nor U3236 (N_3236,N_2421,N_2063);
or U3237 (N_3237,N_2976,N_2842);
or U3238 (N_3238,N_2499,N_2676);
or U3239 (N_3239,N_2665,N_2872);
and U3240 (N_3240,N_2432,N_2661);
nor U3241 (N_3241,N_2356,N_2434);
or U3242 (N_3242,N_2205,N_2201);
xor U3243 (N_3243,N_2708,N_2805);
nand U3244 (N_3244,N_2241,N_2969);
xor U3245 (N_3245,N_2450,N_2613);
xor U3246 (N_3246,N_2885,N_2897);
and U3247 (N_3247,N_2520,N_2245);
and U3248 (N_3248,N_2932,N_2257);
nand U3249 (N_3249,N_2193,N_2816);
or U3250 (N_3250,N_2644,N_2079);
nand U3251 (N_3251,N_2230,N_2259);
or U3252 (N_3252,N_2873,N_2381);
nor U3253 (N_3253,N_2948,N_2190);
nor U3254 (N_3254,N_2777,N_2046);
and U3255 (N_3255,N_2238,N_2917);
nand U3256 (N_3256,N_2184,N_2119);
nor U3257 (N_3257,N_2820,N_2951);
and U3258 (N_3258,N_2022,N_2549);
and U3259 (N_3259,N_2108,N_2617);
xor U3260 (N_3260,N_2307,N_2896);
nand U3261 (N_3261,N_2575,N_2025);
and U3262 (N_3262,N_2480,N_2208);
and U3263 (N_3263,N_2095,N_2700);
xor U3264 (N_3264,N_2783,N_2124);
and U3265 (N_3265,N_2707,N_2226);
and U3266 (N_3266,N_2582,N_2893);
and U3267 (N_3267,N_2804,N_2007);
xnor U3268 (N_3268,N_2720,N_2258);
nand U3269 (N_3269,N_2248,N_2121);
xor U3270 (N_3270,N_2991,N_2142);
xor U3271 (N_3271,N_2548,N_2127);
or U3272 (N_3272,N_2581,N_2547);
nand U3273 (N_3273,N_2511,N_2562);
or U3274 (N_3274,N_2363,N_2425);
nor U3275 (N_3275,N_2650,N_2160);
nand U3276 (N_3276,N_2264,N_2037);
nor U3277 (N_3277,N_2747,N_2021);
nor U3278 (N_3278,N_2981,N_2411);
and U3279 (N_3279,N_2394,N_2831);
nand U3280 (N_3280,N_2325,N_2474);
nand U3281 (N_3281,N_2535,N_2967);
or U3282 (N_3282,N_2851,N_2478);
xnor U3283 (N_3283,N_2811,N_2330);
nor U3284 (N_3284,N_2084,N_2533);
or U3285 (N_3285,N_2289,N_2466);
xnor U3286 (N_3286,N_2672,N_2565);
and U3287 (N_3287,N_2492,N_2623);
or U3288 (N_3288,N_2346,N_2044);
nor U3289 (N_3289,N_2408,N_2455);
and U3290 (N_3290,N_2634,N_2792);
nor U3291 (N_3291,N_2887,N_2781);
or U3292 (N_3292,N_2354,N_2758);
or U3293 (N_3293,N_2462,N_2978);
nand U3294 (N_3294,N_2986,N_2344);
and U3295 (N_3295,N_2646,N_2111);
or U3296 (N_3296,N_2542,N_2435);
nor U3297 (N_3297,N_2563,N_2580);
nand U3298 (N_3298,N_2648,N_2477);
nand U3299 (N_3299,N_2904,N_2888);
xnor U3300 (N_3300,N_2534,N_2195);
and U3301 (N_3301,N_2396,N_2691);
or U3302 (N_3302,N_2604,N_2367);
nand U3303 (N_3303,N_2770,N_2774);
nand U3304 (N_3304,N_2751,N_2794);
and U3305 (N_3305,N_2566,N_2445);
xor U3306 (N_3306,N_2507,N_2135);
nor U3307 (N_3307,N_2336,N_2415);
nand U3308 (N_3308,N_2994,N_2718);
nor U3309 (N_3309,N_2860,N_2235);
nor U3310 (N_3310,N_2830,N_2793);
nor U3311 (N_3311,N_2891,N_2865);
xnor U3312 (N_3312,N_2166,N_2051);
nand U3313 (N_3313,N_2207,N_2357);
or U3314 (N_3314,N_2099,N_2744);
or U3315 (N_3315,N_2149,N_2070);
nand U3316 (N_3316,N_2839,N_2372);
and U3317 (N_3317,N_2558,N_2267);
nand U3318 (N_3318,N_2622,N_2734);
or U3319 (N_3319,N_2403,N_2484);
xor U3320 (N_3320,N_2630,N_2567);
nor U3321 (N_3321,N_2685,N_2692);
xnor U3322 (N_3322,N_2555,N_2847);
nor U3323 (N_3323,N_2523,N_2353);
nand U3324 (N_3324,N_2012,N_2849);
and U3325 (N_3325,N_2171,N_2360);
nor U3326 (N_3326,N_2826,N_2260);
nor U3327 (N_3327,N_2848,N_2402);
xnor U3328 (N_3328,N_2972,N_2778);
xor U3329 (N_3329,N_2427,N_2938);
or U3330 (N_3330,N_2503,N_2468);
xnor U3331 (N_3331,N_2009,N_2027);
and U3332 (N_3332,N_2469,N_2075);
xnor U3333 (N_3333,N_2002,N_2275);
nor U3334 (N_3334,N_2693,N_2824);
or U3335 (N_3335,N_2561,N_2524);
nor U3336 (N_3336,N_2414,N_2610);
xor U3337 (N_3337,N_2030,N_2959);
xnor U3338 (N_3338,N_2324,N_2194);
nor U3339 (N_3339,N_2290,N_2914);
nor U3340 (N_3340,N_2249,N_2626);
nand U3341 (N_3341,N_2168,N_2276);
nand U3342 (N_3342,N_2375,N_2096);
nor U3343 (N_3343,N_2153,N_2681);
and U3344 (N_3344,N_2679,N_2071);
or U3345 (N_3345,N_2799,N_2611);
nand U3346 (N_3346,N_2725,N_2400);
xnor U3347 (N_3347,N_2844,N_2852);
nand U3348 (N_3348,N_2361,N_2080);
and U3349 (N_3349,N_2033,N_2014);
nor U3350 (N_3350,N_2306,N_2922);
and U3351 (N_3351,N_2299,N_2899);
xnor U3352 (N_3352,N_2355,N_2673);
nand U3353 (N_3353,N_2637,N_2608);
xor U3354 (N_3354,N_2090,N_2008);
xor U3355 (N_3355,N_2612,N_2825);
or U3356 (N_3356,N_2105,N_2871);
and U3357 (N_3357,N_2001,N_2192);
nand U3358 (N_3358,N_2074,N_2652);
nor U3359 (N_3359,N_2232,N_2342);
xor U3360 (N_3360,N_2181,N_2754);
or U3361 (N_3361,N_2016,N_2906);
and U3362 (N_3362,N_2690,N_2145);
nor U3363 (N_3363,N_2072,N_2569);
and U3364 (N_3364,N_2748,N_2386);
xnor U3365 (N_3365,N_2058,N_2379);
nor U3366 (N_3366,N_2060,N_2983);
and U3367 (N_3367,N_2179,N_2919);
nor U3368 (N_3368,N_2081,N_2180);
xor U3369 (N_3369,N_2409,N_2815);
nand U3370 (N_3370,N_2550,N_2629);
xor U3371 (N_3371,N_2782,N_2701);
and U3372 (N_3372,N_2894,N_2905);
nand U3373 (N_3373,N_2784,N_2863);
and U3374 (N_3374,N_2141,N_2483);
and U3375 (N_3375,N_2327,N_2268);
xnor U3376 (N_3376,N_2944,N_2495);
nand U3377 (N_3377,N_2771,N_2958);
or U3378 (N_3378,N_2144,N_2527);
nand U3379 (N_3379,N_2531,N_2735);
nor U3380 (N_3380,N_2174,N_2454);
xnor U3381 (N_3381,N_2553,N_2057);
or U3382 (N_3382,N_2609,N_2845);
nand U3383 (N_3383,N_2989,N_2802);
or U3384 (N_3384,N_2931,N_2992);
or U3385 (N_3385,N_2841,N_2422);
or U3386 (N_3386,N_2585,N_2709);
and U3387 (N_3387,N_2588,N_2261);
nor U3388 (N_3388,N_2441,N_2294);
nor U3389 (N_3389,N_2698,N_2322);
nor U3390 (N_3390,N_2216,N_2912);
xor U3391 (N_3391,N_2642,N_2911);
nor U3392 (N_3392,N_2696,N_2559);
nand U3393 (N_3393,N_2577,N_2129);
or U3394 (N_3394,N_2436,N_2320);
or U3395 (N_3395,N_2966,N_2048);
nand U3396 (N_3396,N_2660,N_2628);
or U3397 (N_3397,N_2362,N_2950);
and U3398 (N_3398,N_2413,N_2838);
xnor U3399 (N_3399,N_2463,N_2143);
and U3400 (N_3400,N_2551,N_2514);
nor U3401 (N_3401,N_2817,N_2557);
nand U3402 (N_3402,N_2437,N_2382);
nand U3403 (N_3403,N_2488,N_2923);
nor U3404 (N_3404,N_2733,N_2370);
nand U3405 (N_3405,N_2752,N_2471);
xnor U3406 (N_3406,N_2187,N_2955);
and U3407 (N_3407,N_2619,N_2957);
nor U3408 (N_3408,N_2704,N_2358);
nor U3409 (N_3409,N_2886,N_2295);
nor U3410 (N_3410,N_2982,N_2500);
nor U3411 (N_3411,N_2444,N_2256);
nand U3412 (N_3412,N_2110,N_2940);
or U3413 (N_3413,N_2263,N_2599);
nand U3414 (N_3414,N_2564,N_2285);
or U3415 (N_3415,N_2876,N_2371);
and U3416 (N_3416,N_2594,N_2587);
and U3417 (N_3417,N_2745,N_2443);
and U3418 (N_3418,N_2884,N_2250);
nand U3419 (N_3419,N_2116,N_2508);
and U3420 (N_3420,N_2323,N_2636);
or U3421 (N_3421,N_2485,N_2602);
xor U3422 (N_3422,N_2091,N_2148);
xor U3423 (N_3423,N_2936,N_2658);
xor U3424 (N_3424,N_2595,N_2269);
nand U3425 (N_3425,N_2999,N_2291);
nor U3426 (N_3426,N_2640,N_2389);
nor U3427 (N_3427,N_2391,N_2214);
and U3428 (N_3428,N_2277,N_2487);
nand U3429 (N_3429,N_2977,N_2010);
nand U3430 (N_3430,N_2318,N_2165);
nand U3431 (N_3431,N_2018,N_2239);
or U3432 (N_3432,N_2233,N_2889);
xor U3433 (N_3433,N_2536,N_2423);
or U3434 (N_3434,N_2417,N_2054);
xnor U3435 (N_3435,N_2206,N_2131);
xor U3436 (N_3436,N_2292,N_2255);
xnor U3437 (N_3437,N_2212,N_2571);
and U3438 (N_3438,N_2952,N_2300);
or U3439 (N_3439,N_2498,N_2122);
xnor U3440 (N_3440,N_2668,N_2304);
and U3441 (N_3441,N_2664,N_2868);
and U3442 (N_3442,N_2050,N_2810);
and U3443 (N_3443,N_2169,N_2641);
nand U3444 (N_3444,N_2158,N_2901);
or U3445 (N_3445,N_2252,N_2635);
xor U3446 (N_3446,N_2984,N_2760);
or U3447 (N_3447,N_2759,N_2737);
nor U3448 (N_3448,N_2453,N_2217);
nand U3449 (N_3449,N_2545,N_2407);
xor U3450 (N_3450,N_2251,N_2756);
nor U3451 (N_3451,N_2247,N_2215);
xnor U3452 (N_3452,N_2440,N_2882);
xnor U3453 (N_3453,N_2833,N_2023);
xor U3454 (N_3454,N_2583,N_2157);
or U3455 (N_3455,N_2350,N_2620);
nand U3456 (N_3456,N_2920,N_2159);
nor U3457 (N_3457,N_2776,N_2540);
or U3458 (N_3458,N_2715,N_2651);
nand U3459 (N_3459,N_2303,N_2606);
nand U3460 (N_3460,N_2663,N_2934);
or U3461 (N_3461,N_2004,N_2694);
nor U3462 (N_3462,N_2006,N_2284);
or U3463 (N_3463,N_2589,N_2243);
and U3464 (N_3464,N_2280,N_2862);
nand U3465 (N_3465,N_2341,N_2351);
and U3466 (N_3466,N_2426,N_2947);
nand U3467 (N_3467,N_2475,N_2019);
or U3468 (N_3468,N_2424,N_2814);
nor U3469 (N_3469,N_2898,N_2167);
and U3470 (N_3470,N_2662,N_2519);
xnor U3471 (N_3471,N_2273,N_2073);
and U3472 (N_3472,N_2695,N_2828);
xnor U3473 (N_3473,N_2313,N_2100);
xor U3474 (N_3474,N_2064,N_2960);
nor U3475 (N_3475,N_2031,N_2486);
or U3476 (N_3476,N_2598,N_2076);
nor U3477 (N_3477,N_2506,N_2464);
xnor U3478 (N_3478,N_2832,N_2574);
nand U3479 (N_3479,N_2801,N_2729);
and U3480 (N_3480,N_2902,N_2140);
nand U3481 (N_3481,N_2870,N_2133);
nor U3482 (N_3482,N_2182,N_2120);
and U3483 (N_3483,N_2130,N_2675);
or U3484 (N_3484,N_2036,N_2796);
nand U3485 (N_3485,N_2787,N_2279);
and U3486 (N_3486,N_2597,N_2314);
and U3487 (N_3487,N_2042,N_2786);
nor U3488 (N_3488,N_2504,N_2085);
xor U3489 (N_3489,N_2479,N_2005);
or U3490 (N_3490,N_2593,N_2234);
xor U3491 (N_3491,N_2521,N_2772);
and U3492 (N_3492,N_2034,N_2605);
or U3493 (N_3493,N_2328,N_2657);
nand U3494 (N_3494,N_2618,N_2185);
nand U3495 (N_3495,N_2753,N_2281);
nor U3496 (N_3496,N_2875,N_2686);
nand U3497 (N_3497,N_2419,N_2283);
nor U3498 (N_3498,N_2083,N_2554);
xor U3499 (N_3499,N_2996,N_2442);
and U3500 (N_3500,N_2030,N_2589);
xor U3501 (N_3501,N_2156,N_2334);
xnor U3502 (N_3502,N_2824,N_2887);
or U3503 (N_3503,N_2418,N_2967);
nand U3504 (N_3504,N_2423,N_2612);
xor U3505 (N_3505,N_2762,N_2219);
nor U3506 (N_3506,N_2010,N_2719);
and U3507 (N_3507,N_2818,N_2875);
and U3508 (N_3508,N_2855,N_2913);
nor U3509 (N_3509,N_2610,N_2044);
nand U3510 (N_3510,N_2661,N_2626);
nor U3511 (N_3511,N_2062,N_2143);
or U3512 (N_3512,N_2467,N_2980);
and U3513 (N_3513,N_2440,N_2817);
nand U3514 (N_3514,N_2398,N_2171);
and U3515 (N_3515,N_2432,N_2447);
nand U3516 (N_3516,N_2999,N_2237);
nor U3517 (N_3517,N_2973,N_2142);
xor U3518 (N_3518,N_2561,N_2706);
nor U3519 (N_3519,N_2064,N_2920);
nand U3520 (N_3520,N_2934,N_2380);
xnor U3521 (N_3521,N_2879,N_2515);
nor U3522 (N_3522,N_2860,N_2274);
nand U3523 (N_3523,N_2090,N_2510);
nand U3524 (N_3524,N_2326,N_2749);
or U3525 (N_3525,N_2550,N_2640);
nor U3526 (N_3526,N_2405,N_2558);
xnor U3527 (N_3527,N_2598,N_2496);
and U3528 (N_3528,N_2056,N_2911);
nand U3529 (N_3529,N_2803,N_2990);
xnor U3530 (N_3530,N_2491,N_2141);
nor U3531 (N_3531,N_2406,N_2942);
nor U3532 (N_3532,N_2709,N_2488);
or U3533 (N_3533,N_2430,N_2180);
and U3534 (N_3534,N_2018,N_2442);
and U3535 (N_3535,N_2846,N_2225);
and U3536 (N_3536,N_2200,N_2631);
and U3537 (N_3537,N_2011,N_2345);
or U3538 (N_3538,N_2612,N_2410);
and U3539 (N_3539,N_2856,N_2828);
nand U3540 (N_3540,N_2230,N_2995);
nand U3541 (N_3541,N_2126,N_2474);
and U3542 (N_3542,N_2526,N_2330);
and U3543 (N_3543,N_2681,N_2010);
nand U3544 (N_3544,N_2955,N_2938);
nand U3545 (N_3545,N_2309,N_2873);
and U3546 (N_3546,N_2520,N_2678);
nor U3547 (N_3547,N_2064,N_2175);
or U3548 (N_3548,N_2362,N_2027);
nand U3549 (N_3549,N_2456,N_2185);
nand U3550 (N_3550,N_2694,N_2873);
or U3551 (N_3551,N_2081,N_2221);
and U3552 (N_3552,N_2976,N_2644);
nand U3553 (N_3553,N_2373,N_2363);
or U3554 (N_3554,N_2917,N_2358);
or U3555 (N_3555,N_2279,N_2702);
nor U3556 (N_3556,N_2181,N_2498);
xnor U3557 (N_3557,N_2932,N_2876);
and U3558 (N_3558,N_2926,N_2244);
and U3559 (N_3559,N_2248,N_2565);
and U3560 (N_3560,N_2973,N_2825);
and U3561 (N_3561,N_2944,N_2074);
and U3562 (N_3562,N_2623,N_2526);
nand U3563 (N_3563,N_2158,N_2990);
or U3564 (N_3564,N_2787,N_2033);
xnor U3565 (N_3565,N_2526,N_2160);
nand U3566 (N_3566,N_2934,N_2081);
and U3567 (N_3567,N_2530,N_2318);
and U3568 (N_3568,N_2000,N_2625);
or U3569 (N_3569,N_2471,N_2407);
nand U3570 (N_3570,N_2408,N_2879);
xnor U3571 (N_3571,N_2537,N_2221);
nand U3572 (N_3572,N_2210,N_2642);
nand U3573 (N_3573,N_2064,N_2761);
nor U3574 (N_3574,N_2810,N_2911);
nor U3575 (N_3575,N_2211,N_2142);
xnor U3576 (N_3576,N_2787,N_2458);
nand U3577 (N_3577,N_2705,N_2860);
and U3578 (N_3578,N_2621,N_2273);
or U3579 (N_3579,N_2123,N_2344);
or U3580 (N_3580,N_2948,N_2060);
and U3581 (N_3581,N_2985,N_2194);
nor U3582 (N_3582,N_2392,N_2373);
or U3583 (N_3583,N_2256,N_2583);
nand U3584 (N_3584,N_2775,N_2852);
and U3585 (N_3585,N_2023,N_2870);
nand U3586 (N_3586,N_2275,N_2173);
and U3587 (N_3587,N_2478,N_2777);
nand U3588 (N_3588,N_2156,N_2142);
nand U3589 (N_3589,N_2382,N_2953);
and U3590 (N_3590,N_2778,N_2837);
nand U3591 (N_3591,N_2852,N_2893);
or U3592 (N_3592,N_2753,N_2519);
and U3593 (N_3593,N_2774,N_2321);
nor U3594 (N_3594,N_2510,N_2674);
or U3595 (N_3595,N_2503,N_2206);
or U3596 (N_3596,N_2451,N_2233);
or U3597 (N_3597,N_2371,N_2072);
nand U3598 (N_3598,N_2748,N_2328);
nand U3599 (N_3599,N_2160,N_2473);
xor U3600 (N_3600,N_2266,N_2960);
or U3601 (N_3601,N_2196,N_2370);
or U3602 (N_3602,N_2603,N_2428);
nor U3603 (N_3603,N_2831,N_2227);
xor U3604 (N_3604,N_2496,N_2918);
nor U3605 (N_3605,N_2338,N_2289);
or U3606 (N_3606,N_2959,N_2512);
and U3607 (N_3607,N_2259,N_2858);
nand U3608 (N_3608,N_2805,N_2234);
xor U3609 (N_3609,N_2560,N_2238);
nor U3610 (N_3610,N_2543,N_2246);
xnor U3611 (N_3611,N_2754,N_2037);
nor U3612 (N_3612,N_2716,N_2154);
and U3613 (N_3613,N_2422,N_2391);
xor U3614 (N_3614,N_2274,N_2704);
and U3615 (N_3615,N_2405,N_2495);
nand U3616 (N_3616,N_2483,N_2641);
nand U3617 (N_3617,N_2207,N_2551);
and U3618 (N_3618,N_2581,N_2446);
xnor U3619 (N_3619,N_2240,N_2136);
nor U3620 (N_3620,N_2920,N_2205);
nand U3621 (N_3621,N_2827,N_2237);
nand U3622 (N_3622,N_2946,N_2407);
xor U3623 (N_3623,N_2129,N_2448);
xor U3624 (N_3624,N_2470,N_2528);
nor U3625 (N_3625,N_2990,N_2951);
nor U3626 (N_3626,N_2394,N_2741);
nand U3627 (N_3627,N_2834,N_2935);
or U3628 (N_3628,N_2127,N_2593);
and U3629 (N_3629,N_2983,N_2698);
nand U3630 (N_3630,N_2106,N_2467);
nor U3631 (N_3631,N_2444,N_2580);
and U3632 (N_3632,N_2352,N_2466);
nor U3633 (N_3633,N_2125,N_2874);
nor U3634 (N_3634,N_2537,N_2203);
xor U3635 (N_3635,N_2387,N_2839);
nand U3636 (N_3636,N_2590,N_2548);
nor U3637 (N_3637,N_2487,N_2932);
xnor U3638 (N_3638,N_2308,N_2680);
and U3639 (N_3639,N_2528,N_2501);
or U3640 (N_3640,N_2199,N_2805);
nand U3641 (N_3641,N_2356,N_2853);
nand U3642 (N_3642,N_2150,N_2374);
xnor U3643 (N_3643,N_2926,N_2606);
nor U3644 (N_3644,N_2432,N_2573);
xor U3645 (N_3645,N_2043,N_2338);
and U3646 (N_3646,N_2082,N_2125);
nand U3647 (N_3647,N_2277,N_2187);
and U3648 (N_3648,N_2831,N_2654);
xnor U3649 (N_3649,N_2260,N_2235);
nor U3650 (N_3650,N_2109,N_2224);
nand U3651 (N_3651,N_2926,N_2485);
nor U3652 (N_3652,N_2335,N_2943);
nor U3653 (N_3653,N_2532,N_2662);
or U3654 (N_3654,N_2004,N_2329);
nor U3655 (N_3655,N_2588,N_2355);
xor U3656 (N_3656,N_2588,N_2133);
and U3657 (N_3657,N_2345,N_2012);
xor U3658 (N_3658,N_2092,N_2284);
xnor U3659 (N_3659,N_2004,N_2823);
and U3660 (N_3660,N_2727,N_2161);
and U3661 (N_3661,N_2509,N_2202);
or U3662 (N_3662,N_2180,N_2988);
xor U3663 (N_3663,N_2284,N_2447);
nand U3664 (N_3664,N_2751,N_2558);
and U3665 (N_3665,N_2094,N_2189);
xnor U3666 (N_3666,N_2022,N_2421);
or U3667 (N_3667,N_2911,N_2212);
or U3668 (N_3668,N_2365,N_2912);
and U3669 (N_3669,N_2051,N_2432);
and U3670 (N_3670,N_2417,N_2402);
nor U3671 (N_3671,N_2955,N_2973);
or U3672 (N_3672,N_2164,N_2961);
xnor U3673 (N_3673,N_2854,N_2037);
or U3674 (N_3674,N_2013,N_2333);
nand U3675 (N_3675,N_2448,N_2723);
nor U3676 (N_3676,N_2407,N_2151);
or U3677 (N_3677,N_2004,N_2654);
nor U3678 (N_3678,N_2252,N_2582);
xnor U3679 (N_3679,N_2674,N_2764);
nor U3680 (N_3680,N_2604,N_2421);
nand U3681 (N_3681,N_2398,N_2718);
and U3682 (N_3682,N_2707,N_2877);
and U3683 (N_3683,N_2323,N_2607);
nand U3684 (N_3684,N_2301,N_2581);
xnor U3685 (N_3685,N_2753,N_2685);
nor U3686 (N_3686,N_2662,N_2812);
nand U3687 (N_3687,N_2632,N_2217);
xor U3688 (N_3688,N_2328,N_2887);
and U3689 (N_3689,N_2306,N_2800);
and U3690 (N_3690,N_2245,N_2887);
xnor U3691 (N_3691,N_2390,N_2543);
or U3692 (N_3692,N_2424,N_2857);
xor U3693 (N_3693,N_2767,N_2815);
or U3694 (N_3694,N_2224,N_2879);
or U3695 (N_3695,N_2590,N_2485);
xor U3696 (N_3696,N_2690,N_2142);
and U3697 (N_3697,N_2786,N_2696);
or U3698 (N_3698,N_2195,N_2269);
or U3699 (N_3699,N_2193,N_2512);
xnor U3700 (N_3700,N_2328,N_2860);
and U3701 (N_3701,N_2548,N_2044);
or U3702 (N_3702,N_2042,N_2743);
xor U3703 (N_3703,N_2538,N_2512);
and U3704 (N_3704,N_2154,N_2347);
nor U3705 (N_3705,N_2989,N_2790);
and U3706 (N_3706,N_2890,N_2286);
nor U3707 (N_3707,N_2334,N_2896);
xor U3708 (N_3708,N_2417,N_2707);
nor U3709 (N_3709,N_2311,N_2115);
nand U3710 (N_3710,N_2482,N_2213);
and U3711 (N_3711,N_2488,N_2999);
or U3712 (N_3712,N_2889,N_2347);
and U3713 (N_3713,N_2321,N_2838);
or U3714 (N_3714,N_2152,N_2479);
nor U3715 (N_3715,N_2756,N_2537);
or U3716 (N_3716,N_2010,N_2393);
xnor U3717 (N_3717,N_2948,N_2977);
and U3718 (N_3718,N_2514,N_2645);
xnor U3719 (N_3719,N_2409,N_2906);
nand U3720 (N_3720,N_2604,N_2039);
or U3721 (N_3721,N_2654,N_2900);
nor U3722 (N_3722,N_2222,N_2938);
xor U3723 (N_3723,N_2100,N_2186);
or U3724 (N_3724,N_2063,N_2497);
nor U3725 (N_3725,N_2901,N_2524);
or U3726 (N_3726,N_2128,N_2298);
xor U3727 (N_3727,N_2158,N_2052);
xnor U3728 (N_3728,N_2005,N_2443);
nor U3729 (N_3729,N_2676,N_2776);
and U3730 (N_3730,N_2254,N_2107);
nor U3731 (N_3731,N_2732,N_2894);
xor U3732 (N_3732,N_2260,N_2462);
nand U3733 (N_3733,N_2950,N_2467);
and U3734 (N_3734,N_2674,N_2000);
or U3735 (N_3735,N_2607,N_2989);
or U3736 (N_3736,N_2417,N_2264);
xnor U3737 (N_3737,N_2439,N_2869);
nor U3738 (N_3738,N_2268,N_2692);
nor U3739 (N_3739,N_2889,N_2920);
nor U3740 (N_3740,N_2284,N_2552);
nand U3741 (N_3741,N_2656,N_2626);
xnor U3742 (N_3742,N_2298,N_2898);
or U3743 (N_3743,N_2176,N_2469);
nand U3744 (N_3744,N_2372,N_2574);
or U3745 (N_3745,N_2238,N_2896);
nor U3746 (N_3746,N_2496,N_2025);
xor U3747 (N_3747,N_2104,N_2741);
xnor U3748 (N_3748,N_2268,N_2571);
xor U3749 (N_3749,N_2873,N_2128);
nor U3750 (N_3750,N_2570,N_2932);
nor U3751 (N_3751,N_2660,N_2176);
or U3752 (N_3752,N_2228,N_2815);
nand U3753 (N_3753,N_2379,N_2472);
xor U3754 (N_3754,N_2679,N_2756);
nor U3755 (N_3755,N_2448,N_2488);
xnor U3756 (N_3756,N_2859,N_2495);
and U3757 (N_3757,N_2232,N_2161);
and U3758 (N_3758,N_2698,N_2564);
xor U3759 (N_3759,N_2866,N_2565);
nand U3760 (N_3760,N_2811,N_2944);
xor U3761 (N_3761,N_2253,N_2474);
or U3762 (N_3762,N_2725,N_2642);
nand U3763 (N_3763,N_2107,N_2275);
xnor U3764 (N_3764,N_2298,N_2360);
nor U3765 (N_3765,N_2490,N_2203);
nand U3766 (N_3766,N_2164,N_2659);
or U3767 (N_3767,N_2294,N_2801);
xor U3768 (N_3768,N_2824,N_2665);
nand U3769 (N_3769,N_2366,N_2960);
nand U3770 (N_3770,N_2435,N_2127);
nor U3771 (N_3771,N_2897,N_2450);
nor U3772 (N_3772,N_2366,N_2003);
or U3773 (N_3773,N_2516,N_2600);
and U3774 (N_3774,N_2324,N_2465);
nor U3775 (N_3775,N_2993,N_2527);
xor U3776 (N_3776,N_2623,N_2058);
nor U3777 (N_3777,N_2200,N_2487);
nand U3778 (N_3778,N_2169,N_2555);
xor U3779 (N_3779,N_2623,N_2258);
or U3780 (N_3780,N_2469,N_2442);
nor U3781 (N_3781,N_2245,N_2391);
or U3782 (N_3782,N_2834,N_2906);
and U3783 (N_3783,N_2792,N_2537);
nand U3784 (N_3784,N_2501,N_2134);
or U3785 (N_3785,N_2489,N_2974);
or U3786 (N_3786,N_2798,N_2852);
xnor U3787 (N_3787,N_2316,N_2915);
nand U3788 (N_3788,N_2822,N_2048);
nand U3789 (N_3789,N_2769,N_2567);
xnor U3790 (N_3790,N_2829,N_2946);
nand U3791 (N_3791,N_2784,N_2246);
and U3792 (N_3792,N_2864,N_2322);
xnor U3793 (N_3793,N_2334,N_2793);
xnor U3794 (N_3794,N_2485,N_2878);
nor U3795 (N_3795,N_2484,N_2801);
nor U3796 (N_3796,N_2645,N_2496);
and U3797 (N_3797,N_2003,N_2218);
nand U3798 (N_3798,N_2385,N_2870);
nor U3799 (N_3799,N_2155,N_2479);
or U3800 (N_3800,N_2438,N_2777);
nor U3801 (N_3801,N_2572,N_2848);
nor U3802 (N_3802,N_2862,N_2593);
nor U3803 (N_3803,N_2990,N_2326);
and U3804 (N_3804,N_2340,N_2517);
xor U3805 (N_3805,N_2334,N_2698);
and U3806 (N_3806,N_2046,N_2505);
nand U3807 (N_3807,N_2001,N_2233);
nor U3808 (N_3808,N_2805,N_2212);
xnor U3809 (N_3809,N_2303,N_2513);
nor U3810 (N_3810,N_2172,N_2955);
and U3811 (N_3811,N_2170,N_2596);
nand U3812 (N_3812,N_2979,N_2087);
nor U3813 (N_3813,N_2769,N_2004);
and U3814 (N_3814,N_2614,N_2812);
and U3815 (N_3815,N_2854,N_2992);
or U3816 (N_3816,N_2899,N_2214);
nand U3817 (N_3817,N_2071,N_2470);
nor U3818 (N_3818,N_2469,N_2462);
xor U3819 (N_3819,N_2808,N_2968);
nand U3820 (N_3820,N_2335,N_2286);
nand U3821 (N_3821,N_2701,N_2192);
nor U3822 (N_3822,N_2099,N_2234);
and U3823 (N_3823,N_2764,N_2223);
nor U3824 (N_3824,N_2407,N_2808);
or U3825 (N_3825,N_2693,N_2333);
nor U3826 (N_3826,N_2564,N_2715);
nand U3827 (N_3827,N_2809,N_2567);
nor U3828 (N_3828,N_2767,N_2671);
or U3829 (N_3829,N_2387,N_2984);
or U3830 (N_3830,N_2795,N_2908);
nand U3831 (N_3831,N_2502,N_2084);
or U3832 (N_3832,N_2303,N_2622);
nor U3833 (N_3833,N_2088,N_2072);
and U3834 (N_3834,N_2543,N_2440);
nor U3835 (N_3835,N_2843,N_2601);
or U3836 (N_3836,N_2477,N_2152);
nor U3837 (N_3837,N_2257,N_2304);
xnor U3838 (N_3838,N_2391,N_2574);
or U3839 (N_3839,N_2130,N_2709);
or U3840 (N_3840,N_2392,N_2509);
xor U3841 (N_3841,N_2784,N_2815);
and U3842 (N_3842,N_2306,N_2144);
nand U3843 (N_3843,N_2113,N_2765);
nand U3844 (N_3844,N_2195,N_2600);
nand U3845 (N_3845,N_2928,N_2748);
or U3846 (N_3846,N_2454,N_2932);
or U3847 (N_3847,N_2553,N_2613);
nand U3848 (N_3848,N_2803,N_2456);
nand U3849 (N_3849,N_2166,N_2154);
xnor U3850 (N_3850,N_2741,N_2431);
and U3851 (N_3851,N_2296,N_2395);
or U3852 (N_3852,N_2724,N_2734);
xor U3853 (N_3853,N_2478,N_2084);
nor U3854 (N_3854,N_2981,N_2955);
xor U3855 (N_3855,N_2107,N_2326);
nor U3856 (N_3856,N_2731,N_2940);
or U3857 (N_3857,N_2156,N_2158);
and U3858 (N_3858,N_2620,N_2946);
nand U3859 (N_3859,N_2857,N_2502);
xnor U3860 (N_3860,N_2370,N_2693);
and U3861 (N_3861,N_2756,N_2265);
or U3862 (N_3862,N_2022,N_2218);
nand U3863 (N_3863,N_2749,N_2448);
or U3864 (N_3864,N_2456,N_2213);
and U3865 (N_3865,N_2577,N_2371);
nor U3866 (N_3866,N_2335,N_2691);
and U3867 (N_3867,N_2116,N_2993);
or U3868 (N_3868,N_2950,N_2956);
nand U3869 (N_3869,N_2081,N_2367);
and U3870 (N_3870,N_2652,N_2645);
xor U3871 (N_3871,N_2324,N_2765);
xnor U3872 (N_3872,N_2721,N_2262);
xor U3873 (N_3873,N_2251,N_2927);
or U3874 (N_3874,N_2036,N_2524);
or U3875 (N_3875,N_2501,N_2413);
or U3876 (N_3876,N_2020,N_2148);
or U3877 (N_3877,N_2653,N_2465);
nand U3878 (N_3878,N_2300,N_2517);
and U3879 (N_3879,N_2666,N_2255);
xnor U3880 (N_3880,N_2638,N_2024);
nor U3881 (N_3881,N_2851,N_2263);
or U3882 (N_3882,N_2529,N_2297);
and U3883 (N_3883,N_2371,N_2287);
and U3884 (N_3884,N_2977,N_2806);
and U3885 (N_3885,N_2049,N_2123);
xnor U3886 (N_3886,N_2463,N_2612);
nor U3887 (N_3887,N_2825,N_2980);
and U3888 (N_3888,N_2958,N_2292);
and U3889 (N_3889,N_2296,N_2408);
nor U3890 (N_3890,N_2365,N_2746);
nand U3891 (N_3891,N_2936,N_2091);
or U3892 (N_3892,N_2642,N_2431);
nand U3893 (N_3893,N_2417,N_2213);
or U3894 (N_3894,N_2331,N_2718);
or U3895 (N_3895,N_2567,N_2972);
nand U3896 (N_3896,N_2050,N_2107);
xor U3897 (N_3897,N_2613,N_2565);
and U3898 (N_3898,N_2248,N_2280);
or U3899 (N_3899,N_2834,N_2978);
nor U3900 (N_3900,N_2648,N_2910);
xor U3901 (N_3901,N_2733,N_2533);
and U3902 (N_3902,N_2645,N_2046);
xnor U3903 (N_3903,N_2822,N_2009);
and U3904 (N_3904,N_2535,N_2548);
nor U3905 (N_3905,N_2286,N_2704);
nand U3906 (N_3906,N_2866,N_2346);
and U3907 (N_3907,N_2444,N_2177);
nor U3908 (N_3908,N_2321,N_2247);
nor U3909 (N_3909,N_2569,N_2949);
nand U3910 (N_3910,N_2225,N_2626);
or U3911 (N_3911,N_2091,N_2925);
and U3912 (N_3912,N_2759,N_2895);
nand U3913 (N_3913,N_2916,N_2943);
xnor U3914 (N_3914,N_2859,N_2218);
nor U3915 (N_3915,N_2778,N_2686);
xnor U3916 (N_3916,N_2128,N_2391);
xor U3917 (N_3917,N_2940,N_2797);
and U3918 (N_3918,N_2571,N_2962);
nor U3919 (N_3919,N_2477,N_2679);
nand U3920 (N_3920,N_2981,N_2596);
and U3921 (N_3921,N_2485,N_2476);
nand U3922 (N_3922,N_2301,N_2874);
xnor U3923 (N_3923,N_2112,N_2299);
nor U3924 (N_3924,N_2627,N_2855);
xor U3925 (N_3925,N_2126,N_2067);
or U3926 (N_3926,N_2107,N_2252);
or U3927 (N_3927,N_2337,N_2884);
or U3928 (N_3928,N_2620,N_2343);
and U3929 (N_3929,N_2642,N_2190);
and U3930 (N_3930,N_2484,N_2620);
nand U3931 (N_3931,N_2399,N_2829);
xor U3932 (N_3932,N_2201,N_2979);
and U3933 (N_3933,N_2773,N_2526);
nand U3934 (N_3934,N_2391,N_2554);
xor U3935 (N_3935,N_2624,N_2265);
nand U3936 (N_3936,N_2557,N_2472);
nand U3937 (N_3937,N_2356,N_2457);
or U3938 (N_3938,N_2207,N_2079);
or U3939 (N_3939,N_2666,N_2923);
nor U3940 (N_3940,N_2957,N_2075);
nand U3941 (N_3941,N_2858,N_2734);
nand U3942 (N_3942,N_2935,N_2360);
and U3943 (N_3943,N_2378,N_2358);
or U3944 (N_3944,N_2380,N_2556);
or U3945 (N_3945,N_2201,N_2474);
xor U3946 (N_3946,N_2328,N_2567);
nor U3947 (N_3947,N_2732,N_2328);
or U3948 (N_3948,N_2072,N_2931);
and U3949 (N_3949,N_2112,N_2138);
nand U3950 (N_3950,N_2335,N_2480);
nor U3951 (N_3951,N_2647,N_2729);
nor U3952 (N_3952,N_2783,N_2948);
nor U3953 (N_3953,N_2190,N_2107);
xnor U3954 (N_3954,N_2772,N_2865);
xnor U3955 (N_3955,N_2597,N_2804);
and U3956 (N_3956,N_2688,N_2159);
xor U3957 (N_3957,N_2054,N_2370);
and U3958 (N_3958,N_2492,N_2074);
nor U3959 (N_3959,N_2107,N_2627);
and U3960 (N_3960,N_2921,N_2577);
and U3961 (N_3961,N_2861,N_2073);
or U3962 (N_3962,N_2415,N_2008);
xor U3963 (N_3963,N_2317,N_2988);
and U3964 (N_3964,N_2023,N_2066);
xor U3965 (N_3965,N_2459,N_2300);
nor U3966 (N_3966,N_2905,N_2581);
nor U3967 (N_3967,N_2749,N_2698);
xnor U3968 (N_3968,N_2304,N_2922);
nor U3969 (N_3969,N_2244,N_2768);
and U3970 (N_3970,N_2506,N_2588);
or U3971 (N_3971,N_2420,N_2460);
or U3972 (N_3972,N_2100,N_2638);
or U3973 (N_3973,N_2004,N_2754);
nor U3974 (N_3974,N_2931,N_2670);
and U3975 (N_3975,N_2667,N_2042);
nor U3976 (N_3976,N_2233,N_2565);
and U3977 (N_3977,N_2387,N_2202);
or U3978 (N_3978,N_2074,N_2963);
xor U3979 (N_3979,N_2153,N_2661);
nor U3980 (N_3980,N_2259,N_2607);
and U3981 (N_3981,N_2554,N_2475);
nand U3982 (N_3982,N_2803,N_2580);
nor U3983 (N_3983,N_2689,N_2338);
nand U3984 (N_3984,N_2339,N_2456);
or U3985 (N_3985,N_2529,N_2325);
nor U3986 (N_3986,N_2871,N_2003);
nand U3987 (N_3987,N_2878,N_2614);
nand U3988 (N_3988,N_2382,N_2452);
nor U3989 (N_3989,N_2962,N_2892);
or U3990 (N_3990,N_2655,N_2649);
or U3991 (N_3991,N_2012,N_2321);
nor U3992 (N_3992,N_2202,N_2596);
nand U3993 (N_3993,N_2911,N_2255);
xor U3994 (N_3994,N_2448,N_2261);
or U3995 (N_3995,N_2964,N_2596);
or U3996 (N_3996,N_2725,N_2715);
and U3997 (N_3997,N_2670,N_2159);
xor U3998 (N_3998,N_2303,N_2563);
or U3999 (N_3999,N_2941,N_2623);
xnor U4000 (N_4000,N_3582,N_3046);
and U4001 (N_4001,N_3435,N_3760);
nor U4002 (N_4002,N_3425,N_3681);
or U4003 (N_4003,N_3024,N_3195);
or U4004 (N_4004,N_3336,N_3232);
nand U4005 (N_4005,N_3276,N_3999);
nand U4006 (N_4006,N_3236,N_3190);
xor U4007 (N_4007,N_3152,N_3936);
nor U4008 (N_4008,N_3077,N_3537);
nor U4009 (N_4009,N_3734,N_3436);
nor U4010 (N_4010,N_3587,N_3421);
xor U4011 (N_4011,N_3818,N_3163);
or U4012 (N_4012,N_3676,N_3127);
or U4013 (N_4013,N_3669,N_3738);
nor U4014 (N_4014,N_3072,N_3899);
nor U4015 (N_4015,N_3775,N_3983);
xnor U4016 (N_4016,N_3339,N_3020);
xor U4017 (N_4017,N_3594,N_3591);
nand U4018 (N_4018,N_3275,N_3571);
or U4019 (N_4019,N_3929,N_3352);
nor U4020 (N_4020,N_3419,N_3874);
or U4021 (N_4021,N_3909,N_3688);
or U4022 (N_4022,N_3016,N_3401);
or U4023 (N_4023,N_3757,N_3031);
nand U4024 (N_4024,N_3431,N_3958);
nand U4025 (N_4025,N_3430,N_3846);
nand U4026 (N_4026,N_3870,N_3881);
and U4027 (N_4027,N_3648,N_3674);
and U4028 (N_4028,N_3144,N_3923);
nor U4029 (N_4029,N_3329,N_3735);
and U4030 (N_4030,N_3740,N_3182);
or U4031 (N_4031,N_3231,N_3854);
xor U4032 (N_4032,N_3531,N_3724);
nor U4033 (N_4033,N_3378,N_3322);
nor U4034 (N_4034,N_3529,N_3940);
and U4035 (N_4035,N_3885,N_3301);
nand U4036 (N_4036,N_3203,N_3579);
and U4037 (N_4037,N_3592,N_3604);
nor U4038 (N_4038,N_3570,N_3984);
nand U4039 (N_4039,N_3908,N_3911);
nand U4040 (N_4040,N_3053,N_3943);
xor U4041 (N_4041,N_3883,N_3354);
xnor U4042 (N_4042,N_3776,N_3270);
nand U4043 (N_4043,N_3575,N_3122);
and U4044 (N_4044,N_3222,N_3959);
and U4045 (N_4045,N_3644,N_3337);
nand U4046 (N_4046,N_3777,N_3189);
xor U4047 (N_4047,N_3711,N_3120);
xor U4048 (N_4048,N_3054,N_3710);
nor U4049 (N_4049,N_3827,N_3995);
nand U4050 (N_4050,N_3603,N_3312);
nor U4051 (N_4051,N_3458,N_3910);
nor U4052 (N_4052,N_3461,N_3768);
or U4053 (N_4053,N_3173,N_3493);
nand U4054 (N_4054,N_3765,N_3297);
nand U4055 (N_4055,N_3863,N_3149);
and U4056 (N_4056,N_3832,N_3879);
or U4057 (N_4057,N_3498,N_3573);
xnor U4058 (N_4058,N_3991,N_3460);
nand U4059 (N_4059,N_3761,N_3652);
nor U4060 (N_4060,N_3975,N_3230);
or U4061 (N_4061,N_3141,N_3852);
nand U4062 (N_4062,N_3932,N_3853);
xnor U4063 (N_4063,N_3902,N_3209);
xnor U4064 (N_4064,N_3606,N_3447);
or U4065 (N_4065,N_3081,N_3484);
nor U4066 (N_4066,N_3332,N_3828);
nor U4067 (N_4067,N_3721,N_3264);
nand U4068 (N_4068,N_3891,N_3553);
and U4069 (N_4069,N_3955,N_3471);
or U4070 (N_4070,N_3013,N_3025);
nand U4071 (N_4071,N_3680,N_3810);
nor U4072 (N_4072,N_3219,N_3503);
nor U4073 (N_4073,N_3820,N_3739);
or U4074 (N_4074,N_3366,N_3698);
and U4075 (N_4075,N_3617,N_3894);
and U4076 (N_4076,N_3560,N_3028);
or U4077 (N_4077,N_3248,N_3713);
and U4078 (N_4078,N_3517,N_3340);
or U4079 (N_4079,N_3521,N_3727);
or U4080 (N_4080,N_3186,N_3912);
and U4081 (N_4081,N_3489,N_3041);
xnor U4082 (N_4082,N_3622,N_3183);
nand U4083 (N_4083,N_3801,N_3884);
nor U4084 (N_4084,N_3282,N_3858);
nand U4085 (N_4085,N_3783,N_3930);
or U4086 (N_4086,N_3043,N_3288);
or U4087 (N_4087,N_3831,N_3866);
nor U4088 (N_4088,N_3840,N_3067);
xnor U4089 (N_4089,N_3369,N_3368);
and U4090 (N_4090,N_3245,N_3095);
and U4091 (N_4091,N_3581,N_3974);
xnor U4092 (N_4092,N_3420,N_3205);
nor U4093 (N_4093,N_3821,N_3611);
nor U4094 (N_4094,N_3153,N_3374);
nand U4095 (N_4095,N_3084,N_3961);
nor U4096 (N_4096,N_3422,N_3121);
nand U4097 (N_4097,N_3289,N_3497);
xor U4098 (N_4098,N_3736,N_3226);
or U4099 (N_4099,N_3147,N_3860);
and U4100 (N_4100,N_3628,N_3010);
nand U4101 (N_4101,N_3917,N_3563);
nand U4102 (N_4102,N_3947,N_3459);
nor U4103 (N_4103,N_3962,N_3888);
nand U4104 (N_4104,N_3396,N_3822);
xnor U4105 (N_4105,N_3968,N_3868);
nand U4106 (N_4106,N_3785,N_3310);
nand U4107 (N_4107,N_3706,N_3625);
nand U4108 (N_4108,N_3406,N_3414);
nor U4109 (N_4109,N_3600,N_3439);
nand U4110 (N_4110,N_3371,N_3048);
nand U4111 (N_4111,N_3491,N_3819);
and U4112 (N_4112,N_3725,N_3349);
and U4113 (N_4113,N_3238,N_3382);
or U4114 (N_4114,N_3400,N_3130);
nor U4115 (N_4115,N_3100,N_3705);
xnor U4116 (N_4116,N_3945,N_3500);
nor U4117 (N_4117,N_3265,N_3326);
or U4118 (N_4118,N_3511,N_3823);
xor U4119 (N_4119,N_3426,N_3791);
xnor U4120 (N_4120,N_3809,N_3377);
nor U4121 (N_4121,N_3919,N_3311);
nor U4122 (N_4122,N_3477,N_3770);
xor U4123 (N_4123,N_3399,N_3309);
and U4124 (N_4124,N_3097,N_3159);
or U4125 (N_4125,N_3754,N_3034);
nor U4126 (N_4126,N_3814,N_3508);
xnor U4127 (N_4127,N_3651,N_3085);
nand U4128 (N_4128,N_3428,N_3277);
and U4129 (N_4129,N_3824,N_3254);
xnor U4130 (N_4130,N_3221,N_3807);
xnor U4131 (N_4131,N_3645,N_3880);
nor U4132 (N_4132,N_3825,N_3177);
xor U4133 (N_4133,N_3082,N_3012);
and U4134 (N_4134,N_3403,N_3331);
nor U4135 (N_4135,N_3981,N_3093);
nand U4136 (N_4136,N_3574,N_3679);
nor U4137 (N_4137,N_3344,N_3014);
or U4138 (N_4138,N_3335,N_3675);
nand U4139 (N_4139,N_3812,N_3145);
and U4140 (N_4140,N_3078,N_3715);
or U4141 (N_4141,N_3154,N_3741);
nor U4142 (N_4142,N_3750,N_3000);
xnor U4143 (N_4143,N_3786,N_3049);
or U4144 (N_4144,N_3596,N_3948);
or U4145 (N_4145,N_3532,N_3134);
and U4146 (N_4146,N_3992,N_3616);
xnor U4147 (N_4147,N_3970,N_3779);
nor U4148 (N_4148,N_3623,N_3108);
xor U4149 (N_4149,N_3480,N_3971);
and U4150 (N_4150,N_3583,N_3318);
xor U4151 (N_4151,N_3355,N_3576);
and U4152 (N_4152,N_3045,N_3522);
nand U4153 (N_4153,N_3937,N_3106);
nand U4154 (N_4154,N_3957,N_3844);
nor U4155 (N_4155,N_3607,N_3685);
and U4156 (N_4156,N_3061,N_3193);
nor U4157 (N_4157,N_3638,N_3615);
nor U4158 (N_4158,N_3762,N_3367);
nor U4159 (N_4159,N_3001,N_3898);
and U4160 (N_4160,N_3321,N_3671);
xor U4161 (N_4161,N_3307,N_3811);
nor U4162 (N_4162,N_3683,N_3117);
and U4163 (N_4163,N_3184,N_3548);
nor U4164 (N_4164,N_3720,N_3125);
and U4165 (N_4165,N_3758,N_3677);
or U4166 (N_4166,N_3882,N_3621);
xor U4167 (N_4167,N_3197,N_3561);
nor U4168 (N_4168,N_3637,N_3543);
or U4169 (N_4169,N_3467,N_3386);
or U4170 (N_4170,N_3798,N_3951);
xor U4171 (N_4171,N_3287,N_3328);
or U4172 (N_4172,N_3730,N_3257);
nand U4173 (N_4173,N_3759,N_3080);
or U4174 (N_4174,N_3556,N_3363);
or U4175 (N_4175,N_3742,N_3303);
and U4176 (N_4176,N_3523,N_3901);
nor U4177 (N_4177,N_3552,N_3415);
or U4178 (N_4178,N_3057,N_3502);
nand U4179 (N_4179,N_3389,N_3123);
or U4180 (N_4180,N_3417,N_3073);
or U4181 (N_4181,N_3160,N_3058);
nor U4182 (N_4182,N_3897,N_3906);
nand U4183 (N_4183,N_3052,N_3712);
xor U4184 (N_4184,N_3071,N_3180);
xor U4185 (N_4185,N_3784,N_3550);
or U4186 (N_4186,N_3692,N_3214);
and U4187 (N_4187,N_3364,N_3486);
and U4188 (N_4188,N_3920,N_3124);
nand U4189 (N_4189,N_3345,N_3167);
xnor U4190 (N_4190,N_3250,N_3731);
and U4191 (N_4191,N_3895,N_3797);
or U4192 (N_4192,N_3472,N_3176);
nor U4193 (N_4193,N_3083,N_3572);
and U4194 (N_4194,N_3997,N_3207);
xor U4195 (N_4195,N_3050,N_3719);
and U4196 (N_4196,N_3857,N_3033);
nand U4197 (N_4197,N_3746,N_3808);
xor U4198 (N_4198,N_3562,N_3941);
nor U4199 (N_4199,N_3360,N_3261);
nor U4200 (N_4200,N_3869,N_3004);
or U4201 (N_4201,N_3102,N_3060);
nor U4202 (N_4202,N_3613,N_3589);
or U4203 (N_4203,N_3732,N_3800);
nand U4204 (N_4204,N_3640,N_3068);
nand U4205 (N_4205,N_3567,N_3315);
and U4206 (N_4206,N_3633,N_3475);
or U4207 (N_4207,N_3978,N_3817);
nand U4208 (N_4208,N_3223,N_3593);
xnor U4209 (N_4209,N_3111,N_3952);
nor U4210 (N_4210,N_3836,N_3528);
nor U4211 (N_4211,N_3384,N_3729);
or U4212 (N_4212,N_3136,N_3370);
and U4213 (N_4213,N_3518,N_3285);
or U4214 (N_4214,N_3294,N_3849);
nor U4215 (N_4215,N_3114,N_3158);
xor U4216 (N_4216,N_3717,N_3474);
or U4217 (N_4217,N_3466,N_3404);
and U4218 (N_4218,N_3156,N_3509);
nor U4219 (N_4219,N_3672,N_3977);
xor U4220 (N_4220,N_3172,N_3927);
and U4221 (N_4221,N_3663,N_3632);
or U4222 (N_4222,N_3643,N_3142);
xnor U4223 (N_4223,N_3774,N_3896);
nand U4224 (N_4224,N_3540,N_3707);
nor U4225 (N_4225,N_3185,N_3148);
xor U4226 (N_4226,N_3505,N_3204);
or U4227 (N_4227,N_3216,N_3942);
nor U4228 (N_4228,N_3485,N_3157);
or U4229 (N_4229,N_3639,N_3047);
and U4230 (N_4230,N_3541,N_3026);
or U4231 (N_4231,N_3703,N_3280);
nor U4232 (N_4232,N_3262,N_3056);
xor U4233 (N_4233,N_3383,N_3090);
nor U4234 (N_4234,N_3949,N_3390);
nor U4235 (N_4235,N_3642,N_3059);
and U4236 (N_4236,N_3751,N_3065);
xor U4237 (N_4237,N_3418,N_3094);
xor U4238 (N_4238,N_3969,N_3660);
nor U4239 (N_4239,N_3341,N_3040);
or U4240 (N_4240,N_3027,N_3449);
nor U4241 (N_4241,N_3987,N_3343);
or U4242 (N_4242,N_3653,N_3805);
nand U4243 (N_4243,N_3440,N_3524);
xnor U4244 (N_4244,N_3538,N_3877);
and U4245 (N_4245,N_3551,N_3003);
and U4246 (N_4246,N_3925,N_3922);
nand U4247 (N_4247,N_3842,N_3709);
or U4248 (N_4248,N_3744,N_3423);
nor U4249 (N_4249,N_3782,N_3237);
xor U4250 (N_4250,N_3308,N_3778);
nor U4251 (N_4251,N_3011,N_3533);
xnor U4252 (N_4252,N_3424,N_3602);
nand U4253 (N_4253,N_3075,N_3916);
nor U4254 (N_4254,N_3037,N_3373);
and U4255 (N_4255,N_3728,N_3586);
or U4256 (N_4256,N_3385,N_3848);
xnor U4257 (N_4257,N_3387,N_3333);
and U4258 (N_4258,N_3405,N_3023);
xor U4259 (N_4259,N_3062,N_3259);
nor U4260 (N_4260,N_3224,N_3697);
nand U4261 (N_4261,N_3351,N_3631);
and U4262 (N_4262,N_3789,N_3926);
and U4263 (N_4263,N_3434,N_3446);
xor U4264 (N_4264,N_3166,N_3008);
nand U4265 (N_4265,N_3150,N_3693);
nand U4266 (N_4266,N_3039,N_3269);
or U4267 (N_4267,N_3397,N_3074);
xor U4268 (N_4268,N_3317,N_3687);
nor U4269 (N_4269,N_3989,N_3861);
nor U4270 (N_4270,N_3099,N_3064);
or U4271 (N_4271,N_3833,N_3169);
nor U4272 (N_4272,N_3665,N_3856);
nand U4273 (N_4273,N_3376,N_3772);
xor U4274 (N_4274,N_3859,N_3200);
and U4275 (N_4275,N_3365,N_3361);
nand U4276 (N_4276,N_3678,N_3829);
or U4277 (N_4277,N_3356,N_3752);
or U4278 (N_4278,N_3131,N_3664);
nor U4279 (N_4279,N_3402,N_3855);
and U4280 (N_4280,N_3455,N_3196);
or U4281 (N_4281,N_3412,N_3139);
and U4282 (N_4282,N_3996,N_3716);
and U4283 (N_4283,N_3982,N_3578);
nor U4284 (N_4284,N_3488,N_3771);
nand U4285 (N_4285,N_3965,N_3334);
or U4286 (N_4286,N_3889,N_3601);
xnor U4287 (N_4287,N_3702,N_3267);
xor U4288 (N_4288,N_3875,N_3939);
and U4289 (N_4289,N_3492,N_3626);
nor U4290 (N_4290,N_3577,N_3994);
and U4291 (N_4291,N_3864,N_3164);
and U4292 (N_4292,N_3242,N_3691);
nor U4293 (N_4293,N_3393,N_3605);
or U4294 (N_4294,N_3960,N_3862);
nand U4295 (N_4295,N_3069,N_3300);
nor U4296 (N_4296,N_3661,N_3140);
and U4297 (N_4297,N_3217,N_3465);
xnor U4298 (N_4298,N_3813,N_3499);
xor U4299 (N_4299,N_3281,N_3346);
or U4300 (N_4300,N_3950,N_3161);
nor U4301 (N_4301,N_3769,N_3588);
xnor U4302 (N_4302,N_3441,N_3319);
nor U4303 (N_4303,N_3035,N_3890);
xor U4304 (N_4304,N_3137,N_3608);
nor U4305 (N_4305,N_3564,N_3273);
or U4306 (N_4306,N_3468,N_3380);
or U4307 (N_4307,N_3115,N_3438);
and U4308 (N_4308,N_3295,N_3019);
and U4309 (N_4309,N_3168,N_3079);
or U4310 (N_4310,N_3756,N_3938);
xnor U4311 (N_4311,N_3251,N_3293);
xor U4312 (N_4312,N_3566,N_3747);
and U4313 (N_4313,N_3055,N_3260);
or U4314 (N_4314,N_3298,N_3228);
nor U4315 (N_4315,N_3963,N_3478);
or U4316 (N_4316,N_3568,N_3748);
xnor U4317 (N_4317,N_3513,N_3764);
or U4318 (N_4318,N_3103,N_3456);
and U4319 (N_4319,N_3704,N_3634);
and U4320 (N_4320,N_3347,N_3091);
xnor U4321 (N_4321,N_3520,N_3263);
nor U4322 (N_4322,N_3802,N_3635);
xor U4323 (N_4323,N_3796,N_3448);
or U4324 (N_4324,N_3473,N_3051);
xor U4325 (N_4325,N_3481,N_3444);
or U4326 (N_4326,N_3042,N_3871);
xor U4327 (N_4327,N_3138,N_3525);
and U4328 (N_4328,N_3395,N_3743);
xor U4329 (N_4329,N_3956,N_3029);
nor U4330 (N_4330,N_3504,N_3501);
and U4331 (N_4331,N_3793,N_3787);
or U4332 (N_4332,N_3815,N_3620);
nand U4333 (N_4333,N_3876,N_3530);
nand U4334 (N_4334,N_3650,N_3202);
xor U4335 (N_4335,N_3972,N_3442);
xor U4336 (N_4336,N_3737,N_3443);
or U4337 (N_4337,N_3655,N_3411);
and U4338 (N_4338,N_3580,N_3695);
nor U4339 (N_4339,N_3063,N_3432);
nor U4340 (N_4340,N_3584,N_3116);
nand U4341 (N_4341,N_3476,N_3155);
xor U4342 (N_4342,N_3795,N_3549);
xor U4343 (N_4343,N_3220,N_3954);
nand U4344 (N_4344,N_3656,N_3837);
xnor U4345 (N_4345,N_3194,N_3233);
nor U4346 (N_4346,N_3253,N_3032);
nand U4347 (N_4347,N_3353,N_3865);
nand U4348 (N_4348,N_3171,N_3535);
nand U4349 (N_4349,N_3165,N_3781);
or U4350 (N_4350,N_3658,N_3391);
or U4351 (N_4351,N_3749,N_3437);
nand U4352 (N_4352,N_3595,N_3452);
xor U4353 (N_4353,N_3714,N_3699);
nor U4354 (N_4354,N_3255,N_3279);
xor U4355 (N_4355,N_3700,N_3792);
or U4356 (N_4356,N_3128,N_3118);
nor U4357 (N_4357,N_3913,N_3274);
or U4358 (N_4358,N_3445,N_3305);
xnor U4359 (N_4359,N_3234,N_3694);
xor U4360 (N_4360,N_3998,N_3009);
or U4361 (N_4361,N_3227,N_3174);
nor U4362 (N_4362,N_3208,N_3427);
or U4363 (N_4363,N_3873,N_3753);
and U4364 (N_4364,N_3886,N_3666);
and U4365 (N_4365,N_3838,N_3433);
xnor U4366 (N_4366,N_3038,N_3022);
or U4367 (N_4367,N_3545,N_3271);
or U4368 (N_4368,N_3278,N_3483);
nand U4369 (N_4369,N_3358,N_3187);
nor U4370 (N_4370,N_3244,N_3066);
nor U4371 (N_4371,N_3268,N_3243);
or U4372 (N_4372,N_3018,N_3191);
xnor U4373 (N_4373,N_3469,N_3181);
or U4374 (N_4374,N_3510,N_3088);
nand U4375 (N_4375,N_3211,N_3647);
xor U4376 (N_4376,N_3519,N_3841);
or U4377 (N_4377,N_3636,N_3905);
nand U4378 (N_4378,N_3283,N_3726);
xnor U4379 (N_4379,N_3985,N_3429);
xor U4380 (N_4380,N_3342,N_3496);
and U4381 (N_4381,N_3109,N_3559);
and U4382 (N_4382,N_3931,N_3175);
or U4383 (N_4383,N_3953,N_3935);
nor U4384 (N_4384,N_3372,N_3348);
nand U4385 (N_4385,N_3464,N_3557);
or U4386 (N_4386,N_3002,N_3803);
nor U4387 (N_4387,N_3918,N_3092);
or U4388 (N_4388,N_3199,N_3847);
and U4389 (N_4389,N_3506,N_3629);
nor U4390 (N_4390,N_3104,N_3313);
xor U4391 (N_4391,N_3722,N_3790);
nor U4392 (N_4392,N_3534,N_3087);
nor U4393 (N_4393,N_3398,N_3338);
xor U4394 (N_4394,N_3536,N_3558);
or U4395 (N_4395,N_3667,N_3933);
nor U4396 (N_4396,N_3357,N_3070);
and U4397 (N_4397,N_3215,N_3686);
nand U4398 (N_4398,N_3453,N_3036);
and U4399 (N_4399,N_3907,N_3394);
nor U4400 (N_4400,N_3113,N_3988);
nand U4401 (N_4401,N_3657,N_3089);
or U4402 (N_4402,N_3210,N_3839);
xor U4403 (N_4403,N_3696,N_3733);
or U4404 (N_4404,N_3755,N_3388);
nand U4405 (N_4405,N_3973,N_3105);
and U4406 (N_4406,N_3893,N_3512);
and U4407 (N_4407,N_3590,N_3286);
nor U4408 (N_4408,N_3314,N_3044);
xor U4409 (N_4409,N_3816,N_3964);
xor U4410 (N_4410,N_3599,N_3021);
and U4411 (N_4411,N_3462,N_3585);
xor U4412 (N_4412,N_3381,N_3723);
and U4413 (N_4413,N_3684,N_3835);
and U4414 (N_4414,N_3129,N_3284);
nand U4415 (N_4415,N_3098,N_3872);
xor U4416 (N_4416,N_3296,N_3544);
xnor U4417 (N_4417,N_3976,N_3126);
xnor U4418 (N_4418,N_3851,N_3007);
or U4419 (N_4419,N_3843,N_3773);
nor U4420 (N_4420,N_3213,N_3241);
xnor U4421 (N_4421,N_3229,N_3662);
or U4422 (N_4422,N_3290,N_3457);
nand U4423 (N_4423,N_3554,N_3966);
and U4424 (N_4424,N_3619,N_3246);
nand U4425 (N_4425,N_3304,N_3641);
and U4426 (N_4426,N_3017,N_3515);
and U4427 (N_4427,N_3479,N_3258);
xnor U4428 (N_4428,N_3323,N_3618);
nor U4429 (N_4429,N_3132,N_3627);
nor U4430 (N_4430,N_3006,N_3324);
xor U4431 (N_4431,N_3076,N_3133);
nor U4432 (N_4432,N_3030,N_3979);
and U4433 (N_4433,N_3107,N_3110);
xnor U4434 (N_4434,N_3612,N_3799);
xor U4435 (N_4435,N_3162,N_3101);
xnor U4436 (N_4436,N_3555,N_3850);
nor U4437 (N_4437,N_3198,N_3610);
xnor U4438 (N_4438,N_3410,N_3362);
and U4439 (N_4439,N_3921,N_3654);
nor U4440 (N_4440,N_3516,N_3845);
or U4441 (N_4441,N_3569,N_3507);
and U4442 (N_4442,N_3718,N_3609);
and U4443 (N_4443,N_3766,N_3806);
nor U4444 (N_4444,N_3614,N_3291);
nor U4445 (N_4445,N_3915,N_3413);
or U4446 (N_4446,N_3299,N_3788);
and U4447 (N_4447,N_3892,N_3867);
and U4448 (N_4448,N_3225,N_3526);
or U4449 (N_4449,N_3900,N_3143);
and U4450 (N_4450,N_3247,N_3780);
xnor U4451 (N_4451,N_3212,N_3767);
and U4452 (N_4452,N_3826,N_3670);
or U4453 (N_4453,N_3928,N_3256);
nand U4454 (N_4454,N_3359,N_3763);
nor U4455 (N_4455,N_3542,N_3539);
nand U4456 (N_4456,N_3272,N_3490);
or U4457 (N_4457,N_3914,N_3986);
xor U4458 (N_4458,N_3192,N_3630);
nor U4459 (N_4459,N_3218,N_3330);
nand U4460 (N_4460,N_3993,N_3463);
and U4461 (N_4461,N_3112,N_3392);
and U4462 (N_4462,N_3320,N_3546);
and U4463 (N_4463,N_3235,N_3266);
nand U4464 (N_4464,N_3527,N_3495);
xnor U4465 (N_4465,N_3179,N_3239);
xor U4466 (N_4466,N_3316,N_3514);
or U4467 (N_4467,N_3494,N_3325);
and U4468 (N_4468,N_3450,N_3096);
and U4469 (N_4469,N_3834,N_3454);
or U4470 (N_4470,N_3170,N_3292);
and U4471 (N_4471,N_3804,N_3946);
nand U4472 (N_4472,N_3327,N_3701);
nor U4473 (N_4473,N_3668,N_3887);
or U4474 (N_4474,N_3178,N_3487);
or U4475 (N_4475,N_3005,N_3673);
or U4476 (N_4476,N_3646,N_3980);
xnor U4477 (N_4477,N_3649,N_3302);
nor U4478 (N_4478,N_3682,N_3416);
nand U4479 (N_4479,N_3119,N_3565);
and U4480 (N_4480,N_3689,N_3659);
and U4481 (N_4481,N_3188,N_3934);
or U4482 (N_4482,N_3015,N_3624);
nand U4483 (N_4483,N_3482,N_3708);
nor U4484 (N_4484,N_3201,N_3967);
nand U4485 (N_4485,N_3690,N_3904);
or U4486 (N_4486,N_3990,N_3306);
or U4487 (N_4487,N_3794,N_3924);
nor U4488 (N_4488,N_3350,N_3408);
xor U4489 (N_4489,N_3944,N_3903);
nand U4490 (N_4490,N_3409,N_3249);
nand U4491 (N_4491,N_3451,N_3086);
or U4492 (N_4492,N_3146,N_3470);
xnor U4493 (N_4493,N_3379,N_3151);
nand U4494 (N_4494,N_3407,N_3830);
and U4495 (N_4495,N_3240,N_3597);
or U4496 (N_4496,N_3252,N_3135);
and U4497 (N_4497,N_3206,N_3745);
nor U4498 (N_4498,N_3878,N_3375);
nor U4499 (N_4499,N_3598,N_3547);
xor U4500 (N_4500,N_3060,N_3409);
and U4501 (N_4501,N_3510,N_3697);
nor U4502 (N_4502,N_3041,N_3753);
xnor U4503 (N_4503,N_3181,N_3957);
nor U4504 (N_4504,N_3100,N_3446);
xor U4505 (N_4505,N_3721,N_3809);
or U4506 (N_4506,N_3582,N_3694);
and U4507 (N_4507,N_3642,N_3611);
xor U4508 (N_4508,N_3341,N_3048);
or U4509 (N_4509,N_3751,N_3778);
nor U4510 (N_4510,N_3324,N_3147);
and U4511 (N_4511,N_3123,N_3902);
and U4512 (N_4512,N_3358,N_3646);
or U4513 (N_4513,N_3382,N_3010);
nor U4514 (N_4514,N_3785,N_3833);
and U4515 (N_4515,N_3976,N_3758);
nor U4516 (N_4516,N_3638,N_3288);
xnor U4517 (N_4517,N_3601,N_3456);
nor U4518 (N_4518,N_3568,N_3109);
or U4519 (N_4519,N_3330,N_3103);
and U4520 (N_4520,N_3330,N_3464);
nand U4521 (N_4521,N_3780,N_3291);
or U4522 (N_4522,N_3813,N_3425);
or U4523 (N_4523,N_3066,N_3405);
nand U4524 (N_4524,N_3641,N_3353);
nor U4525 (N_4525,N_3594,N_3246);
or U4526 (N_4526,N_3407,N_3462);
nor U4527 (N_4527,N_3372,N_3045);
nand U4528 (N_4528,N_3812,N_3370);
and U4529 (N_4529,N_3362,N_3561);
and U4530 (N_4530,N_3401,N_3107);
nor U4531 (N_4531,N_3996,N_3136);
xor U4532 (N_4532,N_3059,N_3836);
xor U4533 (N_4533,N_3562,N_3989);
nand U4534 (N_4534,N_3684,N_3590);
or U4535 (N_4535,N_3260,N_3072);
nor U4536 (N_4536,N_3598,N_3710);
and U4537 (N_4537,N_3604,N_3586);
nor U4538 (N_4538,N_3589,N_3757);
and U4539 (N_4539,N_3863,N_3098);
nor U4540 (N_4540,N_3878,N_3021);
or U4541 (N_4541,N_3583,N_3441);
or U4542 (N_4542,N_3485,N_3569);
nor U4543 (N_4543,N_3677,N_3244);
nand U4544 (N_4544,N_3217,N_3588);
and U4545 (N_4545,N_3928,N_3843);
or U4546 (N_4546,N_3197,N_3387);
nor U4547 (N_4547,N_3507,N_3299);
nor U4548 (N_4548,N_3399,N_3910);
or U4549 (N_4549,N_3563,N_3078);
or U4550 (N_4550,N_3844,N_3972);
or U4551 (N_4551,N_3715,N_3704);
or U4552 (N_4552,N_3682,N_3507);
xor U4553 (N_4553,N_3200,N_3714);
nor U4554 (N_4554,N_3976,N_3616);
or U4555 (N_4555,N_3435,N_3638);
nand U4556 (N_4556,N_3546,N_3742);
and U4557 (N_4557,N_3704,N_3909);
and U4558 (N_4558,N_3049,N_3305);
nor U4559 (N_4559,N_3566,N_3281);
nor U4560 (N_4560,N_3659,N_3555);
nand U4561 (N_4561,N_3828,N_3570);
or U4562 (N_4562,N_3237,N_3719);
nand U4563 (N_4563,N_3855,N_3378);
and U4564 (N_4564,N_3008,N_3745);
xor U4565 (N_4565,N_3935,N_3817);
or U4566 (N_4566,N_3056,N_3753);
nor U4567 (N_4567,N_3144,N_3336);
xnor U4568 (N_4568,N_3186,N_3734);
nand U4569 (N_4569,N_3399,N_3136);
nor U4570 (N_4570,N_3878,N_3874);
xnor U4571 (N_4571,N_3689,N_3021);
or U4572 (N_4572,N_3500,N_3608);
and U4573 (N_4573,N_3809,N_3029);
nor U4574 (N_4574,N_3330,N_3474);
and U4575 (N_4575,N_3852,N_3772);
nor U4576 (N_4576,N_3576,N_3020);
or U4577 (N_4577,N_3217,N_3100);
or U4578 (N_4578,N_3692,N_3405);
nor U4579 (N_4579,N_3442,N_3269);
nand U4580 (N_4580,N_3214,N_3494);
nand U4581 (N_4581,N_3406,N_3737);
nor U4582 (N_4582,N_3663,N_3132);
or U4583 (N_4583,N_3610,N_3577);
nand U4584 (N_4584,N_3914,N_3454);
xor U4585 (N_4585,N_3721,N_3196);
nand U4586 (N_4586,N_3523,N_3281);
xnor U4587 (N_4587,N_3707,N_3890);
nand U4588 (N_4588,N_3265,N_3098);
xnor U4589 (N_4589,N_3992,N_3859);
nor U4590 (N_4590,N_3988,N_3678);
nor U4591 (N_4591,N_3501,N_3767);
xor U4592 (N_4592,N_3713,N_3104);
and U4593 (N_4593,N_3292,N_3802);
and U4594 (N_4594,N_3171,N_3282);
nand U4595 (N_4595,N_3896,N_3268);
nand U4596 (N_4596,N_3125,N_3440);
nor U4597 (N_4597,N_3405,N_3234);
nand U4598 (N_4598,N_3857,N_3259);
xor U4599 (N_4599,N_3891,N_3993);
and U4600 (N_4600,N_3054,N_3013);
or U4601 (N_4601,N_3826,N_3988);
and U4602 (N_4602,N_3707,N_3967);
xnor U4603 (N_4603,N_3942,N_3215);
nand U4604 (N_4604,N_3288,N_3145);
and U4605 (N_4605,N_3309,N_3392);
nand U4606 (N_4606,N_3883,N_3197);
xnor U4607 (N_4607,N_3106,N_3100);
nor U4608 (N_4608,N_3776,N_3597);
and U4609 (N_4609,N_3710,N_3923);
nor U4610 (N_4610,N_3325,N_3606);
or U4611 (N_4611,N_3986,N_3719);
and U4612 (N_4612,N_3605,N_3625);
nand U4613 (N_4613,N_3441,N_3485);
or U4614 (N_4614,N_3731,N_3057);
nand U4615 (N_4615,N_3473,N_3205);
and U4616 (N_4616,N_3435,N_3806);
and U4617 (N_4617,N_3130,N_3760);
and U4618 (N_4618,N_3882,N_3040);
xor U4619 (N_4619,N_3804,N_3949);
nor U4620 (N_4620,N_3546,N_3330);
and U4621 (N_4621,N_3122,N_3191);
xnor U4622 (N_4622,N_3851,N_3139);
nand U4623 (N_4623,N_3721,N_3377);
and U4624 (N_4624,N_3680,N_3513);
and U4625 (N_4625,N_3972,N_3717);
nor U4626 (N_4626,N_3720,N_3421);
xor U4627 (N_4627,N_3948,N_3523);
or U4628 (N_4628,N_3697,N_3373);
and U4629 (N_4629,N_3203,N_3041);
nor U4630 (N_4630,N_3891,N_3098);
and U4631 (N_4631,N_3882,N_3011);
nor U4632 (N_4632,N_3408,N_3969);
and U4633 (N_4633,N_3233,N_3396);
and U4634 (N_4634,N_3780,N_3347);
or U4635 (N_4635,N_3525,N_3308);
nand U4636 (N_4636,N_3853,N_3144);
nor U4637 (N_4637,N_3614,N_3896);
or U4638 (N_4638,N_3207,N_3490);
nor U4639 (N_4639,N_3955,N_3213);
nor U4640 (N_4640,N_3344,N_3836);
nand U4641 (N_4641,N_3844,N_3641);
nor U4642 (N_4642,N_3274,N_3057);
nand U4643 (N_4643,N_3378,N_3130);
xor U4644 (N_4644,N_3589,N_3668);
nand U4645 (N_4645,N_3827,N_3882);
and U4646 (N_4646,N_3982,N_3271);
nand U4647 (N_4647,N_3684,N_3838);
nor U4648 (N_4648,N_3779,N_3489);
nor U4649 (N_4649,N_3088,N_3932);
nor U4650 (N_4650,N_3862,N_3024);
or U4651 (N_4651,N_3270,N_3402);
and U4652 (N_4652,N_3815,N_3685);
xnor U4653 (N_4653,N_3547,N_3207);
xnor U4654 (N_4654,N_3301,N_3718);
nor U4655 (N_4655,N_3397,N_3091);
xnor U4656 (N_4656,N_3346,N_3822);
xnor U4657 (N_4657,N_3186,N_3195);
nand U4658 (N_4658,N_3018,N_3176);
nand U4659 (N_4659,N_3758,N_3643);
and U4660 (N_4660,N_3541,N_3640);
or U4661 (N_4661,N_3205,N_3015);
and U4662 (N_4662,N_3319,N_3731);
and U4663 (N_4663,N_3901,N_3069);
nand U4664 (N_4664,N_3834,N_3113);
nor U4665 (N_4665,N_3874,N_3764);
and U4666 (N_4666,N_3185,N_3991);
and U4667 (N_4667,N_3979,N_3898);
nand U4668 (N_4668,N_3315,N_3488);
and U4669 (N_4669,N_3945,N_3311);
and U4670 (N_4670,N_3872,N_3119);
or U4671 (N_4671,N_3026,N_3288);
nor U4672 (N_4672,N_3855,N_3845);
xor U4673 (N_4673,N_3657,N_3992);
nor U4674 (N_4674,N_3371,N_3090);
and U4675 (N_4675,N_3335,N_3984);
xor U4676 (N_4676,N_3314,N_3137);
and U4677 (N_4677,N_3605,N_3056);
xnor U4678 (N_4678,N_3814,N_3706);
nand U4679 (N_4679,N_3821,N_3783);
or U4680 (N_4680,N_3080,N_3430);
xnor U4681 (N_4681,N_3979,N_3457);
nand U4682 (N_4682,N_3032,N_3547);
nand U4683 (N_4683,N_3115,N_3162);
nand U4684 (N_4684,N_3636,N_3963);
or U4685 (N_4685,N_3845,N_3292);
xor U4686 (N_4686,N_3088,N_3596);
nor U4687 (N_4687,N_3857,N_3377);
and U4688 (N_4688,N_3073,N_3531);
nand U4689 (N_4689,N_3028,N_3134);
or U4690 (N_4690,N_3868,N_3476);
or U4691 (N_4691,N_3441,N_3110);
xor U4692 (N_4692,N_3942,N_3529);
xnor U4693 (N_4693,N_3325,N_3692);
nand U4694 (N_4694,N_3607,N_3047);
nor U4695 (N_4695,N_3890,N_3220);
nor U4696 (N_4696,N_3658,N_3384);
nor U4697 (N_4697,N_3442,N_3002);
xnor U4698 (N_4698,N_3188,N_3571);
nand U4699 (N_4699,N_3566,N_3358);
or U4700 (N_4700,N_3273,N_3847);
or U4701 (N_4701,N_3467,N_3435);
nand U4702 (N_4702,N_3995,N_3905);
or U4703 (N_4703,N_3900,N_3825);
xor U4704 (N_4704,N_3434,N_3579);
nand U4705 (N_4705,N_3101,N_3408);
or U4706 (N_4706,N_3426,N_3640);
nand U4707 (N_4707,N_3997,N_3388);
or U4708 (N_4708,N_3606,N_3691);
and U4709 (N_4709,N_3154,N_3966);
nor U4710 (N_4710,N_3614,N_3424);
and U4711 (N_4711,N_3280,N_3692);
and U4712 (N_4712,N_3637,N_3111);
or U4713 (N_4713,N_3897,N_3197);
and U4714 (N_4714,N_3977,N_3734);
or U4715 (N_4715,N_3553,N_3846);
or U4716 (N_4716,N_3285,N_3084);
xor U4717 (N_4717,N_3530,N_3513);
nor U4718 (N_4718,N_3394,N_3498);
nor U4719 (N_4719,N_3436,N_3466);
or U4720 (N_4720,N_3502,N_3660);
nand U4721 (N_4721,N_3651,N_3398);
nor U4722 (N_4722,N_3093,N_3503);
nand U4723 (N_4723,N_3772,N_3311);
xor U4724 (N_4724,N_3776,N_3285);
and U4725 (N_4725,N_3599,N_3400);
xnor U4726 (N_4726,N_3103,N_3499);
and U4727 (N_4727,N_3970,N_3380);
and U4728 (N_4728,N_3817,N_3856);
nand U4729 (N_4729,N_3308,N_3238);
or U4730 (N_4730,N_3143,N_3849);
or U4731 (N_4731,N_3312,N_3000);
and U4732 (N_4732,N_3158,N_3318);
nor U4733 (N_4733,N_3845,N_3389);
or U4734 (N_4734,N_3990,N_3878);
xor U4735 (N_4735,N_3818,N_3518);
xor U4736 (N_4736,N_3752,N_3129);
nand U4737 (N_4737,N_3475,N_3502);
xnor U4738 (N_4738,N_3416,N_3801);
nand U4739 (N_4739,N_3848,N_3085);
nor U4740 (N_4740,N_3970,N_3141);
nor U4741 (N_4741,N_3841,N_3612);
xnor U4742 (N_4742,N_3633,N_3804);
or U4743 (N_4743,N_3644,N_3664);
nor U4744 (N_4744,N_3526,N_3695);
xor U4745 (N_4745,N_3227,N_3616);
or U4746 (N_4746,N_3562,N_3695);
xor U4747 (N_4747,N_3609,N_3150);
xnor U4748 (N_4748,N_3598,N_3189);
or U4749 (N_4749,N_3102,N_3838);
nor U4750 (N_4750,N_3157,N_3289);
or U4751 (N_4751,N_3919,N_3459);
xor U4752 (N_4752,N_3697,N_3263);
nand U4753 (N_4753,N_3803,N_3113);
nor U4754 (N_4754,N_3534,N_3226);
or U4755 (N_4755,N_3388,N_3576);
and U4756 (N_4756,N_3922,N_3267);
nor U4757 (N_4757,N_3175,N_3795);
or U4758 (N_4758,N_3113,N_3372);
xor U4759 (N_4759,N_3955,N_3949);
nand U4760 (N_4760,N_3555,N_3356);
and U4761 (N_4761,N_3008,N_3296);
or U4762 (N_4762,N_3008,N_3780);
or U4763 (N_4763,N_3773,N_3984);
nand U4764 (N_4764,N_3235,N_3178);
nand U4765 (N_4765,N_3206,N_3889);
xnor U4766 (N_4766,N_3767,N_3399);
nor U4767 (N_4767,N_3195,N_3048);
or U4768 (N_4768,N_3815,N_3151);
nor U4769 (N_4769,N_3781,N_3683);
and U4770 (N_4770,N_3663,N_3548);
xor U4771 (N_4771,N_3593,N_3590);
nand U4772 (N_4772,N_3080,N_3344);
or U4773 (N_4773,N_3596,N_3610);
and U4774 (N_4774,N_3586,N_3046);
nand U4775 (N_4775,N_3959,N_3075);
nand U4776 (N_4776,N_3827,N_3585);
xor U4777 (N_4777,N_3806,N_3110);
nor U4778 (N_4778,N_3460,N_3576);
nor U4779 (N_4779,N_3403,N_3928);
nand U4780 (N_4780,N_3841,N_3310);
nand U4781 (N_4781,N_3411,N_3680);
and U4782 (N_4782,N_3254,N_3548);
xnor U4783 (N_4783,N_3449,N_3994);
xor U4784 (N_4784,N_3354,N_3803);
or U4785 (N_4785,N_3513,N_3503);
nor U4786 (N_4786,N_3442,N_3075);
nand U4787 (N_4787,N_3407,N_3580);
nand U4788 (N_4788,N_3427,N_3065);
and U4789 (N_4789,N_3081,N_3382);
and U4790 (N_4790,N_3981,N_3363);
or U4791 (N_4791,N_3956,N_3338);
nand U4792 (N_4792,N_3478,N_3943);
nand U4793 (N_4793,N_3354,N_3263);
and U4794 (N_4794,N_3749,N_3922);
or U4795 (N_4795,N_3579,N_3338);
or U4796 (N_4796,N_3495,N_3136);
or U4797 (N_4797,N_3386,N_3485);
or U4798 (N_4798,N_3586,N_3776);
or U4799 (N_4799,N_3499,N_3243);
and U4800 (N_4800,N_3532,N_3775);
and U4801 (N_4801,N_3185,N_3242);
and U4802 (N_4802,N_3431,N_3683);
nor U4803 (N_4803,N_3164,N_3024);
nand U4804 (N_4804,N_3473,N_3465);
or U4805 (N_4805,N_3392,N_3043);
nor U4806 (N_4806,N_3332,N_3685);
or U4807 (N_4807,N_3218,N_3823);
xnor U4808 (N_4808,N_3359,N_3645);
xor U4809 (N_4809,N_3367,N_3063);
or U4810 (N_4810,N_3835,N_3747);
and U4811 (N_4811,N_3466,N_3353);
and U4812 (N_4812,N_3059,N_3283);
and U4813 (N_4813,N_3342,N_3514);
xnor U4814 (N_4814,N_3843,N_3157);
and U4815 (N_4815,N_3981,N_3684);
xor U4816 (N_4816,N_3280,N_3011);
nor U4817 (N_4817,N_3641,N_3323);
xnor U4818 (N_4818,N_3783,N_3970);
xnor U4819 (N_4819,N_3329,N_3592);
nor U4820 (N_4820,N_3844,N_3958);
or U4821 (N_4821,N_3590,N_3084);
nand U4822 (N_4822,N_3727,N_3620);
xnor U4823 (N_4823,N_3636,N_3573);
nor U4824 (N_4824,N_3554,N_3110);
xor U4825 (N_4825,N_3974,N_3852);
and U4826 (N_4826,N_3663,N_3077);
and U4827 (N_4827,N_3879,N_3406);
or U4828 (N_4828,N_3141,N_3541);
nand U4829 (N_4829,N_3446,N_3811);
and U4830 (N_4830,N_3323,N_3929);
or U4831 (N_4831,N_3986,N_3264);
xnor U4832 (N_4832,N_3523,N_3350);
or U4833 (N_4833,N_3853,N_3272);
nand U4834 (N_4834,N_3843,N_3076);
and U4835 (N_4835,N_3850,N_3375);
xor U4836 (N_4836,N_3297,N_3959);
nand U4837 (N_4837,N_3656,N_3114);
nand U4838 (N_4838,N_3786,N_3563);
or U4839 (N_4839,N_3144,N_3746);
or U4840 (N_4840,N_3756,N_3194);
nor U4841 (N_4841,N_3193,N_3044);
and U4842 (N_4842,N_3807,N_3041);
nand U4843 (N_4843,N_3228,N_3354);
or U4844 (N_4844,N_3612,N_3846);
or U4845 (N_4845,N_3210,N_3981);
and U4846 (N_4846,N_3153,N_3448);
xnor U4847 (N_4847,N_3368,N_3840);
nor U4848 (N_4848,N_3343,N_3349);
nor U4849 (N_4849,N_3160,N_3611);
nand U4850 (N_4850,N_3612,N_3316);
nor U4851 (N_4851,N_3909,N_3420);
or U4852 (N_4852,N_3719,N_3927);
or U4853 (N_4853,N_3148,N_3215);
xor U4854 (N_4854,N_3007,N_3564);
nand U4855 (N_4855,N_3437,N_3763);
nor U4856 (N_4856,N_3073,N_3748);
nor U4857 (N_4857,N_3836,N_3478);
or U4858 (N_4858,N_3952,N_3045);
and U4859 (N_4859,N_3750,N_3094);
and U4860 (N_4860,N_3786,N_3236);
and U4861 (N_4861,N_3505,N_3261);
and U4862 (N_4862,N_3935,N_3741);
nand U4863 (N_4863,N_3642,N_3971);
and U4864 (N_4864,N_3660,N_3312);
or U4865 (N_4865,N_3100,N_3981);
nand U4866 (N_4866,N_3108,N_3294);
and U4867 (N_4867,N_3746,N_3516);
nand U4868 (N_4868,N_3981,N_3140);
nor U4869 (N_4869,N_3980,N_3647);
nor U4870 (N_4870,N_3996,N_3292);
or U4871 (N_4871,N_3657,N_3590);
or U4872 (N_4872,N_3764,N_3498);
or U4873 (N_4873,N_3605,N_3324);
or U4874 (N_4874,N_3026,N_3855);
nand U4875 (N_4875,N_3127,N_3181);
nand U4876 (N_4876,N_3851,N_3610);
xnor U4877 (N_4877,N_3452,N_3500);
and U4878 (N_4878,N_3133,N_3281);
nor U4879 (N_4879,N_3274,N_3694);
xor U4880 (N_4880,N_3950,N_3582);
nor U4881 (N_4881,N_3694,N_3360);
and U4882 (N_4882,N_3546,N_3120);
nor U4883 (N_4883,N_3657,N_3869);
and U4884 (N_4884,N_3017,N_3460);
and U4885 (N_4885,N_3208,N_3130);
nand U4886 (N_4886,N_3771,N_3382);
xnor U4887 (N_4887,N_3431,N_3971);
nand U4888 (N_4888,N_3023,N_3779);
nand U4889 (N_4889,N_3898,N_3308);
or U4890 (N_4890,N_3526,N_3720);
nand U4891 (N_4891,N_3075,N_3362);
and U4892 (N_4892,N_3475,N_3050);
or U4893 (N_4893,N_3708,N_3684);
and U4894 (N_4894,N_3468,N_3196);
nand U4895 (N_4895,N_3571,N_3902);
xnor U4896 (N_4896,N_3619,N_3757);
nor U4897 (N_4897,N_3666,N_3512);
nor U4898 (N_4898,N_3562,N_3771);
nor U4899 (N_4899,N_3597,N_3647);
or U4900 (N_4900,N_3466,N_3528);
and U4901 (N_4901,N_3175,N_3889);
xnor U4902 (N_4902,N_3619,N_3748);
or U4903 (N_4903,N_3439,N_3317);
xor U4904 (N_4904,N_3584,N_3669);
and U4905 (N_4905,N_3724,N_3607);
and U4906 (N_4906,N_3488,N_3189);
nand U4907 (N_4907,N_3451,N_3854);
or U4908 (N_4908,N_3991,N_3281);
nand U4909 (N_4909,N_3805,N_3013);
or U4910 (N_4910,N_3406,N_3489);
nand U4911 (N_4911,N_3375,N_3410);
nand U4912 (N_4912,N_3163,N_3823);
nand U4913 (N_4913,N_3419,N_3059);
nor U4914 (N_4914,N_3534,N_3784);
or U4915 (N_4915,N_3680,N_3787);
and U4916 (N_4916,N_3274,N_3940);
and U4917 (N_4917,N_3241,N_3900);
xor U4918 (N_4918,N_3582,N_3000);
nand U4919 (N_4919,N_3614,N_3315);
and U4920 (N_4920,N_3865,N_3488);
nand U4921 (N_4921,N_3603,N_3269);
and U4922 (N_4922,N_3059,N_3215);
nand U4923 (N_4923,N_3578,N_3761);
nor U4924 (N_4924,N_3437,N_3934);
nand U4925 (N_4925,N_3791,N_3117);
nor U4926 (N_4926,N_3839,N_3466);
or U4927 (N_4927,N_3419,N_3617);
nor U4928 (N_4928,N_3123,N_3376);
xnor U4929 (N_4929,N_3830,N_3561);
xor U4930 (N_4930,N_3169,N_3812);
nand U4931 (N_4931,N_3989,N_3474);
or U4932 (N_4932,N_3716,N_3005);
nand U4933 (N_4933,N_3745,N_3870);
or U4934 (N_4934,N_3623,N_3244);
and U4935 (N_4935,N_3022,N_3511);
and U4936 (N_4936,N_3037,N_3851);
and U4937 (N_4937,N_3839,N_3818);
nand U4938 (N_4938,N_3544,N_3719);
and U4939 (N_4939,N_3937,N_3070);
and U4940 (N_4940,N_3377,N_3464);
nand U4941 (N_4941,N_3438,N_3801);
and U4942 (N_4942,N_3152,N_3280);
and U4943 (N_4943,N_3868,N_3330);
nand U4944 (N_4944,N_3420,N_3827);
nor U4945 (N_4945,N_3241,N_3949);
nor U4946 (N_4946,N_3305,N_3566);
nor U4947 (N_4947,N_3472,N_3321);
or U4948 (N_4948,N_3139,N_3232);
xnor U4949 (N_4949,N_3518,N_3177);
xor U4950 (N_4950,N_3106,N_3787);
nor U4951 (N_4951,N_3574,N_3401);
or U4952 (N_4952,N_3835,N_3783);
nand U4953 (N_4953,N_3342,N_3822);
or U4954 (N_4954,N_3784,N_3351);
nor U4955 (N_4955,N_3566,N_3139);
and U4956 (N_4956,N_3189,N_3931);
xor U4957 (N_4957,N_3074,N_3674);
and U4958 (N_4958,N_3667,N_3226);
or U4959 (N_4959,N_3994,N_3047);
nor U4960 (N_4960,N_3112,N_3345);
or U4961 (N_4961,N_3304,N_3263);
nand U4962 (N_4962,N_3399,N_3151);
and U4963 (N_4963,N_3835,N_3655);
nand U4964 (N_4964,N_3546,N_3400);
xor U4965 (N_4965,N_3990,N_3803);
xor U4966 (N_4966,N_3803,N_3378);
nand U4967 (N_4967,N_3494,N_3359);
nor U4968 (N_4968,N_3819,N_3029);
or U4969 (N_4969,N_3033,N_3137);
nor U4970 (N_4970,N_3440,N_3893);
and U4971 (N_4971,N_3402,N_3651);
nor U4972 (N_4972,N_3112,N_3774);
and U4973 (N_4973,N_3894,N_3884);
and U4974 (N_4974,N_3060,N_3733);
and U4975 (N_4975,N_3135,N_3626);
or U4976 (N_4976,N_3095,N_3756);
or U4977 (N_4977,N_3084,N_3889);
or U4978 (N_4978,N_3226,N_3508);
or U4979 (N_4979,N_3885,N_3538);
xor U4980 (N_4980,N_3707,N_3554);
xnor U4981 (N_4981,N_3191,N_3049);
or U4982 (N_4982,N_3579,N_3576);
nor U4983 (N_4983,N_3969,N_3295);
and U4984 (N_4984,N_3516,N_3345);
or U4985 (N_4985,N_3821,N_3240);
nand U4986 (N_4986,N_3335,N_3436);
nand U4987 (N_4987,N_3115,N_3718);
or U4988 (N_4988,N_3052,N_3545);
or U4989 (N_4989,N_3041,N_3150);
nand U4990 (N_4990,N_3520,N_3951);
nor U4991 (N_4991,N_3254,N_3162);
nor U4992 (N_4992,N_3945,N_3966);
or U4993 (N_4993,N_3038,N_3895);
or U4994 (N_4994,N_3233,N_3855);
or U4995 (N_4995,N_3996,N_3864);
and U4996 (N_4996,N_3551,N_3176);
nand U4997 (N_4997,N_3534,N_3466);
and U4998 (N_4998,N_3899,N_3119);
or U4999 (N_4999,N_3951,N_3072);
nor U5000 (N_5000,N_4623,N_4282);
nand U5001 (N_5001,N_4577,N_4483);
nand U5002 (N_5002,N_4021,N_4436);
and U5003 (N_5003,N_4299,N_4293);
or U5004 (N_5004,N_4074,N_4938);
nand U5005 (N_5005,N_4934,N_4118);
or U5006 (N_5006,N_4472,N_4316);
or U5007 (N_5007,N_4978,N_4538);
nor U5008 (N_5008,N_4261,N_4106);
nor U5009 (N_5009,N_4552,N_4053);
or U5010 (N_5010,N_4831,N_4659);
nand U5011 (N_5011,N_4460,N_4789);
nor U5012 (N_5012,N_4794,N_4433);
xor U5013 (N_5013,N_4264,N_4758);
or U5014 (N_5014,N_4712,N_4802);
nand U5015 (N_5015,N_4543,N_4320);
nor U5016 (N_5016,N_4667,N_4216);
nor U5017 (N_5017,N_4816,N_4829);
and U5018 (N_5018,N_4446,N_4920);
and U5019 (N_5019,N_4176,N_4398);
nor U5020 (N_5020,N_4211,N_4757);
and U5021 (N_5021,N_4926,N_4510);
nand U5022 (N_5022,N_4091,N_4057);
or U5023 (N_5023,N_4513,N_4346);
nor U5024 (N_5024,N_4078,N_4533);
or U5025 (N_5025,N_4677,N_4358);
or U5026 (N_5026,N_4896,N_4917);
nor U5027 (N_5027,N_4050,N_4773);
xor U5028 (N_5028,N_4144,N_4394);
or U5029 (N_5029,N_4471,N_4891);
or U5030 (N_5030,N_4930,N_4806);
xnor U5031 (N_5031,N_4683,N_4412);
nand U5032 (N_5032,N_4991,N_4127);
nand U5033 (N_5033,N_4808,N_4632);
or U5034 (N_5034,N_4355,N_4395);
nand U5035 (N_5035,N_4351,N_4760);
xnor U5036 (N_5036,N_4734,N_4788);
xnor U5037 (N_5037,N_4933,N_4307);
or U5038 (N_5038,N_4912,N_4479);
or U5039 (N_5039,N_4180,N_4588);
nor U5040 (N_5040,N_4907,N_4418);
nand U5041 (N_5041,N_4833,N_4321);
or U5042 (N_5042,N_4646,N_4255);
or U5043 (N_5043,N_4243,N_4855);
or U5044 (N_5044,N_4524,N_4842);
or U5045 (N_5045,N_4849,N_4569);
xnor U5046 (N_5046,N_4288,N_4850);
or U5047 (N_5047,N_4685,N_4182);
xnor U5048 (N_5048,N_4923,N_4553);
and U5049 (N_5049,N_4691,N_4033);
and U5050 (N_5050,N_4694,N_4283);
nor U5051 (N_5051,N_4972,N_4813);
nand U5052 (N_5052,N_4340,N_4408);
nor U5053 (N_5053,N_4751,N_4130);
and U5054 (N_5054,N_4034,N_4464);
xor U5055 (N_5055,N_4109,N_4890);
nor U5056 (N_5056,N_4804,N_4970);
xnor U5057 (N_5057,N_4983,N_4442);
nand U5058 (N_5058,N_4402,N_4542);
nand U5059 (N_5059,N_4413,N_4003);
nor U5060 (N_5060,N_4429,N_4156);
nor U5061 (N_5061,N_4837,N_4603);
nand U5062 (N_5062,N_4946,N_4864);
xor U5063 (N_5063,N_4012,N_4092);
and U5064 (N_5064,N_4810,N_4680);
nand U5065 (N_5065,N_4707,N_4382);
nor U5066 (N_5066,N_4531,N_4690);
or U5067 (N_5067,N_4763,N_4620);
nor U5068 (N_5068,N_4625,N_4766);
nor U5069 (N_5069,N_4624,N_4187);
and U5070 (N_5070,N_4103,N_4207);
nand U5071 (N_5071,N_4304,N_4893);
xor U5072 (N_5072,N_4640,N_4824);
and U5073 (N_5073,N_4771,N_4076);
or U5074 (N_5074,N_4518,N_4090);
xor U5075 (N_5075,N_4517,N_4098);
nor U5076 (N_5076,N_4062,N_4750);
nand U5077 (N_5077,N_4800,N_4753);
nand U5078 (N_5078,N_4449,N_4173);
and U5079 (N_5079,N_4922,N_4245);
nor U5080 (N_5080,N_4140,N_4637);
or U5081 (N_5081,N_4489,N_4242);
nand U5082 (N_5082,N_4055,N_4997);
xnor U5083 (N_5083,N_4452,N_4727);
xor U5084 (N_5084,N_4230,N_4841);
nand U5085 (N_5085,N_4411,N_4966);
or U5086 (N_5086,N_4698,N_4294);
xor U5087 (N_5087,N_4328,N_4882);
xnor U5088 (N_5088,N_4693,N_4768);
and U5089 (N_5089,N_4711,N_4740);
nor U5090 (N_5090,N_4585,N_4780);
xor U5091 (N_5091,N_4819,N_4861);
nand U5092 (N_5092,N_4277,N_4581);
xnor U5093 (N_5093,N_4499,N_4765);
nand U5094 (N_5094,N_4774,N_4183);
xor U5095 (N_5095,N_4713,N_4641);
nand U5096 (N_5096,N_4171,N_4032);
nor U5097 (N_5097,N_4146,N_4086);
xnor U5098 (N_5098,N_4152,N_4404);
xor U5099 (N_5099,N_4291,N_4077);
or U5100 (N_5100,N_4162,N_4611);
nor U5101 (N_5101,N_4338,N_4201);
and U5102 (N_5102,N_4072,N_4224);
and U5103 (N_5103,N_4915,N_4481);
and U5104 (N_5104,N_4593,N_4151);
and U5105 (N_5105,N_4082,N_4035);
nand U5106 (N_5106,N_4018,N_4823);
nor U5107 (N_5107,N_4326,N_4237);
nor U5108 (N_5108,N_4847,N_4700);
and U5109 (N_5109,N_4134,N_4164);
or U5110 (N_5110,N_4105,N_4486);
xor U5111 (N_5111,N_4002,N_4225);
or U5112 (N_5112,N_4633,N_4434);
xnor U5113 (N_5113,N_4631,N_4571);
and U5114 (N_5114,N_4607,N_4403);
and U5115 (N_5115,N_4252,N_4929);
nand U5116 (N_5116,N_4600,N_4276);
or U5117 (N_5117,N_4424,N_4662);
and U5118 (N_5118,N_4107,N_4960);
and U5119 (N_5119,N_4241,N_4166);
xor U5120 (N_5120,N_4254,N_4142);
xnor U5121 (N_5121,N_4303,N_4451);
and U5122 (N_5122,N_4122,N_4781);
and U5123 (N_5123,N_4139,N_4958);
xor U5124 (N_5124,N_4115,N_4535);
nor U5125 (N_5125,N_4016,N_4844);
nor U5126 (N_5126,N_4342,N_4744);
xnor U5127 (N_5127,N_4329,N_4888);
xnor U5128 (N_5128,N_4463,N_4605);
xor U5129 (N_5129,N_4121,N_4526);
nor U5130 (N_5130,N_4557,N_4023);
xnor U5131 (N_5131,N_4423,N_4163);
nor U5132 (N_5132,N_4560,N_4881);
nand U5133 (N_5133,N_4132,N_4634);
and U5134 (N_5134,N_4584,N_4330);
or U5135 (N_5135,N_4809,N_4573);
xor U5136 (N_5136,N_4942,N_4722);
or U5137 (N_5137,N_4879,N_4520);
and U5138 (N_5138,N_4601,N_4537);
or U5139 (N_5139,N_4719,N_4953);
and U5140 (N_5140,N_4515,N_4563);
nor U5141 (N_5141,N_4431,N_4791);
or U5142 (N_5142,N_4678,N_4718);
xnor U5143 (N_5143,N_4961,N_4417);
xnor U5144 (N_5144,N_4393,N_4415);
xor U5145 (N_5145,N_4026,N_4478);
xnor U5146 (N_5146,N_4410,N_4653);
and U5147 (N_5147,N_4370,N_4206);
xnor U5148 (N_5148,N_4660,N_4337);
nand U5149 (N_5149,N_4811,N_4219);
nand U5150 (N_5150,N_4209,N_4046);
xnor U5151 (N_5151,N_4422,N_4948);
xor U5152 (N_5152,N_4143,N_4238);
and U5153 (N_5153,N_4221,N_4854);
xor U5154 (N_5154,N_4188,N_4777);
and U5155 (N_5155,N_4795,N_4742);
nand U5156 (N_5156,N_4281,N_4706);
or U5157 (N_5157,N_4570,N_4544);
nor U5158 (N_5158,N_4014,N_4373);
nand U5159 (N_5159,N_4167,N_4863);
nand U5160 (N_5160,N_4598,N_4709);
nand U5161 (N_5161,N_4636,N_4372);
and U5162 (N_5162,N_4889,N_4582);
nand U5163 (N_5163,N_4686,N_4068);
xnor U5164 (N_5164,N_4285,N_4916);
and U5165 (N_5165,N_4097,N_4903);
and U5166 (N_5166,N_4721,N_4732);
nand U5167 (N_5167,N_4295,N_4250);
or U5168 (N_5168,N_4170,N_4738);
xor U5169 (N_5169,N_4843,N_4583);
nor U5170 (N_5170,N_4733,N_4060);
nand U5171 (N_5171,N_4931,N_4400);
nor U5172 (N_5172,N_4943,N_4967);
or U5173 (N_5173,N_4317,N_4473);
xor U5174 (N_5174,N_4001,N_4739);
and U5175 (N_5175,N_4038,N_4042);
xor U5176 (N_5176,N_4987,N_4749);
xnor U5177 (N_5177,N_4503,N_4214);
or U5178 (N_5178,N_4880,N_4244);
or U5179 (N_5179,N_4939,N_4432);
xnor U5180 (N_5180,N_4703,N_4101);
nor U5181 (N_5181,N_4562,N_4778);
nor U5182 (N_5182,N_4969,N_4704);
and U5183 (N_5183,N_4477,N_4852);
xnor U5184 (N_5184,N_4364,N_4821);
xnor U5185 (N_5185,N_4947,N_4856);
nand U5186 (N_5186,N_4494,N_4131);
and U5187 (N_5187,N_4595,N_4697);
nor U5188 (N_5188,N_4665,N_4755);
or U5189 (N_5189,N_4061,N_4935);
xor U5190 (N_5190,N_4735,N_4249);
nor U5191 (N_5191,N_4487,N_4608);
or U5192 (N_5192,N_4696,N_4671);
or U5193 (N_5193,N_4467,N_4391);
or U5194 (N_5194,N_4007,N_4054);
xor U5195 (N_5195,N_4507,N_4797);
xnor U5196 (N_5196,N_4271,N_4807);
nand U5197 (N_5197,N_4325,N_4482);
or U5198 (N_5198,N_4825,N_4724);
nor U5199 (N_5199,N_4871,N_4799);
xor U5200 (N_5200,N_4558,N_4309);
nand U5201 (N_5201,N_4367,N_4361);
xnor U5202 (N_5202,N_4204,N_4610);
nand U5203 (N_5203,N_4918,N_4009);
or U5204 (N_5204,N_4857,N_4462);
nand U5205 (N_5205,N_4616,N_4664);
nand U5206 (N_5206,N_4450,N_4902);
nand U5207 (N_5207,N_4315,N_4874);
and U5208 (N_5208,N_4123,N_4792);
or U5209 (N_5209,N_4908,N_4215);
xor U5210 (N_5210,N_4318,N_4022);
and U5211 (N_5211,N_4924,N_4530);
and U5212 (N_5212,N_4651,N_4335);
or U5213 (N_5213,N_4070,N_4787);
nand U5214 (N_5214,N_4095,N_4615);
or U5215 (N_5215,N_4897,N_4976);
nor U5216 (N_5216,N_4602,N_4913);
nor U5217 (N_5217,N_4425,N_4622);
nor U5218 (N_5218,N_4154,N_4591);
nand U5219 (N_5219,N_4228,N_4996);
nand U5220 (N_5220,N_4990,N_4617);
nand U5221 (N_5221,N_4561,N_4455);
nor U5222 (N_5222,N_4223,N_4401);
nand U5223 (N_5223,N_4365,N_4812);
nand U5224 (N_5224,N_4521,N_4576);
xnor U5225 (N_5225,N_4292,N_4974);
and U5226 (N_5226,N_4168,N_4748);
and U5227 (N_5227,N_4147,N_4716);
nor U5228 (N_5228,N_4199,N_4392);
or U5229 (N_5229,N_4052,N_4312);
nor U5230 (N_5230,N_4783,N_4975);
nor U5231 (N_5231,N_4165,N_4754);
and U5232 (N_5232,N_4456,N_4347);
or U5233 (N_5233,N_4387,N_4441);
nor U5234 (N_5234,N_4944,N_4084);
xor U5235 (N_5235,N_4759,N_4905);
and U5236 (N_5236,N_4150,N_4246);
nor U5237 (N_5237,N_4448,N_4222);
and U5238 (N_5238,N_4865,N_4957);
nor U5239 (N_5239,N_4604,N_4454);
nor U5240 (N_5240,N_4301,N_4687);
nand U5241 (N_5241,N_4100,N_4005);
nor U5242 (N_5242,N_4772,N_4549);
nor U5243 (N_5243,N_4884,N_4323);
nand U5244 (N_5244,N_4289,N_4803);
nand U5245 (N_5245,N_4814,N_4626);
nand U5246 (N_5246,N_4045,N_4348);
or U5247 (N_5247,N_4087,N_4112);
nand U5248 (N_5248,N_4971,N_4838);
nor U5249 (N_5249,N_4937,N_4159);
nor U5250 (N_5250,N_4419,N_4314);
nor U5251 (N_5251,N_4669,N_4233);
nand U5252 (N_5252,N_4438,N_4149);
xor U5253 (N_5253,N_4786,N_4067);
xnor U5254 (N_5254,N_4208,N_4220);
and U5255 (N_5255,N_4440,N_4037);
or U5256 (N_5256,N_4488,N_4682);
nor U5257 (N_5257,N_4505,N_4073);
nand U5258 (N_5258,N_4259,N_4263);
nand U5259 (N_5259,N_4476,N_4534);
nand U5260 (N_5260,N_4684,N_4927);
nor U5261 (N_5261,N_4267,N_4752);
xnor U5262 (N_5262,N_4430,N_4239);
xor U5263 (N_5263,N_4284,N_4217);
nor U5264 (N_5264,N_4193,N_4555);
or U5265 (N_5265,N_4203,N_4114);
nor U5266 (N_5266,N_4546,N_4426);
nor U5267 (N_5267,N_4652,N_4029);
and U5268 (N_5268,N_4189,N_4240);
or U5269 (N_5269,N_4845,N_4248);
and U5270 (N_5270,N_4491,N_4088);
nand U5271 (N_5271,N_4470,N_4679);
xnor U5272 (N_5272,N_4554,N_4213);
xnor U5273 (N_5273,N_4296,N_4099);
xnor U5274 (N_5274,N_4715,N_4689);
xnor U5275 (N_5275,N_4699,N_4069);
or U5276 (N_5276,N_4185,N_4878);
nor U5277 (N_5277,N_4688,N_4374);
or U5278 (N_5278,N_4195,N_4728);
nor U5279 (N_5279,N_4331,N_4936);
and U5280 (N_5280,N_4859,N_4514);
xor U5281 (N_5281,N_4272,N_4994);
and U5282 (N_5282,N_4117,N_4049);
and U5283 (N_5283,N_4984,N_4258);
or U5284 (N_5284,N_4396,N_4904);
nand U5285 (N_5285,N_4028,N_4349);
xor U5286 (N_5286,N_4275,N_4089);
and U5287 (N_5287,N_4390,N_4172);
xor U5288 (N_5288,N_4319,N_4815);
nor U5289 (N_5289,N_4104,N_4357);
nor U5290 (N_5290,N_4725,N_4059);
nand U5291 (N_5291,N_4663,N_4643);
nand U5292 (N_5292,N_4767,N_4041);
nand U5293 (N_5293,N_4564,N_4369);
nand U5294 (N_5294,N_4359,N_4710);
nand U5295 (N_5295,N_4770,N_4645);
and U5296 (N_5296,N_4898,N_4932);
or U5297 (N_5297,N_4386,N_4895);
or U5298 (N_5298,N_4327,N_4399);
nor U5299 (N_5299,N_4835,N_4036);
nor U5300 (N_5300,N_4899,N_4673);
nand U5301 (N_5301,N_4736,N_4234);
or U5302 (N_5302,N_4305,N_4928);
or U5303 (N_5303,N_4551,N_4614);
nor U5304 (N_5304,N_4981,N_4498);
nand U5305 (N_5305,N_4226,N_4674);
or U5306 (N_5306,N_4366,N_4290);
and U5307 (N_5307,N_4818,N_4043);
xnor U5308 (N_5308,N_4236,N_4579);
and U5309 (N_5309,N_4065,N_4421);
or U5310 (N_5310,N_4726,N_4025);
and U5311 (N_5311,N_4468,N_4108);
or U5312 (N_5312,N_4324,N_4322);
xor U5313 (N_5313,N_4137,N_4385);
nor U5314 (N_5314,N_4894,N_4253);
xor U5315 (N_5315,N_4764,N_4982);
xnor U5316 (N_5316,N_4876,N_4378);
xor U5317 (N_5317,N_4820,N_4790);
or U5318 (N_5318,N_4516,N_4523);
or U5319 (N_5319,N_4145,N_4251);
or U5320 (N_5320,N_4492,N_4302);
nand U5321 (N_5321,N_4497,N_4853);
and U5322 (N_5322,N_4658,N_4247);
and U5323 (N_5323,N_4968,N_4093);
nand U5324 (N_5324,N_4495,N_4020);
xor U5325 (N_5325,N_4031,N_4197);
nor U5326 (N_5326,N_4868,N_4475);
or U5327 (N_5327,N_4177,N_4741);
nor U5328 (N_5328,N_4527,N_4599);
nand U5329 (N_5329,N_4836,N_4407);
xnor U5330 (N_5330,N_4427,N_4877);
and U5331 (N_5331,N_4262,N_4529);
or U5332 (N_5332,N_4039,N_4138);
nor U5333 (N_5333,N_4609,N_4649);
or U5334 (N_5334,N_4414,N_4545);
and U5335 (N_5335,N_4550,N_4509);
xor U5336 (N_5336,N_4071,N_4257);
or U5337 (N_5337,N_4575,N_4175);
and U5338 (N_5338,N_4380,N_4941);
nand U5339 (N_5339,N_4190,N_4962);
and U5340 (N_5340,N_4474,N_4126);
and U5341 (N_5341,N_4278,N_4191);
nand U5342 (N_5342,N_4873,N_4119);
nand U5343 (N_5343,N_4011,N_4504);
and U5344 (N_5344,N_4096,N_4672);
or U5345 (N_5345,N_4532,N_4730);
nor U5346 (N_5346,N_4701,N_4848);
nand U5347 (N_5347,N_4914,N_4024);
or U5348 (N_5348,N_4298,N_4747);
and U5349 (N_5349,N_4959,N_4621);
xor U5350 (N_5350,N_4642,N_4875);
nand U5351 (N_5351,N_4501,N_4592);
xnor U5352 (N_5352,N_4830,N_4169);
xnor U5353 (N_5353,N_4862,N_4428);
and U5354 (N_5354,N_4851,N_4729);
nand U5355 (N_5355,N_4921,N_4784);
or U5356 (N_5356,N_4083,N_4801);
or U5357 (N_5357,N_4695,N_4860);
and U5358 (N_5358,N_4416,N_4574);
nor U5359 (N_5359,N_4120,N_4980);
nand U5360 (N_5360,N_4508,N_4158);
xnor U5361 (N_5361,N_4639,N_4113);
nand U5362 (N_5362,N_4568,N_4619);
and U5363 (N_5363,N_4834,N_4556);
nor U5364 (N_5364,N_4965,N_4827);
and U5365 (N_5365,N_4354,N_4995);
or U5366 (N_5366,N_4629,N_4776);
and U5367 (N_5367,N_4313,N_4040);
or U5368 (N_5368,N_4279,N_4133);
or U5369 (N_5369,N_4080,N_4260);
xnor U5370 (N_5370,N_4157,N_4368);
nor U5371 (N_5371,N_4465,N_4480);
nor U5372 (N_5372,N_4461,N_4332);
xnor U5373 (N_5373,N_4048,N_4128);
nand U5374 (N_5374,N_4940,N_4381);
nor U5375 (N_5375,N_4343,N_4085);
nor U5376 (N_5376,N_4647,N_4989);
or U5377 (N_5377,N_4746,N_4160);
nor U5378 (N_5378,N_4388,N_4883);
xor U5379 (N_5379,N_4435,N_4056);
nand U5380 (N_5380,N_4136,N_4153);
and U5381 (N_5381,N_4951,N_4779);
nand U5382 (N_5382,N_4075,N_4785);
nand U5383 (N_5383,N_4443,N_4900);
and U5384 (N_5384,N_4828,N_4949);
nor U5385 (N_5385,N_4963,N_4867);
or U5386 (N_5386,N_4266,N_4178);
and U5387 (N_5387,N_4596,N_4110);
or U5388 (N_5388,N_4743,N_4079);
or U5389 (N_5389,N_4692,N_4306);
or U5390 (N_5390,N_4397,N_4578);
or U5391 (N_5391,N_4566,N_4384);
and U5392 (N_5392,N_4988,N_4590);
or U5393 (N_5393,N_4998,N_4661);
and U5394 (N_5394,N_4594,N_4184);
or U5395 (N_5395,N_4437,N_4612);
nor U5396 (N_5396,N_4287,N_4270);
and U5397 (N_5397,N_4004,N_4124);
or U5398 (N_5398,N_4511,N_4539);
and U5399 (N_5399,N_4352,N_4606);
nor U5400 (N_5400,N_4027,N_4064);
xnor U5401 (N_5401,N_4447,N_4116);
nor U5402 (N_5402,N_4668,N_4840);
or U5403 (N_5403,N_4453,N_4383);
or U5404 (N_5404,N_4286,N_4227);
or U5405 (N_5405,N_4702,N_4496);
nand U5406 (N_5406,N_4200,N_4565);
xor U5407 (N_5407,N_4015,N_4232);
nand U5408 (N_5408,N_4886,N_4212);
xor U5409 (N_5409,N_4644,N_4363);
nand U5410 (N_5410,N_4058,N_4008);
or U5411 (N_5411,N_4256,N_4376);
and U5412 (N_5412,N_4627,N_4409);
or U5413 (N_5413,N_4310,N_4405);
or U5414 (N_5414,N_4798,N_4648);
nand U5415 (N_5415,N_4141,N_4000);
or U5416 (N_5416,N_4179,N_4181);
or U5417 (N_5417,N_4723,N_4379);
nor U5418 (N_5418,N_4775,N_4512);
xor U5419 (N_5419,N_4051,N_4580);
xnor U5420 (N_5420,N_4375,N_4210);
nor U5421 (N_5421,N_4955,N_4737);
or U5422 (N_5422,N_4300,N_4541);
and U5423 (N_5423,N_4274,N_4506);
or U5424 (N_5424,N_4782,N_4952);
and U5425 (N_5425,N_4638,N_4341);
nor U5426 (N_5426,N_4536,N_4676);
nand U5427 (N_5427,N_4964,N_4796);
nor U5428 (N_5428,N_4666,N_4202);
xnor U5429 (N_5429,N_4125,N_4469);
xnor U5430 (N_5430,N_4192,N_4205);
or U5431 (N_5431,N_4196,N_4635);
and U5432 (N_5432,N_4892,N_4377);
nor U5433 (N_5433,N_4484,N_4013);
or U5434 (N_5434,N_4406,N_4909);
nor U5435 (N_5435,N_4954,N_4458);
nor U5436 (N_5436,N_4589,N_4992);
and U5437 (N_5437,N_4817,N_4044);
nor U5438 (N_5438,N_4597,N_4910);
nor U5439 (N_5439,N_4805,N_4655);
nand U5440 (N_5440,N_4030,N_4887);
and U5441 (N_5441,N_4714,N_4360);
xor U5442 (N_5442,N_4656,N_4986);
and U5443 (N_5443,N_4870,N_4720);
nand U5444 (N_5444,N_4832,N_4650);
nand U5445 (N_5445,N_4102,N_4344);
and U5446 (N_5446,N_4705,N_4756);
or U5447 (N_5447,N_4519,N_4869);
nand U5448 (N_5448,N_4493,N_4280);
nor U5449 (N_5449,N_4528,N_4334);
nor U5450 (N_5450,N_4459,N_4950);
or U5451 (N_5451,N_4885,N_4587);
and U5452 (N_5452,N_4822,N_4135);
nor U5453 (N_5453,N_4567,N_4866);
and U5454 (N_5454,N_4846,N_4762);
and U5455 (N_5455,N_4129,N_4977);
or U5456 (N_5456,N_4457,N_4345);
nand U5457 (N_5457,N_4630,N_4269);
and U5458 (N_5458,N_4362,N_4973);
nand U5459 (N_5459,N_4066,N_4485);
or U5460 (N_5460,N_4444,N_4445);
nand U5461 (N_5461,N_4198,N_4708);
xor U5462 (N_5462,N_4420,N_4006);
xor U5463 (N_5463,N_4047,N_4745);
or U5464 (N_5464,N_4356,N_4613);
or U5465 (N_5465,N_4628,N_4161);
nand U5466 (N_5466,N_4872,N_4502);
xor U5467 (N_5467,N_4063,N_4559);
or U5468 (N_5468,N_4265,N_4731);
nand U5469 (N_5469,N_4229,N_4548);
xor U5470 (N_5470,N_4945,N_4333);
xnor U5471 (N_5471,N_4793,N_4350);
nand U5472 (N_5472,N_4901,N_4094);
and U5473 (N_5473,N_4155,N_4670);
nand U5474 (N_5474,N_4371,N_4081);
nand U5475 (N_5475,N_4389,N_4858);
xnor U5476 (N_5476,N_4769,N_4353);
or U5477 (N_5477,N_4999,N_4906);
nor U5478 (N_5478,N_4311,N_4572);
and U5479 (N_5479,N_4979,N_4231);
xor U5480 (N_5480,N_4174,N_4956);
xnor U5481 (N_5481,N_4268,N_4654);
and U5482 (N_5482,N_4466,N_4235);
xor U5483 (N_5483,N_4993,N_4194);
xnor U5484 (N_5484,N_4540,N_4218);
and U5485 (N_5485,N_4111,N_4911);
nor U5486 (N_5486,N_4826,N_4273);
nor U5487 (N_5487,N_4547,N_4985);
or U5488 (N_5488,N_4308,N_4717);
nand U5489 (N_5489,N_4586,N_4490);
and U5490 (N_5490,N_4525,N_4297);
or U5491 (N_5491,N_4500,N_4919);
or U5492 (N_5492,N_4186,N_4522);
nor U5493 (N_5493,N_4681,N_4010);
xor U5494 (N_5494,N_4761,N_4148);
and U5495 (N_5495,N_4339,N_4019);
xnor U5496 (N_5496,N_4839,N_4657);
or U5497 (N_5497,N_4017,N_4925);
and U5498 (N_5498,N_4618,N_4675);
xnor U5499 (N_5499,N_4336,N_4439);
xnor U5500 (N_5500,N_4635,N_4435);
nand U5501 (N_5501,N_4140,N_4159);
or U5502 (N_5502,N_4889,N_4054);
xor U5503 (N_5503,N_4331,N_4775);
nand U5504 (N_5504,N_4934,N_4935);
and U5505 (N_5505,N_4206,N_4214);
and U5506 (N_5506,N_4426,N_4402);
nor U5507 (N_5507,N_4969,N_4559);
and U5508 (N_5508,N_4329,N_4065);
and U5509 (N_5509,N_4983,N_4626);
or U5510 (N_5510,N_4601,N_4005);
and U5511 (N_5511,N_4689,N_4078);
nand U5512 (N_5512,N_4454,N_4536);
xnor U5513 (N_5513,N_4989,N_4026);
and U5514 (N_5514,N_4690,N_4896);
nand U5515 (N_5515,N_4969,N_4375);
nand U5516 (N_5516,N_4710,N_4580);
and U5517 (N_5517,N_4478,N_4552);
nor U5518 (N_5518,N_4985,N_4663);
nand U5519 (N_5519,N_4047,N_4470);
xor U5520 (N_5520,N_4178,N_4634);
nor U5521 (N_5521,N_4953,N_4246);
xnor U5522 (N_5522,N_4883,N_4343);
or U5523 (N_5523,N_4156,N_4113);
and U5524 (N_5524,N_4766,N_4176);
or U5525 (N_5525,N_4746,N_4698);
nand U5526 (N_5526,N_4189,N_4219);
nand U5527 (N_5527,N_4646,N_4673);
nor U5528 (N_5528,N_4582,N_4011);
xnor U5529 (N_5529,N_4614,N_4401);
nand U5530 (N_5530,N_4772,N_4331);
nand U5531 (N_5531,N_4404,N_4284);
or U5532 (N_5532,N_4085,N_4226);
and U5533 (N_5533,N_4825,N_4488);
xor U5534 (N_5534,N_4186,N_4286);
nand U5535 (N_5535,N_4245,N_4844);
nand U5536 (N_5536,N_4907,N_4332);
and U5537 (N_5537,N_4455,N_4224);
xnor U5538 (N_5538,N_4815,N_4313);
or U5539 (N_5539,N_4331,N_4167);
and U5540 (N_5540,N_4477,N_4108);
nor U5541 (N_5541,N_4134,N_4711);
or U5542 (N_5542,N_4382,N_4179);
nand U5543 (N_5543,N_4743,N_4383);
nor U5544 (N_5544,N_4893,N_4492);
xnor U5545 (N_5545,N_4583,N_4602);
or U5546 (N_5546,N_4577,N_4937);
nor U5547 (N_5547,N_4030,N_4547);
nor U5548 (N_5548,N_4713,N_4945);
nor U5549 (N_5549,N_4864,N_4010);
or U5550 (N_5550,N_4821,N_4949);
xor U5551 (N_5551,N_4601,N_4595);
or U5552 (N_5552,N_4525,N_4441);
xnor U5553 (N_5553,N_4659,N_4098);
nand U5554 (N_5554,N_4319,N_4335);
or U5555 (N_5555,N_4096,N_4517);
and U5556 (N_5556,N_4242,N_4547);
or U5557 (N_5557,N_4113,N_4852);
nand U5558 (N_5558,N_4202,N_4282);
nand U5559 (N_5559,N_4816,N_4759);
nand U5560 (N_5560,N_4693,N_4048);
xnor U5561 (N_5561,N_4361,N_4334);
and U5562 (N_5562,N_4874,N_4813);
nor U5563 (N_5563,N_4646,N_4592);
and U5564 (N_5564,N_4352,N_4965);
or U5565 (N_5565,N_4288,N_4452);
or U5566 (N_5566,N_4344,N_4949);
nand U5567 (N_5567,N_4304,N_4892);
nand U5568 (N_5568,N_4163,N_4739);
nor U5569 (N_5569,N_4273,N_4168);
nand U5570 (N_5570,N_4567,N_4164);
and U5571 (N_5571,N_4606,N_4599);
or U5572 (N_5572,N_4351,N_4148);
nand U5573 (N_5573,N_4689,N_4337);
xnor U5574 (N_5574,N_4653,N_4925);
nor U5575 (N_5575,N_4220,N_4032);
and U5576 (N_5576,N_4123,N_4770);
nor U5577 (N_5577,N_4474,N_4096);
or U5578 (N_5578,N_4729,N_4407);
xnor U5579 (N_5579,N_4449,N_4373);
or U5580 (N_5580,N_4644,N_4987);
or U5581 (N_5581,N_4188,N_4756);
and U5582 (N_5582,N_4508,N_4353);
nor U5583 (N_5583,N_4476,N_4748);
and U5584 (N_5584,N_4089,N_4827);
or U5585 (N_5585,N_4603,N_4509);
xnor U5586 (N_5586,N_4316,N_4665);
xnor U5587 (N_5587,N_4926,N_4196);
xor U5588 (N_5588,N_4968,N_4977);
nand U5589 (N_5589,N_4381,N_4886);
and U5590 (N_5590,N_4688,N_4394);
or U5591 (N_5591,N_4754,N_4331);
and U5592 (N_5592,N_4807,N_4437);
or U5593 (N_5593,N_4829,N_4358);
or U5594 (N_5594,N_4253,N_4531);
or U5595 (N_5595,N_4713,N_4588);
nand U5596 (N_5596,N_4870,N_4196);
xnor U5597 (N_5597,N_4864,N_4772);
nor U5598 (N_5598,N_4265,N_4220);
or U5599 (N_5599,N_4699,N_4123);
xor U5600 (N_5600,N_4288,N_4494);
or U5601 (N_5601,N_4046,N_4416);
nor U5602 (N_5602,N_4204,N_4075);
nand U5603 (N_5603,N_4525,N_4382);
nand U5604 (N_5604,N_4308,N_4213);
or U5605 (N_5605,N_4000,N_4995);
xor U5606 (N_5606,N_4305,N_4030);
and U5607 (N_5607,N_4069,N_4747);
and U5608 (N_5608,N_4867,N_4972);
xnor U5609 (N_5609,N_4956,N_4334);
xor U5610 (N_5610,N_4869,N_4640);
nand U5611 (N_5611,N_4270,N_4074);
nor U5612 (N_5612,N_4591,N_4357);
and U5613 (N_5613,N_4146,N_4849);
xor U5614 (N_5614,N_4923,N_4459);
and U5615 (N_5615,N_4990,N_4348);
and U5616 (N_5616,N_4295,N_4615);
xor U5617 (N_5617,N_4957,N_4166);
or U5618 (N_5618,N_4250,N_4405);
and U5619 (N_5619,N_4079,N_4141);
nor U5620 (N_5620,N_4948,N_4188);
nor U5621 (N_5621,N_4389,N_4830);
nand U5622 (N_5622,N_4829,N_4559);
nor U5623 (N_5623,N_4283,N_4781);
nor U5624 (N_5624,N_4316,N_4918);
and U5625 (N_5625,N_4645,N_4049);
nor U5626 (N_5626,N_4696,N_4402);
and U5627 (N_5627,N_4415,N_4389);
and U5628 (N_5628,N_4678,N_4943);
nand U5629 (N_5629,N_4350,N_4846);
xnor U5630 (N_5630,N_4820,N_4614);
nand U5631 (N_5631,N_4187,N_4629);
nand U5632 (N_5632,N_4745,N_4206);
or U5633 (N_5633,N_4738,N_4903);
xor U5634 (N_5634,N_4257,N_4441);
nor U5635 (N_5635,N_4732,N_4311);
or U5636 (N_5636,N_4039,N_4466);
and U5637 (N_5637,N_4719,N_4304);
xnor U5638 (N_5638,N_4875,N_4575);
nor U5639 (N_5639,N_4394,N_4566);
xor U5640 (N_5640,N_4991,N_4167);
xnor U5641 (N_5641,N_4075,N_4885);
or U5642 (N_5642,N_4141,N_4755);
nor U5643 (N_5643,N_4280,N_4504);
xnor U5644 (N_5644,N_4410,N_4181);
nor U5645 (N_5645,N_4352,N_4059);
nor U5646 (N_5646,N_4863,N_4749);
or U5647 (N_5647,N_4427,N_4846);
and U5648 (N_5648,N_4421,N_4043);
and U5649 (N_5649,N_4543,N_4567);
nor U5650 (N_5650,N_4633,N_4155);
and U5651 (N_5651,N_4123,N_4558);
nand U5652 (N_5652,N_4691,N_4832);
xor U5653 (N_5653,N_4778,N_4255);
or U5654 (N_5654,N_4375,N_4755);
and U5655 (N_5655,N_4033,N_4194);
or U5656 (N_5656,N_4133,N_4959);
nand U5657 (N_5657,N_4074,N_4910);
or U5658 (N_5658,N_4128,N_4652);
and U5659 (N_5659,N_4364,N_4237);
nand U5660 (N_5660,N_4954,N_4867);
or U5661 (N_5661,N_4567,N_4688);
and U5662 (N_5662,N_4674,N_4811);
nor U5663 (N_5663,N_4690,N_4794);
or U5664 (N_5664,N_4808,N_4366);
or U5665 (N_5665,N_4746,N_4705);
and U5666 (N_5666,N_4745,N_4726);
xor U5667 (N_5667,N_4569,N_4431);
or U5668 (N_5668,N_4136,N_4953);
nor U5669 (N_5669,N_4815,N_4054);
and U5670 (N_5670,N_4652,N_4593);
xnor U5671 (N_5671,N_4929,N_4617);
or U5672 (N_5672,N_4541,N_4420);
and U5673 (N_5673,N_4775,N_4976);
nor U5674 (N_5674,N_4320,N_4461);
nand U5675 (N_5675,N_4908,N_4331);
nor U5676 (N_5676,N_4074,N_4043);
or U5677 (N_5677,N_4231,N_4740);
or U5678 (N_5678,N_4790,N_4960);
and U5679 (N_5679,N_4300,N_4354);
and U5680 (N_5680,N_4172,N_4659);
or U5681 (N_5681,N_4204,N_4484);
xor U5682 (N_5682,N_4233,N_4540);
nand U5683 (N_5683,N_4137,N_4519);
and U5684 (N_5684,N_4445,N_4090);
nor U5685 (N_5685,N_4278,N_4157);
and U5686 (N_5686,N_4994,N_4623);
nor U5687 (N_5687,N_4663,N_4463);
nand U5688 (N_5688,N_4118,N_4776);
xnor U5689 (N_5689,N_4537,N_4783);
nor U5690 (N_5690,N_4004,N_4492);
or U5691 (N_5691,N_4904,N_4088);
or U5692 (N_5692,N_4827,N_4651);
or U5693 (N_5693,N_4386,N_4823);
nand U5694 (N_5694,N_4392,N_4962);
xor U5695 (N_5695,N_4232,N_4138);
or U5696 (N_5696,N_4051,N_4009);
nand U5697 (N_5697,N_4766,N_4188);
nand U5698 (N_5698,N_4849,N_4755);
nor U5699 (N_5699,N_4718,N_4275);
or U5700 (N_5700,N_4402,N_4850);
xor U5701 (N_5701,N_4055,N_4475);
nand U5702 (N_5702,N_4572,N_4433);
nor U5703 (N_5703,N_4877,N_4124);
and U5704 (N_5704,N_4576,N_4182);
and U5705 (N_5705,N_4605,N_4062);
nand U5706 (N_5706,N_4572,N_4420);
and U5707 (N_5707,N_4885,N_4892);
and U5708 (N_5708,N_4261,N_4098);
xor U5709 (N_5709,N_4707,N_4767);
xnor U5710 (N_5710,N_4135,N_4401);
xor U5711 (N_5711,N_4933,N_4312);
and U5712 (N_5712,N_4884,N_4972);
xor U5713 (N_5713,N_4790,N_4413);
xor U5714 (N_5714,N_4534,N_4694);
nand U5715 (N_5715,N_4337,N_4658);
nand U5716 (N_5716,N_4582,N_4320);
nand U5717 (N_5717,N_4498,N_4429);
and U5718 (N_5718,N_4545,N_4515);
nor U5719 (N_5719,N_4014,N_4672);
xnor U5720 (N_5720,N_4616,N_4938);
xor U5721 (N_5721,N_4033,N_4283);
nor U5722 (N_5722,N_4067,N_4684);
nor U5723 (N_5723,N_4219,N_4547);
nor U5724 (N_5724,N_4162,N_4151);
or U5725 (N_5725,N_4808,N_4851);
nand U5726 (N_5726,N_4617,N_4958);
or U5727 (N_5727,N_4391,N_4288);
xnor U5728 (N_5728,N_4421,N_4028);
nand U5729 (N_5729,N_4980,N_4677);
or U5730 (N_5730,N_4277,N_4335);
xnor U5731 (N_5731,N_4018,N_4436);
nor U5732 (N_5732,N_4798,N_4970);
or U5733 (N_5733,N_4619,N_4078);
or U5734 (N_5734,N_4474,N_4215);
nor U5735 (N_5735,N_4616,N_4284);
nor U5736 (N_5736,N_4595,N_4573);
or U5737 (N_5737,N_4602,N_4751);
nand U5738 (N_5738,N_4654,N_4397);
xnor U5739 (N_5739,N_4953,N_4137);
nand U5740 (N_5740,N_4605,N_4307);
and U5741 (N_5741,N_4121,N_4246);
and U5742 (N_5742,N_4391,N_4959);
and U5743 (N_5743,N_4952,N_4163);
and U5744 (N_5744,N_4119,N_4517);
nor U5745 (N_5745,N_4530,N_4019);
xor U5746 (N_5746,N_4080,N_4152);
or U5747 (N_5747,N_4639,N_4570);
and U5748 (N_5748,N_4951,N_4078);
or U5749 (N_5749,N_4284,N_4086);
nor U5750 (N_5750,N_4158,N_4595);
nand U5751 (N_5751,N_4570,N_4488);
xnor U5752 (N_5752,N_4357,N_4188);
nand U5753 (N_5753,N_4045,N_4888);
and U5754 (N_5754,N_4338,N_4702);
xor U5755 (N_5755,N_4926,N_4684);
nand U5756 (N_5756,N_4895,N_4029);
or U5757 (N_5757,N_4637,N_4303);
xor U5758 (N_5758,N_4268,N_4805);
and U5759 (N_5759,N_4322,N_4225);
xnor U5760 (N_5760,N_4855,N_4447);
and U5761 (N_5761,N_4223,N_4863);
or U5762 (N_5762,N_4397,N_4006);
nor U5763 (N_5763,N_4325,N_4345);
and U5764 (N_5764,N_4503,N_4527);
nand U5765 (N_5765,N_4908,N_4165);
nor U5766 (N_5766,N_4299,N_4255);
nand U5767 (N_5767,N_4015,N_4827);
and U5768 (N_5768,N_4963,N_4672);
or U5769 (N_5769,N_4179,N_4945);
nor U5770 (N_5770,N_4064,N_4407);
nor U5771 (N_5771,N_4238,N_4151);
or U5772 (N_5772,N_4376,N_4107);
and U5773 (N_5773,N_4644,N_4901);
and U5774 (N_5774,N_4968,N_4888);
or U5775 (N_5775,N_4489,N_4974);
nand U5776 (N_5776,N_4986,N_4526);
or U5777 (N_5777,N_4546,N_4660);
xnor U5778 (N_5778,N_4241,N_4402);
nand U5779 (N_5779,N_4146,N_4658);
nor U5780 (N_5780,N_4478,N_4160);
nor U5781 (N_5781,N_4392,N_4482);
nand U5782 (N_5782,N_4446,N_4847);
or U5783 (N_5783,N_4162,N_4318);
or U5784 (N_5784,N_4366,N_4005);
nand U5785 (N_5785,N_4181,N_4852);
or U5786 (N_5786,N_4430,N_4045);
xor U5787 (N_5787,N_4475,N_4385);
or U5788 (N_5788,N_4277,N_4877);
nor U5789 (N_5789,N_4388,N_4347);
and U5790 (N_5790,N_4982,N_4191);
and U5791 (N_5791,N_4415,N_4826);
nand U5792 (N_5792,N_4820,N_4858);
nand U5793 (N_5793,N_4087,N_4066);
xor U5794 (N_5794,N_4913,N_4072);
or U5795 (N_5795,N_4667,N_4369);
nand U5796 (N_5796,N_4639,N_4579);
nand U5797 (N_5797,N_4303,N_4961);
xor U5798 (N_5798,N_4748,N_4918);
and U5799 (N_5799,N_4554,N_4813);
xnor U5800 (N_5800,N_4791,N_4908);
and U5801 (N_5801,N_4853,N_4064);
xor U5802 (N_5802,N_4152,N_4772);
and U5803 (N_5803,N_4951,N_4568);
xor U5804 (N_5804,N_4465,N_4368);
nor U5805 (N_5805,N_4484,N_4029);
nor U5806 (N_5806,N_4809,N_4617);
and U5807 (N_5807,N_4290,N_4725);
nor U5808 (N_5808,N_4205,N_4795);
nor U5809 (N_5809,N_4563,N_4851);
or U5810 (N_5810,N_4611,N_4858);
nor U5811 (N_5811,N_4961,N_4392);
or U5812 (N_5812,N_4052,N_4617);
or U5813 (N_5813,N_4840,N_4376);
nor U5814 (N_5814,N_4068,N_4118);
or U5815 (N_5815,N_4895,N_4458);
nor U5816 (N_5816,N_4511,N_4475);
or U5817 (N_5817,N_4002,N_4467);
xor U5818 (N_5818,N_4574,N_4609);
xnor U5819 (N_5819,N_4379,N_4060);
nor U5820 (N_5820,N_4234,N_4468);
or U5821 (N_5821,N_4907,N_4479);
nand U5822 (N_5822,N_4447,N_4554);
and U5823 (N_5823,N_4583,N_4604);
or U5824 (N_5824,N_4851,N_4004);
and U5825 (N_5825,N_4676,N_4210);
nor U5826 (N_5826,N_4997,N_4671);
nor U5827 (N_5827,N_4523,N_4793);
nor U5828 (N_5828,N_4714,N_4855);
nor U5829 (N_5829,N_4975,N_4265);
nor U5830 (N_5830,N_4591,N_4249);
nand U5831 (N_5831,N_4740,N_4010);
or U5832 (N_5832,N_4858,N_4793);
and U5833 (N_5833,N_4498,N_4882);
or U5834 (N_5834,N_4140,N_4470);
and U5835 (N_5835,N_4735,N_4746);
and U5836 (N_5836,N_4446,N_4705);
nor U5837 (N_5837,N_4447,N_4596);
and U5838 (N_5838,N_4909,N_4627);
xnor U5839 (N_5839,N_4231,N_4805);
nor U5840 (N_5840,N_4453,N_4964);
and U5841 (N_5841,N_4418,N_4412);
xnor U5842 (N_5842,N_4104,N_4423);
or U5843 (N_5843,N_4309,N_4293);
nand U5844 (N_5844,N_4423,N_4649);
nor U5845 (N_5845,N_4499,N_4944);
nor U5846 (N_5846,N_4944,N_4346);
or U5847 (N_5847,N_4793,N_4047);
and U5848 (N_5848,N_4395,N_4812);
nor U5849 (N_5849,N_4492,N_4129);
or U5850 (N_5850,N_4419,N_4137);
xnor U5851 (N_5851,N_4271,N_4135);
and U5852 (N_5852,N_4059,N_4639);
nor U5853 (N_5853,N_4394,N_4924);
or U5854 (N_5854,N_4605,N_4970);
and U5855 (N_5855,N_4852,N_4856);
nor U5856 (N_5856,N_4135,N_4033);
or U5857 (N_5857,N_4451,N_4834);
or U5858 (N_5858,N_4380,N_4351);
or U5859 (N_5859,N_4077,N_4231);
nand U5860 (N_5860,N_4273,N_4255);
nand U5861 (N_5861,N_4485,N_4245);
and U5862 (N_5862,N_4930,N_4542);
or U5863 (N_5863,N_4770,N_4022);
or U5864 (N_5864,N_4437,N_4904);
xor U5865 (N_5865,N_4720,N_4483);
xnor U5866 (N_5866,N_4424,N_4476);
and U5867 (N_5867,N_4350,N_4742);
and U5868 (N_5868,N_4533,N_4512);
xor U5869 (N_5869,N_4113,N_4752);
nor U5870 (N_5870,N_4359,N_4531);
or U5871 (N_5871,N_4481,N_4204);
nand U5872 (N_5872,N_4910,N_4085);
and U5873 (N_5873,N_4154,N_4891);
and U5874 (N_5874,N_4604,N_4828);
or U5875 (N_5875,N_4563,N_4465);
nor U5876 (N_5876,N_4337,N_4511);
and U5877 (N_5877,N_4961,N_4122);
or U5878 (N_5878,N_4898,N_4601);
nor U5879 (N_5879,N_4074,N_4808);
or U5880 (N_5880,N_4100,N_4838);
nor U5881 (N_5881,N_4265,N_4267);
xor U5882 (N_5882,N_4522,N_4583);
xor U5883 (N_5883,N_4368,N_4703);
xnor U5884 (N_5884,N_4928,N_4722);
or U5885 (N_5885,N_4362,N_4971);
xor U5886 (N_5886,N_4509,N_4269);
or U5887 (N_5887,N_4678,N_4798);
nand U5888 (N_5888,N_4724,N_4071);
nor U5889 (N_5889,N_4824,N_4278);
or U5890 (N_5890,N_4750,N_4937);
xor U5891 (N_5891,N_4659,N_4917);
and U5892 (N_5892,N_4087,N_4417);
or U5893 (N_5893,N_4335,N_4104);
nand U5894 (N_5894,N_4441,N_4748);
xnor U5895 (N_5895,N_4428,N_4139);
nor U5896 (N_5896,N_4124,N_4001);
xor U5897 (N_5897,N_4355,N_4872);
nand U5898 (N_5898,N_4301,N_4669);
and U5899 (N_5899,N_4696,N_4472);
nor U5900 (N_5900,N_4362,N_4725);
nor U5901 (N_5901,N_4786,N_4267);
nand U5902 (N_5902,N_4854,N_4542);
nand U5903 (N_5903,N_4357,N_4960);
nor U5904 (N_5904,N_4641,N_4834);
and U5905 (N_5905,N_4690,N_4985);
or U5906 (N_5906,N_4051,N_4124);
xnor U5907 (N_5907,N_4399,N_4558);
and U5908 (N_5908,N_4257,N_4649);
nand U5909 (N_5909,N_4345,N_4878);
xnor U5910 (N_5910,N_4749,N_4207);
or U5911 (N_5911,N_4434,N_4715);
or U5912 (N_5912,N_4444,N_4876);
nor U5913 (N_5913,N_4609,N_4133);
nor U5914 (N_5914,N_4756,N_4052);
nand U5915 (N_5915,N_4544,N_4773);
xor U5916 (N_5916,N_4451,N_4511);
nand U5917 (N_5917,N_4740,N_4957);
xor U5918 (N_5918,N_4024,N_4068);
or U5919 (N_5919,N_4673,N_4935);
nand U5920 (N_5920,N_4967,N_4604);
xnor U5921 (N_5921,N_4302,N_4848);
or U5922 (N_5922,N_4453,N_4544);
xnor U5923 (N_5923,N_4336,N_4484);
xnor U5924 (N_5924,N_4781,N_4650);
xor U5925 (N_5925,N_4976,N_4115);
and U5926 (N_5926,N_4209,N_4299);
or U5927 (N_5927,N_4801,N_4719);
or U5928 (N_5928,N_4078,N_4387);
nand U5929 (N_5929,N_4656,N_4949);
xnor U5930 (N_5930,N_4000,N_4892);
nand U5931 (N_5931,N_4111,N_4665);
or U5932 (N_5932,N_4554,N_4089);
nor U5933 (N_5933,N_4927,N_4631);
nor U5934 (N_5934,N_4039,N_4007);
nor U5935 (N_5935,N_4074,N_4280);
nand U5936 (N_5936,N_4470,N_4734);
or U5937 (N_5937,N_4819,N_4935);
xor U5938 (N_5938,N_4454,N_4035);
or U5939 (N_5939,N_4154,N_4778);
and U5940 (N_5940,N_4081,N_4781);
and U5941 (N_5941,N_4338,N_4808);
xnor U5942 (N_5942,N_4840,N_4922);
or U5943 (N_5943,N_4239,N_4722);
nor U5944 (N_5944,N_4147,N_4586);
or U5945 (N_5945,N_4742,N_4900);
nand U5946 (N_5946,N_4732,N_4222);
or U5947 (N_5947,N_4325,N_4767);
xnor U5948 (N_5948,N_4764,N_4183);
nand U5949 (N_5949,N_4005,N_4526);
xnor U5950 (N_5950,N_4891,N_4217);
or U5951 (N_5951,N_4597,N_4803);
nand U5952 (N_5952,N_4088,N_4282);
and U5953 (N_5953,N_4073,N_4852);
and U5954 (N_5954,N_4267,N_4568);
nor U5955 (N_5955,N_4998,N_4911);
and U5956 (N_5956,N_4566,N_4547);
or U5957 (N_5957,N_4676,N_4773);
xnor U5958 (N_5958,N_4210,N_4489);
or U5959 (N_5959,N_4217,N_4545);
or U5960 (N_5960,N_4937,N_4354);
or U5961 (N_5961,N_4705,N_4841);
or U5962 (N_5962,N_4461,N_4954);
xor U5963 (N_5963,N_4913,N_4992);
and U5964 (N_5964,N_4297,N_4648);
or U5965 (N_5965,N_4141,N_4749);
and U5966 (N_5966,N_4160,N_4960);
and U5967 (N_5967,N_4844,N_4299);
and U5968 (N_5968,N_4520,N_4935);
or U5969 (N_5969,N_4596,N_4282);
and U5970 (N_5970,N_4445,N_4183);
or U5971 (N_5971,N_4720,N_4105);
or U5972 (N_5972,N_4428,N_4571);
xor U5973 (N_5973,N_4752,N_4670);
or U5974 (N_5974,N_4182,N_4116);
and U5975 (N_5975,N_4971,N_4127);
and U5976 (N_5976,N_4850,N_4148);
or U5977 (N_5977,N_4368,N_4569);
or U5978 (N_5978,N_4966,N_4508);
nand U5979 (N_5979,N_4348,N_4128);
nand U5980 (N_5980,N_4545,N_4423);
nand U5981 (N_5981,N_4541,N_4423);
nand U5982 (N_5982,N_4987,N_4594);
nor U5983 (N_5983,N_4168,N_4393);
or U5984 (N_5984,N_4386,N_4396);
and U5985 (N_5985,N_4290,N_4909);
nor U5986 (N_5986,N_4617,N_4717);
xor U5987 (N_5987,N_4458,N_4910);
xor U5988 (N_5988,N_4538,N_4087);
and U5989 (N_5989,N_4766,N_4930);
and U5990 (N_5990,N_4284,N_4264);
xnor U5991 (N_5991,N_4481,N_4140);
or U5992 (N_5992,N_4334,N_4017);
or U5993 (N_5993,N_4131,N_4622);
xnor U5994 (N_5994,N_4132,N_4867);
xnor U5995 (N_5995,N_4673,N_4347);
or U5996 (N_5996,N_4140,N_4702);
and U5997 (N_5997,N_4052,N_4351);
nand U5998 (N_5998,N_4376,N_4116);
nor U5999 (N_5999,N_4064,N_4475);
or U6000 (N_6000,N_5633,N_5644);
or U6001 (N_6001,N_5865,N_5520);
and U6002 (N_6002,N_5033,N_5091);
and U6003 (N_6003,N_5157,N_5888);
nor U6004 (N_6004,N_5073,N_5743);
nor U6005 (N_6005,N_5626,N_5204);
xnor U6006 (N_6006,N_5110,N_5989);
xnor U6007 (N_6007,N_5828,N_5405);
xnor U6008 (N_6008,N_5312,N_5031);
or U6009 (N_6009,N_5314,N_5666);
xor U6010 (N_6010,N_5253,N_5317);
and U6011 (N_6011,N_5416,N_5257);
xnor U6012 (N_6012,N_5239,N_5118);
and U6013 (N_6013,N_5237,N_5207);
or U6014 (N_6014,N_5211,N_5776);
nor U6015 (N_6015,N_5128,N_5191);
xnor U6016 (N_6016,N_5680,N_5150);
or U6017 (N_6017,N_5451,N_5430);
nand U6018 (N_6018,N_5299,N_5899);
nand U6019 (N_6019,N_5948,N_5876);
or U6020 (N_6020,N_5562,N_5189);
nor U6021 (N_6021,N_5295,N_5821);
xnor U6022 (N_6022,N_5533,N_5918);
nor U6023 (N_6023,N_5111,N_5124);
nand U6024 (N_6024,N_5668,N_5774);
nand U6025 (N_6025,N_5878,N_5014);
and U6026 (N_6026,N_5673,N_5027);
and U6027 (N_6027,N_5275,N_5045);
nor U6028 (N_6028,N_5561,N_5137);
and U6029 (N_6029,N_5374,N_5907);
nand U6030 (N_6030,N_5398,N_5245);
or U6031 (N_6031,N_5811,N_5539);
and U6032 (N_6032,N_5302,N_5143);
xor U6033 (N_6033,N_5351,N_5505);
xor U6034 (N_6034,N_5601,N_5671);
nor U6035 (N_6035,N_5754,N_5762);
nand U6036 (N_6036,N_5264,N_5493);
or U6037 (N_6037,N_5917,N_5650);
and U6038 (N_6038,N_5305,N_5779);
nor U6039 (N_6039,N_5632,N_5690);
or U6040 (N_6040,N_5285,N_5165);
or U6041 (N_6041,N_5062,N_5311);
nand U6042 (N_6042,N_5660,N_5838);
xor U6043 (N_6043,N_5350,N_5467);
xor U6044 (N_6044,N_5476,N_5063);
nand U6045 (N_6045,N_5766,N_5689);
xor U6046 (N_6046,N_5373,N_5786);
or U6047 (N_6047,N_5144,N_5688);
nor U6048 (N_6048,N_5745,N_5997);
nand U6049 (N_6049,N_5117,N_5551);
xnor U6050 (N_6050,N_5453,N_5640);
and U6051 (N_6051,N_5654,N_5103);
and U6052 (N_6052,N_5885,N_5622);
and U6053 (N_6053,N_5837,N_5956);
nor U6054 (N_6054,N_5010,N_5566);
nor U6055 (N_6055,N_5557,N_5658);
nand U6056 (N_6056,N_5517,N_5353);
nand U6057 (N_6057,N_5209,N_5290);
xor U6058 (N_6058,N_5126,N_5094);
or U6059 (N_6059,N_5200,N_5707);
nand U6060 (N_6060,N_5906,N_5621);
or U6061 (N_6061,N_5852,N_5602);
or U6062 (N_6062,N_5716,N_5574);
xnor U6063 (N_6063,N_5459,N_5213);
nand U6064 (N_6064,N_5729,N_5313);
or U6065 (N_6065,N_5278,N_5210);
xnor U6066 (N_6066,N_5342,N_5968);
nor U6067 (N_6067,N_5423,N_5923);
or U6068 (N_6068,N_5482,N_5404);
nor U6069 (N_6069,N_5634,N_5586);
or U6070 (N_6070,N_5319,N_5643);
nor U6071 (N_6071,N_5901,N_5758);
and U6072 (N_6072,N_5347,N_5530);
xnor U6073 (N_6073,N_5034,N_5733);
and U6074 (N_6074,N_5617,N_5366);
xnor U6075 (N_6075,N_5734,N_5882);
nand U6076 (N_6076,N_5233,N_5147);
nor U6077 (N_6077,N_5406,N_5387);
and U6078 (N_6078,N_5502,N_5479);
or U6079 (N_6079,N_5529,N_5006);
nor U6080 (N_6080,N_5785,N_5352);
or U6081 (N_6081,N_5655,N_5125);
nor U6082 (N_6082,N_5470,N_5746);
xor U6083 (N_6083,N_5097,N_5691);
and U6084 (N_6084,N_5518,N_5021);
xor U6085 (N_6085,N_5605,N_5616);
nor U6086 (N_6086,N_5506,N_5166);
and U6087 (N_6087,N_5267,N_5874);
xor U6088 (N_6088,N_5120,N_5130);
nor U6089 (N_6089,N_5362,N_5846);
and U6090 (N_6090,N_5234,N_5383);
nor U6091 (N_6091,N_5256,N_5826);
or U6092 (N_6092,N_5399,N_5265);
nand U6093 (N_6093,N_5364,N_5273);
or U6094 (N_6094,N_5104,N_5061);
xnor U6095 (N_6095,N_5855,N_5148);
nor U6096 (N_6096,N_5296,N_5015);
nand U6097 (N_6097,N_5523,N_5613);
nor U6098 (N_6098,N_5735,N_5537);
xnor U6099 (N_6099,N_5294,N_5829);
xnor U6100 (N_6100,N_5197,N_5077);
and U6101 (N_6101,N_5456,N_5939);
nand U6102 (N_6102,N_5369,N_5844);
or U6103 (N_6103,N_5386,N_5370);
nor U6104 (N_6104,N_5095,N_5921);
or U6105 (N_6105,N_5608,N_5193);
xor U6106 (N_6106,N_5343,N_5934);
nand U6107 (N_6107,N_5935,N_5814);
xnor U6108 (N_6108,N_5646,N_5395);
nor U6109 (N_6109,N_5615,N_5426);
xor U6110 (N_6110,N_5949,N_5903);
and U6111 (N_6111,N_5259,N_5116);
and U6112 (N_6112,N_5262,N_5998);
and U6113 (N_6113,N_5135,N_5411);
or U6114 (N_6114,N_5202,N_5208);
xnor U6115 (N_6115,N_5757,N_5065);
nor U6116 (N_6116,N_5696,N_5565);
nand U6117 (N_6117,N_5967,N_5744);
and U6118 (N_6118,N_5315,N_5136);
and U6119 (N_6119,N_5127,N_5833);
or U6120 (N_6120,N_5986,N_5215);
nand U6121 (N_6121,N_5944,N_5895);
and U6122 (N_6122,N_5408,N_5188);
nand U6123 (N_6123,N_5832,N_5869);
nor U6124 (N_6124,N_5236,N_5752);
nand U6125 (N_6125,N_5330,N_5979);
nor U6126 (N_6126,N_5164,N_5526);
xnor U6127 (N_6127,N_5581,N_5898);
nand U6128 (N_6128,N_5019,N_5791);
nor U6129 (N_6129,N_5804,N_5066);
or U6130 (N_6130,N_5636,N_5618);
or U6131 (N_6131,N_5198,N_5926);
or U6132 (N_6132,N_5071,N_5086);
nor U6133 (N_6133,N_5925,N_5805);
or U6134 (N_6134,N_5108,N_5464);
nor U6135 (N_6135,N_5985,N_5790);
xnor U6136 (N_6136,N_5683,N_5401);
nor U6137 (N_6137,N_5721,N_5775);
xnor U6138 (N_6138,N_5331,N_5220);
nor U6139 (N_6139,N_5971,N_5235);
and U6140 (N_6140,N_5559,N_5810);
xor U6141 (N_6141,N_5079,N_5175);
xnor U6142 (N_6142,N_5339,N_5276);
nand U6143 (N_6143,N_5549,N_5185);
and U6144 (N_6144,N_5932,N_5981);
nand U6145 (N_6145,N_5830,N_5485);
and U6146 (N_6146,N_5146,N_5912);
nand U6147 (N_6147,N_5571,N_5902);
and U6148 (N_6148,N_5114,N_5623);
or U6149 (N_6149,N_5867,N_5280);
and U6150 (N_6150,N_5454,N_5794);
or U6151 (N_6151,N_5609,N_5109);
nor U6152 (N_6152,N_5064,N_5717);
nor U6153 (N_6153,N_5772,N_5291);
or U6154 (N_6154,N_5349,N_5229);
nor U6155 (N_6155,N_5227,N_5977);
nor U6156 (N_6156,N_5797,N_5345);
xnor U6157 (N_6157,N_5060,N_5699);
nand U6158 (N_6158,N_5324,N_5011);
xnor U6159 (N_6159,N_5528,N_5879);
nand U6160 (N_6160,N_5684,N_5871);
and U6161 (N_6161,N_5667,N_5022);
xor U6162 (N_6162,N_5041,N_5793);
xnor U6163 (N_6163,N_5008,N_5085);
or U6164 (N_6164,N_5192,N_5444);
xnor U6165 (N_6165,N_5473,N_5681);
or U6166 (N_6166,N_5067,N_5242);
or U6167 (N_6167,N_5412,N_5069);
or U6168 (N_6168,N_5788,N_5142);
nand U6169 (N_6169,N_5983,N_5051);
nand U6170 (N_6170,N_5122,N_5099);
and U6171 (N_6171,N_5897,N_5807);
and U6172 (N_6172,N_5836,N_5354);
and U6173 (N_6173,N_5297,N_5980);
xor U6174 (N_6174,N_5472,N_5230);
nor U6175 (N_6175,N_5449,N_5372);
or U6176 (N_6176,N_5709,N_5875);
or U6177 (N_6177,N_5536,N_5145);
and U6178 (N_6178,N_5138,N_5205);
nor U6179 (N_6179,N_5945,N_5823);
and U6180 (N_6180,N_5947,N_5271);
and U6181 (N_6181,N_5820,N_5252);
nor U6182 (N_6182,N_5162,N_5083);
nor U6183 (N_6183,N_5808,N_5216);
or U6184 (N_6184,N_5403,N_5089);
xnor U6185 (N_6185,N_5740,N_5892);
nand U6186 (N_6186,N_5381,N_5139);
nor U6187 (N_6187,N_5627,N_5570);
nand U6188 (N_6188,N_5475,N_5219);
nor U6189 (N_6189,N_5163,N_5554);
and U6190 (N_6190,N_5186,N_5973);
xnor U6191 (N_6191,N_5555,N_5507);
xnor U6192 (N_6192,N_5853,N_5665);
nor U6193 (N_6193,N_5864,N_5910);
or U6194 (N_6194,N_5760,N_5751);
or U6195 (N_6195,N_5240,N_5129);
nor U6196 (N_6196,N_5556,N_5438);
nor U6197 (N_6197,N_5904,N_5327);
nand U6198 (N_6198,N_5346,N_5038);
xnor U6199 (N_6199,N_5877,N_5883);
and U6200 (N_6200,N_5248,N_5440);
or U6201 (N_6201,N_5418,N_5052);
nand U6202 (N_6202,N_5577,N_5687);
or U6203 (N_6203,N_5427,N_5677);
nor U6204 (N_6204,N_5742,N_5042);
xnor U6205 (N_6205,N_5669,N_5462);
xnor U6206 (N_6206,N_5471,N_5706);
or U6207 (N_6207,N_5787,N_5357);
and U6208 (N_6208,N_5950,N_5579);
or U6209 (N_6209,N_5886,N_5084);
or U6210 (N_6210,N_5784,N_5318);
or U6211 (N_6211,N_5310,N_5203);
and U6212 (N_6212,N_5516,N_5726);
nor U6213 (N_6213,N_5670,N_5196);
nor U6214 (N_6214,N_5035,N_5806);
nor U6215 (N_6215,N_5963,N_5379);
xnor U6216 (N_6216,N_5719,N_5504);
xor U6217 (N_6217,N_5737,N_5780);
xnor U6218 (N_6218,N_5802,N_5488);
and U6219 (N_6219,N_5777,N_5951);
or U6220 (N_6220,N_5873,N_5771);
and U6221 (N_6221,N_5238,N_5954);
nor U6222 (N_6222,N_5004,N_5450);
nor U6223 (N_6223,N_5619,N_5016);
xnor U6224 (N_6224,N_5891,N_5141);
and U6225 (N_6225,N_5739,N_5704);
nor U6226 (N_6226,N_5422,N_5512);
xor U6227 (N_6227,N_5323,N_5563);
nor U6228 (N_6228,N_5712,N_5160);
xnor U6229 (N_6229,N_5039,N_5705);
xor U6230 (N_6230,N_5380,N_5113);
nor U6231 (N_6231,N_5999,N_5585);
nand U6232 (N_6232,N_5708,N_5856);
nor U6233 (N_6233,N_5552,N_5753);
nand U6234 (N_6234,N_5348,N_5458);
and U6235 (N_6235,N_5550,N_5920);
nor U6236 (N_6236,N_5172,N_5840);
and U6237 (N_6237,N_5631,N_5007);
and U6238 (N_6238,N_5417,N_5761);
and U6239 (N_6239,N_5937,N_5952);
nor U6240 (N_6240,N_5941,N_5635);
nor U6241 (N_6241,N_5942,N_5976);
and U6242 (N_6242,N_5121,N_5657);
nand U6243 (N_6243,N_5268,N_5419);
and U6244 (N_6244,N_5431,N_5272);
nand U6245 (N_6245,N_5604,N_5720);
and U6246 (N_6246,N_5896,N_5599);
nor U6247 (N_6247,N_5298,N_5152);
nor U6248 (N_6248,N_5088,N_5541);
xor U6249 (N_6249,N_5663,N_5994);
xor U6250 (N_6250,N_5629,N_5843);
and U6251 (N_6251,N_5970,N_5445);
nand U6252 (N_6252,N_5914,N_5106);
xor U6253 (N_6253,N_5773,N_5591);
xnor U6254 (N_6254,N_5569,N_5491);
nor U6255 (N_6255,N_5965,N_5567);
xor U6256 (N_6256,N_5410,N_5212);
and U6257 (N_6257,N_5222,N_5492);
and U6258 (N_6258,N_5661,N_5819);
nand U6259 (N_6259,N_5960,N_5560);
or U6260 (N_6260,N_5589,N_5490);
nor U6261 (N_6261,N_5281,N_5076);
and U6262 (N_6262,N_5070,N_5538);
and U6263 (N_6263,N_5170,N_5218);
xor U6264 (N_6264,N_5649,N_5659);
xnor U6265 (N_6265,N_5044,N_5258);
nor U6266 (N_6266,N_5055,N_5483);
nand U6267 (N_6267,N_5795,N_5713);
nor U6268 (N_6268,N_5698,N_5815);
nand U6269 (N_6269,N_5260,N_5159);
xor U6270 (N_6270,N_5090,N_5024);
nor U6271 (N_6271,N_5301,N_5226);
and U6272 (N_6272,N_5940,N_5769);
nor U6273 (N_6273,N_5176,N_5749);
nor U6274 (N_6274,N_5862,N_5368);
nand U6275 (N_6275,N_5582,N_5587);
nor U6276 (N_6276,N_5376,N_5755);
or U6277 (N_6277,N_5005,N_5724);
nor U6278 (N_6278,N_5511,N_5723);
and U6279 (N_6279,N_5767,N_5792);
xor U6280 (N_6280,N_5286,N_5214);
or U6281 (N_6281,N_5887,N_5283);
and U6282 (N_6282,N_5964,N_5221);
nand U6283 (N_6283,N_5382,N_5307);
nor U6284 (N_6284,N_5012,N_5182);
nand U6285 (N_6285,N_5481,N_5452);
and U6286 (N_6286,N_5715,N_5328);
nor U6287 (N_6287,N_5572,N_5857);
and U6288 (N_6288,N_5580,N_5595);
nand U6289 (N_6289,N_5390,N_5881);
or U6290 (N_6290,N_5420,N_5187);
xor U6291 (N_6291,N_5375,N_5993);
nor U6292 (N_6292,N_5763,N_5421);
nor U6293 (N_6293,N_5335,N_5756);
nand U6294 (N_6294,N_5023,N_5527);
or U6295 (N_6295,N_5255,N_5000);
xnor U6296 (N_6296,N_5289,N_5924);
xor U6297 (N_6297,N_5782,N_5020);
or U6298 (N_6298,N_5468,N_5812);
or U6299 (N_6299,N_5075,N_5149);
or U6300 (N_6300,N_5266,N_5850);
nor U6301 (N_6301,N_5072,N_5013);
nand U6302 (N_6302,N_5741,N_5603);
nand U6303 (N_6303,N_5831,N_5269);
or U6304 (N_6304,N_5645,N_5893);
nor U6305 (N_6305,N_5036,N_5890);
xor U6306 (N_6306,N_5499,N_5974);
and U6307 (N_6307,N_5540,N_5393);
nor U6308 (N_6308,N_5816,N_5694);
and U6309 (N_6309,N_5322,N_5057);
xnor U6310 (N_6310,N_5714,N_5478);
nand U6311 (N_6311,N_5053,N_5783);
nor U6312 (N_6312,N_5858,N_5101);
nand U6313 (N_6313,N_5630,N_5402);
and U6314 (N_6314,N_5930,N_5702);
and U6315 (N_6315,N_5725,N_5448);
xnor U6316 (N_6316,N_5461,N_5880);
nor U6317 (N_6317,N_5338,N_5839);
or U6318 (N_6318,N_5277,N_5849);
nand U6319 (N_6319,N_5542,N_5336);
or U6320 (N_6320,N_5710,N_5080);
and U6321 (N_6321,N_5524,N_5119);
and U6322 (N_6322,N_5279,N_5610);
xnor U6323 (N_6323,N_5025,N_5415);
nand U6324 (N_6324,N_5340,N_5534);
nand U6325 (N_6325,N_5432,N_5486);
or U6326 (N_6326,N_5732,N_5588);
and U6327 (N_6327,N_5384,N_5046);
nand U6328 (N_6328,N_5962,N_5394);
or U6329 (N_6329,N_5442,N_5261);
or U6330 (N_6330,N_5711,N_5446);
nor U6331 (N_6331,N_5274,N_5824);
and U6332 (N_6332,N_5600,N_5778);
xor U6333 (N_6333,N_5508,N_5341);
nand U6334 (N_6334,N_5465,N_5428);
xnor U6335 (N_6335,N_5597,N_5848);
or U6336 (N_6336,N_5624,N_5397);
nand U6337 (N_6337,N_5466,N_5391);
and U6338 (N_6338,N_5140,N_5407);
xor U6339 (N_6339,N_5672,N_5969);
or U6340 (N_6340,N_5984,N_5484);
nand U6341 (N_6341,N_5333,N_5593);
or U6342 (N_6342,N_5544,N_5747);
and U6343 (N_6343,N_5731,N_5360);
and U6344 (N_6344,N_5435,N_5463);
nand U6345 (N_6345,N_5953,N_5532);
nor U6346 (N_6346,N_5522,N_5361);
or U6347 (N_6347,N_5915,N_5800);
nor U6348 (N_6348,N_5596,N_5332);
or U6349 (N_6349,N_5992,N_5612);
and U6350 (N_6350,N_5987,N_5048);
nand U6351 (N_6351,N_5851,N_5329);
nor U6352 (N_6352,N_5058,N_5115);
or U6353 (N_6353,N_5292,N_5548);
and U6354 (N_6354,N_5497,N_5513);
or U6355 (N_6355,N_5909,N_5841);
and U6356 (N_6356,N_5798,N_5183);
nand U6357 (N_6357,N_5501,N_5558);
nand U6358 (N_6358,N_5938,N_5223);
and U6359 (N_6359,N_5047,N_5889);
nand U6360 (N_6360,N_5433,N_5913);
and U6361 (N_6361,N_5845,N_5653);
or U6362 (N_6362,N_5098,N_5325);
nor U6363 (N_6363,N_5096,N_5441);
or U6364 (N_6364,N_5133,N_5206);
xor U6365 (N_6365,N_5662,N_5575);
xnor U6366 (N_6366,N_5409,N_5378);
nor U6367 (N_6367,N_5817,N_5975);
xnor U6368 (N_6368,N_5727,N_5525);
nor U6369 (N_6369,N_5371,N_5972);
and U6370 (N_6370,N_5509,N_5982);
nor U6371 (N_6371,N_5181,N_5447);
or U6372 (N_6372,N_5676,N_5358);
xor U6373 (N_6373,N_5151,N_5102);
nor U6374 (N_6374,N_5781,N_5009);
nand U6375 (N_6375,N_5642,N_5990);
nor U6376 (N_6376,N_5573,N_5400);
and U6377 (N_6377,N_5225,N_5978);
xor U6378 (N_6378,N_5545,N_5764);
nand U6379 (N_6379,N_5576,N_5614);
nor U6380 (N_6380,N_5243,N_5620);
xnor U6381 (N_6381,N_5736,N_5693);
or U6382 (N_6382,N_5946,N_5543);
nand U6383 (N_6383,N_5270,N_5173);
nor U6384 (N_6384,N_5241,N_5232);
xor U6385 (N_6385,N_5639,N_5195);
or U6386 (N_6386,N_5303,N_5199);
nor U6387 (N_6387,N_5703,N_5487);
nor U6388 (N_6388,N_5510,N_5425);
and U6389 (N_6389,N_5933,N_5583);
or U6390 (N_6390,N_5796,N_5123);
nand U6391 (N_6391,N_5607,N_5474);
and U6392 (N_6392,N_5592,N_5469);
or U6393 (N_6393,N_5457,N_5413);
nor U6394 (N_6394,N_5789,N_5988);
nor U6395 (N_6395,N_5578,N_5553);
xnor U6396 (N_6396,N_5228,N_5078);
xor U6397 (N_6397,N_5872,N_5201);
nand U6398 (N_6398,N_5718,N_5911);
or U6399 (N_6399,N_5300,N_5799);
and U6400 (N_6400,N_5894,N_5955);
or U6401 (N_6401,N_5489,N_5167);
xnor U6402 (N_6402,N_5822,N_5682);
nor U6403 (N_6403,N_5641,N_5040);
and U6404 (N_6404,N_5590,N_5652);
nand U6405 (N_6405,N_5304,N_5584);
nand U6406 (N_6406,N_5958,N_5943);
or U6407 (N_6407,N_5246,N_5087);
or U6408 (N_6408,N_5648,N_5647);
nand U6409 (N_6409,N_5168,N_5870);
or U6410 (N_6410,N_5037,N_5498);
and U6411 (N_6411,N_5460,N_5931);
nor U6412 (N_6412,N_5177,N_5434);
and U6413 (N_6413,N_5344,N_5959);
nand U6414 (N_6414,N_5293,N_5367);
and U6415 (N_6415,N_5919,N_5834);
nand U6416 (N_6416,N_5770,N_5217);
xnor U6417 (N_6417,N_5813,N_5847);
nand U6418 (N_6418,N_5679,N_5363);
nand U6419 (N_6419,N_5685,N_5134);
or U6420 (N_6420,N_5564,N_5519);
nor U6421 (N_6421,N_5594,N_5026);
xor U6422 (N_6422,N_5863,N_5827);
xor U6423 (N_6423,N_5436,N_5675);
or U6424 (N_6424,N_5029,N_5309);
and U6425 (N_6425,N_5054,N_5455);
xnor U6426 (N_6426,N_5100,N_5697);
nand U6427 (N_6427,N_5477,N_5287);
nand U6428 (N_6428,N_5153,N_5598);
nand U6429 (N_6429,N_5759,N_5768);
xnor U6430 (N_6430,N_5611,N_5535);
nor U6431 (N_6431,N_5105,N_5927);
xnor U6432 (N_6432,N_5443,N_5859);
and U6433 (N_6433,N_5625,N_5835);
nand U6434 (N_6434,N_5818,N_5396);
or U6435 (N_6435,N_5437,N_5161);
or U6436 (N_6436,N_5651,N_5001);
nand U6437 (N_6437,N_5765,N_5178);
xor U6438 (N_6438,N_5308,N_5359);
or U6439 (N_6439,N_5628,N_5002);
or U6440 (N_6440,N_5154,N_5184);
nand U6441 (N_6441,N_5049,N_5606);
nand U6442 (N_6442,N_5179,N_5730);
or U6443 (N_6443,N_5503,N_5017);
or U6444 (N_6444,N_5320,N_5695);
and U6445 (N_6445,N_5132,N_5686);
xnor U6446 (N_6446,N_5250,N_5638);
nor U6447 (N_6447,N_5500,N_5355);
xor U6448 (N_6448,N_5018,N_5429);
nand U6449 (N_6449,N_5169,N_5356);
or U6450 (N_6450,N_5092,N_5546);
xor U6451 (N_6451,N_5748,N_5112);
nand U6452 (N_6452,N_5547,N_5326);
or U6453 (N_6453,N_5231,N_5905);
and U6454 (N_6454,N_5247,N_5496);
nor U6455 (N_6455,N_5388,N_5068);
nor U6456 (N_6456,N_5531,N_5809);
nor U6457 (N_6457,N_5568,N_5254);
nand U6458 (N_6458,N_5392,N_5996);
nand U6459 (N_6459,N_5263,N_5722);
xor U6460 (N_6460,N_5916,N_5656);
nor U6461 (N_6461,N_5059,N_5190);
xor U6462 (N_6462,N_5334,N_5043);
and U6463 (N_6463,N_5074,N_5174);
or U6464 (N_6464,N_5854,N_5728);
and U6465 (N_6465,N_5171,N_5900);
xnor U6466 (N_6466,N_5032,N_5093);
xor U6467 (N_6467,N_5082,N_5158);
nor U6468 (N_6468,N_5480,N_5389);
nand U6469 (N_6469,N_5155,N_5936);
and U6470 (N_6470,N_5107,N_5385);
or U6471 (N_6471,N_5929,N_5282);
xor U6472 (N_6472,N_5494,N_5028);
and U6473 (N_6473,N_5424,N_5249);
nor U6474 (N_6474,N_5316,N_5365);
and U6475 (N_6475,N_5514,N_5674);
and U6476 (N_6476,N_5180,N_5056);
nor U6477 (N_6477,N_5922,N_5801);
and U6478 (N_6478,N_5521,N_5884);
or U6479 (N_6479,N_5700,N_5081);
nand U6480 (N_6480,N_5803,N_5337);
nand U6481 (N_6481,N_5738,N_5991);
and U6482 (N_6482,N_5961,N_5957);
or U6483 (N_6483,N_5860,N_5678);
and U6484 (N_6484,N_5131,N_5495);
and U6485 (N_6485,N_5750,N_5637);
xnor U6486 (N_6486,N_5284,N_5244);
xnor U6487 (N_6487,N_5306,N_5321);
nand U6488 (N_6488,N_5030,N_5003);
and U6489 (N_6489,N_5825,N_5908);
xnor U6490 (N_6490,N_5515,N_5701);
or U6491 (N_6491,N_5866,N_5050);
nand U6492 (N_6492,N_5224,N_5439);
nor U6493 (N_6493,N_5928,N_5377);
or U6494 (N_6494,N_5156,N_5868);
xnor U6495 (N_6495,N_5194,N_5664);
nor U6496 (N_6496,N_5995,N_5966);
and U6497 (N_6497,N_5288,N_5861);
and U6498 (N_6498,N_5251,N_5842);
nand U6499 (N_6499,N_5692,N_5414);
xnor U6500 (N_6500,N_5847,N_5016);
or U6501 (N_6501,N_5777,N_5674);
xnor U6502 (N_6502,N_5512,N_5902);
nand U6503 (N_6503,N_5321,N_5421);
xor U6504 (N_6504,N_5707,N_5157);
or U6505 (N_6505,N_5770,N_5081);
and U6506 (N_6506,N_5863,N_5610);
and U6507 (N_6507,N_5369,N_5653);
nand U6508 (N_6508,N_5620,N_5455);
xor U6509 (N_6509,N_5033,N_5343);
or U6510 (N_6510,N_5050,N_5562);
xnor U6511 (N_6511,N_5122,N_5279);
or U6512 (N_6512,N_5418,N_5475);
nor U6513 (N_6513,N_5784,N_5885);
or U6514 (N_6514,N_5130,N_5036);
xor U6515 (N_6515,N_5841,N_5756);
nand U6516 (N_6516,N_5318,N_5638);
nor U6517 (N_6517,N_5450,N_5729);
nor U6518 (N_6518,N_5965,N_5041);
nor U6519 (N_6519,N_5654,N_5432);
or U6520 (N_6520,N_5875,N_5306);
nor U6521 (N_6521,N_5288,N_5533);
nand U6522 (N_6522,N_5056,N_5586);
nor U6523 (N_6523,N_5758,N_5217);
xor U6524 (N_6524,N_5526,N_5690);
or U6525 (N_6525,N_5684,N_5700);
xnor U6526 (N_6526,N_5930,N_5183);
nand U6527 (N_6527,N_5177,N_5585);
nor U6528 (N_6528,N_5372,N_5416);
or U6529 (N_6529,N_5705,N_5427);
xor U6530 (N_6530,N_5197,N_5464);
nand U6531 (N_6531,N_5279,N_5315);
or U6532 (N_6532,N_5620,N_5196);
nand U6533 (N_6533,N_5942,N_5477);
nor U6534 (N_6534,N_5220,N_5939);
and U6535 (N_6535,N_5484,N_5165);
xor U6536 (N_6536,N_5954,N_5790);
nand U6537 (N_6537,N_5105,N_5296);
or U6538 (N_6538,N_5705,N_5935);
nor U6539 (N_6539,N_5443,N_5520);
nand U6540 (N_6540,N_5194,N_5703);
nor U6541 (N_6541,N_5324,N_5163);
nand U6542 (N_6542,N_5265,N_5338);
nor U6543 (N_6543,N_5105,N_5686);
and U6544 (N_6544,N_5804,N_5286);
nor U6545 (N_6545,N_5095,N_5621);
or U6546 (N_6546,N_5314,N_5241);
xor U6547 (N_6547,N_5311,N_5243);
nand U6548 (N_6548,N_5052,N_5806);
nor U6549 (N_6549,N_5938,N_5510);
nand U6550 (N_6550,N_5880,N_5058);
nor U6551 (N_6551,N_5855,N_5610);
and U6552 (N_6552,N_5002,N_5109);
nor U6553 (N_6553,N_5007,N_5549);
nor U6554 (N_6554,N_5359,N_5819);
nor U6555 (N_6555,N_5471,N_5181);
nand U6556 (N_6556,N_5045,N_5715);
or U6557 (N_6557,N_5838,N_5474);
xnor U6558 (N_6558,N_5005,N_5295);
and U6559 (N_6559,N_5273,N_5836);
nor U6560 (N_6560,N_5415,N_5238);
xor U6561 (N_6561,N_5476,N_5814);
or U6562 (N_6562,N_5690,N_5721);
or U6563 (N_6563,N_5633,N_5145);
nor U6564 (N_6564,N_5338,N_5462);
xor U6565 (N_6565,N_5476,N_5317);
nand U6566 (N_6566,N_5348,N_5800);
xnor U6567 (N_6567,N_5402,N_5368);
or U6568 (N_6568,N_5179,N_5959);
and U6569 (N_6569,N_5926,N_5468);
or U6570 (N_6570,N_5754,N_5408);
xnor U6571 (N_6571,N_5879,N_5606);
and U6572 (N_6572,N_5636,N_5874);
nor U6573 (N_6573,N_5208,N_5465);
xor U6574 (N_6574,N_5181,N_5998);
xnor U6575 (N_6575,N_5103,N_5777);
nand U6576 (N_6576,N_5291,N_5145);
xor U6577 (N_6577,N_5206,N_5084);
xnor U6578 (N_6578,N_5847,N_5644);
nand U6579 (N_6579,N_5727,N_5286);
nand U6580 (N_6580,N_5987,N_5487);
nor U6581 (N_6581,N_5373,N_5590);
and U6582 (N_6582,N_5525,N_5855);
xor U6583 (N_6583,N_5180,N_5017);
or U6584 (N_6584,N_5764,N_5058);
nor U6585 (N_6585,N_5682,N_5702);
and U6586 (N_6586,N_5041,N_5536);
xnor U6587 (N_6587,N_5941,N_5091);
or U6588 (N_6588,N_5382,N_5330);
xnor U6589 (N_6589,N_5511,N_5252);
xor U6590 (N_6590,N_5647,N_5940);
xor U6591 (N_6591,N_5020,N_5105);
nor U6592 (N_6592,N_5111,N_5603);
nor U6593 (N_6593,N_5832,N_5787);
nor U6594 (N_6594,N_5602,N_5730);
nand U6595 (N_6595,N_5217,N_5197);
nor U6596 (N_6596,N_5143,N_5539);
nor U6597 (N_6597,N_5801,N_5023);
xnor U6598 (N_6598,N_5975,N_5857);
and U6599 (N_6599,N_5655,N_5576);
and U6600 (N_6600,N_5272,N_5070);
xnor U6601 (N_6601,N_5875,N_5189);
or U6602 (N_6602,N_5688,N_5846);
nor U6603 (N_6603,N_5300,N_5235);
xnor U6604 (N_6604,N_5030,N_5821);
or U6605 (N_6605,N_5491,N_5688);
and U6606 (N_6606,N_5221,N_5611);
or U6607 (N_6607,N_5513,N_5072);
or U6608 (N_6608,N_5495,N_5072);
and U6609 (N_6609,N_5319,N_5577);
and U6610 (N_6610,N_5298,N_5624);
nor U6611 (N_6611,N_5418,N_5415);
xor U6612 (N_6612,N_5695,N_5547);
xnor U6613 (N_6613,N_5577,N_5891);
xnor U6614 (N_6614,N_5107,N_5664);
nor U6615 (N_6615,N_5020,N_5066);
nand U6616 (N_6616,N_5202,N_5817);
xor U6617 (N_6617,N_5358,N_5855);
or U6618 (N_6618,N_5989,N_5096);
and U6619 (N_6619,N_5219,N_5954);
nor U6620 (N_6620,N_5742,N_5781);
and U6621 (N_6621,N_5949,N_5758);
nand U6622 (N_6622,N_5010,N_5645);
and U6623 (N_6623,N_5720,N_5735);
or U6624 (N_6624,N_5245,N_5970);
xnor U6625 (N_6625,N_5681,N_5009);
nor U6626 (N_6626,N_5561,N_5580);
nor U6627 (N_6627,N_5729,N_5008);
or U6628 (N_6628,N_5135,N_5034);
and U6629 (N_6629,N_5054,N_5579);
and U6630 (N_6630,N_5192,N_5662);
and U6631 (N_6631,N_5632,N_5915);
and U6632 (N_6632,N_5975,N_5970);
or U6633 (N_6633,N_5354,N_5380);
nand U6634 (N_6634,N_5101,N_5455);
or U6635 (N_6635,N_5939,N_5421);
or U6636 (N_6636,N_5625,N_5250);
nor U6637 (N_6637,N_5687,N_5156);
nor U6638 (N_6638,N_5265,N_5313);
nand U6639 (N_6639,N_5693,N_5073);
or U6640 (N_6640,N_5658,N_5156);
and U6641 (N_6641,N_5449,N_5053);
and U6642 (N_6642,N_5830,N_5560);
xor U6643 (N_6643,N_5059,N_5136);
and U6644 (N_6644,N_5339,N_5036);
xnor U6645 (N_6645,N_5210,N_5622);
xor U6646 (N_6646,N_5226,N_5191);
nand U6647 (N_6647,N_5433,N_5039);
nand U6648 (N_6648,N_5987,N_5954);
or U6649 (N_6649,N_5669,N_5227);
and U6650 (N_6650,N_5958,N_5156);
or U6651 (N_6651,N_5142,N_5651);
nor U6652 (N_6652,N_5959,N_5439);
or U6653 (N_6653,N_5837,N_5122);
nand U6654 (N_6654,N_5002,N_5407);
and U6655 (N_6655,N_5731,N_5680);
or U6656 (N_6656,N_5578,N_5673);
and U6657 (N_6657,N_5435,N_5534);
xnor U6658 (N_6658,N_5936,N_5315);
and U6659 (N_6659,N_5166,N_5981);
and U6660 (N_6660,N_5628,N_5667);
and U6661 (N_6661,N_5216,N_5104);
xor U6662 (N_6662,N_5603,N_5533);
or U6663 (N_6663,N_5644,N_5663);
or U6664 (N_6664,N_5700,N_5206);
xnor U6665 (N_6665,N_5867,N_5923);
xor U6666 (N_6666,N_5192,N_5504);
or U6667 (N_6667,N_5254,N_5330);
nand U6668 (N_6668,N_5435,N_5788);
xnor U6669 (N_6669,N_5090,N_5750);
xor U6670 (N_6670,N_5607,N_5658);
or U6671 (N_6671,N_5213,N_5644);
nand U6672 (N_6672,N_5571,N_5789);
and U6673 (N_6673,N_5666,N_5564);
and U6674 (N_6674,N_5031,N_5363);
nand U6675 (N_6675,N_5601,N_5500);
and U6676 (N_6676,N_5592,N_5761);
or U6677 (N_6677,N_5257,N_5104);
nor U6678 (N_6678,N_5272,N_5209);
xor U6679 (N_6679,N_5810,N_5807);
and U6680 (N_6680,N_5332,N_5198);
nor U6681 (N_6681,N_5202,N_5935);
nand U6682 (N_6682,N_5551,N_5689);
and U6683 (N_6683,N_5520,N_5945);
nand U6684 (N_6684,N_5295,N_5176);
and U6685 (N_6685,N_5652,N_5723);
nand U6686 (N_6686,N_5347,N_5079);
nand U6687 (N_6687,N_5774,N_5103);
nor U6688 (N_6688,N_5643,N_5078);
or U6689 (N_6689,N_5903,N_5124);
nand U6690 (N_6690,N_5672,N_5915);
nor U6691 (N_6691,N_5569,N_5319);
or U6692 (N_6692,N_5587,N_5100);
nand U6693 (N_6693,N_5115,N_5923);
nand U6694 (N_6694,N_5247,N_5973);
nand U6695 (N_6695,N_5842,N_5789);
nand U6696 (N_6696,N_5418,N_5796);
xor U6697 (N_6697,N_5101,N_5321);
nor U6698 (N_6698,N_5004,N_5860);
and U6699 (N_6699,N_5245,N_5032);
xor U6700 (N_6700,N_5125,N_5818);
nor U6701 (N_6701,N_5893,N_5381);
xnor U6702 (N_6702,N_5967,N_5175);
or U6703 (N_6703,N_5151,N_5827);
xnor U6704 (N_6704,N_5918,N_5586);
nand U6705 (N_6705,N_5475,N_5287);
xnor U6706 (N_6706,N_5144,N_5047);
nor U6707 (N_6707,N_5112,N_5639);
or U6708 (N_6708,N_5729,N_5500);
xor U6709 (N_6709,N_5205,N_5079);
xor U6710 (N_6710,N_5486,N_5246);
and U6711 (N_6711,N_5280,N_5933);
or U6712 (N_6712,N_5926,N_5564);
nand U6713 (N_6713,N_5993,N_5807);
and U6714 (N_6714,N_5056,N_5306);
and U6715 (N_6715,N_5429,N_5044);
xnor U6716 (N_6716,N_5186,N_5829);
and U6717 (N_6717,N_5129,N_5101);
xnor U6718 (N_6718,N_5778,N_5148);
xnor U6719 (N_6719,N_5991,N_5748);
nor U6720 (N_6720,N_5837,N_5078);
and U6721 (N_6721,N_5763,N_5813);
nor U6722 (N_6722,N_5211,N_5210);
nor U6723 (N_6723,N_5119,N_5530);
and U6724 (N_6724,N_5042,N_5441);
nand U6725 (N_6725,N_5170,N_5390);
or U6726 (N_6726,N_5343,N_5960);
and U6727 (N_6727,N_5631,N_5032);
nor U6728 (N_6728,N_5653,N_5243);
nor U6729 (N_6729,N_5106,N_5187);
or U6730 (N_6730,N_5357,N_5163);
nor U6731 (N_6731,N_5237,N_5786);
and U6732 (N_6732,N_5015,N_5325);
xor U6733 (N_6733,N_5938,N_5144);
nor U6734 (N_6734,N_5106,N_5345);
or U6735 (N_6735,N_5562,N_5076);
xor U6736 (N_6736,N_5809,N_5893);
or U6737 (N_6737,N_5848,N_5912);
or U6738 (N_6738,N_5305,N_5926);
or U6739 (N_6739,N_5719,N_5576);
nand U6740 (N_6740,N_5287,N_5949);
or U6741 (N_6741,N_5787,N_5081);
nand U6742 (N_6742,N_5610,N_5111);
nand U6743 (N_6743,N_5981,N_5556);
or U6744 (N_6744,N_5344,N_5008);
nand U6745 (N_6745,N_5711,N_5629);
nand U6746 (N_6746,N_5969,N_5560);
nand U6747 (N_6747,N_5287,N_5622);
nand U6748 (N_6748,N_5900,N_5524);
and U6749 (N_6749,N_5613,N_5078);
nor U6750 (N_6750,N_5632,N_5245);
or U6751 (N_6751,N_5038,N_5724);
nand U6752 (N_6752,N_5014,N_5609);
xor U6753 (N_6753,N_5778,N_5674);
xor U6754 (N_6754,N_5247,N_5744);
and U6755 (N_6755,N_5816,N_5411);
and U6756 (N_6756,N_5404,N_5986);
nor U6757 (N_6757,N_5948,N_5460);
and U6758 (N_6758,N_5141,N_5794);
nand U6759 (N_6759,N_5182,N_5341);
or U6760 (N_6760,N_5746,N_5623);
nor U6761 (N_6761,N_5372,N_5337);
or U6762 (N_6762,N_5303,N_5454);
and U6763 (N_6763,N_5118,N_5265);
or U6764 (N_6764,N_5762,N_5874);
nor U6765 (N_6765,N_5901,N_5314);
nand U6766 (N_6766,N_5432,N_5460);
xor U6767 (N_6767,N_5387,N_5921);
nor U6768 (N_6768,N_5380,N_5452);
nor U6769 (N_6769,N_5516,N_5717);
and U6770 (N_6770,N_5515,N_5858);
or U6771 (N_6771,N_5367,N_5038);
or U6772 (N_6772,N_5257,N_5611);
or U6773 (N_6773,N_5047,N_5820);
nand U6774 (N_6774,N_5140,N_5039);
or U6775 (N_6775,N_5099,N_5354);
nor U6776 (N_6776,N_5634,N_5641);
or U6777 (N_6777,N_5638,N_5202);
or U6778 (N_6778,N_5669,N_5819);
or U6779 (N_6779,N_5217,N_5398);
nand U6780 (N_6780,N_5688,N_5690);
and U6781 (N_6781,N_5211,N_5061);
xnor U6782 (N_6782,N_5161,N_5141);
nor U6783 (N_6783,N_5434,N_5162);
or U6784 (N_6784,N_5401,N_5216);
nand U6785 (N_6785,N_5359,N_5253);
nor U6786 (N_6786,N_5593,N_5709);
xnor U6787 (N_6787,N_5075,N_5332);
nor U6788 (N_6788,N_5214,N_5196);
and U6789 (N_6789,N_5822,N_5543);
nor U6790 (N_6790,N_5742,N_5514);
nor U6791 (N_6791,N_5044,N_5053);
nor U6792 (N_6792,N_5854,N_5551);
nand U6793 (N_6793,N_5623,N_5278);
or U6794 (N_6794,N_5475,N_5436);
or U6795 (N_6795,N_5981,N_5474);
nand U6796 (N_6796,N_5135,N_5663);
or U6797 (N_6797,N_5200,N_5224);
nand U6798 (N_6798,N_5943,N_5590);
or U6799 (N_6799,N_5520,N_5232);
and U6800 (N_6800,N_5794,N_5845);
nand U6801 (N_6801,N_5112,N_5657);
and U6802 (N_6802,N_5823,N_5184);
nand U6803 (N_6803,N_5799,N_5521);
xnor U6804 (N_6804,N_5280,N_5614);
and U6805 (N_6805,N_5091,N_5076);
and U6806 (N_6806,N_5202,N_5940);
nor U6807 (N_6807,N_5213,N_5916);
nand U6808 (N_6808,N_5366,N_5525);
nand U6809 (N_6809,N_5405,N_5258);
or U6810 (N_6810,N_5424,N_5747);
nand U6811 (N_6811,N_5094,N_5874);
or U6812 (N_6812,N_5621,N_5945);
nand U6813 (N_6813,N_5753,N_5402);
nor U6814 (N_6814,N_5337,N_5949);
or U6815 (N_6815,N_5041,N_5509);
nand U6816 (N_6816,N_5513,N_5936);
or U6817 (N_6817,N_5726,N_5590);
nor U6818 (N_6818,N_5795,N_5731);
xor U6819 (N_6819,N_5642,N_5203);
and U6820 (N_6820,N_5547,N_5258);
nand U6821 (N_6821,N_5624,N_5426);
xnor U6822 (N_6822,N_5605,N_5110);
nor U6823 (N_6823,N_5960,N_5591);
nand U6824 (N_6824,N_5408,N_5694);
or U6825 (N_6825,N_5761,N_5560);
nand U6826 (N_6826,N_5840,N_5894);
and U6827 (N_6827,N_5836,N_5428);
or U6828 (N_6828,N_5742,N_5389);
nor U6829 (N_6829,N_5395,N_5565);
and U6830 (N_6830,N_5010,N_5070);
xnor U6831 (N_6831,N_5919,N_5601);
or U6832 (N_6832,N_5663,N_5372);
xor U6833 (N_6833,N_5301,N_5709);
xor U6834 (N_6834,N_5090,N_5801);
xor U6835 (N_6835,N_5786,N_5796);
xor U6836 (N_6836,N_5902,N_5175);
xor U6837 (N_6837,N_5889,N_5948);
nand U6838 (N_6838,N_5526,N_5920);
or U6839 (N_6839,N_5022,N_5548);
nand U6840 (N_6840,N_5226,N_5216);
or U6841 (N_6841,N_5921,N_5620);
nand U6842 (N_6842,N_5158,N_5973);
or U6843 (N_6843,N_5303,N_5227);
nand U6844 (N_6844,N_5466,N_5798);
nand U6845 (N_6845,N_5066,N_5415);
or U6846 (N_6846,N_5983,N_5565);
nor U6847 (N_6847,N_5383,N_5836);
nand U6848 (N_6848,N_5955,N_5364);
or U6849 (N_6849,N_5038,N_5106);
nand U6850 (N_6850,N_5562,N_5831);
xnor U6851 (N_6851,N_5479,N_5020);
or U6852 (N_6852,N_5183,N_5766);
nor U6853 (N_6853,N_5439,N_5207);
nand U6854 (N_6854,N_5969,N_5847);
or U6855 (N_6855,N_5302,N_5899);
nor U6856 (N_6856,N_5071,N_5116);
and U6857 (N_6857,N_5555,N_5498);
xnor U6858 (N_6858,N_5968,N_5742);
nor U6859 (N_6859,N_5275,N_5158);
or U6860 (N_6860,N_5305,N_5918);
nand U6861 (N_6861,N_5515,N_5183);
xor U6862 (N_6862,N_5254,N_5835);
or U6863 (N_6863,N_5454,N_5428);
nor U6864 (N_6864,N_5568,N_5446);
or U6865 (N_6865,N_5483,N_5731);
xnor U6866 (N_6866,N_5421,N_5042);
xnor U6867 (N_6867,N_5094,N_5919);
nand U6868 (N_6868,N_5442,N_5219);
nand U6869 (N_6869,N_5951,N_5708);
nor U6870 (N_6870,N_5586,N_5676);
or U6871 (N_6871,N_5551,N_5213);
or U6872 (N_6872,N_5532,N_5713);
and U6873 (N_6873,N_5293,N_5794);
and U6874 (N_6874,N_5374,N_5497);
xnor U6875 (N_6875,N_5540,N_5292);
nor U6876 (N_6876,N_5233,N_5231);
nor U6877 (N_6877,N_5130,N_5236);
xnor U6878 (N_6878,N_5075,N_5058);
and U6879 (N_6879,N_5196,N_5638);
nand U6880 (N_6880,N_5083,N_5248);
nand U6881 (N_6881,N_5849,N_5869);
nand U6882 (N_6882,N_5092,N_5653);
nand U6883 (N_6883,N_5090,N_5069);
nand U6884 (N_6884,N_5239,N_5775);
nand U6885 (N_6885,N_5334,N_5466);
nor U6886 (N_6886,N_5881,N_5330);
nor U6887 (N_6887,N_5522,N_5338);
xor U6888 (N_6888,N_5539,N_5287);
and U6889 (N_6889,N_5840,N_5022);
nor U6890 (N_6890,N_5175,N_5227);
nor U6891 (N_6891,N_5393,N_5973);
or U6892 (N_6892,N_5639,N_5046);
xnor U6893 (N_6893,N_5391,N_5424);
and U6894 (N_6894,N_5231,N_5225);
xor U6895 (N_6895,N_5742,N_5010);
nor U6896 (N_6896,N_5435,N_5785);
nand U6897 (N_6897,N_5393,N_5565);
or U6898 (N_6898,N_5954,N_5670);
nor U6899 (N_6899,N_5868,N_5201);
xnor U6900 (N_6900,N_5757,N_5694);
or U6901 (N_6901,N_5904,N_5461);
nor U6902 (N_6902,N_5498,N_5116);
nand U6903 (N_6903,N_5952,N_5922);
nand U6904 (N_6904,N_5183,N_5009);
or U6905 (N_6905,N_5242,N_5178);
or U6906 (N_6906,N_5524,N_5554);
xnor U6907 (N_6907,N_5972,N_5711);
and U6908 (N_6908,N_5665,N_5523);
or U6909 (N_6909,N_5354,N_5304);
nor U6910 (N_6910,N_5934,N_5128);
or U6911 (N_6911,N_5723,N_5434);
and U6912 (N_6912,N_5438,N_5929);
and U6913 (N_6913,N_5049,N_5824);
or U6914 (N_6914,N_5298,N_5422);
xor U6915 (N_6915,N_5556,N_5459);
nand U6916 (N_6916,N_5221,N_5788);
nor U6917 (N_6917,N_5902,N_5748);
or U6918 (N_6918,N_5892,N_5943);
nand U6919 (N_6919,N_5285,N_5029);
or U6920 (N_6920,N_5156,N_5364);
nor U6921 (N_6921,N_5152,N_5904);
nor U6922 (N_6922,N_5119,N_5978);
nand U6923 (N_6923,N_5673,N_5947);
or U6924 (N_6924,N_5049,N_5214);
nor U6925 (N_6925,N_5960,N_5479);
xor U6926 (N_6926,N_5696,N_5314);
and U6927 (N_6927,N_5680,N_5547);
or U6928 (N_6928,N_5699,N_5537);
and U6929 (N_6929,N_5663,N_5583);
xor U6930 (N_6930,N_5620,N_5639);
or U6931 (N_6931,N_5694,N_5613);
nor U6932 (N_6932,N_5750,N_5277);
nor U6933 (N_6933,N_5929,N_5232);
nor U6934 (N_6934,N_5070,N_5786);
and U6935 (N_6935,N_5904,N_5263);
nor U6936 (N_6936,N_5572,N_5294);
nor U6937 (N_6937,N_5952,N_5248);
xnor U6938 (N_6938,N_5959,N_5273);
nand U6939 (N_6939,N_5550,N_5000);
or U6940 (N_6940,N_5049,N_5787);
or U6941 (N_6941,N_5861,N_5882);
xnor U6942 (N_6942,N_5124,N_5608);
nor U6943 (N_6943,N_5718,N_5059);
and U6944 (N_6944,N_5841,N_5382);
xnor U6945 (N_6945,N_5655,N_5023);
and U6946 (N_6946,N_5097,N_5435);
or U6947 (N_6947,N_5556,N_5570);
and U6948 (N_6948,N_5244,N_5627);
xor U6949 (N_6949,N_5253,N_5871);
nor U6950 (N_6950,N_5409,N_5887);
and U6951 (N_6951,N_5716,N_5606);
or U6952 (N_6952,N_5711,N_5927);
xor U6953 (N_6953,N_5740,N_5273);
nor U6954 (N_6954,N_5043,N_5460);
or U6955 (N_6955,N_5002,N_5561);
xnor U6956 (N_6956,N_5942,N_5052);
nand U6957 (N_6957,N_5565,N_5037);
nand U6958 (N_6958,N_5754,N_5991);
xor U6959 (N_6959,N_5068,N_5009);
nand U6960 (N_6960,N_5961,N_5256);
and U6961 (N_6961,N_5773,N_5365);
xor U6962 (N_6962,N_5479,N_5016);
xnor U6963 (N_6963,N_5790,N_5907);
and U6964 (N_6964,N_5718,N_5428);
nor U6965 (N_6965,N_5368,N_5790);
nor U6966 (N_6966,N_5366,N_5596);
nor U6967 (N_6967,N_5711,N_5609);
nand U6968 (N_6968,N_5861,N_5712);
or U6969 (N_6969,N_5383,N_5029);
and U6970 (N_6970,N_5723,N_5701);
nor U6971 (N_6971,N_5998,N_5056);
nor U6972 (N_6972,N_5948,N_5212);
or U6973 (N_6973,N_5653,N_5672);
nand U6974 (N_6974,N_5684,N_5393);
nand U6975 (N_6975,N_5447,N_5193);
xor U6976 (N_6976,N_5738,N_5413);
and U6977 (N_6977,N_5530,N_5172);
xor U6978 (N_6978,N_5816,N_5132);
nand U6979 (N_6979,N_5009,N_5330);
or U6980 (N_6980,N_5190,N_5910);
and U6981 (N_6981,N_5325,N_5495);
nand U6982 (N_6982,N_5561,N_5562);
and U6983 (N_6983,N_5867,N_5953);
or U6984 (N_6984,N_5036,N_5976);
nor U6985 (N_6985,N_5903,N_5543);
or U6986 (N_6986,N_5223,N_5876);
xnor U6987 (N_6987,N_5718,N_5135);
xor U6988 (N_6988,N_5274,N_5529);
nor U6989 (N_6989,N_5827,N_5156);
nor U6990 (N_6990,N_5181,N_5018);
or U6991 (N_6991,N_5004,N_5818);
nor U6992 (N_6992,N_5231,N_5047);
xnor U6993 (N_6993,N_5232,N_5973);
xor U6994 (N_6994,N_5877,N_5783);
nand U6995 (N_6995,N_5118,N_5298);
xnor U6996 (N_6996,N_5856,N_5772);
xnor U6997 (N_6997,N_5163,N_5164);
nand U6998 (N_6998,N_5340,N_5027);
xnor U6999 (N_6999,N_5936,N_5468);
nand U7000 (N_7000,N_6621,N_6587);
or U7001 (N_7001,N_6726,N_6592);
xor U7002 (N_7002,N_6523,N_6835);
or U7003 (N_7003,N_6073,N_6636);
xnor U7004 (N_7004,N_6371,N_6915);
and U7005 (N_7005,N_6275,N_6402);
nor U7006 (N_7006,N_6808,N_6454);
nand U7007 (N_7007,N_6052,N_6833);
nor U7008 (N_7008,N_6158,N_6113);
or U7009 (N_7009,N_6686,N_6432);
nand U7010 (N_7010,N_6382,N_6099);
nand U7011 (N_7011,N_6519,N_6150);
xnor U7012 (N_7012,N_6561,N_6663);
nand U7013 (N_7013,N_6579,N_6873);
and U7014 (N_7014,N_6784,N_6023);
nor U7015 (N_7015,N_6494,N_6968);
xor U7016 (N_7016,N_6600,N_6548);
and U7017 (N_7017,N_6672,N_6474);
and U7018 (N_7018,N_6377,N_6249);
xnor U7019 (N_7019,N_6864,N_6811);
and U7020 (N_7020,N_6842,N_6146);
nor U7021 (N_7021,N_6353,N_6963);
nand U7022 (N_7022,N_6263,N_6043);
nor U7023 (N_7023,N_6450,N_6568);
nand U7024 (N_7024,N_6834,N_6143);
xor U7025 (N_7025,N_6046,N_6491);
xnor U7026 (N_7026,N_6197,N_6040);
xor U7027 (N_7027,N_6566,N_6651);
nand U7028 (N_7028,N_6274,N_6369);
nand U7029 (N_7029,N_6209,N_6329);
nor U7030 (N_7030,N_6313,N_6222);
nand U7031 (N_7031,N_6528,N_6221);
xor U7032 (N_7032,N_6495,N_6928);
xor U7033 (N_7033,N_6298,N_6089);
nor U7034 (N_7034,N_6166,N_6152);
or U7035 (N_7035,N_6612,N_6986);
xnor U7036 (N_7036,N_6945,N_6542);
nand U7037 (N_7037,N_6799,N_6302);
nor U7038 (N_7038,N_6457,N_6848);
and U7039 (N_7039,N_6057,N_6169);
nor U7040 (N_7040,N_6220,N_6822);
or U7041 (N_7041,N_6095,N_6085);
xor U7042 (N_7042,N_6815,N_6713);
xnor U7043 (N_7043,N_6892,N_6324);
nor U7044 (N_7044,N_6829,N_6712);
and U7045 (N_7045,N_6747,N_6859);
nor U7046 (N_7046,N_6678,N_6756);
nand U7047 (N_7047,N_6002,N_6477);
and U7048 (N_7048,N_6593,N_6479);
nand U7049 (N_7049,N_6845,N_6520);
nor U7050 (N_7050,N_6252,N_6708);
or U7051 (N_7051,N_6826,N_6164);
nand U7052 (N_7052,N_6530,N_6465);
xor U7053 (N_7053,N_6237,N_6108);
and U7054 (N_7054,N_6696,N_6047);
or U7055 (N_7055,N_6422,N_6580);
nor U7056 (N_7056,N_6656,N_6508);
nor U7057 (N_7057,N_6137,N_6946);
or U7058 (N_7058,N_6412,N_6130);
nor U7059 (N_7059,N_6261,N_6549);
or U7060 (N_7060,N_6832,N_6200);
xnor U7061 (N_7061,N_6560,N_6206);
nor U7062 (N_7062,N_6694,N_6724);
nor U7063 (N_7063,N_6638,N_6644);
and U7064 (N_7064,N_6781,N_6637);
or U7065 (N_7065,N_6253,N_6846);
xnor U7066 (N_7066,N_6414,N_6437);
and U7067 (N_7067,N_6420,N_6155);
or U7068 (N_7068,N_6788,N_6762);
and U7069 (N_7069,N_6987,N_6758);
nor U7070 (N_7070,N_6075,N_6856);
xor U7071 (N_7071,N_6148,N_6136);
nand U7072 (N_7072,N_6468,N_6339);
nand U7073 (N_7073,N_6405,N_6559);
and U7074 (N_7074,N_6092,N_6486);
nand U7075 (N_7075,N_6213,N_6994);
nand U7076 (N_7076,N_6081,N_6004);
nand U7077 (N_7077,N_6105,N_6289);
xnor U7078 (N_7078,N_6322,N_6596);
nor U7079 (N_7079,N_6721,N_6199);
nor U7080 (N_7080,N_6080,N_6719);
or U7081 (N_7081,N_6993,N_6424);
or U7082 (N_7082,N_6373,N_6086);
or U7083 (N_7083,N_6122,N_6731);
and U7084 (N_7084,N_6647,N_6769);
nand U7085 (N_7085,N_6436,N_6916);
or U7086 (N_7086,N_6957,N_6456);
and U7087 (N_7087,N_6540,N_6078);
xnor U7088 (N_7088,N_6074,N_6140);
xnor U7089 (N_7089,N_6624,N_6677);
nor U7090 (N_7090,N_6818,N_6665);
and U7091 (N_7091,N_6959,N_6445);
xnor U7092 (N_7092,N_6506,N_6408);
and U7093 (N_7093,N_6443,N_6648);
nor U7094 (N_7094,N_6689,N_6397);
or U7095 (N_7095,N_6502,N_6280);
nand U7096 (N_7096,N_6933,N_6386);
or U7097 (N_7097,N_6279,N_6425);
and U7098 (N_7098,N_6861,N_6489);
nor U7099 (N_7099,N_6463,N_6783);
xnor U7100 (N_7100,N_6055,N_6983);
nor U7101 (N_7101,N_6490,N_6179);
xnor U7102 (N_7102,N_6910,N_6662);
nand U7103 (N_7103,N_6168,N_6746);
nor U7104 (N_7104,N_6258,N_6673);
xnor U7105 (N_7105,N_6557,N_6773);
and U7106 (N_7106,N_6028,N_6904);
xor U7107 (N_7107,N_6035,N_6185);
nand U7108 (N_7108,N_6884,N_6666);
nor U7109 (N_7109,N_6188,N_6899);
xor U7110 (N_7110,N_6699,N_6021);
and U7111 (N_7111,N_6934,N_6905);
or U7112 (N_7112,N_6416,N_6650);
nor U7113 (N_7113,N_6307,N_6922);
nand U7114 (N_7114,N_6190,N_6142);
nor U7115 (N_7115,N_6608,N_6157);
xor U7116 (N_7116,N_6435,N_6558);
and U7117 (N_7117,N_6367,N_6356);
or U7118 (N_7118,N_6024,N_6501);
nor U7119 (N_7119,N_6332,N_6428);
and U7120 (N_7120,N_6093,N_6124);
nor U7121 (N_7121,N_6334,N_6552);
nand U7122 (N_7122,N_6964,N_6698);
xor U7123 (N_7123,N_6882,N_6544);
or U7124 (N_7124,N_6738,N_6151);
nor U7125 (N_7125,N_6704,N_6399);
xnor U7126 (N_7126,N_6639,N_6238);
xnor U7127 (N_7127,N_6867,N_6452);
xnor U7128 (N_7128,N_6620,N_6264);
or U7129 (N_7129,N_6553,N_6091);
nand U7130 (N_7130,N_6734,N_6088);
nor U7131 (N_7131,N_6740,N_6145);
nor U7132 (N_7132,N_6999,N_6935);
nand U7133 (N_7133,N_6067,N_6281);
or U7134 (N_7134,N_6326,N_6603);
nor U7135 (N_7135,N_6855,N_6215);
and U7136 (N_7136,N_6260,N_6998);
nand U7137 (N_7137,N_6295,N_6819);
nor U7138 (N_7138,N_6582,N_6017);
and U7139 (N_7139,N_6574,N_6655);
xnor U7140 (N_7140,N_6243,N_6676);
nor U7141 (N_7141,N_6201,N_6907);
or U7142 (N_7142,N_6913,N_6615);
or U7143 (N_7143,N_6265,N_6059);
nor U7144 (N_7144,N_6276,N_6966);
and U7145 (N_7145,N_6393,N_6606);
xor U7146 (N_7146,N_6288,N_6908);
xnor U7147 (N_7147,N_6887,N_6730);
and U7148 (N_7148,N_6268,N_6387);
or U7149 (N_7149,N_6446,N_6975);
xnor U7150 (N_7150,N_6352,N_6550);
nor U7151 (N_7151,N_6919,N_6011);
and U7152 (N_7152,N_6785,N_6051);
or U7153 (N_7153,N_6359,N_6466);
or U7154 (N_7154,N_6044,N_6601);
and U7155 (N_7155,N_6009,N_6453);
xor U7156 (N_7156,N_6283,N_6898);
or U7157 (N_7157,N_6400,N_6459);
xnor U7158 (N_7158,N_6187,N_6180);
nor U7159 (N_7159,N_6034,N_6618);
nand U7160 (N_7160,N_6375,N_6320);
nand U7161 (N_7161,N_6880,N_6522);
and U7162 (N_7162,N_6310,N_6628);
and U7163 (N_7163,N_6707,N_6172);
and U7164 (N_7164,N_6690,N_6803);
and U7165 (N_7165,N_6363,N_6054);
and U7166 (N_7166,N_6404,N_6364);
nand U7167 (N_7167,N_6248,N_6349);
or U7168 (N_7168,N_6537,N_6100);
nor U7169 (N_7169,N_6485,N_6003);
and U7170 (N_7170,N_6451,N_6094);
nand U7171 (N_7171,N_6077,N_6189);
nor U7172 (N_7172,N_6555,N_6029);
or U7173 (N_7173,N_6809,N_6792);
or U7174 (N_7174,N_6497,N_6132);
nor U7175 (N_7175,N_6763,N_6000);
nor U7176 (N_7176,N_6695,N_6267);
nand U7177 (N_7177,N_6764,N_6604);
or U7178 (N_7178,N_6160,N_6256);
or U7179 (N_7179,N_6737,N_6729);
or U7180 (N_7180,N_6936,N_6609);
or U7181 (N_7181,N_6970,N_6355);
nand U7182 (N_7182,N_6810,N_6617);
nand U7183 (N_7183,N_6259,N_6346);
xor U7184 (N_7184,N_6794,N_6623);
nand U7185 (N_7185,N_6126,N_6817);
xnor U7186 (N_7186,N_6976,N_6162);
nand U7187 (N_7187,N_6223,N_6217);
xnor U7188 (N_7188,N_6991,N_6610);
and U7189 (N_7189,N_6433,N_6667);
nand U7190 (N_7190,N_6296,N_6039);
nand U7191 (N_7191,N_6571,N_6447);
nor U7192 (N_7192,N_6509,N_6943);
xor U7193 (N_7193,N_6480,N_6594);
xnor U7194 (N_7194,N_6337,N_6518);
or U7195 (N_7195,N_6431,N_6038);
or U7196 (N_7196,N_6183,N_6900);
nor U7197 (N_7197,N_6083,N_6379);
xor U7198 (N_7198,N_6455,N_6374);
or U7199 (N_7199,N_6728,N_6037);
xor U7200 (N_7200,N_6761,N_6668);
or U7201 (N_7201,N_6354,N_6865);
or U7202 (N_7202,N_6875,N_6458);
nor U7203 (N_7203,N_6777,N_6068);
or U7204 (N_7204,N_6564,N_6851);
and U7205 (N_7205,N_6331,N_6210);
xor U7206 (N_7206,N_6025,N_6406);
xor U7207 (N_7207,N_6551,N_6780);
and U7208 (N_7208,N_6026,N_6144);
and U7209 (N_7209,N_6333,N_6543);
nand U7210 (N_7210,N_6242,N_6066);
or U7211 (N_7211,N_6565,N_6679);
and U7212 (N_7212,N_6671,N_6942);
or U7213 (N_7213,N_6498,N_6710);
nor U7214 (N_7214,N_6891,N_6939);
xnor U7215 (N_7215,N_6635,N_6309);
or U7216 (N_7216,N_6511,N_6583);
and U7217 (N_7217,N_6415,N_6335);
and U7218 (N_7218,N_6239,N_6419);
nor U7219 (N_7219,N_6921,N_6972);
xor U7220 (N_7220,N_6717,N_6988);
nand U7221 (N_7221,N_6286,N_6343);
or U7222 (N_7222,N_6653,N_6700);
and U7223 (N_7223,N_6722,N_6439);
xnor U7224 (N_7224,N_6076,N_6643);
xnor U7225 (N_7225,N_6409,N_6982);
or U7226 (N_7226,N_6850,N_6438);
or U7227 (N_7227,N_6049,N_6174);
xnor U7228 (N_7228,N_6351,N_6996);
nor U7229 (N_7229,N_6303,N_6167);
nand U7230 (N_7230,N_6563,N_6484);
or U7231 (N_7231,N_6901,N_6478);
nor U7232 (N_7232,N_6366,N_6545);
xnor U7233 (N_7233,N_6526,N_6849);
and U7234 (N_7234,N_6599,N_6370);
and U7235 (N_7235,N_6546,N_6423);
or U7236 (N_7236,N_6793,N_6954);
nand U7237 (N_7237,N_6776,N_6036);
nor U7238 (N_7238,N_6118,N_6929);
or U7239 (N_7239,N_6398,N_6013);
or U7240 (N_7240,N_6410,N_6119);
xor U7241 (N_7241,N_6517,N_6103);
nand U7242 (N_7242,N_6997,N_6765);
and U7243 (N_7243,N_6585,N_6814);
nor U7244 (N_7244,N_6109,N_6311);
nand U7245 (N_7245,N_6018,N_6874);
xor U7246 (N_7246,N_6471,N_6971);
xor U7247 (N_7247,N_6853,N_6902);
or U7248 (N_7248,N_6175,N_6031);
and U7249 (N_7249,N_6634,N_6225);
nor U7250 (N_7250,N_6787,N_6247);
or U7251 (N_7251,N_6056,N_6828);
and U7252 (N_7252,N_6362,N_6766);
nor U7253 (N_7253,N_6470,N_6589);
xor U7254 (N_7254,N_6607,N_6125);
and U7255 (N_7255,N_6529,N_6595);
nand U7256 (N_7256,N_6032,N_6461);
or U7257 (N_7257,N_6736,N_6858);
nand U7258 (N_7258,N_6981,N_6531);
and U7259 (N_7259,N_6755,N_6821);
and U7260 (N_7260,N_6318,N_6319);
or U7261 (N_7261,N_6956,N_6990);
and U7262 (N_7262,N_6228,N_6868);
or U7263 (N_7263,N_6779,N_6961);
or U7264 (N_7264,N_6840,N_6927);
and U7265 (N_7265,N_6512,N_6652);
or U7266 (N_7266,N_6016,N_6820);
xnor U7267 (N_7267,N_6178,N_6448);
and U7268 (N_7268,N_6232,N_6196);
and U7269 (N_7269,N_6147,N_6503);
xnor U7270 (N_7270,N_6205,N_6951);
xor U7271 (N_7271,N_6872,N_6460);
nor U7272 (N_7272,N_6926,N_6413);
nor U7273 (N_7273,N_6345,N_6467);
and U7274 (N_7274,N_6616,N_6812);
nor U7275 (N_7275,N_6064,N_6277);
nor U7276 (N_7276,N_6775,N_6577);
nand U7277 (N_7277,N_6597,N_6154);
nand U7278 (N_7278,N_6866,N_6153);
nand U7279 (N_7279,N_6058,N_6920);
and U7280 (N_7280,N_6684,N_6930);
or U7281 (N_7281,N_6715,N_6115);
xor U7282 (N_7282,N_6012,N_6824);
or U7283 (N_7283,N_6847,N_6019);
xnor U7284 (N_7284,N_6973,N_6500);
or U7285 (N_7285,N_6360,N_6208);
nor U7286 (N_7286,N_6072,N_6429);
xor U7287 (N_7287,N_6316,N_6378);
nand U7288 (N_7288,N_6321,N_6925);
xor U7289 (N_7289,N_6245,N_6692);
nor U7290 (N_7290,N_6294,N_6590);
and U7291 (N_7291,N_6182,N_6576);
xor U7292 (N_7292,N_6348,N_6389);
nor U7293 (N_7293,N_6657,N_6212);
xor U7294 (N_7294,N_6706,N_6687);
nand U7295 (N_7295,N_6863,N_6805);
or U7296 (N_7296,N_6030,N_6202);
nor U7297 (N_7297,N_6739,N_6895);
nand U7298 (N_7298,N_6417,N_6978);
or U7299 (N_7299,N_6837,N_6640);
or U7300 (N_7300,N_6001,N_6204);
or U7301 (N_7301,N_6266,N_6883);
nand U7302 (N_7302,N_6368,N_6444);
xnor U7303 (N_7303,N_6135,N_6969);
and U7304 (N_7304,N_6149,N_6536);
or U7305 (N_7305,N_6641,N_6790);
and U7306 (N_7306,N_6101,N_6693);
nand U7307 (N_7307,N_6116,N_6312);
or U7308 (N_7308,N_6314,N_6768);
nor U7309 (N_7309,N_6234,N_6984);
nor U7310 (N_7310,N_6723,N_6427);
and U7311 (N_7311,N_6629,N_6795);
and U7312 (N_7312,N_6931,N_6173);
nor U7313 (N_7313,N_6938,N_6513);
and U7314 (N_7314,N_6754,N_6507);
xor U7315 (N_7315,N_6195,N_6669);
or U7316 (N_7316,N_6390,N_6096);
and U7317 (N_7317,N_6749,N_6469);
nand U7318 (N_7318,N_6732,N_6660);
and U7319 (N_7319,N_6308,N_6838);
or U7320 (N_7320,N_6914,N_6060);
or U7321 (N_7321,N_6207,N_6211);
nor U7322 (N_7322,N_6006,N_6575);
nor U7323 (N_7323,N_6798,N_6163);
nand U7324 (N_7324,N_6114,N_6664);
nor U7325 (N_7325,N_6071,N_6952);
or U7326 (N_7326,N_6770,N_6005);
xor U7327 (N_7327,N_6381,N_6138);
nor U7328 (N_7328,N_6654,N_6069);
or U7329 (N_7329,N_6293,N_6789);
or U7330 (N_7330,N_6361,N_6924);
nor U7331 (N_7331,N_6886,N_6889);
and U7332 (N_7332,N_6483,N_6102);
nor U7333 (N_7333,N_6940,N_6284);
and U7334 (N_7334,N_6515,N_6906);
xnor U7335 (N_7335,N_6745,N_6878);
xor U7336 (N_7336,N_6649,N_6744);
xor U7337 (N_7337,N_6133,N_6569);
xor U7338 (N_7338,N_6421,N_6586);
or U7339 (N_7339,N_6801,N_6227);
or U7340 (N_7340,N_6750,N_6807);
or U7341 (N_7341,N_6464,N_6711);
nand U7342 (N_7342,N_6441,N_6688);
and U7343 (N_7343,N_6980,N_6434);
nor U7344 (N_7344,N_6062,N_6918);
or U7345 (N_7345,N_6357,N_6514);
nor U7346 (N_7346,N_6358,N_6287);
xor U7347 (N_7347,N_6462,N_6989);
xnor U7348 (N_7348,N_6584,N_6090);
nor U7349 (N_7349,N_6752,N_6977);
nand U7350 (N_7350,N_6979,N_6893);
nor U7351 (N_7351,N_6767,N_6219);
and U7352 (N_7352,N_6831,N_6107);
xor U7353 (N_7353,N_6251,N_6128);
or U7354 (N_7354,N_6301,N_6341);
xor U7355 (N_7355,N_6282,N_6020);
xor U7356 (N_7356,N_6338,N_6879);
nor U7357 (N_7357,N_6725,N_6186);
or U7358 (N_7358,N_6937,N_6254);
and U7359 (N_7359,N_6087,N_6622);
nand U7360 (N_7360,N_6944,N_6112);
or U7361 (N_7361,N_6097,N_6014);
and U7362 (N_7362,N_6547,N_6860);
and U7363 (N_7363,N_6129,N_6521);
or U7364 (N_7364,N_6554,N_6198);
nor U7365 (N_7365,N_6701,N_6176);
xnor U7366 (N_7366,N_6475,N_6658);
nor U7367 (N_7367,N_6631,N_6403);
nor U7368 (N_7368,N_6246,N_6022);
nor U7369 (N_7369,N_6297,N_6958);
nor U7370 (N_7370,N_6141,N_6401);
or U7371 (N_7371,N_6852,N_6917);
and U7372 (N_7372,N_6830,N_6045);
nand U7373 (N_7373,N_6203,N_6110);
and U7374 (N_7374,N_6953,N_6327);
nand U7375 (N_7375,N_6816,N_6292);
xnor U7376 (N_7376,N_6825,N_6159);
nand U7377 (N_7377,N_6170,N_6082);
nor U7378 (N_7378,N_6778,N_6659);
nand U7379 (N_7379,N_6449,N_6748);
nand U7380 (N_7380,N_6870,N_6800);
nand U7381 (N_7381,N_6236,N_6300);
or U7382 (N_7382,N_6534,N_6941);
nand U7383 (N_7383,N_6562,N_6836);
and U7384 (N_7384,N_6588,N_6131);
nor U7385 (N_7385,N_6070,N_6877);
xor U7386 (N_7386,N_6702,N_6705);
or U7387 (N_7387,N_6079,N_6241);
and U7388 (N_7388,N_6235,N_6304);
nand U7389 (N_7389,N_6048,N_6255);
or U7390 (N_7390,N_6985,N_6084);
xor U7391 (N_7391,N_6912,N_6974);
xnor U7392 (N_7392,N_6797,N_6123);
xnor U7393 (N_7393,N_6675,N_6504);
nor U7394 (N_7394,N_6697,N_6121);
xor U7395 (N_7395,N_6139,N_6871);
nand U7396 (N_7396,N_6890,N_6008);
and U7397 (N_7397,N_6720,N_6718);
or U7398 (N_7398,N_6573,N_6473);
and U7399 (N_7399,N_6661,N_6796);
nand U7400 (N_7400,N_6909,N_6733);
nor U7401 (N_7401,N_6857,N_6193);
and U7402 (N_7402,N_6535,N_6336);
xnor U7403 (N_7403,N_6226,N_6372);
or U7404 (N_7404,N_6407,N_6010);
xor U7405 (N_7405,N_6960,N_6120);
nor U7406 (N_7406,N_6299,N_6743);
nor U7407 (N_7407,N_6098,N_6156);
and U7408 (N_7408,N_6218,N_6053);
and U7409 (N_7409,N_6041,N_6315);
xor U7410 (N_7410,N_6290,N_6325);
and U7411 (N_7411,N_6802,N_6330);
xnor U7412 (N_7412,N_6365,N_6772);
or U7413 (N_7413,N_6903,N_6224);
xor U7414 (N_7414,N_6305,N_6727);
nor U7415 (N_7415,N_6488,N_6556);
xnor U7416 (N_7416,N_6625,N_6681);
nand U7417 (N_7417,N_6760,N_6626);
and U7418 (N_7418,N_6385,N_6843);
and U7419 (N_7419,N_6033,N_6394);
or U7420 (N_7420,N_6442,N_6955);
or U7421 (N_7421,N_6632,N_6881);
and U7422 (N_7422,N_6806,N_6876);
nor U7423 (N_7423,N_6496,N_6683);
xor U7424 (N_7424,N_6630,N_6177);
nor U7425 (N_7425,N_6347,N_6841);
nand U7426 (N_7426,N_6418,N_6194);
xor U7427 (N_7427,N_6257,N_6104);
or U7428 (N_7428,N_6380,N_6392);
nor U7429 (N_7429,N_6613,N_6680);
or U7430 (N_7430,N_6813,N_6965);
nor U7431 (N_7431,N_6962,N_6525);
nor U7432 (N_7432,N_6476,N_6932);
xor U7433 (N_7433,N_6804,N_6230);
xnor U7434 (N_7434,N_6244,N_6757);
nor U7435 (N_7435,N_6703,N_6714);
xor U7436 (N_7436,N_6685,N_6527);
nor U7437 (N_7437,N_6627,N_6165);
nor U7438 (N_7438,N_6869,N_6578);
xnor U7439 (N_7439,N_6161,N_6950);
nor U7440 (N_7440,N_6278,N_6383);
xor U7441 (N_7441,N_6516,N_6645);
nand U7442 (N_7442,N_6250,N_6581);
nand U7443 (N_7443,N_6591,N_6317);
nor U7444 (N_7444,N_6328,N_6134);
nand U7445 (N_7445,N_6481,N_6396);
xor U7446 (N_7446,N_6751,N_6273);
and U7447 (N_7447,N_6742,N_6063);
nor U7448 (N_7448,N_6117,N_6472);
nand U7449 (N_7449,N_6839,N_6342);
and U7450 (N_7450,N_6716,N_6533);
and U7451 (N_7451,N_6395,N_6426);
or U7452 (N_7452,N_6269,N_6532);
nand U7453 (N_7453,N_6539,N_6633);
xor U7454 (N_7454,N_6759,N_6376);
xnor U7455 (N_7455,N_6262,N_6388);
nand U7456 (N_7456,N_6570,N_6691);
xor U7457 (N_7457,N_6911,N_6791);
xor U7458 (N_7458,N_6614,N_6323);
and U7459 (N_7459,N_6541,N_6192);
xor U7460 (N_7460,N_6042,N_6440);
nor U7461 (N_7461,N_6181,N_6050);
and U7462 (N_7462,N_6674,N_6106);
or U7463 (N_7463,N_6487,N_6505);
xor U7464 (N_7464,N_6854,N_6231);
or U7465 (N_7465,N_6611,N_6007);
xor U7466 (N_7466,N_6344,N_6619);
nor U7467 (N_7467,N_6786,N_6888);
or U7468 (N_7468,N_6897,N_6240);
and U7469 (N_7469,N_6923,N_6285);
and U7470 (N_7470,N_6430,N_6524);
or U7471 (N_7471,N_6306,N_6229);
xnor U7472 (N_7472,N_6538,N_6670);
and U7473 (N_7473,N_6844,N_6741);
nor U7474 (N_7474,N_6642,N_6572);
xnor U7475 (N_7475,N_6065,N_6992);
nor U7476 (N_7476,N_6827,N_6482);
or U7477 (N_7477,N_6271,N_6027);
or U7478 (N_7478,N_6184,N_6602);
or U7479 (N_7479,N_6270,N_6015);
nor U7480 (N_7480,N_6391,N_6171);
or U7481 (N_7481,N_6111,N_6949);
and U7482 (N_7482,N_6567,N_6272);
or U7483 (N_7483,N_6340,N_6646);
and U7484 (N_7484,N_6862,N_6885);
nor U7485 (N_7485,N_6191,N_6291);
and U7486 (N_7486,N_6127,N_6598);
and U7487 (N_7487,N_6947,N_6384);
xor U7488 (N_7488,N_6948,N_6753);
or U7489 (N_7489,N_6709,N_6493);
nor U7490 (N_7490,N_6735,N_6216);
or U7491 (N_7491,N_6350,N_6995);
nor U7492 (N_7492,N_6499,N_6967);
nor U7493 (N_7493,N_6774,N_6782);
and U7494 (N_7494,N_6510,N_6894);
or U7495 (N_7495,N_6411,N_6605);
or U7496 (N_7496,N_6061,N_6214);
nand U7497 (N_7497,N_6823,N_6771);
nand U7498 (N_7498,N_6896,N_6682);
and U7499 (N_7499,N_6492,N_6233);
or U7500 (N_7500,N_6807,N_6074);
and U7501 (N_7501,N_6675,N_6940);
nand U7502 (N_7502,N_6179,N_6234);
nor U7503 (N_7503,N_6657,N_6184);
nor U7504 (N_7504,N_6296,N_6461);
nor U7505 (N_7505,N_6169,N_6314);
or U7506 (N_7506,N_6011,N_6162);
and U7507 (N_7507,N_6733,N_6103);
nor U7508 (N_7508,N_6601,N_6046);
and U7509 (N_7509,N_6485,N_6879);
nand U7510 (N_7510,N_6861,N_6510);
xor U7511 (N_7511,N_6180,N_6267);
nand U7512 (N_7512,N_6299,N_6715);
xnor U7513 (N_7513,N_6715,N_6822);
nor U7514 (N_7514,N_6012,N_6266);
nor U7515 (N_7515,N_6447,N_6810);
xor U7516 (N_7516,N_6393,N_6294);
or U7517 (N_7517,N_6994,N_6579);
nor U7518 (N_7518,N_6724,N_6620);
and U7519 (N_7519,N_6517,N_6079);
nand U7520 (N_7520,N_6284,N_6583);
nand U7521 (N_7521,N_6545,N_6173);
nor U7522 (N_7522,N_6853,N_6528);
xor U7523 (N_7523,N_6671,N_6545);
nand U7524 (N_7524,N_6532,N_6488);
nand U7525 (N_7525,N_6119,N_6199);
nand U7526 (N_7526,N_6868,N_6382);
xnor U7527 (N_7527,N_6270,N_6701);
xnor U7528 (N_7528,N_6228,N_6135);
nand U7529 (N_7529,N_6381,N_6834);
and U7530 (N_7530,N_6133,N_6150);
and U7531 (N_7531,N_6667,N_6471);
and U7532 (N_7532,N_6535,N_6265);
nor U7533 (N_7533,N_6166,N_6625);
or U7534 (N_7534,N_6070,N_6241);
xor U7535 (N_7535,N_6586,N_6673);
nor U7536 (N_7536,N_6751,N_6115);
xnor U7537 (N_7537,N_6913,N_6161);
or U7538 (N_7538,N_6137,N_6466);
and U7539 (N_7539,N_6585,N_6643);
nor U7540 (N_7540,N_6975,N_6082);
or U7541 (N_7541,N_6943,N_6811);
and U7542 (N_7542,N_6216,N_6150);
nand U7543 (N_7543,N_6062,N_6183);
nand U7544 (N_7544,N_6407,N_6864);
or U7545 (N_7545,N_6877,N_6917);
and U7546 (N_7546,N_6984,N_6926);
xnor U7547 (N_7547,N_6709,N_6742);
xnor U7548 (N_7548,N_6853,N_6578);
nor U7549 (N_7549,N_6672,N_6571);
nand U7550 (N_7550,N_6931,N_6671);
xor U7551 (N_7551,N_6294,N_6905);
and U7552 (N_7552,N_6008,N_6193);
and U7553 (N_7553,N_6785,N_6260);
xor U7554 (N_7554,N_6011,N_6553);
and U7555 (N_7555,N_6971,N_6505);
or U7556 (N_7556,N_6635,N_6448);
nand U7557 (N_7557,N_6035,N_6553);
xor U7558 (N_7558,N_6103,N_6499);
and U7559 (N_7559,N_6962,N_6202);
nor U7560 (N_7560,N_6706,N_6160);
and U7561 (N_7561,N_6034,N_6479);
and U7562 (N_7562,N_6797,N_6851);
and U7563 (N_7563,N_6718,N_6676);
and U7564 (N_7564,N_6306,N_6155);
or U7565 (N_7565,N_6450,N_6624);
xor U7566 (N_7566,N_6419,N_6655);
and U7567 (N_7567,N_6921,N_6132);
or U7568 (N_7568,N_6632,N_6128);
nand U7569 (N_7569,N_6044,N_6109);
and U7570 (N_7570,N_6795,N_6972);
nand U7571 (N_7571,N_6445,N_6325);
nand U7572 (N_7572,N_6781,N_6595);
xnor U7573 (N_7573,N_6304,N_6789);
and U7574 (N_7574,N_6077,N_6823);
or U7575 (N_7575,N_6931,N_6868);
nor U7576 (N_7576,N_6825,N_6118);
xor U7577 (N_7577,N_6304,N_6595);
nand U7578 (N_7578,N_6453,N_6548);
xor U7579 (N_7579,N_6340,N_6072);
and U7580 (N_7580,N_6463,N_6393);
nand U7581 (N_7581,N_6605,N_6307);
nor U7582 (N_7582,N_6542,N_6130);
and U7583 (N_7583,N_6788,N_6979);
nand U7584 (N_7584,N_6219,N_6800);
and U7585 (N_7585,N_6350,N_6957);
or U7586 (N_7586,N_6487,N_6320);
or U7587 (N_7587,N_6546,N_6967);
xnor U7588 (N_7588,N_6165,N_6251);
xnor U7589 (N_7589,N_6537,N_6195);
xnor U7590 (N_7590,N_6476,N_6166);
or U7591 (N_7591,N_6618,N_6534);
and U7592 (N_7592,N_6332,N_6596);
nand U7593 (N_7593,N_6338,N_6399);
xor U7594 (N_7594,N_6025,N_6335);
and U7595 (N_7595,N_6091,N_6364);
or U7596 (N_7596,N_6727,N_6884);
nor U7597 (N_7597,N_6247,N_6376);
and U7598 (N_7598,N_6845,N_6333);
and U7599 (N_7599,N_6061,N_6891);
or U7600 (N_7600,N_6979,N_6846);
or U7601 (N_7601,N_6216,N_6685);
nand U7602 (N_7602,N_6627,N_6222);
and U7603 (N_7603,N_6628,N_6906);
xnor U7604 (N_7604,N_6300,N_6984);
and U7605 (N_7605,N_6105,N_6674);
nand U7606 (N_7606,N_6553,N_6359);
nand U7607 (N_7607,N_6222,N_6781);
or U7608 (N_7608,N_6021,N_6020);
xnor U7609 (N_7609,N_6321,N_6162);
or U7610 (N_7610,N_6426,N_6425);
or U7611 (N_7611,N_6145,N_6753);
nand U7612 (N_7612,N_6379,N_6337);
xnor U7613 (N_7613,N_6274,N_6676);
xor U7614 (N_7614,N_6339,N_6599);
or U7615 (N_7615,N_6570,N_6110);
nor U7616 (N_7616,N_6477,N_6762);
xor U7617 (N_7617,N_6285,N_6827);
xnor U7618 (N_7618,N_6939,N_6907);
nor U7619 (N_7619,N_6227,N_6241);
nand U7620 (N_7620,N_6182,N_6701);
xnor U7621 (N_7621,N_6771,N_6765);
xor U7622 (N_7622,N_6610,N_6315);
xor U7623 (N_7623,N_6374,N_6567);
nand U7624 (N_7624,N_6457,N_6911);
nand U7625 (N_7625,N_6808,N_6828);
nor U7626 (N_7626,N_6248,N_6716);
nor U7627 (N_7627,N_6398,N_6613);
and U7628 (N_7628,N_6213,N_6723);
xor U7629 (N_7629,N_6853,N_6754);
xor U7630 (N_7630,N_6460,N_6297);
and U7631 (N_7631,N_6241,N_6465);
or U7632 (N_7632,N_6827,N_6593);
and U7633 (N_7633,N_6876,N_6074);
nand U7634 (N_7634,N_6376,N_6920);
and U7635 (N_7635,N_6248,N_6300);
nor U7636 (N_7636,N_6969,N_6893);
or U7637 (N_7637,N_6076,N_6584);
and U7638 (N_7638,N_6980,N_6480);
and U7639 (N_7639,N_6336,N_6475);
or U7640 (N_7640,N_6005,N_6467);
xor U7641 (N_7641,N_6908,N_6935);
or U7642 (N_7642,N_6418,N_6701);
and U7643 (N_7643,N_6773,N_6643);
nand U7644 (N_7644,N_6370,N_6110);
nor U7645 (N_7645,N_6202,N_6930);
xnor U7646 (N_7646,N_6422,N_6607);
and U7647 (N_7647,N_6933,N_6598);
xor U7648 (N_7648,N_6996,N_6055);
and U7649 (N_7649,N_6406,N_6907);
or U7650 (N_7650,N_6815,N_6456);
and U7651 (N_7651,N_6099,N_6867);
xor U7652 (N_7652,N_6807,N_6784);
xnor U7653 (N_7653,N_6955,N_6276);
or U7654 (N_7654,N_6523,N_6164);
or U7655 (N_7655,N_6480,N_6697);
nand U7656 (N_7656,N_6797,N_6866);
and U7657 (N_7657,N_6316,N_6469);
xor U7658 (N_7658,N_6475,N_6201);
or U7659 (N_7659,N_6129,N_6669);
and U7660 (N_7660,N_6243,N_6498);
xor U7661 (N_7661,N_6238,N_6789);
xor U7662 (N_7662,N_6232,N_6221);
or U7663 (N_7663,N_6637,N_6257);
xor U7664 (N_7664,N_6468,N_6747);
nand U7665 (N_7665,N_6081,N_6478);
and U7666 (N_7666,N_6735,N_6725);
xnor U7667 (N_7667,N_6671,N_6412);
xor U7668 (N_7668,N_6643,N_6757);
and U7669 (N_7669,N_6775,N_6167);
nand U7670 (N_7670,N_6723,N_6211);
and U7671 (N_7671,N_6356,N_6028);
xor U7672 (N_7672,N_6115,N_6934);
nand U7673 (N_7673,N_6168,N_6552);
and U7674 (N_7674,N_6834,N_6060);
xor U7675 (N_7675,N_6813,N_6003);
or U7676 (N_7676,N_6168,N_6081);
nor U7677 (N_7677,N_6843,N_6882);
nor U7678 (N_7678,N_6683,N_6230);
xnor U7679 (N_7679,N_6255,N_6202);
nor U7680 (N_7680,N_6938,N_6308);
or U7681 (N_7681,N_6413,N_6365);
or U7682 (N_7682,N_6503,N_6204);
and U7683 (N_7683,N_6774,N_6085);
or U7684 (N_7684,N_6291,N_6549);
nor U7685 (N_7685,N_6585,N_6782);
and U7686 (N_7686,N_6169,N_6665);
xnor U7687 (N_7687,N_6782,N_6299);
xor U7688 (N_7688,N_6793,N_6801);
xnor U7689 (N_7689,N_6534,N_6200);
or U7690 (N_7690,N_6982,N_6331);
xor U7691 (N_7691,N_6314,N_6905);
or U7692 (N_7692,N_6592,N_6218);
nand U7693 (N_7693,N_6475,N_6649);
xnor U7694 (N_7694,N_6079,N_6151);
and U7695 (N_7695,N_6749,N_6697);
and U7696 (N_7696,N_6948,N_6412);
xor U7697 (N_7697,N_6847,N_6100);
xnor U7698 (N_7698,N_6470,N_6158);
nor U7699 (N_7699,N_6890,N_6498);
or U7700 (N_7700,N_6568,N_6578);
xor U7701 (N_7701,N_6691,N_6242);
xnor U7702 (N_7702,N_6284,N_6991);
nor U7703 (N_7703,N_6969,N_6895);
xor U7704 (N_7704,N_6807,N_6686);
nor U7705 (N_7705,N_6393,N_6759);
or U7706 (N_7706,N_6195,N_6822);
xor U7707 (N_7707,N_6956,N_6008);
and U7708 (N_7708,N_6838,N_6214);
xnor U7709 (N_7709,N_6087,N_6534);
nand U7710 (N_7710,N_6314,N_6758);
nor U7711 (N_7711,N_6396,N_6595);
xor U7712 (N_7712,N_6516,N_6758);
and U7713 (N_7713,N_6251,N_6269);
nor U7714 (N_7714,N_6348,N_6337);
xnor U7715 (N_7715,N_6268,N_6106);
and U7716 (N_7716,N_6451,N_6148);
or U7717 (N_7717,N_6598,N_6310);
and U7718 (N_7718,N_6764,N_6107);
nand U7719 (N_7719,N_6663,N_6063);
or U7720 (N_7720,N_6165,N_6746);
nor U7721 (N_7721,N_6946,N_6362);
or U7722 (N_7722,N_6822,N_6051);
or U7723 (N_7723,N_6656,N_6678);
and U7724 (N_7724,N_6051,N_6430);
xnor U7725 (N_7725,N_6267,N_6298);
xor U7726 (N_7726,N_6083,N_6790);
nand U7727 (N_7727,N_6271,N_6352);
nor U7728 (N_7728,N_6685,N_6783);
or U7729 (N_7729,N_6654,N_6968);
nand U7730 (N_7730,N_6939,N_6916);
xor U7731 (N_7731,N_6773,N_6075);
nand U7732 (N_7732,N_6838,N_6145);
or U7733 (N_7733,N_6215,N_6847);
xor U7734 (N_7734,N_6609,N_6453);
and U7735 (N_7735,N_6756,N_6270);
or U7736 (N_7736,N_6638,N_6360);
nor U7737 (N_7737,N_6678,N_6701);
or U7738 (N_7738,N_6712,N_6612);
nand U7739 (N_7739,N_6873,N_6823);
nand U7740 (N_7740,N_6526,N_6926);
nand U7741 (N_7741,N_6733,N_6127);
nor U7742 (N_7742,N_6800,N_6807);
or U7743 (N_7743,N_6511,N_6654);
or U7744 (N_7744,N_6830,N_6398);
nor U7745 (N_7745,N_6517,N_6676);
xor U7746 (N_7746,N_6328,N_6866);
or U7747 (N_7747,N_6451,N_6962);
or U7748 (N_7748,N_6485,N_6928);
nand U7749 (N_7749,N_6403,N_6124);
and U7750 (N_7750,N_6993,N_6920);
nand U7751 (N_7751,N_6877,N_6323);
nand U7752 (N_7752,N_6512,N_6972);
and U7753 (N_7753,N_6604,N_6388);
xor U7754 (N_7754,N_6008,N_6285);
xor U7755 (N_7755,N_6000,N_6274);
xnor U7756 (N_7756,N_6671,N_6659);
or U7757 (N_7757,N_6869,N_6720);
xor U7758 (N_7758,N_6389,N_6983);
or U7759 (N_7759,N_6445,N_6838);
nor U7760 (N_7760,N_6692,N_6824);
nor U7761 (N_7761,N_6768,N_6007);
or U7762 (N_7762,N_6487,N_6008);
xnor U7763 (N_7763,N_6062,N_6362);
nand U7764 (N_7764,N_6445,N_6289);
xor U7765 (N_7765,N_6813,N_6529);
nor U7766 (N_7766,N_6214,N_6473);
or U7767 (N_7767,N_6117,N_6103);
or U7768 (N_7768,N_6865,N_6273);
or U7769 (N_7769,N_6655,N_6615);
nand U7770 (N_7770,N_6652,N_6555);
xor U7771 (N_7771,N_6159,N_6275);
nor U7772 (N_7772,N_6913,N_6077);
nor U7773 (N_7773,N_6227,N_6554);
and U7774 (N_7774,N_6861,N_6103);
and U7775 (N_7775,N_6350,N_6440);
or U7776 (N_7776,N_6664,N_6037);
or U7777 (N_7777,N_6269,N_6000);
nand U7778 (N_7778,N_6404,N_6760);
and U7779 (N_7779,N_6698,N_6093);
or U7780 (N_7780,N_6229,N_6760);
nand U7781 (N_7781,N_6819,N_6570);
nor U7782 (N_7782,N_6604,N_6852);
xnor U7783 (N_7783,N_6473,N_6882);
and U7784 (N_7784,N_6740,N_6244);
xnor U7785 (N_7785,N_6252,N_6665);
nor U7786 (N_7786,N_6455,N_6187);
xor U7787 (N_7787,N_6731,N_6507);
nor U7788 (N_7788,N_6796,N_6056);
or U7789 (N_7789,N_6042,N_6345);
and U7790 (N_7790,N_6111,N_6410);
nand U7791 (N_7791,N_6661,N_6321);
and U7792 (N_7792,N_6086,N_6589);
nor U7793 (N_7793,N_6642,N_6963);
or U7794 (N_7794,N_6848,N_6500);
or U7795 (N_7795,N_6570,N_6251);
nand U7796 (N_7796,N_6870,N_6041);
and U7797 (N_7797,N_6761,N_6346);
or U7798 (N_7798,N_6093,N_6572);
or U7799 (N_7799,N_6734,N_6159);
xor U7800 (N_7800,N_6673,N_6110);
and U7801 (N_7801,N_6382,N_6618);
nor U7802 (N_7802,N_6826,N_6119);
xnor U7803 (N_7803,N_6619,N_6397);
or U7804 (N_7804,N_6053,N_6654);
and U7805 (N_7805,N_6890,N_6477);
xnor U7806 (N_7806,N_6702,N_6966);
nor U7807 (N_7807,N_6073,N_6327);
xor U7808 (N_7808,N_6710,N_6242);
nand U7809 (N_7809,N_6951,N_6107);
nor U7810 (N_7810,N_6123,N_6085);
xor U7811 (N_7811,N_6213,N_6227);
and U7812 (N_7812,N_6903,N_6259);
and U7813 (N_7813,N_6470,N_6299);
and U7814 (N_7814,N_6883,N_6857);
nand U7815 (N_7815,N_6886,N_6635);
xnor U7816 (N_7816,N_6526,N_6477);
nand U7817 (N_7817,N_6358,N_6627);
nor U7818 (N_7818,N_6646,N_6521);
nor U7819 (N_7819,N_6426,N_6583);
xor U7820 (N_7820,N_6844,N_6998);
nor U7821 (N_7821,N_6100,N_6482);
nor U7822 (N_7822,N_6093,N_6237);
and U7823 (N_7823,N_6415,N_6235);
nand U7824 (N_7824,N_6649,N_6890);
nand U7825 (N_7825,N_6538,N_6373);
or U7826 (N_7826,N_6059,N_6411);
or U7827 (N_7827,N_6130,N_6755);
and U7828 (N_7828,N_6394,N_6953);
nor U7829 (N_7829,N_6259,N_6543);
or U7830 (N_7830,N_6862,N_6927);
and U7831 (N_7831,N_6666,N_6109);
and U7832 (N_7832,N_6512,N_6654);
nand U7833 (N_7833,N_6885,N_6594);
nor U7834 (N_7834,N_6806,N_6558);
xor U7835 (N_7835,N_6709,N_6157);
nand U7836 (N_7836,N_6117,N_6751);
xnor U7837 (N_7837,N_6463,N_6996);
nor U7838 (N_7838,N_6291,N_6762);
nand U7839 (N_7839,N_6799,N_6600);
nor U7840 (N_7840,N_6129,N_6960);
nor U7841 (N_7841,N_6282,N_6211);
and U7842 (N_7842,N_6382,N_6051);
and U7843 (N_7843,N_6067,N_6782);
nor U7844 (N_7844,N_6791,N_6772);
xor U7845 (N_7845,N_6345,N_6041);
or U7846 (N_7846,N_6203,N_6771);
or U7847 (N_7847,N_6405,N_6402);
or U7848 (N_7848,N_6929,N_6414);
or U7849 (N_7849,N_6839,N_6800);
nor U7850 (N_7850,N_6781,N_6406);
nor U7851 (N_7851,N_6260,N_6040);
nand U7852 (N_7852,N_6274,N_6700);
or U7853 (N_7853,N_6847,N_6464);
and U7854 (N_7854,N_6744,N_6463);
xor U7855 (N_7855,N_6527,N_6706);
nand U7856 (N_7856,N_6346,N_6410);
xor U7857 (N_7857,N_6309,N_6408);
and U7858 (N_7858,N_6692,N_6554);
xor U7859 (N_7859,N_6108,N_6593);
nand U7860 (N_7860,N_6706,N_6690);
xnor U7861 (N_7861,N_6283,N_6928);
nand U7862 (N_7862,N_6096,N_6619);
xor U7863 (N_7863,N_6883,N_6572);
or U7864 (N_7864,N_6689,N_6051);
or U7865 (N_7865,N_6078,N_6030);
xnor U7866 (N_7866,N_6468,N_6974);
xnor U7867 (N_7867,N_6249,N_6191);
nor U7868 (N_7868,N_6265,N_6595);
or U7869 (N_7869,N_6712,N_6656);
xnor U7870 (N_7870,N_6121,N_6783);
xor U7871 (N_7871,N_6493,N_6664);
nand U7872 (N_7872,N_6737,N_6164);
or U7873 (N_7873,N_6575,N_6465);
xor U7874 (N_7874,N_6351,N_6712);
nor U7875 (N_7875,N_6550,N_6759);
or U7876 (N_7876,N_6693,N_6726);
nand U7877 (N_7877,N_6765,N_6525);
nand U7878 (N_7878,N_6096,N_6873);
xnor U7879 (N_7879,N_6411,N_6659);
nor U7880 (N_7880,N_6911,N_6013);
xnor U7881 (N_7881,N_6965,N_6778);
nand U7882 (N_7882,N_6352,N_6525);
nand U7883 (N_7883,N_6832,N_6779);
xnor U7884 (N_7884,N_6005,N_6339);
or U7885 (N_7885,N_6414,N_6738);
nor U7886 (N_7886,N_6968,N_6677);
xor U7887 (N_7887,N_6583,N_6011);
and U7888 (N_7888,N_6261,N_6310);
nand U7889 (N_7889,N_6038,N_6822);
or U7890 (N_7890,N_6420,N_6888);
nand U7891 (N_7891,N_6731,N_6844);
nand U7892 (N_7892,N_6888,N_6077);
nor U7893 (N_7893,N_6023,N_6081);
nor U7894 (N_7894,N_6479,N_6639);
or U7895 (N_7895,N_6498,N_6322);
nor U7896 (N_7896,N_6738,N_6017);
and U7897 (N_7897,N_6612,N_6902);
nand U7898 (N_7898,N_6415,N_6283);
nand U7899 (N_7899,N_6029,N_6725);
xnor U7900 (N_7900,N_6461,N_6795);
xor U7901 (N_7901,N_6825,N_6274);
nor U7902 (N_7902,N_6752,N_6715);
nand U7903 (N_7903,N_6286,N_6767);
xor U7904 (N_7904,N_6342,N_6966);
xnor U7905 (N_7905,N_6206,N_6136);
nand U7906 (N_7906,N_6828,N_6019);
or U7907 (N_7907,N_6731,N_6839);
and U7908 (N_7908,N_6705,N_6731);
nor U7909 (N_7909,N_6943,N_6278);
nand U7910 (N_7910,N_6888,N_6834);
xnor U7911 (N_7911,N_6189,N_6630);
nand U7912 (N_7912,N_6654,N_6296);
and U7913 (N_7913,N_6368,N_6883);
or U7914 (N_7914,N_6053,N_6569);
nand U7915 (N_7915,N_6298,N_6294);
xor U7916 (N_7916,N_6253,N_6330);
xor U7917 (N_7917,N_6693,N_6518);
nand U7918 (N_7918,N_6640,N_6875);
xnor U7919 (N_7919,N_6702,N_6221);
and U7920 (N_7920,N_6820,N_6229);
nand U7921 (N_7921,N_6560,N_6493);
nand U7922 (N_7922,N_6677,N_6159);
nor U7923 (N_7923,N_6239,N_6256);
nor U7924 (N_7924,N_6410,N_6332);
and U7925 (N_7925,N_6889,N_6715);
or U7926 (N_7926,N_6400,N_6769);
xnor U7927 (N_7927,N_6624,N_6956);
or U7928 (N_7928,N_6950,N_6655);
nor U7929 (N_7929,N_6519,N_6864);
nor U7930 (N_7930,N_6450,N_6670);
nor U7931 (N_7931,N_6190,N_6660);
or U7932 (N_7932,N_6738,N_6580);
or U7933 (N_7933,N_6859,N_6491);
xor U7934 (N_7934,N_6625,N_6616);
or U7935 (N_7935,N_6501,N_6551);
xnor U7936 (N_7936,N_6864,N_6066);
or U7937 (N_7937,N_6542,N_6076);
nor U7938 (N_7938,N_6219,N_6157);
xor U7939 (N_7939,N_6153,N_6273);
or U7940 (N_7940,N_6326,N_6655);
nor U7941 (N_7941,N_6811,N_6835);
nand U7942 (N_7942,N_6084,N_6534);
and U7943 (N_7943,N_6115,N_6547);
xnor U7944 (N_7944,N_6720,N_6864);
or U7945 (N_7945,N_6456,N_6472);
nand U7946 (N_7946,N_6480,N_6351);
xor U7947 (N_7947,N_6697,N_6082);
xor U7948 (N_7948,N_6310,N_6843);
and U7949 (N_7949,N_6499,N_6740);
and U7950 (N_7950,N_6842,N_6585);
xor U7951 (N_7951,N_6727,N_6329);
nor U7952 (N_7952,N_6223,N_6255);
xnor U7953 (N_7953,N_6304,N_6243);
xor U7954 (N_7954,N_6099,N_6462);
nand U7955 (N_7955,N_6555,N_6162);
or U7956 (N_7956,N_6687,N_6331);
nand U7957 (N_7957,N_6185,N_6652);
nor U7958 (N_7958,N_6184,N_6914);
and U7959 (N_7959,N_6987,N_6049);
nand U7960 (N_7960,N_6967,N_6733);
xnor U7961 (N_7961,N_6208,N_6413);
and U7962 (N_7962,N_6775,N_6079);
or U7963 (N_7963,N_6291,N_6879);
nor U7964 (N_7964,N_6097,N_6308);
xnor U7965 (N_7965,N_6023,N_6352);
or U7966 (N_7966,N_6024,N_6215);
nand U7967 (N_7967,N_6636,N_6865);
xnor U7968 (N_7968,N_6519,N_6863);
nand U7969 (N_7969,N_6703,N_6559);
nor U7970 (N_7970,N_6202,N_6824);
xnor U7971 (N_7971,N_6039,N_6720);
xnor U7972 (N_7972,N_6933,N_6238);
and U7973 (N_7973,N_6297,N_6452);
xor U7974 (N_7974,N_6374,N_6444);
nand U7975 (N_7975,N_6131,N_6120);
or U7976 (N_7976,N_6971,N_6782);
and U7977 (N_7977,N_6186,N_6794);
and U7978 (N_7978,N_6712,N_6653);
xor U7979 (N_7979,N_6944,N_6213);
and U7980 (N_7980,N_6185,N_6512);
and U7981 (N_7981,N_6021,N_6221);
xnor U7982 (N_7982,N_6320,N_6597);
and U7983 (N_7983,N_6062,N_6478);
xnor U7984 (N_7984,N_6101,N_6095);
nor U7985 (N_7985,N_6173,N_6314);
nand U7986 (N_7986,N_6995,N_6856);
xor U7987 (N_7987,N_6302,N_6373);
xnor U7988 (N_7988,N_6644,N_6813);
xnor U7989 (N_7989,N_6835,N_6504);
or U7990 (N_7990,N_6067,N_6028);
nor U7991 (N_7991,N_6711,N_6134);
xor U7992 (N_7992,N_6707,N_6462);
nand U7993 (N_7993,N_6843,N_6609);
nand U7994 (N_7994,N_6254,N_6614);
or U7995 (N_7995,N_6276,N_6778);
nor U7996 (N_7996,N_6964,N_6904);
and U7997 (N_7997,N_6005,N_6266);
xor U7998 (N_7998,N_6337,N_6190);
nor U7999 (N_7999,N_6021,N_6115);
nand U8000 (N_8000,N_7075,N_7328);
or U8001 (N_8001,N_7629,N_7275);
nor U8002 (N_8002,N_7253,N_7968);
nor U8003 (N_8003,N_7477,N_7585);
or U8004 (N_8004,N_7244,N_7559);
and U8005 (N_8005,N_7219,N_7911);
nor U8006 (N_8006,N_7535,N_7442);
nand U8007 (N_8007,N_7106,N_7138);
or U8008 (N_8008,N_7603,N_7386);
and U8009 (N_8009,N_7992,N_7870);
or U8010 (N_8010,N_7425,N_7670);
xnor U8011 (N_8011,N_7286,N_7861);
xnor U8012 (N_8012,N_7793,N_7375);
nor U8013 (N_8013,N_7692,N_7744);
nor U8014 (N_8014,N_7979,N_7239);
or U8015 (N_8015,N_7107,N_7536);
and U8016 (N_8016,N_7834,N_7272);
nand U8017 (N_8017,N_7767,N_7482);
nor U8018 (N_8018,N_7056,N_7925);
xor U8019 (N_8019,N_7080,N_7248);
nor U8020 (N_8020,N_7921,N_7489);
or U8021 (N_8021,N_7246,N_7616);
xnor U8022 (N_8022,N_7532,N_7418);
xor U8023 (N_8023,N_7894,N_7833);
xor U8024 (N_8024,N_7913,N_7415);
or U8025 (N_8025,N_7524,N_7513);
xnor U8026 (N_8026,N_7078,N_7654);
nor U8027 (N_8027,N_7070,N_7311);
or U8028 (N_8028,N_7020,N_7452);
xnor U8029 (N_8029,N_7416,N_7940);
nand U8030 (N_8030,N_7096,N_7684);
nor U8031 (N_8031,N_7475,N_7389);
or U8032 (N_8032,N_7326,N_7145);
xnor U8033 (N_8033,N_7666,N_7617);
xor U8034 (N_8034,N_7218,N_7486);
or U8035 (N_8035,N_7731,N_7174);
or U8036 (N_8036,N_7079,N_7976);
nor U8037 (N_8037,N_7095,N_7885);
and U8038 (N_8038,N_7234,N_7615);
or U8039 (N_8039,N_7517,N_7108);
or U8040 (N_8040,N_7050,N_7178);
xnor U8041 (N_8041,N_7689,N_7790);
nor U8042 (N_8042,N_7010,N_7072);
xnor U8043 (N_8043,N_7278,N_7928);
or U8044 (N_8044,N_7539,N_7951);
or U8045 (N_8045,N_7057,N_7573);
nand U8046 (N_8046,N_7268,N_7185);
nor U8047 (N_8047,N_7414,N_7060);
and U8048 (N_8048,N_7284,N_7969);
nor U8049 (N_8049,N_7069,N_7224);
or U8050 (N_8050,N_7267,N_7303);
or U8051 (N_8051,N_7128,N_7022);
nor U8052 (N_8052,N_7453,N_7619);
xor U8053 (N_8053,N_7454,N_7871);
or U8054 (N_8054,N_7896,N_7635);
or U8055 (N_8055,N_7848,N_7238);
xor U8056 (N_8056,N_7537,N_7953);
or U8057 (N_8057,N_7518,N_7903);
xor U8058 (N_8058,N_7351,N_7154);
and U8059 (N_8059,N_7212,N_7592);
and U8060 (N_8060,N_7726,N_7383);
xor U8061 (N_8061,N_7958,N_7538);
nor U8062 (N_8062,N_7643,N_7741);
xor U8063 (N_8063,N_7051,N_7942);
nor U8064 (N_8064,N_7710,N_7166);
nand U8065 (N_8065,N_7490,N_7352);
xor U8066 (N_8066,N_7484,N_7388);
or U8067 (N_8067,N_7739,N_7467);
or U8068 (N_8068,N_7608,N_7909);
or U8069 (N_8069,N_7024,N_7378);
or U8070 (N_8070,N_7465,N_7748);
or U8071 (N_8071,N_7498,N_7655);
and U8072 (N_8072,N_7881,N_7829);
nor U8073 (N_8073,N_7269,N_7437);
nand U8074 (N_8074,N_7485,N_7204);
and U8075 (N_8075,N_7973,N_7799);
and U8076 (N_8076,N_7402,N_7180);
or U8077 (N_8077,N_7541,N_7751);
and U8078 (N_8078,N_7952,N_7830);
and U8079 (N_8079,N_7926,N_7716);
xor U8080 (N_8080,N_7946,N_7408);
and U8081 (N_8081,N_7296,N_7674);
xnor U8082 (N_8082,N_7620,N_7657);
nor U8083 (N_8083,N_7758,N_7695);
nand U8084 (N_8084,N_7165,N_7409);
nand U8085 (N_8085,N_7314,N_7345);
xnor U8086 (N_8086,N_7583,N_7337);
and U8087 (N_8087,N_7675,N_7718);
nand U8088 (N_8088,N_7826,N_7937);
and U8089 (N_8089,N_7124,N_7175);
nand U8090 (N_8090,N_7343,N_7686);
xnor U8091 (N_8091,N_7529,N_7274);
nand U8092 (N_8092,N_7542,N_7957);
xnor U8093 (N_8093,N_7062,N_7333);
nand U8094 (N_8094,N_7419,N_7562);
and U8095 (N_8095,N_7316,N_7971);
and U8096 (N_8096,N_7836,N_7161);
xnor U8097 (N_8097,N_7797,N_7318);
nand U8098 (N_8098,N_7636,N_7281);
nand U8099 (N_8099,N_7480,N_7077);
xor U8100 (N_8100,N_7195,N_7985);
nand U8101 (N_8101,N_7801,N_7504);
or U8102 (N_8102,N_7664,N_7033);
nand U8103 (N_8103,N_7029,N_7914);
or U8104 (N_8104,N_7143,N_7198);
nand U8105 (N_8105,N_7982,N_7663);
nand U8106 (N_8106,N_7858,N_7993);
nand U8107 (N_8107,N_7099,N_7661);
nor U8108 (N_8108,N_7939,N_7354);
and U8109 (N_8109,N_7737,N_7407);
nor U8110 (N_8110,N_7427,N_7956);
nand U8111 (N_8111,N_7397,N_7713);
or U8112 (N_8112,N_7882,N_7468);
nand U8113 (N_8113,N_7508,N_7450);
nand U8114 (N_8114,N_7091,N_7420);
nor U8115 (N_8115,N_7247,N_7747);
or U8116 (N_8116,N_7040,N_7034);
and U8117 (N_8117,N_7647,N_7067);
nand U8118 (N_8118,N_7012,N_7054);
nor U8119 (N_8119,N_7900,N_7796);
and U8120 (N_8120,N_7832,N_7100);
or U8121 (N_8121,N_7152,N_7950);
and U8122 (N_8122,N_7217,N_7488);
nor U8123 (N_8123,N_7941,N_7791);
nand U8124 (N_8124,N_7544,N_7363);
nor U8125 (N_8125,N_7551,N_7089);
xnor U8126 (N_8126,N_7546,N_7644);
or U8127 (N_8127,N_7395,N_7305);
nand U8128 (N_8128,N_7111,N_7358);
xor U8129 (N_8129,N_7349,N_7736);
or U8130 (N_8130,N_7360,N_7630);
nor U8131 (N_8131,N_7340,N_7875);
or U8132 (N_8132,N_7240,N_7851);
xnor U8133 (N_8133,N_7252,N_7859);
and U8134 (N_8134,N_7413,N_7001);
or U8135 (N_8135,N_7819,N_7135);
and U8136 (N_8136,N_7039,N_7564);
nor U8137 (N_8137,N_7260,N_7197);
and U8138 (N_8138,N_7827,N_7458);
xnor U8139 (N_8139,N_7892,N_7464);
nand U8140 (N_8140,N_7313,N_7765);
nor U8141 (N_8141,N_7860,N_7373);
or U8142 (N_8142,N_7769,N_7220);
or U8143 (N_8143,N_7960,N_7552);
xor U8144 (N_8144,N_7474,N_7018);
nand U8145 (N_8145,N_7846,N_7906);
nor U8146 (N_8146,N_7129,N_7182);
nor U8147 (N_8147,N_7706,N_7639);
or U8148 (N_8148,N_7954,N_7599);
and U8149 (N_8149,N_7707,N_7582);
or U8150 (N_8150,N_7778,N_7678);
or U8151 (N_8151,N_7759,N_7614);
or U8152 (N_8152,N_7738,N_7729);
and U8153 (N_8153,N_7591,N_7379);
xnor U8154 (N_8154,N_7249,N_7377);
and U8155 (N_8155,N_7422,N_7622);
nor U8156 (N_8156,N_7624,N_7553);
nor U8157 (N_8157,N_7978,N_7865);
nor U8158 (N_8158,N_7866,N_7203);
nor U8159 (N_8159,N_7857,N_7502);
nor U8160 (N_8160,N_7510,N_7030);
nor U8161 (N_8161,N_7139,N_7642);
and U8162 (N_8162,N_7514,N_7927);
xor U8163 (N_8163,N_7365,N_7595);
xor U8164 (N_8164,N_7336,N_7816);
nor U8165 (N_8165,N_7173,N_7200);
and U8166 (N_8166,N_7507,N_7776);
nor U8167 (N_8167,N_7986,N_7496);
nor U8168 (N_8168,N_7899,N_7523);
or U8169 (N_8169,N_7476,N_7168);
nor U8170 (N_8170,N_7988,N_7715);
nand U8171 (N_8171,N_7322,N_7962);
or U8172 (N_8172,N_7053,N_7558);
and U8173 (N_8173,N_7850,N_7396);
nand U8174 (N_8174,N_7671,N_7646);
nand U8175 (N_8175,N_7821,N_7071);
and U8176 (N_8176,N_7890,N_7501);
nand U8177 (N_8177,N_7259,N_7805);
and U8178 (N_8178,N_7392,N_7688);
nand U8179 (N_8179,N_7121,N_7368);
or U8180 (N_8180,N_7136,N_7901);
nor U8181 (N_8181,N_7719,N_7785);
and U8182 (N_8182,N_7817,N_7123);
nor U8183 (N_8183,N_7183,N_7021);
or U8184 (N_8184,N_7840,N_7459);
nand U8185 (N_8185,N_7170,N_7724);
and U8186 (N_8186,N_7680,N_7932);
nor U8187 (N_8187,N_7561,N_7522);
nor U8188 (N_8188,N_7638,N_7947);
nand U8189 (N_8189,N_7237,N_7366);
and U8190 (N_8190,N_7632,N_7114);
nand U8191 (N_8191,N_7059,N_7110);
nand U8192 (N_8192,N_7245,N_7505);
xnor U8193 (N_8193,N_7933,N_7627);
or U8194 (N_8194,N_7594,N_7186);
nand U8195 (N_8195,N_7660,N_7586);
xnor U8196 (N_8196,N_7527,N_7795);
and U8197 (N_8197,N_7134,N_7261);
and U8198 (N_8198,N_7362,N_7289);
or U8199 (N_8199,N_7086,N_7783);
xor U8200 (N_8200,N_7665,N_7356);
and U8201 (N_8201,N_7478,N_7658);
and U8202 (N_8202,N_7772,N_7779);
and U8203 (N_8203,N_7271,N_7235);
xor U8204 (N_8204,N_7007,N_7633);
xnor U8205 (N_8205,N_7126,N_7216);
nor U8206 (N_8206,N_7812,N_7081);
xor U8207 (N_8207,N_7854,N_7446);
and U8208 (N_8208,N_7109,N_7566);
nand U8209 (N_8209,N_7604,N_7749);
nand U8210 (N_8210,N_7525,N_7317);
and U8211 (N_8211,N_7307,N_7436);
nor U8212 (N_8212,N_7723,N_7277);
xor U8213 (N_8213,N_7412,N_7031);
nor U8214 (N_8214,N_7456,N_7555);
nand U8215 (N_8215,N_7818,N_7290);
and U8216 (N_8216,N_7651,N_7334);
and U8217 (N_8217,N_7530,N_7387);
or U8218 (N_8218,N_7722,N_7005);
nand U8219 (N_8219,N_7043,N_7727);
and U8220 (N_8220,N_7302,N_7210);
nor U8221 (N_8221,N_7883,N_7445);
and U8222 (N_8222,N_7098,N_7983);
or U8223 (N_8223,N_7677,N_7338);
xor U8224 (N_8224,N_7872,N_7667);
and U8225 (N_8225,N_7798,N_7058);
and U8226 (N_8226,N_7920,N_7656);
nor U8227 (N_8227,N_7803,N_7308);
nand U8228 (N_8228,N_7084,N_7807);
or U8229 (N_8229,N_7082,N_7972);
nor U8230 (N_8230,N_7435,N_7970);
nor U8231 (N_8231,N_7626,N_7384);
nand U8232 (N_8232,N_7831,N_7399);
nor U8233 (N_8233,N_7980,N_7550);
and U8234 (N_8234,N_7994,N_7038);
nand U8235 (N_8235,N_7966,N_7721);
or U8236 (N_8236,N_7215,N_7009);
xnor U8237 (N_8237,N_7584,N_7487);
nor U8238 (N_8238,N_7873,N_7199);
xor U8239 (N_8239,N_7090,N_7754);
xnor U8240 (N_8240,N_7519,N_7179);
xnor U8241 (N_8241,N_7087,N_7725);
xnor U8242 (N_8242,N_7142,N_7867);
xor U8243 (N_8243,N_7967,N_7898);
or U8244 (N_8244,N_7232,N_7481);
and U8245 (N_8245,N_7493,N_7015);
nand U8246 (N_8246,N_7549,N_7406);
xnor U8247 (N_8247,N_7499,N_7843);
nor U8248 (N_8248,N_7568,N_7348);
or U8249 (N_8249,N_7405,N_7230);
xnor U8250 (N_8250,N_7611,N_7600);
nor U8251 (N_8251,N_7229,N_7227);
nor U8252 (N_8252,N_7181,N_7113);
nor U8253 (N_8253,N_7528,N_7837);
xor U8254 (N_8254,N_7746,N_7809);
nand U8255 (N_8255,N_7959,N_7006);
and U8256 (N_8256,N_7641,N_7888);
or U8257 (N_8257,N_7158,N_7516);
or U8258 (N_8258,N_7878,N_7623);
nand U8259 (N_8259,N_7662,N_7787);
nor U8260 (N_8260,N_7118,N_7576);
and U8261 (N_8261,N_7825,N_7162);
nand U8262 (N_8262,N_7382,N_7367);
xor U8263 (N_8263,N_7222,N_7441);
or U8264 (N_8264,N_7285,N_7169);
nor U8265 (N_8265,N_7699,N_7364);
xor U8266 (N_8266,N_7961,N_7208);
and U8267 (N_8267,N_7596,N_7000);
xor U8268 (N_8268,N_7391,N_7279);
xor U8269 (N_8269,N_7443,N_7140);
nand U8270 (N_8270,N_7580,N_7008);
or U8271 (N_8271,N_7672,N_7652);
xnor U8272 (N_8272,N_7880,N_7401);
or U8273 (N_8273,N_7922,N_7804);
or U8274 (N_8274,N_7097,N_7172);
xnor U8275 (N_8275,N_7984,N_7189);
and U8276 (N_8276,N_7905,N_7424);
or U8277 (N_8277,N_7262,N_7404);
and U8278 (N_8278,N_7844,N_7579);
nor U8279 (N_8279,N_7815,N_7730);
nand U8280 (N_8280,N_7841,N_7104);
or U8281 (N_8281,N_7634,N_7255);
nor U8282 (N_8282,N_7125,N_7187);
and U8283 (N_8283,N_7207,N_7293);
xor U8284 (N_8284,N_7828,N_7449);
xor U8285 (N_8285,N_7612,N_7511);
nand U8286 (N_8286,N_7254,N_7711);
nor U8287 (N_8287,N_7842,N_7701);
and U8288 (N_8288,N_7673,N_7046);
nand U8289 (N_8289,N_7241,N_7431);
nor U8290 (N_8290,N_7910,N_7534);
and U8291 (N_8291,N_7270,N_7694);
xnor U8292 (N_8292,N_7370,N_7280);
nand U8293 (N_8293,N_7775,N_7587);
or U8294 (N_8294,N_7974,N_7575);
and U8295 (N_8295,N_7588,N_7512);
nor U8296 (N_8296,N_7133,N_7495);
nand U8297 (N_8297,N_7037,N_7800);
nand U8298 (N_8298,N_7963,N_7891);
or U8299 (N_8299,N_7201,N_7202);
nand U8300 (N_8300,N_7073,N_7112);
or U8301 (N_8301,N_7155,N_7088);
xnor U8302 (N_8302,N_7410,N_7917);
nand U8303 (N_8303,N_7451,N_7417);
xor U8304 (N_8304,N_7466,N_7621);
nand U8305 (N_8305,N_7734,N_7390);
nand U8306 (N_8306,N_7810,N_7120);
and U8307 (N_8307,N_7064,N_7342);
nand U8308 (N_8308,N_7766,N_7117);
and U8309 (N_8309,N_7794,N_7889);
nand U8310 (N_8310,N_7045,N_7223);
nand U8311 (N_8311,N_7374,N_7601);
xnor U8312 (N_8312,N_7945,N_7886);
or U8313 (N_8313,N_7188,N_7026);
and U8314 (N_8314,N_7457,N_7789);
or U8315 (N_8315,N_7931,N_7225);
or U8316 (N_8316,N_7036,N_7742);
and U8317 (N_8317,N_7631,N_7915);
nand U8318 (N_8318,N_7243,N_7668);
nand U8319 (N_8319,N_7101,N_7548);
nor U8320 (N_8320,N_7565,N_7845);
nand U8321 (N_8321,N_7292,N_7792);
or U8322 (N_8322,N_7863,N_7160);
nor U8323 (N_8323,N_7304,N_7531);
xor U8324 (N_8324,N_7315,N_7572);
nor U8325 (N_8325,N_7288,N_7209);
nor U8326 (N_8326,N_7426,N_7609);
or U8327 (N_8327,N_7211,N_7017);
or U8328 (N_8328,N_7720,N_7421);
and U8329 (N_8329,N_7049,N_7753);
and U8330 (N_8330,N_7864,N_7700);
xor U8331 (N_8331,N_7042,N_7439);
nor U8332 (N_8332,N_7214,N_7773);
or U8333 (N_8333,N_7717,N_7256);
or U8334 (N_8334,N_7589,N_7003);
nor U8335 (N_8335,N_7907,N_7306);
or U8336 (N_8336,N_7690,N_7335);
nor U8337 (N_8337,N_7545,N_7132);
nor U8338 (N_8338,N_7869,N_7141);
nand U8339 (N_8339,N_7811,N_7163);
xnor U8340 (N_8340,N_7704,N_7462);
nand U8341 (N_8341,N_7990,N_7159);
nor U8342 (N_8342,N_7813,N_7618);
nand U8343 (N_8343,N_7788,N_7897);
xnor U8344 (N_8344,N_7774,N_7902);
nand U8345 (N_8345,N_7023,N_7428);
nand U8346 (N_8346,N_7273,N_7697);
nand U8347 (N_8347,N_7369,N_7471);
nor U8348 (N_8348,N_7226,N_7849);
nand U8349 (N_8349,N_7102,N_7693);
and U8350 (N_8350,N_7300,N_7838);
nor U8351 (N_8351,N_7411,N_7835);
and U8352 (N_8352,N_7743,N_7563);
nand U8353 (N_8353,N_7301,N_7784);
nand U8354 (N_8354,N_7782,N_7590);
nor U8355 (N_8355,N_7068,N_7887);
and U8356 (N_8356,N_7709,N_7578);
xnor U8357 (N_8357,N_7148,N_7332);
and U8358 (N_8358,N_7061,N_7085);
nor U8359 (N_8359,N_7287,N_7506);
nand U8360 (N_8360,N_7757,N_7176);
and U8361 (N_8361,N_7597,N_7035);
and U8362 (N_8362,N_7122,N_7761);
or U8363 (N_8363,N_7492,N_7004);
xor U8364 (N_8364,N_7503,N_7698);
or U8365 (N_8365,N_7105,N_7606);
xor U8366 (N_8366,N_7066,N_7157);
and U8367 (N_8367,N_7092,N_7093);
nor U8368 (N_8368,N_7987,N_7177);
nand U8369 (N_8369,N_7919,N_7756);
nor U8370 (N_8370,N_7802,N_7372);
nor U8371 (N_8371,N_7236,N_7310);
nand U8372 (N_8372,N_7598,N_7344);
xor U8373 (N_8373,N_7814,N_7027);
xor U8374 (N_8374,N_7242,N_7137);
and U8375 (N_8375,N_7119,N_7904);
nor U8376 (N_8376,N_7014,N_7533);
or U8377 (N_8377,N_7461,N_7312);
xor U8378 (N_8378,N_7577,N_7650);
and U8379 (N_8379,N_7607,N_7327);
or U8380 (N_8380,N_7297,N_7052);
and U8381 (N_8381,N_7771,N_7221);
nor U8382 (N_8382,N_7497,N_7679);
and U8383 (N_8383,N_7291,N_7028);
nor U8384 (N_8384,N_7329,N_7924);
nand U8385 (N_8385,N_7127,N_7824);
or U8386 (N_8386,N_7041,N_7822);
xor U8387 (N_8387,N_7380,N_7936);
xnor U8388 (N_8388,N_7044,N_7393);
and U8389 (N_8389,N_7321,N_7628);
xnor U8390 (N_8390,N_7944,N_7683);
xor U8391 (N_8391,N_7299,N_7196);
and U8392 (N_8392,N_7013,N_7320);
nor U8393 (N_8393,N_7324,N_7434);
nand U8394 (N_8394,N_7470,N_7991);
nor U8395 (N_8395,N_7032,N_7786);
and U8396 (N_8396,N_7965,N_7912);
and U8397 (N_8397,N_7923,N_7750);
xnor U8398 (N_8398,N_7687,N_7648);
xnor U8399 (N_8399,N_7948,N_7341);
nor U8400 (N_8400,N_7977,N_7076);
xor U8401 (N_8401,N_7808,N_7153);
nor U8402 (N_8402,N_7964,N_7515);
nand U8403 (N_8403,N_7862,N_7011);
nor U8404 (N_8404,N_7856,N_7649);
xnor U8405 (N_8405,N_7130,N_7055);
xor U8406 (N_8406,N_7433,N_7781);
or U8407 (N_8407,N_7521,N_7547);
nand U8408 (N_8408,N_7949,N_7463);
nand U8409 (N_8409,N_7429,N_7171);
and U8410 (N_8410,N_7653,N_7567);
nor U8411 (N_8411,N_7935,N_7876);
nor U8412 (N_8412,N_7613,N_7884);
nand U8413 (N_8413,N_7473,N_7560);
and U8414 (N_8414,N_7602,N_7194);
and U8415 (N_8415,N_7989,N_7908);
nor U8416 (N_8416,N_7479,N_7581);
nand U8417 (N_8417,N_7893,N_7371);
and U8418 (N_8418,N_7570,N_7877);
nor U8419 (N_8419,N_7571,N_7147);
xor U8420 (N_8420,N_7400,N_7150);
xor U8421 (N_8421,N_7509,N_7762);
xnor U8422 (N_8422,N_7430,N_7556);
nand U8423 (N_8423,N_7025,N_7266);
and U8424 (N_8424,N_7184,N_7852);
and U8425 (N_8425,N_7353,N_7346);
or U8426 (N_8426,N_7895,N_7676);
xnor U8427 (N_8427,N_7019,N_7156);
nand U8428 (N_8428,N_7806,N_7998);
and U8429 (N_8429,N_7361,N_7943);
xor U8430 (N_8430,N_7625,N_7447);
nor U8431 (N_8431,N_7500,N_7325);
and U8432 (N_8432,N_7712,N_7703);
and U8433 (N_8433,N_7146,N_7440);
and U8434 (N_8434,N_7659,N_7526);
xor U8435 (N_8435,N_7733,N_7997);
xnor U8436 (N_8436,N_7491,N_7282);
nand U8437 (N_8437,N_7745,N_7460);
nor U8438 (N_8438,N_7444,N_7637);
and U8439 (N_8439,N_7438,N_7191);
and U8440 (N_8440,N_7394,N_7839);
and U8441 (N_8441,N_7995,N_7640);
nor U8442 (N_8442,N_7192,N_7755);
nor U8443 (N_8443,N_7257,N_7116);
xor U8444 (N_8444,N_7131,N_7855);
nand U8445 (N_8445,N_7376,N_7853);
and U8446 (N_8446,N_7265,N_7494);
xnor U8447 (N_8447,N_7540,N_7339);
nor U8448 (N_8448,N_7151,N_7016);
or U8449 (N_8449,N_7251,N_7359);
and U8450 (N_8450,N_7263,N_7669);
nand U8451 (N_8451,N_7520,N_7103);
nand U8452 (N_8452,N_7065,N_7764);
xor U8453 (N_8453,N_7323,N_7295);
xnor U8454 (N_8454,N_7735,N_7981);
and U8455 (N_8455,N_7543,N_7728);
and U8456 (N_8456,N_7398,N_7763);
nand U8457 (N_8457,N_7708,N_7593);
or U8458 (N_8458,N_7283,N_7879);
nand U8459 (N_8459,N_7385,N_7975);
nor U8460 (N_8460,N_7206,N_7752);
or U8461 (N_8461,N_7645,N_7760);
nand U8462 (N_8462,N_7469,N_7847);
xor U8463 (N_8463,N_7298,N_7696);
xnor U8464 (N_8464,N_7823,N_7357);
or U8465 (N_8465,N_7610,N_7918);
xor U8466 (N_8466,N_7205,N_7350);
or U8467 (N_8467,N_7403,N_7002);
nor U8468 (N_8468,N_7929,N_7740);
nand U8469 (N_8469,N_7231,N_7455);
xnor U8470 (N_8470,N_7448,N_7574);
nand U8471 (N_8471,N_7294,N_7714);
or U8472 (N_8472,N_7780,N_7094);
nor U8473 (N_8473,N_7432,N_7331);
nand U8474 (N_8474,N_7355,N_7319);
nand U8475 (N_8475,N_7258,N_7554);
nand U8476 (N_8476,N_7276,N_7938);
nand U8477 (N_8477,N_7347,N_7702);
nand U8478 (N_8478,N_7472,N_7048);
or U8479 (N_8479,N_7228,N_7213);
nand U8480 (N_8480,N_7930,N_7777);
or U8481 (N_8481,N_7955,N_7557);
xnor U8482 (N_8482,N_7233,N_7770);
nor U8483 (N_8483,N_7083,N_7047);
nor U8484 (N_8484,N_7999,N_7115);
nor U8485 (N_8485,N_7063,N_7682);
or U8486 (N_8486,N_7264,N_7934);
xnor U8487 (N_8487,N_7916,N_7167);
and U8488 (N_8488,N_7996,N_7483);
or U8489 (N_8489,N_7381,N_7193);
nand U8490 (N_8490,N_7691,N_7144);
and U8491 (N_8491,N_7190,N_7685);
nand U8492 (N_8492,N_7250,N_7309);
and U8493 (N_8493,N_7164,N_7330);
xnor U8494 (N_8494,N_7149,N_7423);
and U8495 (N_8495,N_7074,N_7681);
xor U8496 (N_8496,N_7874,N_7820);
or U8497 (N_8497,N_7605,N_7569);
nor U8498 (N_8498,N_7705,N_7868);
nand U8499 (N_8499,N_7732,N_7768);
or U8500 (N_8500,N_7462,N_7016);
nand U8501 (N_8501,N_7934,N_7982);
and U8502 (N_8502,N_7418,N_7634);
nand U8503 (N_8503,N_7337,N_7022);
and U8504 (N_8504,N_7598,N_7906);
and U8505 (N_8505,N_7149,N_7858);
nor U8506 (N_8506,N_7855,N_7651);
and U8507 (N_8507,N_7913,N_7789);
and U8508 (N_8508,N_7435,N_7168);
and U8509 (N_8509,N_7426,N_7054);
or U8510 (N_8510,N_7607,N_7763);
nor U8511 (N_8511,N_7420,N_7233);
nor U8512 (N_8512,N_7321,N_7614);
nor U8513 (N_8513,N_7592,N_7700);
and U8514 (N_8514,N_7941,N_7196);
and U8515 (N_8515,N_7266,N_7534);
nor U8516 (N_8516,N_7563,N_7168);
or U8517 (N_8517,N_7237,N_7201);
nand U8518 (N_8518,N_7021,N_7612);
and U8519 (N_8519,N_7596,N_7235);
or U8520 (N_8520,N_7465,N_7547);
nand U8521 (N_8521,N_7193,N_7488);
nor U8522 (N_8522,N_7506,N_7499);
and U8523 (N_8523,N_7273,N_7381);
nand U8524 (N_8524,N_7139,N_7852);
or U8525 (N_8525,N_7239,N_7096);
xor U8526 (N_8526,N_7350,N_7127);
nand U8527 (N_8527,N_7016,N_7017);
xnor U8528 (N_8528,N_7117,N_7004);
nor U8529 (N_8529,N_7683,N_7359);
or U8530 (N_8530,N_7441,N_7531);
or U8531 (N_8531,N_7573,N_7182);
and U8532 (N_8532,N_7589,N_7324);
and U8533 (N_8533,N_7765,N_7340);
and U8534 (N_8534,N_7277,N_7801);
xnor U8535 (N_8535,N_7781,N_7191);
nand U8536 (N_8536,N_7924,N_7766);
nor U8537 (N_8537,N_7634,N_7022);
xnor U8538 (N_8538,N_7050,N_7699);
and U8539 (N_8539,N_7665,N_7399);
or U8540 (N_8540,N_7696,N_7334);
nand U8541 (N_8541,N_7719,N_7198);
nand U8542 (N_8542,N_7060,N_7966);
xor U8543 (N_8543,N_7189,N_7385);
nor U8544 (N_8544,N_7628,N_7275);
xor U8545 (N_8545,N_7724,N_7092);
nor U8546 (N_8546,N_7792,N_7937);
and U8547 (N_8547,N_7960,N_7827);
and U8548 (N_8548,N_7202,N_7462);
nand U8549 (N_8549,N_7873,N_7984);
and U8550 (N_8550,N_7423,N_7263);
nor U8551 (N_8551,N_7029,N_7516);
or U8552 (N_8552,N_7045,N_7364);
and U8553 (N_8553,N_7328,N_7448);
xor U8554 (N_8554,N_7079,N_7784);
xnor U8555 (N_8555,N_7188,N_7541);
and U8556 (N_8556,N_7870,N_7595);
nand U8557 (N_8557,N_7368,N_7983);
nor U8558 (N_8558,N_7865,N_7485);
xnor U8559 (N_8559,N_7290,N_7903);
xor U8560 (N_8560,N_7926,N_7445);
xnor U8561 (N_8561,N_7154,N_7051);
and U8562 (N_8562,N_7312,N_7606);
nor U8563 (N_8563,N_7940,N_7661);
and U8564 (N_8564,N_7645,N_7300);
nand U8565 (N_8565,N_7950,N_7880);
and U8566 (N_8566,N_7797,N_7781);
nor U8567 (N_8567,N_7468,N_7875);
or U8568 (N_8568,N_7085,N_7112);
nand U8569 (N_8569,N_7453,N_7294);
xnor U8570 (N_8570,N_7898,N_7864);
and U8571 (N_8571,N_7981,N_7214);
or U8572 (N_8572,N_7909,N_7525);
and U8573 (N_8573,N_7466,N_7487);
xor U8574 (N_8574,N_7441,N_7978);
nor U8575 (N_8575,N_7434,N_7023);
xor U8576 (N_8576,N_7544,N_7812);
and U8577 (N_8577,N_7983,N_7234);
xnor U8578 (N_8578,N_7092,N_7243);
xnor U8579 (N_8579,N_7076,N_7392);
nor U8580 (N_8580,N_7946,N_7691);
nor U8581 (N_8581,N_7323,N_7205);
and U8582 (N_8582,N_7225,N_7835);
nand U8583 (N_8583,N_7854,N_7635);
nor U8584 (N_8584,N_7035,N_7465);
nand U8585 (N_8585,N_7194,N_7003);
nor U8586 (N_8586,N_7159,N_7689);
or U8587 (N_8587,N_7522,N_7874);
and U8588 (N_8588,N_7129,N_7030);
or U8589 (N_8589,N_7694,N_7102);
or U8590 (N_8590,N_7496,N_7661);
xnor U8591 (N_8591,N_7759,N_7398);
xnor U8592 (N_8592,N_7898,N_7074);
nor U8593 (N_8593,N_7203,N_7737);
nor U8594 (N_8594,N_7678,N_7181);
nand U8595 (N_8595,N_7115,N_7626);
or U8596 (N_8596,N_7250,N_7016);
nor U8597 (N_8597,N_7662,N_7762);
nor U8598 (N_8598,N_7719,N_7376);
nand U8599 (N_8599,N_7451,N_7980);
xnor U8600 (N_8600,N_7716,N_7063);
xnor U8601 (N_8601,N_7596,N_7739);
nand U8602 (N_8602,N_7870,N_7773);
or U8603 (N_8603,N_7921,N_7588);
or U8604 (N_8604,N_7498,N_7376);
or U8605 (N_8605,N_7554,N_7876);
and U8606 (N_8606,N_7662,N_7193);
xor U8607 (N_8607,N_7017,N_7571);
or U8608 (N_8608,N_7400,N_7732);
and U8609 (N_8609,N_7954,N_7423);
nor U8610 (N_8610,N_7258,N_7007);
or U8611 (N_8611,N_7560,N_7159);
xor U8612 (N_8612,N_7473,N_7637);
and U8613 (N_8613,N_7453,N_7522);
nor U8614 (N_8614,N_7710,N_7953);
or U8615 (N_8615,N_7359,N_7111);
or U8616 (N_8616,N_7617,N_7622);
xnor U8617 (N_8617,N_7035,N_7903);
xor U8618 (N_8618,N_7676,N_7962);
and U8619 (N_8619,N_7052,N_7338);
and U8620 (N_8620,N_7002,N_7605);
or U8621 (N_8621,N_7910,N_7412);
xnor U8622 (N_8622,N_7861,N_7390);
nand U8623 (N_8623,N_7742,N_7959);
nand U8624 (N_8624,N_7816,N_7815);
xnor U8625 (N_8625,N_7961,N_7182);
xnor U8626 (N_8626,N_7871,N_7730);
nand U8627 (N_8627,N_7750,N_7588);
nor U8628 (N_8628,N_7995,N_7528);
and U8629 (N_8629,N_7215,N_7537);
xor U8630 (N_8630,N_7694,N_7550);
xnor U8631 (N_8631,N_7051,N_7395);
xor U8632 (N_8632,N_7896,N_7351);
or U8633 (N_8633,N_7870,N_7986);
nand U8634 (N_8634,N_7338,N_7144);
xnor U8635 (N_8635,N_7137,N_7064);
or U8636 (N_8636,N_7777,N_7538);
or U8637 (N_8637,N_7116,N_7606);
xnor U8638 (N_8638,N_7014,N_7462);
or U8639 (N_8639,N_7780,N_7983);
or U8640 (N_8640,N_7062,N_7745);
nor U8641 (N_8641,N_7142,N_7271);
nor U8642 (N_8642,N_7054,N_7253);
xnor U8643 (N_8643,N_7921,N_7923);
or U8644 (N_8644,N_7648,N_7495);
and U8645 (N_8645,N_7008,N_7867);
xnor U8646 (N_8646,N_7819,N_7290);
xnor U8647 (N_8647,N_7654,N_7107);
and U8648 (N_8648,N_7266,N_7359);
nand U8649 (N_8649,N_7523,N_7160);
or U8650 (N_8650,N_7061,N_7739);
nand U8651 (N_8651,N_7206,N_7078);
xnor U8652 (N_8652,N_7315,N_7012);
or U8653 (N_8653,N_7246,N_7904);
or U8654 (N_8654,N_7025,N_7589);
xor U8655 (N_8655,N_7117,N_7086);
xor U8656 (N_8656,N_7336,N_7692);
or U8657 (N_8657,N_7259,N_7495);
and U8658 (N_8658,N_7868,N_7933);
nor U8659 (N_8659,N_7395,N_7753);
or U8660 (N_8660,N_7869,N_7892);
and U8661 (N_8661,N_7605,N_7595);
or U8662 (N_8662,N_7039,N_7109);
xnor U8663 (N_8663,N_7325,N_7415);
nor U8664 (N_8664,N_7295,N_7740);
xnor U8665 (N_8665,N_7919,N_7315);
nor U8666 (N_8666,N_7240,N_7884);
xnor U8667 (N_8667,N_7939,N_7807);
and U8668 (N_8668,N_7092,N_7438);
xor U8669 (N_8669,N_7797,N_7304);
nand U8670 (N_8670,N_7138,N_7434);
xor U8671 (N_8671,N_7809,N_7485);
nor U8672 (N_8672,N_7127,N_7603);
and U8673 (N_8673,N_7590,N_7325);
nand U8674 (N_8674,N_7057,N_7728);
and U8675 (N_8675,N_7716,N_7310);
nor U8676 (N_8676,N_7097,N_7656);
nor U8677 (N_8677,N_7318,N_7122);
and U8678 (N_8678,N_7030,N_7020);
and U8679 (N_8679,N_7501,N_7140);
xnor U8680 (N_8680,N_7818,N_7825);
or U8681 (N_8681,N_7360,N_7982);
xnor U8682 (N_8682,N_7562,N_7561);
nand U8683 (N_8683,N_7383,N_7672);
xnor U8684 (N_8684,N_7457,N_7682);
or U8685 (N_8685,N_7664,N_7547);
nand U8686 (N_8686,N_7334,N_7949);
and U8687 (N_8687,N_7033,N_7440);
and U8688 (N_8688,N_7400,N_7124);
or U8689 (N_8689,N_7793,N_7786);
nand U8690 (N_8690,N_7141,N_7143);
xnor U8691 (N_8691,N_7241,N_7769);
or U8692 (N_8692,N_7526,N_7960);
nor U8693 (N_8693,N_7066,N_7487);
nand U8694 (N_8694,N_7332,N_7998);
or U8695 (N_8695,N_7866,N_7124);
xor U8696 (N_8696,N_7464,N_7266);
and U8697 (N_8697,N_7497,N_7849);
nand U8698 (N_8698,N_7232,N_7078);
and U8699 (N_8699,N_7644,N_7044);
nand U8700 (N_8700,N_7476,N_7327);
or U8701 (N_8701,N_7772,N_7403);
nor U8702 (N_8702,N_7912,N_7453);
nand U8703 (N_8703,N_7826,N_7426);
or U8704 (N_8704,N_7605,N_7536);
nor U8705 (N_8705,N_7831,N_7342);
nand U8706 (N_8706,N_7714,N_7355);
xor U8707 (N_8707,N_7950,N_7278);
nand U8708 (N_8708,N_7246,N_7707);
and U8709 (N_8709,N_7094,N_7855);
or U8710 (N_8710,N_7397,N_7715);
or U8711 (N_8711,N_7724,N_7927);
or U8712 (N_8712,N_7587,N_7469);
xnor U8713 (N_8713,N_7526,N_7066);
nor U8714 (N_8714,N_7458,N_7810);
and U8715 (N_8715,N_7961,N_7344);
or U8716 (N_8716,N_7512,N_7777);
nand U8717 (N_8717,N_7050,N_7924);
xnor U8718 (N_8718,N_7178,N_7815);
nor U8719 (N_8719,N_7897,N_7893);
or U8720 (N_8720,N_7081,N_7490);
nand U8721 (N_8721,N_7534,N_7442);
nand U8722 (N_8722,N_7900,N_7193);
nand U8723 (N_8723,N_7523,N_7710);
xnor U8724 (N_8724,N_7566,N_7121);
and U8725 (N_8725,N_7049,N_7052);
nor U8726 (N_8726,N_7165,N_7955);
or U8727 (N_8727,N_7723,N_7865);
nand U8728 (N_8728,N_7653,N_7818);
and U8729 (N_8729,N_7115,N_7198);
nand U8730 (N_8730,N_7713,N_7180);
and U8731 (N_8731,N_7607,N_7317);
or U8732 (N_8732,N_7772,N_7523);
and U8733 (N_8733,N_7077,N_7498);
or U8734 (N_8734,N_7800,N_7660);
or U8735 (N_8735,N_7063,N_7880);
nor U8736 (N_8736,N_7405,N_7603);
or U8737 (N_8737,N_7939,N_7593);
and U8738 (N_8738,N_7571,N_7927);
and U8739 (N_8739,N_7078,N_7774);
nor U8740 (N_8740,N_7353,N_7418);
xor U8741 (N_8741,N_7325,N_7266);
nor U8742 (N_8742,N_7852,N_7576);
nand U8743 (N_8743,N_7571,N_7363);
xnor U8744 (N_8744,N_7531,N_7549);
nor U8745 (N_8745,N_7769,N_7046);
nand U8746 (N_8746,N_7748,N_7078);
nor U8747 (N_8747,N_7459,N_7061);
nor U8748 (N_8748,N_7960,N_7841);
nor U8749 (N_8749,N_7303,N_7128);
nor U8750 (N_8750,N_7934,N_7654);
and U8751 (N_8751,N_7386,N_7829);
nand U8752 (N_8752,N_7876,N_7670);
xor U8753 (N_8753,N_7835,N_7735);
nor U8754 (N_8754,N_7912,N_7589);
nor U8755 (N_8755,N_7407,N_7551);
nor U8756 (N_8756,N_7901,N_7208);
nand U8757 (N_8757,N_7806,N_7501);
nor U8758 (N_8758,N_7105,N_7203);
nor U8759 (N_8759,N_7499,N_7037);
xnor U8760 (N_8760,N_7375,N_7022);
xnor U8761 (N_8761,N_7866,N_7093);
nor U8762 (N_8762,N_7124,N_7021);
xnor U8763 (N_8763,N_7449,N_7685);
nor U8764 (N_8764,N_7286,N_7476);
nor U8765 (N_8765,N_7771,N_7241);
nand U8766 (N_8766,N_7609,N_7920);
nor U8767 (N_8767,N_7752,N_7775);
and U8768 (N_8768,N_7506,N_7257);
and U8769 (N_8769,N_7944,N_7266);
xor U8770 (N_8770,N_7228,N_7638);
nor U8771 (N_8771,N_7904,N_7641);
nand U8772 (N_8772,N_7522,N_7083);
or U8773 (N_8773,N_7489,N_7420);
xnor U8774 (N_8774,N_7736,N_7234);
nor U8775 (N_8775,N_7255,N_7090);
nor U8776 (N_8776,N_7711,N_7640);
or U8777 (N_8777,N_7351,N_7137);
xnor U8778 (N_8778,N_7016,N_7348);
and U8779 (N_8779,N_7752,N_7350);
and U8780 (N_8780,N_7428,N_7369);
nand U8781 (N_8781,N_7788,N_7427);
xor U8782 (N_8782,N_7146,N_7391);
or U8783 (N_8783,N_7077,N_7135);
xor U8784 (N_8784,N_7608,N_7146);
nand U8785 (N_8785,N_7569,N_7382);
nor U8786 (N_8786,N_7685,N_7045);
nor U8787 (N_8787,N_7320,N_7006);
nor U8788 (N_8788,N_7997,N_7893);
nor U8789 (N_8789,N_7004,N_7116);
nand U8790 (N_8790,N_7773,N_7638);
or U8791 (N_8791,N_7911,N_7446);
or U8792 (N_8792,N_7561,N_7926);
and U8793 (N_8793,N_7155,N_7255);
and U8794 (N_8794,N_7214,N_7975);
or U8795 (N_8795,N_7876,N_7564);
or U8796 (N_8796,N_7582,N_7759);
nor U8797 (N_8797,N_7107,N_7590);
nand U8798 (N_8798,N_7416,N_7316);
nand U8799 (N_8799,N_7805,N_7084);
xnor U8800 (N_8800,N_7517,N_7037);
xnor U8801 (N_8801,N_7848,N_7028);
xnor U8802 (N_8802,N_7865,N_7966);
nand U8803 (N_8803,N_7304,N_7318);
and U8804 (N_8804,N_7912,N_7406);
nor U8805 (N_8805,N_7509,N_7465);
nor U8806 (N_8806,N_7089,N_7115);
nand U8807 (N_8807,N_7551,N_7093);
nor U8808 (N_8808,N_7098,N_7752);
nand U8809 (N_8809,N_7582,N_7300);
nor U8810 (N_8810,N_7498,N_7956);
and U8811 (N_8811,N_7818,N_7204);
xor U8812 (N_8812,N_7033,N_7773);
nor U8813 (N_8813,N_7087,N_7954);
nor U8814 (N_8814,N_7401,N_7775);
or U8815 (N_8815,N_7948,N_7807);
and U8816 (N_8816,N_7378,N_7016);
or U8817 (N_8817,N_7387,N_7785);
xnor U8818 (N_8818,N_7737,N_7977);
nand U8819 (N_8819,N_7651,N_7445);
and U8820 (N_8820,N_7928,N_7160);
or U8821 (N_8821,N_7323,N_7791);
and U8822 (N_8822,N_7200,N_7825);
nand U8823 (N_8823,N_7804,N_7571);
nand U8824 (N_8824,N_7680,N_7496);
or U8825 (N_8825,N_7965,N_7843);
xnor U8826 (N_8826,N_7664,N_7565);
and U8827 (N_8827,N_7881,N_7297);
nand U8828 (N_8828,N_7424,N_7725);
nand U8829 (N_8829,N_7541,N_7756);
nand U8830 (N_8830,N_7077,N_7921);
nand U8831 (N_8831,N_7125,N_7580);
and U8832 (N_8832,N_7015,N_7531);
or U8833 (N_8833,N_7049,N_7614);
nor U8834 (N_8834,N_7370,N_7770);
or U8835 (N_8835,N_7099,N_7995);
and U8836 (N_8836,N_7503,N_7181);
nor U8837 (N_8837,N_7306,N_7584);
nor U8838 (N_8838,N_7186,N_7603);
and U8839 (N_8839,N_7312,N_7218);
and U8840 (N_8840,N_7124,N_7861);
nand U8841 (N_8841,N_7559,N_7714);
nor U8842 (N_8842,N_7668,N_7203);
xor U8843 (N_8843,N_7865,N_7764);
nand U8844 (N_8844,N_7864,N_7107);
nor U8845 (N_8845,N_7698,N_7847);
or U8846 (N_8846,N_7020,N_7384);
and U8847 (N_8847,N_7059,N_7237);
nand U8848 (N_8848,N_7164,N_7573);
nor U8849 (N_8849,N_7033,N_7678);
and U8850 (N_8850,N_7256,N_7388);
xor U8851 (N_8851,N_7964,N_7231);
nand U8852 (N_8852,N_7756,N_7885);
or U8853 (N_8853,N_7921,N_7421);
or U8854 (N_8854,N_7995,N_7719);
or U8855 (N_8855,N_7321,N_7329);
nand U8856 (N_8856,N_7687,N_7545);
and U8857 (N_8857,N_7090,N_7349);
and U8858 (N_8858,N_7432,N_7165);
nor U8859 (N_8859,N_7883,N_7421);
xnor U8860 (N_8860,N_7471,N_7144);
xnor U8861 (N_8861,N_7561,N_7787);
nand U8862 (N_8862,N_7640,N_7291);
xor U8863 (N_8863,N_7918,N_7632);
nand U8864 (N_8864,N_7123,N_7187);
or U8865 (N_8865,N_7173,N_7607);
nand U8866 (N_8866,N_7580,N_7052);
or U8867 (N_8867,N_7822,N_7085);
and U8868 (N_8868,N_7060,N_7194);
nor U8869 (N_8869,N_7155,N_7753);
and U8870 (N_8870,N_7779,N_7281);
and U8871 (N_8871,N_7042,N_7138);
nand U8872 (N_8872,N_7236,N_7328);
nor U8873 (N_8873,N_7979,N_7615);
and U8874 (N_8874,N_7219,N_7591);
and U8875 (N_8875,N_7309,N_7061);
or U8876 (N_8876,N_7468,N_7490);
and U8877 (N_8877,N_7726,N_7598);
xnor U8878 (N_8878,N_7715,N_7486);
nor U8879 (N_8879,N_7615,N_7656);
xnor U8880 (N_8880,N_7401,N_7598);
nand U8881 (N_8881,N_7052,N_7206);
or U8882 (N_8882,N_7961,N_7459);
or U8883 (N_8883,N_7574,N_7052);
nand U8884 (N_8884,N_7585,N_7757);
nand U8885 (N_8885,N_7596,N_7793);
or U8886 (N_8886,N_7130,N_7519);
or U8887 (N_8887,N_7092,N_7844);
nor U8888 (N_8888,N_7265,N_7423);
nor U8889 (N_8889,N_7884,N_7388);
and U8890 (N_8890,N_7925,N_7064);
or U8891 (N_8891,N_7043,N_7014);
nor U8892 (N_8892,N_7177,N_7653);
and U8893 (N_8893,N_7878,N_7012);
nand U8894 (N_8894,N_7125,N_7582);
or U8895 (N_8895,N_7407,N_7499);
nand U8896 (N_8896,N_7310,N_7063);
xnor U8897 (N_8897,N_7697,N_7558);
and U8898 (N_8898,N_7503,N_7379);
nor U8899 (N_8899,N_7271,N_7619);
or U8900 (N_8900,N_7593,N_7888);
xor U8901 (N_8901,N_7111,N_7844);
xnor U8902 (N_8902,N_7542,N_7267);
nor U8903 (N_8903,N_7456,N_7070);
or U8904 (N_8904,N_7950,N_7928);
xnor U8905 (N_8905,N_7561,N_7978);
nor U8906 (N_8906,N_7189,N_7248);
nand U8907 (N_8907,N_7912,N_7103);
xnor U8908 (N_8908,N_7250,N_7428);
and U8909 (N_8909,N_7730,N_7758);
and U8910 (N_8910,N_7569,N_7099);
nand U8911 (N_8911,N_7143,N_7897);
nor U8912 (N_8912,N_7787,N_7962);
xnor U8913 (N_8913,N_7202,N_7081);
nor U8914 (N_8914,N_7727,N_7856);
nand U8915 (N_8915,N_7974,N_7019);
nor U8916 (N_8916,N_7834,N_7593);
nor U8917 (N_8917,N_7769,N_7943);
or U8918 (N_8918,N_7099,N_7391);
xor U8919 (N_8919,N_7351,N_7970);
and U8920 (N_8920,N_7148,N_7550);
and U8921 (N_8921,N_7694,N_7571);
nor U8922 (N_8922,N_7902,N_7705);
and U8923 (N_8923,N_7414,N_7590);
nand U8924 (N_8924,N_7913,N_7983);
xor U8925 (N_8925,N_7663,N_7437);
nand U8926 (N_8926,N_7118,N_7790);
and U8927 (N_8927,N_7772,N_7977);
and U8928 (N_8928,N_7972,N_7099);
and U8929 (N_8929,N_7807,N_7042);
nand U8930 (N_8930,N_7702,N_7739);
nor U8931 (N_8931,N_7262,N_7975);
and U8932 (N_8932,N_7786,N_7043);
xnor U8933 (N_8933,N_7106,N_7934);
and U8934 (N_8934,N_7173,N_7450);
xor U8935 (N_8935,N_7105,N_7614);
nor U8936 (N_8936,N_7899,N_7159);
nor U8937 (N_8937,N_7018,N_7143);
nor U8938 (N_8938,N_7796,N_7603);
nor U8939 (N_8939,N_7842,N_7969);
nor U8940 (N_8940,N_7902,N_7613);
nand U8941 (N_8941,N_7591,N_7895);
and U8942 (N_8942,N_7296,N_7136);
and U8943 (N_8943,N_7630,N_7378);
xor U8944 (N_8944,N_7359,N_7992);
and U8945 (N_8945,N_7354,N_7611);
nand U8946 (N_8946,N_7499,N_7712);
xor U8947 (N_8947,N_7801,N_7939);
or U8948 (N_8948,N_7577,N_7957);
or U8949 (N_8949,N_7872,N_7633);
nor U8950 (N_8950,N_7590,N_7020);
or U8951 (N_8951,N_7227,N_7258);
xnor U8952 (N_8952,N_7046,N_7566);
nor U8953 (N_8953,N_7713,N_7491);
and U8954 (N_8954,N_7479,N_7257);
or U8955 (N_8955,N_7977,N_7696);
nor U8956 (N_8956,N_7699,N_7533);
nand U8957 (N_8957,N_7265,N_7477);
nor U8958 (N_8958,N_7571,N_7469);
xor U8959 (N_8959,N_7951,N_7691);
nand U8960 (N_8960,N_7698,N_7712);
xnor U8961 (N_8961,N_7274,N_7533);
xor U8962 (N_8962,N_7223,N_7404);
nor U8963 (N_8963,N_7522,N_7040);
xnor U8964 (N_8964,N_7481,N_7476);
and U8965 (N_8965,N_7675,N_7372);
xor U8966 (N_8966,N_7818,N_7392);
nor U8967 (N_8967,N_7189,N_7834);
nor U8968 (N_8968,N_7033,N_7363);
nand U8969 (N_8969,N_7478,N_7670);
and U8970 (N_8970,N_7227,N_7148);
nand U8971 (N_8971,N_7037,N_7956);
and U8972 (N_8972,N_7679,N_7522);
nor U8973 (N_8973,N_7260,N_7934);
xor U8974 (N_8974,N_7189,N_7943);
nor U8975 (N_8975,N_7367,N_7547);
or U8976 (N_8976,N_7653,N_7878);
nor U8977 (N_8977,N_7043,N_7478);
or U8978 (N_8978,N_7213,N_7878);
nor U8979 (N_8979,N_7488,N_7594);
nand U8980 (N_8980,N_7787,N_7578);
or U8981 (N_8981,N_7063,N_7935);
nand U8982 (N_8982,N_7996,N_7295);
xor U8983 (N_8983,N_7844,N_7240);
nand U8984 (N_8984,N_7522,N_7892);
xnor U8985 (N_8985,N_7885,N_7495);
nand U8986 (N_8986,N_7993,N_7589);
or U8987 (N_8987,N_7179,N_7293);
nor U8988 (N_8988,N_7535,N_7208);
or U8989 (N_8989,N_7117,N_7298);
nand U8990 (N_8990,N_7872,N_7723);
xor U8991 (N_8991,N_7213,N_7165);
nor U8992 (N_8992,N_7345,N_7394);
nor U8993 (N_8993,N_7691,N_7155);
and U8994 (N_8994,N_7233,N_7342);
and U8995 (N_8995,N_7689,N_7493);
nor U8996 (N_8996,N_7093,N_7780);
xnor U8997 (N_8997,N_7719,N_7799);
or U8998 (N_8998,N_7353,N_7277);
xor U8999 (N_8999,N_7219,N_7899);
nor U9000 (N_9000,N_8478,N_8028);
or U9001 (N_9001,N_8457,N_8200);
or U9002 (N_9002,N_8448,N_8105);
or U9003 (N_9003,N_8760,N_8694);
and U9004 (N_9004,N_8249,N_8787);
xnor U9005 (N_9005,N_8469,N_8503);
nand U9006 (N_9006,N_8012,N_8711);
nor U9007 (N_9007,N_8312,N_8133);
xor U9008 (N_9008,N_8776,N_8464);
xnor U9009 (N_9009,N_8961,N_8553);
or U9010 (N_9010,N_8538,N_8391);
nor U9011 (N_9011,N_8686,N_8543);
nor U9012 (N_9012,N_8955,N_8534);
xnor U9013 (N_9013,N_8284,N_8832);
or U9014 (N_9014,N_8178,N_8299);
or U9015 (N_9015,N_8705,N_8993);
nand U9016 (N_9016,N_8870,N_8680);
xor U9017 (N_9017,N_8821,N_8468);
xnor U9018 (N_9018,N_8096,N_8772);
nand U9019 (N_9019,N_8229,N_8631);
nand U9020 (N_9020,N_8412,N_8640);
nor U9021 (N_9021,N_8591,N_8514);
or U9022 (N_9022,N_8668,N_8794);
xnor U9023 (N_9023,N_8283,N_8988);
nor U9024 (N_9024,N_8084,N_8564);
or U9025 (N_9025,N_8806,N_8756);
nor U9026 (N_9026,N_8195,N_8098);
and U9027 (N_9027,N_8739,N_8318);
or U9028 (N_9028,N_8052,N_8279);
nor U9029 (N_9029,N_8759,N_8777);
nor U9030 (N_9030,N_8629,N_8292);
or U9031 (N_9031,N_8859,N_8966);
and U9032 (N_9032,N_8264,N_8723);
xnor U9033 (N_9033,N_8823,N_8928);
or U9034 (N_9034,N_8883,N_8311);
xor U9035 (N_9035,N_8519,N_8903);
xor U9036 (N_9036,N_8344,N_8143);
nor U9037 (N_9037,N_8878,N_8490);
or U9038 (N_9038,N_8493,N_8377);
nor U9039 (N_9039,N_8453,N_8313);
nor U9040 (N_9040,N_8471,N_8071);
nand U9041 (N_9041,N_8994,N_8511);
xnor U9042 (N_9042,N_8207,N_8697);
nor U9043 (N_9043,N_8527,N_8358);
nor U9044 (N_9044,N_8745,N_8325);
or U9045 (N_9045,N_8150,N_8803);
xor U9046 (N_9046,N_8065,N_8274);
nor U9047 (N_9047,N_8288,N_8792);
nor U9048 (N_9048,N_8417,N_8039);
nand U9049 (N_9049,N_8350,N_8339);
nor U9050 (N_9050,N_8376,N_8996);
nor U9051 (N_9051,N_8450,N_8671);
nand U9052 (N_9052,N_8634,N_8428);
nand U9053 (N_9053,N_8060,N_8969);
nor U9054 (N_9054,N_8851,N_8778);
nand U9055 (N_9055,N_8086,N_8338);
or U9056 (N_9056,N_8191,N_8384);
nor U9057 (N_9057,N_8819,N_8854);
xnor U9058 (N_9058,N_8702,N_8751);
xnor U9059 (N_9059,N_8943,N_8425);
or U9060 (N_9060,N_8517,N_8183);
nor U9061 (N_9061,N_8965,N_8773);
xnor U9062 (N_9062,N_8922,N_8612);
or U9063 (N_9063,N_8542,N_8979);
nand U9064 (N_9064,N_8816,N_8923);
nor U9065 (N_9065,N_8132,N_8390);
nor U9066 (N_9066,N_8822,N_8306);
and U9067 (N_9067,N_8622,N_8891);
nor U9068 (N_9068,N_8092,N_8704);
nand U9069 (N_9069,N_8246,N_8151);
nand U9070 (N_9070,N_8693,N_8364);
or U9071 (N_9071,N_8407,N_8103);
nor U9072 (N_9072,N_8186,N_8304);
xor U9073 (N_9073,N_8985,N_8775);
and U9074 (N_9074,N_8930,N_8418);
and U9075 (N_9075,N_8203,N_8477);
or U9076 (N_9076,N_8952,N_8333);
or U9077 (N_9077,N_8341,N_8526);
and U9078 (N_9078,N_8245,N_8633);
xor U9079 (N_9079,N_8408,N_8995);
or U9080 (N_9080,N_8545,N_8804);
nor U9081 (N_9081,N_8653,N_8649);
or U9082 (N_9082,N_8992,N_8427);
nor U9083 (N_9083,N_8958,N_8608);
and U9084 (N_9084,N_8076,N_8467);
nand U9085 (N_9085,N_8416,N_8480);
or U9086 (N_9086,N_8244,N_8395);
xor U9087 (N_9087,N_8434,N_8415);
or U9088 (N_9088,N_8379,N_8632);
xor U9089 (N_9089,N_8546,N_8072);
or U9090 (N_9090,N_8647,N_8555);
or U9091 (N_9091,N_8253,N_8691);
nor U9092 (N_9092,N_8316,N_8826);
xor U9093 (N_9093,N_8446,N_8662);
xor U9094 (N_9094,N_8894,N_8753);
nand U9095 (N_9095,N_8242,N_8815);
and U9096 (N_9096,N_8199,N_8127);
nor U9097 (N_9097,N_8025,N_8232);
xnor U9098 (N_9098,N_8366,N_8795);
nand U9099 (N_9099,N_8948,N_8205);
nor U9100 (N_9100,N_8524,N_8860);
or U9101 (N_9101,N_8607,N_8830);
or U9102 (N_9102,N_8682,N_8677);
nand U9103 (N_9103,N_8611,N_8257);
xor U9104 (N_9104,N_8474,N_8675);
or U9105 (N_9105,N_8699,N_8411);
nand U9106 (N_9106,N_8053,N_8362);
nand U9107 (N_9107,N_8315,N_8125);
or U9108 (N_9108,N_8650,N_8241);
or U9109 (N_9109,N_8354,N_8398);
or U9110 (N_9110,N_8042,N_8939);
nand U9111 (N_9111,N_8101,N_8626);
xor U9112 (N_9112,N_8004,N_8472);
and U9113 (N_9113,N_8569,N_8820);
or U9114 (N_9114,N_8655,N_8637);
or U9115 (N_9115,N_8960,N_8858);
or U9116 (N_9116,N_8134,N_8404);
or U9117 (N_9117,N_8018,N_8678);
nor U9118 (N_9118,N_8485,N_8188);
nand U9119 (N_9119,N_8309,N_8214);
xnor U9120 (N_9120,N_8443,N_8347);
or U9121 (N_9121,N_8173,N_8145);
nand U9122 (N_9122,N_8095,N_8920);
xnor U9123 (N_9123,N_8642,N_8837);
or U9124 (N_9124,N_8862,N_8849);
nor U9125 (N_9125,N_8610,N_8159);
xnor U9126 (N_9126,N_8267,N_8005);
nand U9127 (N_9127,N_8951,N_8378);
nand U9128 (N_9128,N_8077,N_8964);
and U9129 (N_9129,N_8360,N_8314);
xnor U9130 (N_9130,N_8152,N_8209);
xor U9131 (N_9131,N_8281,N_8556);
or U9132 (N_9132,N_8067,N_8164);
nand U9133 (N_9133,N_8847,N_8954);
xor U9134 (N_9134,N_8196,N_8409);
and U9135 (N_9135,N_8630,N_8603);
xnor U9136 (N_9136,N_8654,N_8153);
xor U9137 (N_9137,N_8783,N_8268);
nor U9138 (N_9138,N_8648,N_8031);
and U9139 (N_9139,N_8117,N_8400);
xor U9140 (N_9140,N_8158,N_8522);
nand U9141 (N_9141,N_8373,N_8447);
nor U9142 (N_9142,N_8997,N_8334);
xor U9143 (N_9143,N_8836,N_8540);
or U9144 (N_9144,N_8547,N_8405);
and U9145 (N_9145,N_8124,N_8714);
or U9146 (N_9146,N_8601,N_8710);
and U9147 (N_9147,N_8614,N_8352);
nor U9148 (N_9148,N_8827,N_8104);
nor U9149 (N_9149,N_8029,N_8303);
nor U9150 (N_9150,N_8768,N_8566);
xnor U9151 (N_9151,N_8718,N_8818);
or U9152 (N_9152,N_8643,N_8459);
nand U9153 (N_9153,N_8070,N_8831);
or U9154 (N_9154,N_8509,N_8280);
and U9155 (N_9155,N_8687,N_8009);
xnor U9156 (N_9156,N_8536,N_8278);
and U9157 (N_9157,N_8500,N_8208);
nor U9158 (N_9158,N_8893,N_8646);
nor U9159 (N_9159,N_8496,N_8735);
or U9160 (N_9160,N_8436,N_8110);
and U9161 (N_9161,N_8737,N_8866);
or U9162 (N_9162,N_8238,N_8658);
and U9163 (N_9163,N_8355,N_8666);
or U9164 (N_9164,N_8984,N_8224);
xor U9165 (N_9165,N_8684,N_8030);
nand U9166 (N_9166,N_8275,N_8872);
and U9167 (N_9167,N_8627,N_8982);
nor U9168 (N_9168,N_8329,N_8709);
or U9169 (N_9169,N_8880,N_8290);
nand U9170 (N_9170,N_8285,N_8703);
xnor U9171 (N_9171,N_8081,N_8736);
and U9172 (N_9172,N_8064,N_8906);
and U9173 (N_9173,N_8106,N_8482);
nand U9174 (N_9174,N_8027,N_8618);
and U9175 (N_9175,N_8613,N_8841);
or U9176 (N_9176,N_8990,N_8911);
nand U9177 (N_9177,N_8380,N_8825);
nand U9178 (N_9178,N_8215,N_8864);
and U9179 (N_9179,N_8237,N_8730);
xor U9180 (N_9180,N_8506,N_8925);
nand U9181 (N_9181,N_8410,N_8382);
or U9182 (N_9182,N_8879,N_8754);
or U9183 (N_9183,N_8424,N_8824);
and U9184 (N_9184,N_8273,N_8094);
and U9185 (N_9185,N_8321,N_8367);
or U9186 (N_9186,N_8896,N_8790);
nand U9187 (N_9187,N_8057,N_8796);
nor U9188 (N_9188,N_8763,N_8091);
and U9189 (N_9189,N_8596,N_8577);
nor U9190 (N_9190,N_8359,N_8904);
xnor U9191 (N_9191,N_8024,N_8912);
or U9192 (N_9192,N_8293,N_8075);
and U9193 (N_9193,N_8585,N_8583);
and U9194 (N_9194,N_8243,N_8270);
nor U9195 (N_9195,N_8959,N_8010);
or U9196 (N_9196,N_8255,N_8254);
nor U9197 (N_9197,N_8659,N_8115);
nor U9198 (N_9198,N_8073,N_8497);
or U9199 (N_9199,N_8889,N_8144);
nand U9200 (N_9200,N_8219,N_8038);
or U9201 (N_9201,N_8122,N_8840);
xor U9202 (N_9202,N_8797,N_8296);
nand U9203 (N_9203,N_8251,N_8119);
nand U9204 (N_9204,N_8698,N_8843);
nor U9205 (N_9205,N_8138,N_8910);
or U9206 (N_9206,N_8015,N_8570);
nand U9207 (N_9207,N_8907,N_8058);
and U9208 (N_9208,N_8863,N_8037);
nor U9209 (N_9209,N_8989,N_8456);
nand U9210 (N_9210,N_8580,N_8240);
xor U9211 (N_9211,N_8636,N_8234);
xor U9212 (N_9212,N_8738,N_8676);
or U9213 (N_9213,N_8701,N_8599);
nand U9214 (N_9214,N_8180,N_8833);
xnor U9215 (N_9215,N_8850,N_8892);
or U9216 (N_9216,N_8324,N_8908);
and U9217 (N_9217,N_8828,N_8844);
nand U9218 (N_9218,N_8998,N_8078);
nor U9219 (N_9219,N_8043,N_8929);
nand U9220 (N_9220,N_8048,N_8166);
xor U9221 (N_9221,N_8351,N_8802);
xor U9222 (N_9222,N_8541,N_8715);
nand U9223 (N_9223,N_8041,N_8017);
or U9224 (N_9224,N_8857,N_8807);
xor U9225 (N_9225,N_8431,N_8635);
and U9226 (N_9226,N_8089,N_8848);
and U9227 (N_9227,N_8898,N_8445);
xnor U9228 (N_9228,N_8574,N_8721);
nor U9229 (N_9229,N_8387,N_8558);
nand U9230 (N_9230,N_8269,N_8176);
xnor U9231 (N_9231,N_8227,N_8663);
xnor U9232 (N_9232,N_8973,N_8933);
or U9233 (N_9233,N_8512,N_8349);
and U9234 (N_9234,N_8976,N_8032);
nor U9235 (N_9235,N_8924,N_8707);
or U9236 (N_9236,N_8758,N_8672);
xnor U9237 (N_9237,N_8971,N_8050);
xor U9238 (N_9238,N_8236,N_8728);
xnor U9239 (N_9239,N_8157,N_8770);
nor U9240 (N_9240,N_8462,N_8135);
xor U9241 (N_9241,N_8940,N_8090);
xnor U9242 (N_9242,N_8495,N_8926);
nor U9243 (N_9243,N_8099,N_8869);
xnor U9244 (N_9244,N_8126,N_8054);
and U9245 (N_9245,N_8085,N_8810);
nor U9246 (N_9246,N_8320,N_8949);
nor U9247 (N_9247,N_8720,N_8544);
and U9248 (N_9248,N_8897,N_8800);
xnor U9249 (N_9249,N_8141,N_8455);
nor U9250 (N_9250,N_8520,N_8179);
and U9251 (N_9251,N_8375,N_8323);
nor U9252 (N_9252,N_8838,N_8483);
or U9253 (N_9253,N_8155,N_8968);
and U9254 (N_9254,N_8597,N_8740);
nor U9255 (N_9255,N_8107,N_8835);
nand U9256 (N_9256,N_8036,N_8046);
nor U9257 (N_9257,N_8741,N_8559);
nor U9258 (N_9258,N_8116,N_8584);
nand U9259 (N_9259,N_8248,N_8890);
nand U9260 (N_9260,N_8221,N_8148);
and U9261 (N_9261,N_8888,N_8494);
nand U9262 (N_9262,N_8369,N_8276);
xnor U9263 (N_9263,N_8749,N_8342);
or U9264 (N_9264,N_8689,N_8491);
nor U9265 (N_9265,N_8426,N_8441);
or U9266 (N_9266,N_8172,N_8154);
xnor U9267 (N_9267,N_8045,N_8080);
nand U9268 (N_9268,N_8972,N_8291);
nor U9269 (N_9269,N_8970,N_8801);
nand U9270 (N_9270,N_8732,N_8327);
and U9271 (N_9271,N_8561,N_8282);
nor U9272 (N_9272,N_8147,N_8811);
and U9273 (N_9273,N_8983,N_8228);
nand U9274 (N_9274,N_8330,N_8717);
xor U9275 (N_9275,N_8814,N_8385);
and U9276 (N_9276,N_8146,N_8149);
or U9277 (N_9277,N_8182,N_8656);
and U9278 (N_9278,N_8537,N_8239);
and U9279 (N_9279,N_8393,N_8579);
nor U9280 (N_9280,N_8286,N_8724);
xnor U9281 (N_9281,N_8439,N_8383);
and U9282 (N_9282,N_8565,N_8492);
nand U9283 (N_9283,N_8213,N_8595);
nand U9284 (N_9284,N_8919,N_8747);
nand U9285 (N_9285,N_8729,N_8414);
or U9286 (N_9286,N_8479,N_8220);
nand U9287 (N_9287,N_8013,N_8055);
nand U9288 (N_9288,N_8000,N_8160);
nand U9289 (N_9289,N_8809,N_8808);
and U9290 (N_9290,N_8433,N_8340);
or U9291 (N_9291,N_8389,N_8429);
xnor U9292 (N_9292,N_8999,N_8548);
and U9293 (N_9293,N_8706,N_8442);
or U9294 (N_9294,N_8727,N_8744);
and U9295 (N_9295,N_8136,N_8171);
xor U9296 (N_9296,N_8118,N_8093);
xor U9297 (N_9297,N_8696,N_8513);
xor U9298 (N_9298,N_8163,N_8567);
nor U9299 (N_9299,N_8137,N_8217);
xor U9300 (N_9300,N_8392,N_8295);
nand U9301 (N_9301,N_8957,N_8813);
xor U9302 (N_9302,N_8733,N_8562);
xor U9303 (N_9303,N_8946,N_8805);
nand U9304 (N_9304,N_8665,N_8308);
nand U9305 (N_9305,N_8128,N_8082);
and U9306 (N_9306,N_8980,N_8170);
xor U9307 (N_9307,N_8252,N_8007);
xnor U9308 (N_9308,N_8839,N_8430);
and U9309 (N_9309,N_8936,N_8034);
and U9310 (N_9310,N_8619,N_8616);
or U9311 (N_9311,N_8573,N_8123);
xnor U9312 (N_9312,N_8343,N_8003);
and U9313 (N_9313,N_8162,N_8001);
xnor U9314 (N_9314,N_8165,N_8300);
xor U9315 (N_9315,N_8363,N_8184);
and U9316 (N_9316,N_8865,N_8793);
and U9317 (N_9317,N_8307,N_8109);
nand U9318 (N_9318,N_8921,N_8868);
or U9319 (N_9319,N_8780,N_8481);
nand U9320 (N_9320,N_8197,N_8235);
xor U9321 (N_9321,N_8683,N_8593);
or U9322 (N_9322,N_8586,N_8470);
nand U9323 (N_9323,N_8765,N_8218);
and U9324 (N_9324,N_8401,N_8088);
xnor U9325 (N_9325,N_8575,N_8233);
or U9326 (N_9326,N_8396,N_8069);
and U9327 (N_9327,N_8287,N_8681);
nand U9328 (N_9328,N_8139,N_8917);
nor U9329 (N_9329,N_8909,N_8750);
nor U9330 (N_9330,N_8589,N_8578);
or U9331 (N_9331,N_8552,N_8263);
and U9332 (N_9332,N_8621,N_8531);
or U9333 (N_9333,N_8047,N_8774);
or U9334 (N_9334,N_8590,N_8421);
xnor U9335 (N_9335,N_8515,N_8399);
nor U9336 (N_9336,N_8016,N_8023);
nor U9337 (N_9337,N_8761,N_8247);
nor U9338 (N_9338,N_8956,N_8068);
and U9339 (N_9339,N_8317,N_8365);
nor U9340 (N_9340,N_8189,N_8167);
xor U9341 (N_9341,N_8033,N_8097);
nor U9342 (N_9342,N_8679,N_8554);
and U9343 (N_9343,N_8855,N_8769);
or U9344 (N_9344,N_8420,N_8059);
and U9345 (N_9345,N_8346,N_8690);
xnor U9346 (N_9346,N_8598,N_8782);
and U9347 (N_9347,N_8916,N_8371);
and U9348 (N_9348,N_8402,N_8791);
xor U9349 (N_9349,N_8461,N_8074);
xnor U9350 (N_9350,N_8617,N_8652);
or U9351 (N_9351,N_8061,N_8168);
and U9352 (N_9352,N_8353,N_8265);
nor U9353 (N_9353,N_8661,N_8882);
or U9354 (N_9354,N_8193,N_8669);
xnor U9355 (N_9355,N_8987,N_8615);
nand U9356 (N_9356,N_8322,N_8386);
xnor U9357 (N_9357,N_8489,N_8877);
or U9358 (N_9358,N_8298,N_8206);
nor U9359 (N_9359,N_8931,N_8963);
nand U9360 (N_9360,N_8660,N_8438);
or U9361 (N_9361,N_8845,N_8044);
nand U9362 (N_9362,N_8842,N_8111);
nand U9363 (N_9363,N_8201,N_8934);
nand U9364 (N_9364,N_8035,N_8087);
nor U9365 (N_9365,N_8798,N_8852);
xor U9366 (N_9366,N_8521,N_8011);
or U9367 (N_9367,N_8938,N_8901);
and U9368 (N_9368,N_8177,N_8670);
and U9369 (N_9369,N_8465,N_8731);
xor U9370 (N_9370,N_8222,N_8915);
xor U9371 (N_9371,N_8799,N_8700);
nor U9372 (N_9372,N_8887,N_8625);
or U9373 (N_9373,N_8326,N_8576);
or U9374 (N_9374,N_8572,N_8764);
or U9375 (N_9375,N_8458,N_8505);
xnor U9376 (N_9376,N_8673,N_8927);
xor U9377 (N_9377,N_8602,N_8476);
nand U9378 (N_9378,N_8140,N_8991);
nand U9379 (N_9379,N_8454,N_8331);
nor U9380 (N_9380,N_8156,N_8752);
nor U9381 (N_9381,N_8947,N_8600);
xor U9382 (N_9382,N_8260,N_8726);
or U9383 (N_9383,N_8962,N_8722);
nor U9384 (N_9384,N_8624,N_8685);
or U9385 (N_9385,N_8743,N_8781);
or U9386 (N_9386,N_8876,N_8210);
nand U9387 (N_9387,N_8422,N_8530);
xor U9388 (N_9388,N_8834,N_8337);
and U9389 (N_9389,N_8895,N_8937);
xor U9390 (N_9390,N_8504,N_8757);
nor U9391 (N_9391,N_8120,N_8645);
nor U9392 (N_9392,N_8594,N_8786);
and U9393 (N_9393,N_8006,N_8488);
and U9394 (N_9394,N_8432,N_8551);
nor U9395 (N_9395,N_8008,N_8112);
xor U9396 (N_9396,N_8435,N_8049);
or U9397 (N_9397,N_8950,N_8609);
nor U9398 (N_9398,N_8767,N_8846);
and U9399 (N_9399,N_8368,N_8040);
nand U9400 (N_9400,N_8692,N_8905);
or U9401 (N_9401,N_8664,N_8529);
nand U9402 (N_9402,N_8762,N_8528);
xnor U9403 (N_9403,N_8974,N_8657);
xor U9404 (N_9404,N_8169,N_8535);
xor U9405 (N_9405,N_8190,N_8066);
nor U9406 (N_9406,N_8230,N_8725);
xor U9407 (N_9407,N_8397,N_8114);
xnor U9408 (N_9408,N_8463,N_8277);
or U9409 (N_9409,N_8022,N_8319);
nand U9410 (N_9410,N_8305,N_8861);
or U9411 (N_9411,N_8486,N_8867);
and U9412 (N_9412,N_8871,N_8582);
nor U9413 (N_9413,N_8539,N_8026);
xor U9414 (N_9414,N_8019,N_8550);
nor U9415 (N_9415,N_8262,N_8002);
or U9416 (N_9416,N_8560,N_8563);
xnor U9417 (N_9417,N_8370,N_8620);
nor U9418 (N_9418,N_8674,N_8204);
xnor U9419 (N_9419,N_8328,N_8746);
and U9420 (N_9420,N_8419,N_8473);
xor U9421 (N_9421,N_8185,N_8161);
and U9422 (N_9422,N_8986,N_8131);
or U9423 (N_9423,N_8708,N_8935);
and U9424 (N_9424,N_8639,N_8516);
or U9425 (N_9425,N_8523,N_8638);
xor U9426 (N_9426,N_8102,N_8605);
and U9427 (N_9427,N_8272,N_8261);
nand U9428 (N_9428,N_8348,N_8604);
and U9429 (N_9429,N_8449,N_8335);
or U9430 (N_9430,N_8587,N_8256);
nand U9431 (N_9431,N_8977,N_8651);
xor U9432 (N_9432,N_8571,N_8444);
or U9433 (N_9433,N_8734,N_8357);
or U9434 (N_9434,N_8113,N_8748);
and U9435 (N_9435,N_8216,N_8533);
or U9436 (N_9436,N_8223,N_8902);
xor U9437 (N_9437,N_8817,N_8079);
or U9438 (N_9438,N_8266,N_8388);
and U9439 (N_9439,N_8932,N_8142);
and U9440 (N_9440,N_8423,N_8588);
xnor U9441 (N_9441,N_8785,N_8225);
nand U9442 (N_9442,N_8374,N_8381);
and U9443 (N_9443,N_8451,N_8755);
or U9444 (N_9444,N_8062,N_8944);
nor U9445 (N_9445,N_8507,N_8881);
nor U9446 (N_9446,N_8302,N_8406);
xnor U9447 (N_9447,N_8695,N_8644);
nor U9448 (N_9448,N_8198,N_8899);
and U9449 (N_9449,N_8581,N_8310);
nor U9450 (N_9450,N_8100,N_8942);
xor U9451 (N_9451,N_8766,N_8475);
or U9452 (N_9452,N_8501,N_8413);
xnor U9453 (N_9453,N_8914,N_8975);
xor U9454 (N_9454,N_8174,N_8231);
nand U9455 (N_9455,N_8742,N_8083);
or U9456 (N_9456,N_8063,N_8784);
and U9457 (N_9457,N_8981,N_8211);
and U9458 (N_9458,N_8121,N_8372);
or U9459 (N_9459,N_8918,N_8623);
nor U9460 (N_9460,N_8688,N_8532);
and U9461 (N_9461,N_8886,N_8549);
xnor U9462 (N_9462,N_8884,N_8771);
nor U9463 (N_9463,N_8874,N_8297);
and U9464 (N_9464,N_8192,N_8345);
xnor U9465 (N_9465,N_8466,N_8258);
xnor U9466 (N_9466,N_8719,N_8332);
nand U9467 (N_9467,N_8194,N_8394);
nand U9468 (N_9468,N_8789,N_8667);
nor U9469 (N_9469,N_8020,N_8301);
or U9470 (N_9470,N_8606,N_8187);
nand U9471 (N_9471,N_8641,N_8978);
nand U9472 (N_9472,N_8294,N_8557);
and U9473 (N_9473,N_8452,N_8856);
and U9474 (N_9474,N_8788,N_8525);
nand U9475 (N_9475,N_8181,N_8437);
or U9476 (N_9476,N_8250,N_8403);
nor U9477 (N_9477,N_8945,N_8885);
xor U9478 (N_9478,N_8051,N_8484);
nor U9479 (N_9479,N_8628,N_8289);
xor U9480 (N_9480,N_8853,N_8014);
and U9481 (N_9481,N_8130,N_8226);
nand U9482 (N_9482,N_8175,N_8900);
and U9483 (N_9483,N_8913,N_8498);
nor U9484 (N_9484,N_8129,N_8568);
and U9485 (N_9485,N_8592,N_8361);
and U9486 (N_9486,N_8440,N_8875);
or U9487 (N_9487,N_8953,N_8499);
nand U9488 (N_9488,N_8487,N_8212);
xor U9489 (N_9489,N_8873,N_8713);
or U9490 (N_9490,N_8779,N_8967);
nor U9491 (N_9491,N_8829,N_8716);
and U9492 (N_9492,N_8202,N_8259);
nand U9493 (N_9493,N_8518,N_8356);
nand U9494 (N_9494,N_8941,N_8712);
xnor U9495 (N_9495,N_8056,N_8271);
or U9496 (N_9496,N_8812,N_8510);
and U9497 (N_9497,N_8508,N_8460);
nand U9498 (N_9498,N_8336,N_8021);
or U9499 (N_9499,N_8502,N_8108);
xor U9500 (N_9500,N_8336,N_8558);
nand U9501 (N_9501,N_8907,N_8162);
and U9502 (N_9502,N_8878,N_8180);
nand U9503 (N_9503,N_8527,N_8223);
nor U9504 (N_9504,N_8286,N_8030);
nor U9505 (N_9505,N_8215,N_8177);
nand U9506 (N_9506,N_8634,N_8311);
and U9507 (N_9507,N_8314,N_8732);
nand U9508 (N_9508,N_8210,N_8911);
nor U9509 (N_9509,N_8336,N_8981);
nor U9510 (N_9510,N_8693,N_8714);
xor U9511 (N_9511,N_8077,N_8194);
xor U9512 (N_9512,N_8414,N_8200);
xnor U9513 (N_9513,N_8635,N_8825);
nand U9514 (N_9514,N_8054,N_8519);
or U9515 (N_9515,N_8155,N_8705);
and U9516 (N_9516,N_8496,N_8113);
xor U9517 (N_9517,N_8074,N_8963);
nand U9518 (N_9518,N_8736,N_8091);
xor U9519 (N_9519,N_8289,N_8627);
nor U9520 (N_9520,N_8269,N_8865);
nor U9521 (N_9521,N_8054,N_8206);
nand U9522 (N_9522,N_8573,N_8843);
nor U9523 (N_9523,N_8934,N_8472);
nor U9524 (N_9524,N_8490,N_8350);
xnor U9525 (N_9525,N_8236,N_8569);
xor U9526 (N_9526,N_8911,N_8714);
nand U9527 (N_9527,N_8569,N_8689);
or U9528 (N_9528,N_8478,N_8900);
nor U9529 (N_9529,N_8574,N_8760);
xnor U9530 (N_9530,N_8963,N_8702);
nor U9531 (N_9531,N_8300,N_8735);
or U9532 (N_9532,N_8709,N_8143);
or U9533 (N_9533,N_8768,N_8387);
nor U9534 (N_9534,N_8290,N_8123);
nor U9535 (N_9535,N_8797,N_8585);
xnor U9536 (N_9536,N_8603,N_8851);
xnor U9537 (N_9537,N_8034,N_8610);
nor U9538 (N_9538,N_8404,N_8534);
nor U9539 (N_9539,N_8431,N_8384);
and U9540 (N_9540,N_8227,N_8489);
or U9541 (N_9541,N_8978,N_8849);
or U9542 (N_9542,N_8975,N_8610);
or U9543 (N_9543,N_8456,N_8441);
nand U9544 (N_9544,N_8710,N_8860);
xnor U9545 (N_9545,N_8847,N_8763);
and U9546 (N_9546,N_8960,N_8433);
nor U9547 (N_9547,N_8482,N_8979);
nand U9548 (N_9548,N_8210,N_8546);
nand U9549 (N_9549,N_8229,N_8798);
xor U9550 (N_9550,N_8129,N_8575);
nand U9551 (N_9551,N_8940,N_8497);
or U9552 (N_9552,N_8472,N_8192);
nand U9553 (N_9553,N_8826,N_8195);
or U9554 (N_9554,N_8253,N_8535);
or U9555 (N_9555,N_8029,N_8847);
and U9556 (N_9556,N_8627,N_8613);
xnor U9557 (N_9557,N_8067,N_8964);
xnor U9558 (N_9558,N_8168,N_8119);
nor U9559 (N_9559,N_8026,N_8130);
xnor U9560 (N_9560,N_8404,N_8563);
and U9561 (N_9561,N_8743,N_8975);
nand U9562 (N_9562,N_8806,N_8455);
nand U9563 (N_9563,N_8455,N_8654);
nor U9564 (N_9564,N_8496,N_8421);
nand U9565 (N_9565,N_8492,N_8987);
nand U9566 (N_9566,N_8460,N_8254);
nand U9567 (N_9567,N_8554,N_8740);
and U9568 (N_9568,N_8505,N_8896);
xor U9569 (N_9569,N_8607,N_8453);
or U9570 (N_9570,N_8117,N_8901);
nand U9571 (N_9571,N_8405,N_8331);
or U9572 (N_9572,N_8645,N_8071);
and U9573 (N_9573,N_8575,N_8671);
xnor U9574 (N_9574,N_8240,N_8046);
nor U9575 (N_9575,N_8630,N_8706);
nand U9576 (N_9576,N_8050,N_8587);
nand U9577 (N_9577,N_8104,N_8276);
xor U9578 (N_9578,N_8326,N_8743);
nor U9579 (N_9579,N_8541,N_8651);
nor U9580 (N_9580,N_8316,N_8426);
nor U9581 (N_9581,N_8842,N_8557);
and U9582 (N_9582,N_8987,N_8253);
nor U9583 (N_9583,N_8147,N_8655);
and U9584 (N_9584,N_8190,N_8129);
xnor U9585 (N_9585,N_8942,N_8736);
xor U9586 (N_9586,N_8321,N_8207);
or U9587 (N_9587,N_8829,N_8752);
or U9588 (N_9588,N_8289,N_8610);
nand U9589 (N_9589,N_8003,N_8372);
xor U9590 (N_9590,N_8013,N_8551);
nand U9591 (N_9591,N_8940,N_8160);
nand U9592 (N_9592,N_8179,N_8082);
nand U9593 (N_9593,N_8588,N_8516);
nand U9594 (N_9594,N_8615,N_8322);
nor U9595 (N_9595,N_8447,N_8193);
nand U9596 (N_9596,N_8278,N_8495);
xnor U9597 (N_9597,N_8453,N_8916);
xnor U9598 (N_9598,N_8854,N_8550);
nor U9599 (N_9599,N_8205,N_8628);
nand U9600 (N_9600,N_8427,N_8354);
or U9601 (N_9601,N_8147,N_8553);
or U9602 (N_9602,N_8189,N_8935);
nand U9603 (N_9603,N_8472,N_8385);
nor U9604 (N_9604,N_8067,N_8872);
nand U9605 (N_9605,N_8256,N_8046);
or U9606 (N_9606,N_8307,N_8878);
or U9607 (N_9607,N_8277,N_8450);
and U9608 (N_9608,N_8135,N_8540);
and U9609 (N_9609,N_8674,N_8248);
xor U9610 (N_9610,N_8916,N_8154);
or U9611 (N_9611,N_8837,N_8930);
nand U9612 (N_9612,N_8692,N_8406);
or U9613 (N_9613,N_8907,N_8808);
xnor U9614 (N_9614,N_8589,N_8180);
nor U9615 (N_9615,N_8592,N_8218);
nand U9616 (N_9616,N_8979,N_8018);
or U9617 (N_9617,N_8214,N_8454);
and U9618 (N_9618,N_8967,N_8912);
and U9619 (N_9619,N_8122,N_8423);
nand U9620 (N_9620,N_8680,N_8776);
xnor U9621 (N_9621,N_8855,N_8763);
xnor U9622 (N_9622,N_8515,N_8348);
nand U9623 (N_9623,N_8164,N_8970);
xor U9624 (N_9624,N_8289,N_8968);
and U9625 (N_9625,N_8951,N_8264);
or U9626 (N_9626,N_8486,N_8779);
nand U9627 (N_9627,N_8579,N_8729);
xnor U9628 (N_9628,N_8684,N_8236);
nand U9629 (N_9629,N_8496,N_8625);
xnor U9630 (N_9630,N_8327,N_8780);
nor U9631 (N_9631,N_8066,N_8747);
xor U9632 (N_9632,N_8293,N_8759);
xor U9633 (N_9633,N_8119,N_8678);
nor U9634 (N_9634,N_8859,N_8570);
or U9635 (N_9635,N_8199,N_8310);
or U9636 (N_9636,N_8228,N_8077);
nor U9637 (N_9637,N_8859,N_8971);
xnor U9638 (N_9638,N_8121,N_8256);
nor U9639 (N_9639,N_8406,N_8156);
and U9640 (N_9640,N_8754,N_8762);
xnor U9641 (N_9641,N_8142,N_8841);
or U9642 (N_9642,N_8542,N_8151);
or U9643 (N_9643,N_8698,N_8705);
xor U9644 (N_9644,N_8778,N_8179);
xnor U9645 (N_9645,N_8305,N_8633);
xnor U9646 (N_9646,N_8048,N_8694);
xor U9647 (N_9647,N_8850,N_8417);
xnor U9648 (N_9648,N_8027,N_8388);
xnor U9649 (N_9649,N_8604,N_8745);
or U9650 (N_9650,N_8991,N_8576);
or U9651 (N_9651,N_8192,N_8057);
and U9652 (N_9652,N_8564,N_8684);
nor U9653 (N_9653,N_8803,N_8075);
xor U9654 (N_9654,N_8149,N_8542);
xnor U9655 (N_9655,N_8346,N_8384);
or U9656 (N_9656,N_8536,N_8214);
and U9657 (N_9657,N_8600,N_8589);
nor U9658 (N_9658,N_8251,N_8596);
nor U9659 (N_9659,N_8898,N_8134);
nor U9660 (N_9660,N_8286,N_8705);
nor U9661 (N_9661,N_8131,N_8766);
or U9662 (N_9662,N_8053,N_8281);
and U9663 (N_9663,N_8591,N_8741);
and U9664 (N_9664,N_8486,N_8665);
and U9665 (N_9665,N_8883,N_8546);
xor U9666 (N_9666,N_8614,N_8784);
and U9667 (N_9667,N_8415,N_8731);
nor U9668 (N_9668,N_8507,N_8690);
and U9669 (N_9669,N_8158,N_8835);
xor U9670 (N_9670,N_8450,N_8577);
nor U9671 (N_9671,N_8118,N_8217);
nand U9672 (N_9672,N_8783,N_8254);
or U9673 (N_9673,N_8569,N_8020);
and U9674 (N_9674,N_8433,N_8234);
nand U9675 (N_9675,N_8258,N_8105);
xor U9676 (N_9676,N_8253,N_8452);
nor U9677 (N_9677,N_8684,N_8703);
nor U9678 (N_9678,N_8986,N_8182);
nand U9679 (N_9679,N_8372,N_8939);
or U9680 (N_9680,N_8985,N_8860);
nor U9681 (N_9681,N_8381,N_8395);
and U9682 (N_9682,N_8030,N_8082);
or U9683 (N_9683,N_8581,N_8244);
nand U9684 (N_9684,N_8247,N_8167);
nand U9685 (N_9685,N_8999,N_8227);
nand U9686 (N_9686,N_8951,N_8132);
or U9687 (N_9687,N_8473,N_8555);
xnor U9688 (N_9688,N_8006,N_8569);
nand U9689 (N_9689,N_8643,N_8886);
nor U9690 (N_9690,N_8806,N_8920);
xnor U9691 (N_9691,N_8355,N_8893);
nand U9692 (N_9692,N_8866,N_8070);
and U9693 (N_9693,N_8071,N_8457);
nand U9694 (N_9694,N_8679,N_8832);
xor U9695 (N_9695,N_8008,N_8646);
nor U9696 (N_9696,N_8268,N_8049);
nor U9697 (N_9697,N_8865,N_8781);
xor U9698 (N_9698,N_8382,N_8823);
xor U9699 (N_9699,N_8395,N_8147);
nand U9700 (N_9700,N_8815,N_8336);
nor U9701 (N_9701,N_8148,N_8810);
nand U9702 (N_9702,N_8462,N_8380);
or U9703 (N_9703,N_8039,N_8944);
and U9704 (N_9704,N_8986,N_8152);
or U9705 (N_9705,N_8888,N_8022);
nor U9706 (N_9706,N_8451,N_8599);
xor U9707 (N_9707,N_8548,N_8464);
and U9708 (N_9708,N_8433,N_8368);
and U9709 (N_9709,N_8630,N_8436);
nand U9710 (N_9710,N_8135,N_8703);
xor U9711 (N_9711,N_8483,N_8736);
and U9712 (N_9712,N_8496,N_8028);
or U9713 (N_9713,N_8594,N_8462);
nand U9714 (N_9714,N_8556,N_8379);
or U9715 (N_9715,N_8181,N_8015);
nand U9716 (N_9716,N_8484,N_8985);
and U9717 (N_9717,N_8003,N_8704);
nand U9718 (N_9718,N_8934,N_8073);
nand U9719 (N_9719,N_8091,N_8310);
nand U9720 (N_9720,N_8250,N_8835);
nor U9721 (N_9721,N_8821,N_8657);
nor U9722 (N_9722,N_8093,N_8647);
nor U9723 (N_9723,N_8770,N_8208);
or U9724 (N_9724,N_8781,N_8634);
xor U9725 (N_9725,N_8065,N_8105);
and U9726 (N_9726,N_8169,N_8827);
nand U9727 (N_9727,N_8043,N_8152);
or U9728 (N_9728,N_8395,N_8827);
xor U9729 (N_9729,N_8920,N_8189);
nor U9730 (N_9730,N_8981,N_8848);
or U9731 (N_9731,N_8565,N_8295);
and U9732 (N_9732,N_8342,N_8327);
or U9733 (N_9733,N_8987,N_8119);
and U9734 (N_9734,N_8053,N_8883);
nand U9735 (N_9735,N_8951,N_8193);
nor U9736 (N_9736,N_8282,N_8161);
or U9737 (N_9737,N_8301,N_8017);
nand U9738 (N_9738,N_8636,N_8837);
nand U9739 (N_9739,N_8703,N_8600);
and U9740 (N_9740,N_8959,N_8127);
xnor U9741 (N_9741,N_8312,N_8784);
and U9742 (N_9742,N_8813,N_8394);
and U9743 (N_9743,N_8164,N_8495);
nand U9744 (N_9744,N_8308,N_8464);
or U9745 (N_9745,N_8082,N_8048);
xor U9746 (N_9746,N_8220,N_8031);
nor U9747 (N_9747,N_8146,N_8016);
nor U9748 (N_9748,N_8812,N_8034);
nor U9749 (N_9749,N_8377,N_8582);
and U9750 (N_9750,N_8881,N_8912);
xor U9751 (N_9751,N_8400,N_8039);
nor U9752 (N_9752,N_8510,N_8140);
xnor U9753 (N_9753,N_8048,N_8852);
nor U9754 (N_9754,N_8795,N_8198);
and U9755 (N_9755,N_8748,N_8536);
and U9756 (N_9756,N_8456,N_8516);
and U9757 (N_9757,N_8307,N_8143);
or U9758 (N_9758,N_8347,N_8942);
nand U9759 (N_9759,N_8625,N_8169);
nor U9760 (N_9760,N_8062,N_8060);
or U9761 (N_9761,N_8306,N_8655);
nand U9762 (N_9762,N_8933,N_8450);
xnor U9763 (N_9763,N_8743,N_8953);
xnor U9764 (N_9764,N_8856,N_8458);
nand U9765 (N_9765,N_8247,N_8031);
nand U9766 (N_9766,N_8894,N_8695);
and U9767 (N_9767,N_8654,N_8017);
nand U9768 (N_9768,N_8230,N_8105);
nand U9769 (N_9769,N_8795,N_8423);
nor U9770 (N_9770,N_8022,N_8876);
nor U9771 (N_9771,N_8753,N_8170);
nand U9772 (N_9772,N_8671,N_8407);
and U9773 (N_9773,N_8855,N_8875);
or U9774 (N_9774,N_8650,N_8444);
and U9775 (N_9775,N_8589,N_8863);
and U9776 (N_9776,N_8297,N_8141);
nor U9777 (N_9777,N_8375,N_8754);
nor U9778 (N_9778,N_8730,N_8272);
or U9779 (N_9779,N_8267,N_8626);
and U9780 (N_9780,N_8673,N_8506);
xnor U9781 (N_9781,N_8002,N_8062);
xor U9782 (N_9782,N_8601,N_8800);
xor U9783 (N_9783,N_8762,N_8262);
xnor U9784 (N_9784,N_8921,N_8149);
xor U9785 (N_9785,N_8051,N_8863);
and U9786 (N_9786,N_8797,N_8246);
or U9787 (N_9787,N_8204,N_8000);
xor U9788 (N_9788,N_8706,N_8346);
and U9789 (N_9789,N_8664,N_8221);
nor U9790 (N_9790,N_8908,N_8343);
nand U9791 (N_9791,N_8207,N_8890);
and U9792 (N_9792,N_8563,N_8726);
xor U9793 (N_9793,N_8054,N_8417);
or U9794 (N_9794,N_8663,N_8701);
and U9795 (N_9795,N_8213,N_8766);
and U9796 (N_9796,N_8824,N_8079);
and U9797 (N_9797,N_8729,N_8635);
or U9798 (N_9798,N_8115,N_8737);
and U9799 (N_9799,N_8106,N_8925);
and U9800 (N_9800,N_8046,N_8936);
nor U9801 (N_9801,N_8845,N_8216);
and U9802 (N_9802,N_8885,N_8613);
and U9803 (N_9803,N_8314,N_8356);
nor U9804 (N_9804,N_8074,N_8634);
xnor U9805 (N_9805,N_8476,N_8276);
and U9806 (N_9806,N_8935,N_8661);
or U9807 (N_9807,N_8471,N_8956);
nand U9808 (N_9808,N_8537,N_8055);
xnor U9809 (N_9809,N_8185,N_8142);
and U9810 (N_9810,N_8509,N_8893);
and U9811 (N_9811,N_8010,N_8600);
and U9812 (N_9812,N_8475,N_8720);
nand U9813 (N_9813,N_8303,N_8464);
nor U9814 (N_9814,N_8687,N_8042);
or U9815 (N_9815,N_8830,N_8165);
xnor U9816 (N_9816,N_8906,N_8364);
nand U9817 (N_9817,N_8485,N_8687);
nand U9818 (N_9818,N_8504,N_8222);
nand U9819 (N_9819,N_8753,N_8650);
and U9820 (N_9820,N_8423,N_8394);
xnor U9821 (N_9821,N_8527,N_8626);
nor U9822 (N_9822,N_8128,N_8470);
and U9823 (N_9823,N_8446,N_8631);
or U9824 (N_9824,N_8719,N_8439);
and U9825 (N_9825,N_8483,N_8814);
or U9826 (N_9826,N_8922,N_8569);
nand U9827 (N_9827,N_8039,N_8536);
nor U9828 (N_9828,N_8989,N_8397);
and U9829 (N_9829,N_8825,N_8374);
or U9830 (N_9830,N_8654,N_8942);
nor U9831 (N_9831,N_8599,N_8885);
nand U9832 (N_9832,N_8284,N_8017);
nand U9833 (N_9833,N_8688,N_8917);
nor U9834 (N_9834,N_8227,N_8542);
nand U9835 (N_9835,N_8282,N_8381);
xnor U9836 (N_9836,N_8529,N_8776);
or U9837 (N_9837,N_8854,N_8837);
nand U9838 (N_9838,N_8584,N_8394);
xnor U9839 (N_9839,N_8672,N_8276);
xor U9840 (N_9840,N_8512,N_8274);
xnor U9841 (N_9841,N_8291,N_8552);
xnor U9842 (N_9842,N_8441,N_8876);
nor U9843 (N_9843,N_8585,N_8795);
and U9844 (N_9844,N_8139,N_8672);
nor U9845 (N_9845,N_8220,N_8836);
nor U9846 (N_9846,N_8879,N_8458);
nor U9847 (N_9847,N_8847,N_8257);
or U9848 (N_9848,N_8167,N_8265);
xor U9849 (N_9849,N_8360,N_8254);
nor U9850 (N_9850,N_8469,N_8717);
and U9851 (N_9851,N_8136,N_8335);
nor U9852 (N_9852,N_8377,N_8752);
nand U9853 (N_9853,N_8901,N_8716);
nand U9854 (N_9854,N_8576,N_8566);
xor U9855 (N_9855,N_8164,N_8113);
xnor U9856 (N_9856,N_8388,N_8690);
xor U9857 (N_9857,N_8390,N_8851);
and U9858 (N_9858,N_8005,N_8432);
nand U9859 (N_9859,N_8447,N_8928);
or U9860 (N_9860,N_8440,N_8496);
xnor U9861 (N_9861,N_8292,N_8174);
and U9862 (N_9862,N_8305,N_8257);
xor U9863 (N_9863,N_8658,N_8659);
nand U9864 (N_9864,N_8267,N_8476);
xor U9865 (N_9865,N_8784,N_8886);
xnor U9866 (N_9866,N_8663,N_8294);
nor U9867 (N_9867,N_8812,N_8299);
or U9868 (N_9868,N_8557,N_8009);
or U9869 (N_9869,N_8099,N_8820);
xor U9870 (N_9870,N_8593,N_8698);
or U9871 (N_9871,N_8787,N_8794);
xnor U9872 (N_9872,N_8926,N_8272);
or U9873 (N_9873,N_8255,N_8595);
or U9874 (N_9874,N_8458,N_8886);
or U9875 (N_9875,N_8479,N_8488);
xnor U9876 (N_9876,N_8736,N_8879);
xor U9877 (N_9877,N_8874,N_8026);
xor U9878 (N_9878,N_8536,N_8395);
nor U9879 (N_9879,N_8301,N_8048);
and U9880 (N_9880,N_8190,N_8885);
nand U9881 (N_9881,N_8316,N_8282);
and U9882 (N_9882,N_8853,N_8357);
xnor U9883 (N_9883,N_8419,N_8956);
and U9884 (N_9884,N_8847,N_8332);
nand U9885 (N_9885,N_8222,N_8556);
nor U9886 (N_9886,N_8534,N_8952);
nor U9887 (N_9887,N_8172,N_8416);
xnor U9888 (N_9888,N_8592,N_8388);
or U9889 (N_9889,N_8866,N_8493);
or U9890 (N_9890,N_8435,N_8192);
xor U9891 (N_9891,N_8807,N_8983);
or U9892 (N_9892,N_8861,N_8629);
nand U9893 (N_9893,N_8627,N_8737);
xor U9894 (N_9894,N_8259,N_8788);
or U9895 (N_9895,N_8498,N_8307);
xnor U9896 (N_9896,N_8992,N_8746);
xor U9897 (N_9897,N_8373,N_8781);
and U9898 (N_9898,N_8535,N_8600);
or U9899 (N_9899,N_8599,N_8490);
and U9900 (N_9900,N_8303,N_8732);
or U9901 (N_9901,N_8888,N_8949);
or U9902 (N_9902,N_8377,N_8289);
and U9903 (N_9903,N_8963,N_8437);
nor U9904 (N_9904,N_8264,N_8566);
or U9905 (N_9905,N_8773,N_8520);
xor U9906 (N_9906,N_8141,N_8803);
nor U9907 (N_9907,N_8368,N_8641);
or U9908 (N_9908,N_8474,N_8103);
and U9909 (N_9909,N_8392,N_8283);
nor U9910 (N_9910,N_8771,N_8113);
and U9911 (N_9911,N_8153,N_8930);
or U9912 (N_9912,N_8800,N_8951);
nand U9913 (N_9913,N_8619,N_8162);
and U9914 (N_9914,N_8791,N_8502);
nand U9915 (N_9915,N_8055,N_8104);
or U9916 (N_9916,N_8200,N_8421);
xor U9917 (N_9917,N_8164,N_8734);
xnor U9918 (N_9918,N_8186,N_8836);
and U9919 (N_9919,N_8741,N_8867);
nor U9920 (N_9920,N_8707,N_8672);
and U9921 (N_9921,N_8643,N_8555);
or U9922 (N_9922,N_8731,N_8159);
xnor U9923 (N_9923,N_8403,N_8485);
and U9924 (N_9924,N_8502,N_8621);
xor U9925 (N_9925,N_8383,N_8971);
nor U9926 (N_9926,N_8784,N_8699);
or U9927 (N_9927,N_8915,N_8331);
or U9928 (N_9928,N_8827,N_8769);
or U9929 (N_9929,N_8177,N_8740);
and U9930 (N_9930,N_8378,N_8802);
xor U9931 (N_9931,N_8768,N_8707);
nor U9932 (N_9932,N_8261,N_8668);
nor U9933 (N_9933,N_8969,N_8808);
or U9934 (N_9934,N_8876,N_8857);
nand U9935 (N_9935,N_8060,N_8064);
and U9936 (N_9936,N_8508,N_8966);
nand U9937 (N_9937,N_8989,N_8785);
xnor U9938 (N_9938,N_8137,N_8142);
nand U9939 (N_9939,N_8654,N_8744);
or U9940 (N_9940,N_8305,N_8157);
xnor U9941 (N_9941,N_8081,N_8195);
and U9942 (N_9942,N_8314,N_8188);
nand U9943 (N_9943,N_8643,N_8507);
xnor U9944 (N_9944,N_8904,N_8377);
nand U9945 (N_9945,N_8067,N_8564);
xnor U9946 (N_9946,N_8026,N_8138);
nand U9947 (N_9947,N_8289,N_8245);
xnor U9948 (N_9948,N_8897,N_8146);
xor U9949 (N_9949,N_8355,N_8444);
nor U9950 (N_9950,N_8466,N_8105);
xnor U9951 (N_9951,N_8785,N_8291);
or U9952 (N_9952,N_8527,N_8492);
xnor U9953 (N_9953,N_8557,N_8194);
and U9954 (N_9954,N_8372,N_8040);
and U9955 (N_9955,N_8098,N_8649);
nor U9956 (N_9956,N_8607,N_8437);
xnor U9957 (N_9957,N_8437,N_8639);
nor U9958 (N_9958,N_8664,N_8307);
nor U9959 (N_9959,N_8904,N_8656);
nand U9960 (N_9960,N_8022,N_8406);
or U9961 (N_9961,N_8229,N_8819);
nand U9962 (N_9962,N_8228,N_8387);
and U9963 (N_9963,N_8552,N_8629);
xor U9964 (N_9964,N_8160,N_8761);
or U9965 (N_9965,N_8065,N_8378);
nand U9966 (N_9966,N_8849,N_8936);
nand U9967 (N_9967,N_8383,N_8190);
nor U9968 (N_9968,N_8967,N_8804);
nand U9969 (N_9969,N_8563,N_8356);
nor U9970 (N_9970,N_8931,N_8328);
nand U9971 (N_9971,N_8579,N_8921);
nand U9972 (N_9972,N_8790,N_8472);
nand U9973 (N_9973,N_8152,N_8967);
and U9974 (N_9974,N_8554,N_8313);
and U9975 (N_9975,N_8567,N_8812);
and U9976 (N_9976,N_8169,N_8498);
nand U9977 (N_9977,N_8474,N_8789);
nor U9978 (N_9978,N_8490,N_8655);
xnor U9979 (N_9979,N_8599,N_8787);
or U9980 (N_9980,N_8603,N_8577);
nor U9981 (N_9981,N_8197,N_8648);
or U9982 (N_9982,N_8536,N_8741);
nor U9983 (N_9983,N_8420,N_8243);
or U9984 (N_9984,N_8282,N_8579);
nor U9985 (N_9985,N_8226,N_8044);
or U9986 (N_9986,N_8498,N_8242);
nor U9987 (N_9987,N_8189,N_8376);
nor U9988 (N_9988,N_8903,N_8505);
nand U9989 (N_9989,N_8823,N_8617);
and U9990 (N_9990,N_8811,N_8916);
xor U9991 (N_9991,N_8304,N_8353);
xor U9992 (N_9992,N_8412,N_8248);
nand U9993 (N_9993,N_8455,N_8919);
nand U9994 (N_9994,N_8721,N_8520);
nor U9995 (N_9995,N_8617,N_8587);
nand U9996 (N_9996,N_8807,N_8818);
xor U9997 (N_9997,N_8071,N_8976);
nor U9998 (N_9998,N_8725,N_8957);
nand U9999 (N_9999,N_8039,N_8593);
xor U10000 (N_10000,N_9390,N_9750);
or U10001 (N_10001,N_9803,N_9552);
or U10002 (N_10002,N_9460,N_9828);
nand U10003 (N_10003,N_9616,N_9222);
and U10004 (N_10004,N_9225,N_9626);
and U10005 (N_10005,N_9804,N_9637);
xnor U10006 (N_10006,N_9685,N_9125);
nor U10007 (N_10007,N_9530,N_9009);
nand U10008 (N_10008,N_9364,N_9712);
or U10009 (N_10009,N_9705,N_9501);
or U10010 (N_10010,N_9141,N_9055);
nor U10011 (N_10011,N_9696,N_9752);
nand U10012 (N_10012,N_9150,N_9057);
nor U10013 (N_10013,N_9094,N_9149);
or U10014 (N_10014,N_9076,N_9972);
or U10015 (N_10015,N_9519,N_9349);
xnor U10016 (N_10016,N_9904,N_9682);
or U10017 (N_10017,N_9264,N_9909);
xnor U10018 (N_10018,N_9516,N_9002);
nand U10019 (N_10019,N_9678,N_9158);
or U10020 (N_10020,N_9433,N_9013);
or U10021 (N_10021,N_9117,N_9343);
or U10022 (N_10022,N_9533,N_9048);
nor U10023 (N_10023,N_9618,N_9858);
xnor U10024 (N_10024,N_9274,N_9469);
and U10025 (N_10025,N_9554,N_9262);
and U10026 (N_10026,N_9140,N_9820);
nor U10027 (N_10027,N_9593,N_9236);
nand U10028 (N_10028,N_9760,N_9755);
nand U10029 (N_10029,N_9913,N_9352);
nor U10030 (N_10030,N_9346,N_9537);
xnor U10031 (N_10031,N_9454,N_9894);
and U10032 (N_10032,N_9553,N_9765);
nand U10033 (N_10033,N_9170,N_9890);
xor U10034 (N_10034,N_9216,N_9463);
and U10035 (N_10035,N_9590,N_9490);
or U10036 (N_10036,N_9511,N_9413);
xor U10037 (N_10037,N_9322,N_9353);
or U10038 (N_10038,N_9132,N_9059);
or U10039 (N_10039,N_9987,N_9947);
and U10040 (N_10040,N_9266,N_9676);
nor U10041 (N_10041,N_9321,N_9428);
nor U10042 (N_10042,N_9694,N_9611);
or U10043 (N_10043,N_9237,N_9697);
and U10044 (N_10044,N_9974,N_9869);
nand U10045 (N_10045,N_9500,N_9597);
and U10046 (N_10046,N_9394,N_9914);
or U10047 (N_10047,N_9699,N_9587);
or U10048 (N_10048,N_9206,N_9186);
and U10049 (N_10049,N_9456,N_9050);
xnor U10050 (N_10050,N_9415,N_9317);
and U10051 (N_10051,N_9453,N_9448);
nand U10052 (N_10052,N_9328,N_9998);
or U10053 (N_10053,N_9212,N_9984);
or U10054 (N_10054,N_9153,N_9856);
nand U10055 (N_10055,N_9534,N_9101);
and U10056 (N_10056,N_9208,N_9794);
nor U10057 (N_10057,N_9019,N_9444);
xnor U10058 (N_10058,N_9806,N_9323);
or U10059 (N_10059,N_9548,N_9562);
or U10060 (N_10060,N_9224,N_9205);
or U10061 (N_10061,N_9066,N_9639);
or U10062 (N_10062,N_9931,N_9635);
nor U10063 (N_10063,N_9812,N_9690);
nor U10064 (N_10064,N_9768,N_9598);
xor U10065 (N_10065,N_9591,N_9811);
nand U10066 (N_10066,N_9991,N_9831);
nor U10067 (N_10067,N_9793,N_9217);
or U10068 (N_10068,N_9333,N_9753);
nand U10069 (N_10069,N_9367,N_9119);
nand U10070 (N_10070,N_9350,N_9619);
xnor U10071 (N_10071,N_9289,N_9403);
nor U10072 (N_10072,N_9508,N_9852);
and U10073 (N_10073,N_9195,N_9502);
or U10074 (N_10074,N_9551,N_9324);
or U10075 (N_10075,N_9443,N_9191);
nor U10076 (N_10076,N_9853,N_9997);
nor U10077 (N_10077,N_9392,N_9848);
or U10078 (N_10078,N_9484,N_9065);
or U10079 (N_10079,N_9020,N_9418);
xor U10080 (N_10080,N_9666,N_9044);
or U10081 (N_10081,N_9097,N_9371);
xor U10082 (N_10082,N_9389,N_9800);
nor U10083 (N_10083,N_9067,N_9201);
nand U10084 (N_10084,N_9429,N_9681);
xnor U10085 (N_10085,N_9139,N_9994);
nand U10086 (N_10086,N_9198,N_9467);
nand U10087 (N_10087,N_9046,N_9992);
and U10088 (N_10088,N_9640,N_9409);
xnor U10089 (N_10089,N_9383,N_9190);
and U10090 (N_10090,N_9609,N_9646);
and U10091 (N_10091,N_9246,N_9315);
or U10092 (N_10092,N_9393,N_9340);
xnor U10093 (N_10093,N_9620,N_9568);
or U10094 (N_10094,N_9900,N_9683);
xor U10095 (N_10095,N_9007,N_9129);
and U10096 (N_10096,N_9575,N_9870);
nand U10097 (N_10097,N_9218,N_9247);
or U10098 (N_10098,N_9263,N_9532);
or U10099 (N_10099,N_9165,N_9301);
nor U10100 (N_10100,N_9729,N_9245);
or U10101 (N_10101,N_9868,N_9993);
and U10102 (N_10102,N_9033,N_9585);
and U10103 (N_10103,N_9041,N_9926);
and U10104 (N_10104,N_9632,N_9505);
nand U10105 (N_10105,N_9691,N_9507);
nand U10106 (N_10106,N_9572,N_9095);
and U10107 (N_10107,N_9298,N_9475);
xor U10108 (N_10108,N_9331,N_9819);
xor U10109 (N_10109,N_9897,N_9813);
nor U10110 (N_10110,N_9608,N_9614);
nor U10111 (N_10111,N_9335,N_9010);
xnor U10112 (N_10112,N_9024,N_9173);
or U10113 (N_10113,N_9157,N_9910);
or U10114 (N_10114,N_9178,N_9847);
nor U10115 (N_10115,N_9134,N_9946);
or U10116 (N_10116,N_9399,N_9580);
xor U10117 (N_10117,N_9151,N_9907);
and U10118 (N_10118,N_9908,N_9951);
nand U10119 (N_10119,N_9288,N_9079);
or U10120 (N_10120,N_9130,N_9113);
xnor U10121 (N_10121,N_9872,N_9215);
nand U10122 (N_10122,N_9928,N_9492);
and U10123 (N_10123,N_9145,N_9365);
nor U10124 (N_10124,N_9612,N_9665);
and U10125 (N_10125,N_9769,N_9625);
nand U10126 (N_10126,N_9949,N_9885);
nand U10127 (N_10127,N_9647,N_9146);
nor U10128 (N_10128,N_9362,N_9523);
nand U10129 (N_10129,N_9960,N_9782);
and U10130 (N_10130,N_9829,N_9630);
nor U10131 (N_10131,N_9498,N_9796);
or U10132 (N_10132,N_9588,N_9051);
and U10133 (N_10133,N_9242,N_9999);
or U10134 (N_10134,N_9180,N_9849);
and U10135 (N_10135,N_9571,N_9358);
nor U10136 (N_10136,N_9083,N_9496);
xnor U10137 (N_10137,N_9172,N_9012);
nor U10138 (N_10138,N_9027,N_9486);
and U10139 (N_10139,N_9772,N_9701);
and U10140 (N_10140,N_9862,N_9105);
nand U10141 (N_10141,N_9293,N_9382);
xor U10142 (N_10142,N_9159,N_9574);
xnor U10143 (N_10143,N_9470,N_9834);
and U10144 (N_10144,N_9092,N_9169);
or U10145 (N_10145,N_9014,N_9751);
xnor U10146 (N_10146,N_9713,N_9808);
nor U10147 (N_10147,N_9404,N_9600);
and U10148 (N_10148,N_9886,N_9396);
and U10149 (N_10149,N_9108,N_9329);
or U10150 (N_10150,N_9927,N_9643);
and U10151 (N_10151,N_9940,N_9074);
nand U10152 (N_10152,N_9981,N_9969);
nor U10153 (N_10153,N_9096,N_9749);
xor U10154 (N_10154,N_9451,N_9260);
nand U10155 (N_10155,N_9662,N_9202);
or U10156 (N_10156,N_9361,N_9311);
xnor U10157 (N_10157,N_9589,N_9265);
nand U10158 (N_10158,N_9356,N_9162);
or U10159 (N_10159,N_9442,N_9287);
and U10160 (N_10160,N_9269,N_9354);
xor U10161 (N_10161,N_9080,N_9702);
or U10162 (N_10162,N_9320,N_9545);
nor U10163 (N_10163,N_9512,N_9986);
xor U10164 (N_10164,N_9915,N_9836);
xor U10165 (N_10165,N_9430,N_9745);
nor U10166 (N_10166,N_9219,N_9494);
nor U10167 (N_10167,N_9727,N_9474);
xor U10168 (N_10168,N_9156,N_9607);
nor U10169 (N_10169,N_9283,N_9835);
xnor U10170 (N_10170,N_9837,N_9838);
nor U10171 (N_10171,N_9226,N_9957);
nand U10172 (N_10172,N_9045,N_9672);
nor U10173 (N_10173,N_9491,N_9670);
or U10174 (N_10174,N_9982,N_9115);
and U10175 (N_10175,N_9728,N_9517);
nand U10176 (N_10176,N_9944,N_9684);
nand U10177 (N_10177,N_9503,N_9733);
nand U10178 (N_10178,N_9922,N_9419);
nor U10179 (N_10179,N_9121,N_9565);
nor U10180 (N_10180,N_9155,N_9434);
xor U10181 (N_10181,N_9642,N_9735);
or U10182 (N_10182,N_9717,N_9864);
nor U10183 (N_10183,N_9372,N_9763);
nand U10184 (N_10184,N_9230,N_9595);
nor U10185 (N_10185,N_9584,N_9823);
xor U10186 (N_10186,N_9388,N_9114);
xnor U10187 (N_10187,N_9704,N_9310);
or U10188 (N_10188,N_9558,N_9111);
or U10189 (N_10189,N_9304,N_9976);
xnor U10190 (N_10190,N_9197,N_9978);
nand U10191 (N_10191,N_9878,N_9061);
and U10192 (N_10192,N_9290,N_9499);
nor U10193 (N_10193,N_9259,N_9790);
nor U10194 (N_10194,N_9305,N_9000);
nor U10195 (N_10195,N_9905,N_9039);
and U10196 (N_10196,N_9770,N_9325);
xor U10197 (N_10197,N_9090,N_9477);
nor U10198 (N_10198,N_9968,N_9663);
or U10199 (N_10199,N_9303,N_9017);
and U10200 (N_10200,N_9762,N_9996);
xnor U10201 (N_10201,N_9495,N_9743);
and U10202 (N_10202,N_9255,N_9327);
xnor U10203 (N_10203,N_9416,N_9240);
xor U10204 (N_10204,N_9203,N_9406);
and U10205 (N_10205,N_9673,N_9556);
and U10206 (N_10206,N_9714,N_9857);
or U10207 (N_10207,N_9398,N_9137);
xnor U10208 (N_10208,N_9211,N_9192);
nor U10209 (N_10209,N_9881,N_9344);
xor U10210 (N_10210,N_9380,N_9522);
nand U10211 (N_10211,N_9531,N_9815);
nand U10212 (N_10212,N_9307,N_9510);
or U10213 (N_10213,N_9243,N_9777);
or U10214 (N_10214,N_9747,N_9104);
and U10215 (N_10215,N_9131,N_9866);
and U10216 (N_10216,N_9802,N_9824);
nand U10217 (N_10217,N_9623,N_9720);
or U10218 (N_10218,N_9932,N_9238);
xnor U10219 (N_10219,N_9648,N_9979);
nand U10220 (N_10220,N_9730,N_9319);
and U10221 (N_10221,N_9042,N_9459);
xor U10222 (N_10222,N_9724,N_9817);
nor U10223 (N_10223,N_9883,N_9592);
and U10224 (N_10224,N_9441,N_9493);
and U10225 (N_10225,N_9970,N_9711);
nor U10226 (N_10226,N_9291,N_9420);
xor U10227 (N_10227,N_9576,N_9624);
or U10228 (N_10228,N_9488,N_9267);
and U10229 (N_10229,N_9166,N_9379);
or U10230 (N_10230,N_9052,N_9110);
nand U10231 (N_10231,N_9445,N_9309);
xor U10232 (N_10232,N_9843,N_9895);
or U10233 (N_10233,N_9988,N_9543);
or U10234 (N_10234,N_9359,N_9830);
nor U10235 (N_10235,N_9995,N_9641);
and U10236 (N_10236,N_9147,N_9368);
xor U10237 (N_10237,N_9515,N_9069);
or U10238 (N_10238,N_9839,N_9845);
nor U10239 (N_10239,N_9877,N_9478);
nand U10240 (N_10240,N_9275,N_9773);
or U10241 (N_10241,N_9629,N_9832);
nor U10242 (N_10242,N_9314,N_9082);
or U10243 (N_10243,N_9708,N_9758);
or U10244 (N_10244,N_9177,N_9464);
and U10245 (N_10245,N_9468,N_9040);
and U10246 (N_10246,N_9529,N_9391);
xnor U10247 (N_10247,N_9606,N_9422);
nand U10248 (N_10248,N_9355,N_9435);
xor U10249 (N_10249,N_9937,N_9844);
or U10250 (N_10250,N_9058,N_9893);
nand U10251 (N_10251,N_9933,N_9414);
or U10252 (N_10252,N_9249,N_9351);
nand U10253 (N_10253,N_9136,N_9450);
nor U10254 (N_10254,N_9071,N_9043);
and U10255 (N_10255,N_9892,N_9654);
or U10256 (N_10256,N_9652,N_9805);
nand U10257 (N_10257,N_9687,N_9882);
nor U10258 (N_10258,N_9068,N_9138);
xnor U10259 (N_10259,N_9342,N_9457);
nand U10260 (N_10260,N_9360,N_9506);
and U10261 (N_10261,N_9308,N_9603);
or U10262 (N_10262,N_9075,N_9721);
xnor U10263 (N_10263,N_9761,N_9959);
nand U10264 (N_10264,N_9405,N_9655);
nand U10265 (N_10265,N_9254,N_9658);
nand U10266 (N_10266,N_9731,N_9659);
and U10267 (N_10267,N_9471,N_9462);
xor U10268 (N_10268,N_9193,N_9248);
or U10269 (N_10269,N_9792,N_9601);
nand U10270 (N_10270,N_9054,N_9759);
nand U10271 (N_10271,N_9476,N_9566);
nor U10272 (N_10272,N_9966,N_9161);
nand U10273 (N_10273,N_9707,N_9221);
xnor U10274 (N_10274,N_9481,N_9235);
nor U10275 (N_10275,N_9182,N_9022);
nor U10276 (N_10276,N_9898,N_9816);
nor U10277 (N_10277,N_9653,N_9906);
nand U10278 (N_10278,N_9889,N_9480);
or U10279 (N_10279,N_9840,N_9871);
or U10280 (N_10280,N_9188,N_9581);
nand U10281 (N_10281,N_9446,N_9967);
and U10282 (N_10282,N_9376,N_9410);
xnor U10283 (N_10283,N_9272,N_9073);
xnor U10284 (N_10284,N_9294,N_9783);
and U10285 (N_10285,N_9497,N_9809);
nand U10286 (N_10286,N_9473,N_9229);
and U10287 (N_10287,N_9089,N_9313);
nor U10288 (N_10288,N_9723,N_9424);
nor U10289 (N_10289,N_9561,N_9271);
nor U10290 (N_10290,N_9440,N_9417);
and U10291 (N_10291,N_9776,N_9650);
nor U10292 (N_10292,N_9163,N_9718);
and U10293 (N_10293,N_9879,N_9030);
and U10294 (N_10294,N_9525,N_9789);
or U10295 (N_10295,N_9936,N_9295);
nand U10296 (N_10296,N_9370,N_9807);
or U10297 (N_10297,N_9021,N_9023);
or U10298 (N_10298,N_9855,N_9397);
xor U10299 (N_10299,N_9739,N_9377);
nand U10300 (N_10300,N_9144,N_9700);
or U10301 (N_10301,N_9431,N_9479);
or U10302 (N_10302,N_9920,N_9078);
nand U10303 (N_10303,N_9357,N_9680);
nor U10304 (N_10304,N_9689,N_9621);
and U10305 (N_10305,N_9764,N_9175);
or U10306 (N_10306,N_9706,N_9942);
xnor U10307 (N_10307,N_9081,N_9306);
xor U10308 (N_10308,N_9535,N_9189);
or U10309 (N_10309,N_9634,N_9636);
and U10310 (N_10310,N_9774,N_9207);
and U10311 (N_10311,N_9771,N_9651);
and U10312 (N_10312,N_9945,N_9087);
or U10313 (N_10313,N_9228,N_9160);
nor U10314 (N_10314,N_9250,N_9958);
nor U10315 (N_10315,N_9261,N_9656);
nand U10316 (N_10316,N_9550,N_9077);
and U10317 (N_10317,N_9559,N_9126);
nor U10318 (N_10318,N_9003,N_9318);
or U10319 (N_10319,N_9911,N_9709);
nor U10320 (N_10320,N_9780,N_9302);
xor U10321 (N_10321,N_9693,N_9722);
xor U10322 (N_10322,N_9276,N_9513);
nand U10323 (N_10323,N_9638,N_9661);
and U10324 (N_10324,N_9123,N_9567);
nor U10325 (N_10325,N_9466,N_9381);
nor U10326 (N_10326,N_9887,N_9547);
xnor U10327 (N_10327,N_9569,N_9810);
or U10328 (N_10328,N_9427,N_9899);
nand U10329 (N_10329,N_9846,N_9546);
nor U10330 (N_10330,N_9983,N_9004);
nor U10331 (N_10331,N_9439,N_9099);
xnor U10332 (N_10332,N_9120,N_9112);
nand U10333 (N_10333,N_9231,N_9256);
or U10334 (N_10334,N_9710,N_9280);
nor U10335 (N_10335,N_9411,N_9395);
and U10336 (N_10336,N_9387,N_9692);
and U10337 (N_10337,N_9018,N_9924);
xor U10338 (N_10338,N_9859,N_9093);
or U10339 (N_10339,N_9686,N_9677);
nor U10340 (N_10340,N_9179,N_9461);
or U10341 (N_10341,N_9032,N_9176);
and U10342 (N_10342,N_9985,N_9756);
xnor U10343 (N_10343,N_9223,N_9818);
nand U10344 (N_10344,N_9366,N_9929);
and U10345 (N_10345,N_9107,N_9826);
nor U10346 (N_10346,N_9671,N_9605);
and U10347 (N_10347,N_9602,N_9965);
or U10348 (N_10348,N_9627,N_9599);
or U10349 (N_10349,N_9421,N_9766);
xor U10350 (N_10350,N_9742,N_9746);
nor U10351 (N_10351,N_9268,N_9785);
nor U10352 (N_10352,N_9253,N_9821);
or U10353 (N_10353,N_9633,N_9977);
nor U10354 (N_10354,N_9948,N_9423);
and U10355 (N_10355,N_9028,N_9369);
nor U10356 (N_10356,N_9901,N_9085);
or U10357 (N_10357,N_9719,N_9363);
xor U10358 (N_10358,N_9649,N_9918);
nor U10359 (N_10359,N_9016,N_9233);
nand U10360 (N_10360,N_9674,N_9282);
nor U10361 (N_10361,N_9549,N_9458);
xnor U10362 (N_10362,N_9934,N_9675);
and U10363 (N_10363,N_9152,N_9436);
xnor U10364 (N_10364,N_9337,N_9098);
nand U10365 (N_10365,N_9164,N_9784);
and U10366 (N_10366,N_9876,N_9084);
nor U10367 (N_10367,N_9822,N_9989);
or U10368 (N_10368,N_9827,N_9312);
xor U10369 (N_10369,N_9278,N_9564);
or U10370 (N_10370,N_9286,N_9181);
nand U10371 (N_10371,N_9336,N_9912);
or U10372 (N_10372,N_9524,N_9594);
and U10373 (N_10373,N_9025,N_9669);
nor U10374 (N_10374,N_9124,N_9698);
xnor U10375 (N_10375,N_9888,N_9432);
nand U10376 (N_10376,N_9873,N_9005);
nand U10377 (N_10377,N_9127,N_9962);
nand U10378 (N_10378,N_9292,N_9091);
and U10379 (N_10379,N_9174,N_9374);
and U10380 (N_10380,N_9296,N_9171);
nand U10381 (N_10381,N_9106,N_9825);
or U10382 (N_10382,N_9854,N_9521);
xor U10383 (N_10383,N_9916,N_9386);
nor U10384 (N_10384,N_9273,N_9241);
xnor U10385 (N_10385,N_9896,N_9833);
nand U10386 (N_10386,N_9412,N_9540);
nor U10387 (N_10387,N_9875,N_9865);
nor U10388 (N_10388,N_9520,N_9798);
xor U10389 (N_10389,N_9026,N_9187);
xnor U10390 (N_10390,N_9384,N_9064);
or U10391 (N_10391,N_9891,N_9570);
xnor U10392 (N_10392,N_9037,N_9330);
nand U10393 (N_10393,N_9518,N_9257);
xnor U10394 (N_10394,N_9167,N_9788);
xnor U10395 (N_10395,N_9644,N_9631);
nor U10396 (N_10396,N_9465,N_9526);
and U10397 (N_10397,N_9281,N_9034);
or U10398 (N_10398,N_9950,N_9767);
nand U10399 (N_10399,N_9485,N_9741);
or U10400 (N_10400,N_9487,N_9400);
nor U10401 (N_10401,N_9408,N_9143);
nor U10402 (N_10402,N_9199,N_9128);
nand U10403 (N_10403,N_9973,N_9941);
xnor U10404 (N_10404,N_9861,N_9244);
nor U10405 (N_10405,N_9577,N_9482);
or U10406 (N_10406,N_9736,N_9200);
and U10407 (N_10407,N_9285,N_9015);
nor U10408 (N_10408,N_9695,N_9943);
nor U10409 (N_10409,N_9851,N_9006);
nor U10410 (N_10410,N_9483,N_9116);
and U10411 (N_10411,N_9316,N_9557);
xnor U10412 (N_10412,N_9781,N_9667);
xor U10413 (N_10413,N_9063,N_9645);
or U10414 (N_10414,N_9715,N_9196);
xor U10415 (N_10415,N_9514,N_9596);
xor U10416 (N_10416,N_9220,N_9657);
and U10417 (N_10417,N_9622,N_9339);
nand U10418 (N_10418,N_9031,N_9338);
or U10419 (N_10419,N_9185,N_9573);
xor U10420 (N_10420,N_9194,N_9716);
and U10421 (N_10421,N_9449,N_9438);
or U10422 (N_10422,N_9258,N_9072);
nor U10423 (N_10423,N_9437,N_9011);
nand U10424 (N_10424,N_9118,N_9345);
nor U10425 (N_10425,N_9542,N_9279);
nor U10426 (N_10426,N_9679,N_9841);
or U10427 (N_10427,N_9668,N_9053);
and U10428 (N_10428,N_9086,N_9001);
xor U10429 (N_10429,N_9509,N_9921);
or U10430 (N_10430,N_9961,N_9930);
xor U10431 (N_10431,N_9252,N_9541);
or U10432 (N_10432,N_9029,N_9604);
nand U10433 (N_10433,N_9660,N_9903);
xor U10434 (N_10434,N_9953,N_9210);
or U10435 (N_10435,N_9334,N_9232);
nand U10436 (N_10436,N_9504,N_9725);
nor U10437 (N_10437,N_9284,N_9582);
and U10438 (N_10438,N_9975,N_9956);
and U10439 (N_10439,N_9347,N_9555);
or U10440 (N_10440,N_9787,N_9863);
xor U10441 (N_10441,N_9884,N_9938);
xnor U10442 (N_10442,N_9579,N_9239);
xor U10443 (N_10443,N_9425,N_9939);
nor U10444 (N_10444,N_9214,N_9726);
and U10445 (N_10445,N_9860,N_9527);
or U10446 (N_10446,N_9775,N_9234);
or U10447 (N_10447,N_9613,N_9748);
xnor U10448 (N_10448,N_9786,N_9952);
nand U10449 (N_10449,N_9332,N_9122);
nor U10450 (N_10450,N_9737,N_9204);
nand U10451 (N_10451,N_9135,N_9341);
xor U10452 (N_10452,N_9452,N_9183);
nor U10453 (N_10453,N_9056,N_9732);
xor U10454 (N_10454,N_9270,N_9744);
xor U10455 (N_10455,N_9047,N_9277);
or U10456 (N_10456,N_9154,N_9348);
nor U10457 (N_10457,N_9925,N_9610);
xor U10458 (N_10458,N_9935,N_9209);
or U10459 (N_10459,N_9563,N_9740);
and U10460 (N_10460,N_9586,N_9955);
nor U10461 (N_10461,N_9738,N_9954);
nand U10462 (N_10462,N_9734,N_9980);
xnor U10463 (N_10463,N_9227,N_9797);
nor U10464 (N_10464,N_9536,N_9035);
nand U10465 (N_10465,N_9300,N_9902);
nand U10466 (N_10466,N_9791,N_9880);
nand U10467 (N_10467,N_9923,N_9795);
or U10468 (N_10468,N_9528,N_9036);
xnor U10469 (N_10469,N_9299,N_9814);
xor U10470 (N_10470,N_9628,N_9917);
nor U10471 (N_10471,N_9688,N_9990);
and U10472 (N_10472,N_9874,N_9375);
and U10473 (N_10473,N_9060,N_9407);
nor U10474 (N_10474,N_9008,N_9385);
nor U10475 (N_10475,N_9088,N_9401);
or U10476 (N_10476,N_9062,N_9455);
nand U10477 (N_10477,N_9378,N_9297);
and U10478 (N_10478,N_9447,N_9971);
nand U10479 (N_10479,N_9109,N_9251);
nor U10480 (N_10480,N_9213,N_9617);
and U10481 (N_10481,N_9472,N_9919);
nor U10482 (N_10482,N_9489,N_9779);
nor U10483 (N_10483,N_9373,N_9102);
or U10484 (N_10484,N_9038,N_9799);
and U10485 (N_10485,N_9402,N_9964);
xor U10486 (N_10486,N_9426,N_9703);
or U10487 (N_10487,N_9578,N_9539);
and U10488 (N_10488,N_9850,N_9326);
nand U10489 (N_10489,N_9148,N_9142);
nand U10490 (N_10490,N_9583,N_9801);
nand U10491 (N_10491,N_9842,N_9757);
nand U10492 (N_10492,N_9049,N_9778);
xnor U10493 (N_10493,N_9538,N_9168);
xnor U10494 (N_10494,N_9754,N_9133);
nand U10495 (N_10495,N_9184,N_9070);
and U10496 (N_10496,N_9544,N_9615);
nor U10497 (N_10497,N_9664,N_9100);
or U10498 (N_10498,N_9867,N_9963);
nand U10499 (N_10499,N_9103,N_9560);
nor U10500 (N_10500,N_9613,N_9089);
nand U10501 (N_10501,N_9451,N_9114);
nand U10502 (N_10502,N_9865,N_9449);
nor U10503 (N_10503,N_9338,N_9747);
nand U10504 (N_10504,N_9554,N_9451);
xnor U10505 (N_10505,N_9582,N_9295);
nand U10506 (N_10506,N_9742,N_9052);
nand U10507 (N_10507,N_9306,N_9632);
nand U10508 (N_10508,N_9959,N_9469);
or U10509 (N_10509,N_9434,N_9435);
and U10510 (N_10510,N_9342,N_9626);
nor U10511 (N_10511,N_9868,N_9882);
nor U10512 (N_10512,N_9788,N_9681);
or U10513 (N_10513,N_9709,N_9022);
or U10514 (N_10514,N_9099,N_9798);
nor U10515 (N_10515,N_9543,N_9029);
or U10516 (N_10516,N_9346,N_9937);
and U10517 (N_10517,N_9916,N_9951);
xor U10518 (N_10518,N_9511,N_9865);
or U10519 (N_10519,N_9129,N_9903);
or U10520 (N_10520,N_9484,N_9464);
and U10521 (N_10521,N_9056,N_9522);
nand U10522 (N_10522,N_9728,N_9611);
xor U10523 (N_10523,N_9335,N_9098);
nand U10524 (N_10524,N_9897,N_9651);
or U10525 (N_10525,N_9871,N_9387);
nor U10526 (N_10526,N_9332,N_9246);
or U10527 (N_10527,N_9904,N_9686);
nand U10528 (N_10528,N_9582,N_9547);
nand U10529 (N_10529,N_9903,N_9874);
nand U10530 (N_10530,N_9485,N_9522);
or U10531 (N_10531,N_9079,N_9207);
nor U10532 (N_10532,N_9505,N_9595);
xnor U10533 (N_10533,N_9518,N_9009);
xnor U10534 (N_10534,N_9091,N_9601);
or U10535 (N_10535,N_9684,N_9501);
or U10536 (N_10536,N_9802,N_9151);
and U10537 (N_10537,N_9503,N_9465);
nand U10538 (N_10538,N_9896,N_9349);
xor U10539 (N_10539,N_9144,N_9777);
nor U10540 (N_10540,N_9222,N_9413);
and U10541 (N_10541,N_9574,N_9412);
or U10542 (N_10542,N_9249,N_9649);
xnor U10543 (N_10543,N_9434,N_9473);
nand U10544 (N_10544,N_9683,N_9022);
xnor U10545 (N_10545,N_9365,N_9090);
nand U10546 (N_10546,N_9493,N_9964);
or U10547 (N_10547,N_9163,N_9040);
and U10548 (N_10548,N_9733,N_9557);
or U10549 (N_10549,N_9804,N_9304);
nor U10550 (N_10550,N_9428,N_9988);
nor U10551 (N_10551,N_9029,N_9040);
nand U10552 (N_10552,N_9092,N_9750);
xor U10553 (N_10553,N_9166,N_9888);
xnor U10554 (N_10554,N_9418,N_9081);
nor U10555 (N_10555,N_9274,N_9354);
and U10556 (N_10556,N_9080,N_9934);
nor U10557 (N_10557,N_9753,N_9846);
and U10558 (N_10558,N_9972,N_9228);
and U10559 (N_10559,N_9168,N_9256);
and U10560 (N_10560,N_9072,N_9148);
and U10561 (N_10561,N_9251,N_9957);
nand U10562 (N_10562,N_9316,N_9364);
nor U10563 (N_10563,N_9179,N_9560);
and U10564 (N_10564,N_9291,N_9087);
xor U10565 (N_10565,N_9248,N_9370);
nor U10566 (N_10566,N_9678,N_9103);
xnor U10567 (N_10567,N_9343,N_9635);
nand U10568 (N_10568,N_9890,N_9501);
nand U10569 (N_10569,N_9061,N_9397);
nand U10570 (N_10570,N_9589,N_9489);
and U10571 (N_10571,N_9598,N_9101);
nor U10572 (N_10572,N_9053,N_9561);
or U10573 (N_10573,N_9837,N_9394);
xor U10574 (N_10574,N_9074,N_9662);
nand U10575 (N_10575,N_9070,N_9449);
nor U10576 (N_10576,N_9926,N_9431);
or U10577 (N_10577,N_9412,N_9041);
or U10578 (N_10578,N_9242,N_9140);
nand U10579 (N_10579,N_9374,N_9223);
nand U10580 (N_10580,N_9106,N_9276);
nor U10581 (N_10581,N_9365,N_9624);
or U10582 (N_10582,N_9784,N_9608);
nor U10583 (N_10583,N_9014,N_9133);
nand U10584 (N_10584,N_9107,N_9034);
xnor U10585 (N_10585,N_9417,N_9935);
and U10586 (N_10586,N_9544,N_9387);
xor U10587 (N_10587,N_9208,N_9064);
nor U10588 (N_10588,N_9523,N_9277);
nor U10589 (N_10589,N_9231,N_9745);
and U10590 (N_10590,N_9117,N_9254);
or U10591 (N_10591,N_9390,N_9630);
xor U10592 (N_10592,N_9660,N_9760);
and U10593 (N_10593,N_9163,N_9702);
and U10594 (N_10594,N_9946,N_9887);
nand U10595 (N_10595,N_9064,N_9491);
xnor U10596 (N_10596,N_9529,N_9192);
and U10597 (N_10597,N_9288,N_9392);
nand U10598 (N_10598,N_9003,N_9087);
and U10599 (N_10599,N_9229,N_9237);
nand U10600 (N_10600,N_9258,N_9401);
and U10601 (N_10601,N_9596,N_9708);
xnor U10602 (N_10602,N_9040,N_9134);
nand U10603 (N_10603,N_9837,N_9953);
nand U10604 (N_10604,N_9980,N_9923);
nand U10605 (N_10605,N_9602,N_9473);
or U10606 (N_10606,N_9705,N_9649);
or U10607 (N_10607,N_9885,N_9901);
and U10608 (N_10608,N_9536,N_9931);
nand U10609 (N_10609,N_9287,N_9757);
and U10610 (N_10610,N_9189,N_9936);
or U10611 (N_10611,N_9041,N_9640);
nor U10612 (N_10612,N_9682,N_9781);
or U10613 (N_10613,N_9505,N_9652);
or U10614 (N_10614,N_9950,N_9202);
nand U10615 (N_10615,N_9390,N_9462);
and U10616 (N_10616,N_9778,N_9524);
and U10617 (N_10617,N_9414,N_9321);
nor U10618 (N_10618,N_9447,N_9777);
and U10619 (N_10619,N_9972,N_9370);
xnor U10620 (N_10620,N_9088,N_9922);
xnor U10621 (N_10621,N_9205,N_9219);
xnor U10622 (N_10622,N_9627,N_9249);
xnor U10623 (N_10623,N_9835,N_9710);
and U10624 (N_10624,N_9017,N_9151);
or U10625 (N_10625,N_9053,N_9656);
xor U10626 (N_10626,N_9722,N_9088);
nor U10627 (N_10627,N_9009,N_9663);
or U10628 (N_10628,N_9936,N_9514);
nand U10629 (N_10629,N_9898,N_9142);
and U10630 (N_10630,N_9971,N_9273);
nor U10631 (N_10631,N_9862,N_9357);
and U10632 (N_10632,N_9847,N_9062);
or U10633 (N_10633,N_9486,N_9283);
nor U10634 (N_10634,N_9087,N_9698);
nand U10635 (N_10635,N_9098,N_9762);
or U10636 (N_10636,N_9574,N_9442);
nor U10637 (N_10637,N_9582,N_9364);
nor U10638 (N_10638,N_9786,N_9852);
nor U10639 (N_10639,N_9919,N_9264);
xnor U10640 (N_10640,N_9942,N_9873);
and U10641 (N_10641,N_9525,N_9567);
xor U10642 (N_10642,N_9647,N_9249);
nor U10643 (N_10643,N_9170,N_9839);
or U10644 (N_10644,N_9086,N_9661);
nor U10645 (N_10645,N_9972,N_9961);
or U10646 (N_10646,N_9607,N_9525);
or U10647 (N_10647,N_9285,N_9159);
and U10648 (N_10648,N_9804,N_9652);
nand U10649 (N_10649,N_9952,N_9338);
nor U10650 (N_10650,N_9915,N_9695);
and U10651 (N_10651,N_9268,N_9241);
or U10652 (N_10652,N_9046,N_9636);
nand U10653 (N_10653,N_9569,N_9021);
nand U10654 (N_10654,N_9253,N_9741);
nand U10655 (N_10655,N_9244,N_9636);
xnor U10656 (N_10656,N_9879,N_9207);
or U10657 (N_10657,N_9256,N_9850);
or U10658 (N_10658,N_9943,N_9671);
nand U10659 (N_10659,N_9475,N_9842);
or U10660 (N_10660,N_9027,N_9632);
xor U10661 (N_10661,N_9622,N_9831);
nor U10662 (N_10662,N_9445,N_9393);
or U10663 (N_10663,N_9630,N_9022);
or U10664 (N_10664,N_9897,N_9173);
or U10665 (N_10665,N_9751,N_9194);
and U10666 (N_10666,N_9657,N_9656);
and U10667 (N_10667,N_9384,N_9838);
nand U10668 (N_10668,N_9514,N_9639);
or U10669 (N_10669,N_9570,N_9680);
or U10670 (N_10670,N_9923,N_9267);
nor U10671 (N_10671,N_9190,N_9438);
nand U10672 (N_10672,N_9589,N_9413);
nand U10673 (N_10673,N_9340,N_9494);
xnor U10674 (N_10674,N_9645,N_9242);
nand U10675 (N_10675,N_9776,N_9723);
nand U10676 (N_10676,N_9494,N_9500);
nand U10677 (N_10677,N_9040,N_9586);
nor U10678 (N_10678,N_9991,N_9077);
and U10679 (N_10679,N_9603,N_9056);
or U10680 (N_10680,N_9158,N_9724);
nand U10681 (N_10681,N_9971,N_9005);
and U10682 (N_10682,N_9706,N_9233);
nand U10683 (N_10683,N_9292,N_9678);
or U10684 (N_10684,N_9456,N_9572);
nand U10685 (N_10685,N_9257,N_9264);
or U10686 (N_10686,N_9071,N_9369);
nor U10687 (N_10687,N_9816,N_9832);
nand U10688 (N_10688,N_9140,N_9617);
nand U10689 (N_10689,N_9939,N_9101);
and U10690 (N_10690,N_9902,N_9892);
xor U10691 (N_10691,N_9860,N_9491);
or U10692 (N_10692,N_9098,N_9728);
or U10693 (N_10693,N_9763,N_9639);
xnor U10694 (N_10694,N_9046,N_9963);
or U10695 (N_10695,N_9857,N_9186);
xnor U10696 (N_10696,N_9323,N_9170);
nand U10697 (N_10697,N_9488,N_9133);
nor U10698 (N_10698,N_9514,N_9767);
nand U10699 (N_10699,N_9036,N_9554);
nand U10700 (N_10700,N_9607,N_9078);
nor U10701 (N_10701,N_9643,N_9678);
nand U10702 (N_10702,N_9372,N_9183);
or U10703 (N_10703,N_9770,N_9674);
nor U10704 (N_10704,N_9592,N_9104);
and U10705 (N_10705,N_9560,N_9702);
nand U10706 (N_10706,N_9279,N_9995);
and U10707 (N_10707,N_9221,N_9858);
nor U10708 (N_10708,N_9221,N_9806);
nor U10709 (N_10709,N_9339,N_9799);
xor U10710 (N_10710,N_9154,N_9860);
xor U10711 (N_10711,N_9770,N_9754);
nand U10712 (N_10712,N_9846,N_9100);
and U10713 (N_10713,N_9295,N_9820);
nand U10714 (N_10714,N_9015,N_9039);
nand U10715 (N_10715,N_9769,N_9944);
nand U10716 (N_10716,N_9538,N_9514);
nor U10717 (N_10717,N_9219,N_9649);
nor U10718 (N_10718,N_9343,N_9366);
nor U10719 (N_10719,N_9263,N_9186);
xor U10720 (N_10720,N_9430,N_9507);
and U10721 (N_10721,N_9728,N_9991);
and U10722 (N_10722,N_9496,N_9588);
nor U10723 (N_10723,N_9241,N_9966);
nor U10724 (N_10724,N_9334,N_9012);
and U10725 (N_10725,N_9024,N_9958);
and U10726 (N_10726,N_9020,N_9142);
nand U10727 (N_10727,N_9771,N_9820);
nor U10728 (N_10728,N_9939,N_9340);
xnor U10729 (N_10729,N_9201,N_9463);
and U10730 (N_10730,N_9984,N_9442);
or U10731 (N_10731,N_9990,N_9777);
or U10732 (N_10732,N_9440,N_9256);
xnor U10733 (N_10733,N_9501,N_9675);
xor U10734 (N_10734,N_9740,N_9629);
or U10735 (N_10735,N_9317,N_9817);
or U10736 (N_10736,N_9925,N_9644);
and U10737 (N_10737,N_9792,N_9958);
nand U10738 (N_10738,N_9491,N_9529);
nand U10739 (N_10739,N_9833,N_9616);
xor U10740 (N_10740,N_9467,N_9645);
nand U10741 (N_10741,N_9775,N_9854);
and U10742 (N_10742,N_9877,N_9789);
and U10743 (N_10743,N_9953,N_9840);
or U10744 (N_10744,N_9976,N_9044);
or U10745 (N_10745,N_9552,N_9769);
xnor U10746 (N_10746,N_9473,N_9833);
or U10747 (N_10747,N_9856,N_9168);
and U10748 (N_10748,N_9553,N_9378);
nand U10749 (N_10749,N_9803,N_9935);
nor U10750 (N_10750,N_9994,N_9129);
and U10751 (N_10751,N_9171,N_9161);
nor U10752 (N_10752,N_9478,N_9917);
xor U10753 (N_10753,N_9421,N_9663);
and U10754 (N_10754,N_9418,N_9052);
or U10755 (N_10755,N_9951,N_9805);
or U10756 (N_10756,N_9379,N_9418);
nor U10757 (N_10757,N_9554,N_9906);
and U10758 (N_10758,N_9661,N_9489);
xnor U10759 (N_10759,N_9436,N_9030);
or U10760 (N_10760,N_9449,N_9225);
xnor U10761 (N_10761,N_9329,N_9828);
nor U10762 (N_10762,N_9717,N_9756);
nand U10763 (N_10763,N_9639,N_9948);
nor U10764 (N_10764,N_9676,N_9628);
nor U10765 (N_10765,N_9028,N_9669);
or U10766 (N_10766,N_9219,N_9634);
nor U10767 (N_10767,N_9591,N_9686);
nand U10768 (N_10768,N_9396,N_9076);
and U10769 (N_10769,N_9249,N_9231);
nand U10770 (N_10770,N_9720,N_9189);
and U10771 (N_10771,N_9203,N_9955);
xnor U10772 (N_10772,N_9313,N_9516);
xnor U10773 (N_10773,N_9256,N_9581);
and U10774 (N_10774,N_9336,N_9847);
nand U10775 (N_10775,N_9041,N_9828);
nand U10776 (N_10776,N_9082,N_9124);
or U10777 (N_10777,N_9711,N_9085);
xnor U10778 (N_10778,N_9543,N_9778);
nand U10779 (N_10779,N_9807,N_9030);
nor U10780 (N_10780,N_9787,N_9699);
nor U10781 (N_10781,N_9608,N_9235);
nor U10782 (N_10782,N_9112,N_9843);
or U10783 (N_10783,N_9734,N_9581);
nor U10784 (N_10784,N_9184,N_9848);
nor U10785 (N_10785,N_9263,N_9103);
nor U10786 (N_10786,N_9754,N_9173);
or U10787 (N_10787,N_9927,N_9033);
or U10788 (N_10788,N_9554,N_9138);
or U10789 (N_10789,N_9378,N_9576);
nor U10790 (N_10790,N_9795,N_9546);
nor U10791 (N_10791,N_9487,N_9433);
and U10792 (N_10792,N_9171,N_9263);
or U10793 (N_10793,N_9476,N_9420);
nand U10794 (N_10794,N_9688,N_9915);
or U10795 (N_10795,N_9623,N_9718);
nor U10796 (N_10796,N_9662,N_9549);
xnor U10797 (N_10797,N_9171,N_9398);
or U10798 (N_10798,N_9312,N_9973);
and U10799 (N_10799,N_9562,N_9202);
or U10800 (N_10800,N_9862,N_9844);
xor U10801 (N_10801,N_9638,N_9202);
or U10802 (N_10802,N_9819,N_9778);
nor U10803 (N_10803,N_9623,N_9076);
xor U10804 (N_10804,N_9172,N_9877);
xor U10805 (N_10805,N_9768,N_9995);
or U10806 (N_10806,N_9881,N_9180);
nand U10807 (N_10807,N_9201,N_9014);
or U10808 (N_10808,N_9448,N_9960);
xnor U10809 (N_10809,N_9769,N_9737);
xor U10810 (N_10810,N_9322,N_9196);
or U10811 (N_10811,N_9561,N_9729);
and U10812 (N_10812,N_9530,N_9801);
xnor U10813 (N_10813,N_9079,N_9942);
or U10814 (N_10814,N_9324,N_9449);
and U10815 (N_10815,N_9521,N_9343);
and U10816 (N_10816,N_9861,N_9919);
or U10817 (N_10817,N_9820,N_9065);
and U10818 (N_10818,N_9527,N_9813);
and U10819 (N_10819,N_9526,N_9829);
xor U10820 (N_10820,N_9811,N_9040);
or U10821 (N_10821,N_9197,N_9348);
or U10822 (N_10822,N_9954,N_9337);
nor U10823 (N_10823,N_9235,N_9494);
nor U10824 (N_10824,N_9378,N_9612);
xor U10825 (N_10825,N_9176,N_9022);
nor U10826 (N_10826,N_9907,N_9453);
or U10827 (N_10827,N_9330,N_9503);
nand U10828 (N_10828,N_9183,N_9461);
nor U10829 (N_10829,N_9582,N_9596);
nand U10830 (N_10830,N_9219,N_9117);
or U10831 (N_10831,N_9946,N_9442);
nor U10832 (N_10832,N_9810,N_9557);
xnor U10833 (N_10833,N_9658,N_9533);
nand U10834 (N_10834,N_9033,N_9147);
nor U10835 (N_10835,N_9574,N_9019);
nor U10836 (N_10836,N_9309,N_9167);
nand U10837 (N_10837,N_9874,N_9045);
and U10838 (N_10838,N_9147,N_9664);
nand U10839 (N_10839,N_9029,N_9579);
or U10840 (N_10840,N_9156,N_9479);
xor U10841 (N_10841,N_9428,N_9921);
xnor U10842 (N_10842,N_9089,N_9623);
xor U10843 (N_10843,N_9157,N_9232);
xnor U10844 (N_10844,N_9827,N_9611);
and U10845 (N_10845,N_9071,N_9822);
and U10846 (N_10846,N_9037,N_9798);
nand U10847 (N_10847,N_9884,N_9347);
nand U10848 (N_10848,N_9233,N_9214);
or U10849 (N_10849,N_9636,N_9456);
or U10850 (N_10850,N_9648,N_9974);
and U10851 (N_10851,N_9613,N_9625);
xor U10852 (N_10852,N_9290,N_9004);
or U10853 (N_10853,N_9723,N_9854);
nor U10854 (N_10854,N_9201,N_9066);
nand U10855 (N_10855,N_9832,N_9073);
or U10856 (N_10856,N_9232,N_9010);
or U10857 (N_10857,N_9637,N_9190);
nand U10858 (N_10858,N_9096,N_9621);
nand U10859 (N_10859,N_9351,N_9280);
nand U10860 (N_10860,N_9460,N_9302);
nand U10861 (N_10861,N_9971,N_9160);
xnor U10862 (N_10862,N_9251,N_9879);
or U10863 (N_10863,N_9608,N_9910);
or U10864 (N_10864,N_9103,N_9123);
or U10865 (N_10865,N_9908,N_9883);
or U10866 (N_10866,N_9680,N_9500);
or U10867 (N_10867,N_9758,N_9501);
xnor U10868 (N_10868,N_9043,N_9084);
and U10869 (N_10869,N_9174,N_9848);
xor U10870 (N_10870,N_9643,N_9139);
nand U10871 (N_10871,N_9001,N_9991);
xnor U10872 (N_10872,N_9436,N_9794);
xnor U10873 (N_10873,N_9111,N_9385);
and U10874 (N_10874,N_9591,N_9735);
xnor U10875 (N_10875,N_9006,N_9980);
nand U10876 (N_10876,N_9285,N_9424);
nand U10877 (N_10877,N_9670,N_9407);
xnor U10878 (N_10878,N_9343,N_9460);
nand U10879 (N_10879,N_9584,N_9261);
nand U10880 (N_10880,N_9315,N_9127);
nand U10881 (N_10881,N_9275,N_9491);
or U10882 (N_10882,N_9655,N_9677);
nand U10883 (N_10883,N_9651,N_9777);
nor U10884 (N_10884,N_9680,N_9203);
xnor U10885 (N_10885,N_9397,N_9942);
xor U10886 (N_10886,N_9279,N_9039);
nor U10887 (N_10887,N_9229,N_9704);
nor U10888 (N_10888,N_9946,N_9535);
nor U10889 (N_10889,N_9918,N_9958);
and U10890 (N_10890,N_9097,N_9664);
xor U10891 (N_10891,N_9799,N_9926);
nand U10892 (N_10892,N_9600,N_9614);
nand U10893 (N_10893,N_9395,N_9686);
nand U10894 (N_10894,N_9194,N_9105);
nor U10895 (N_10895,N_9730,N_9605);
or U10896 (N_10896,N_9881,N_9898);
nand U10897 (N_10897,N_9519,N_9041);
or U10898 (N_10898,N_9881,N_9681);
nand U10899 (N_10899,N_9170,N_9085);
or U10900 (N_10900,N_9842,N_9415);
nand U10901 (N_10901,N_9508,N_9257);
xor U10902 (N_10902,N_9443,N_9832);
xnor U10903 (N_10903,N_9508,N_9160);
xor U10904 (N_10904,N_9506,N_9244);
nand U10905 (N_10905,N_9393,N_9802);
xor U10906 (N_10906,N_9038,N_9180);
or U10907 (N_10907,N_9656,N_9076);
nand U10908 (N_10908,N_9270,N_9305);
and U10909 (N_10909,N_9712,N_9734);
and U10910 (N_10910,N_9523,N_9708);
and U10911 (N_10911,N_9583,N_9719);
or U10912 (N_10912,N_9395,N_9214);
or U10913 (N_10913,N_9784,N_9955);
or U10914 (N_10914,N_9368,N_9788);
or U10915 (N_10915,N_9367,N_9222);
nor U10916 (N_10916,N_9742,N_9805);
and U10917 (N_10917,N_9759,N_9986);
and U10918 (N_10918,N_9657,N_9224);
nor U10919 (N_10919,N_9742,N_9006);
xor U10920 (N_10920,N_9577,N_9918);
xnor U10921 (N_10921,N_9394,N_9310);
xnor U10922 (N_10922,N_9639,N_9073);
or U10923 (N_10923,N_9173,N_9193);
or U10924 (N_10924,N_9125,N_9909);
nand U10925 (N_10925,N_9684,N_9664);
or U10926 (N_10926,N_9528,N_9536);
nor U10927 (N_10927,N_9267,N_9482);
xor U10928 (N_10928,N_9942,N_9644);
or U10929 (N_10929,N_9059,N_9668);
nand U10930 (N_10930,N_9568,N_9681);
and U10931 (N_10931,N_9041,N_9324);
xnor U10932 (N_10932,N_9653,N_9071);
or U10933 (N_10933,N_9353,N_9612);
and U10934 (N_10934,N_9882,N_9096);
nand U10935 (N_10935,N_9555,N_9562);
xor U10936 (N_10936,N_9781,N_9287);
nor U10937 (N_10937,N_9129,N_9297);
and U10938 (N_10938,N_9805,N_9454);
xnor U10939 (N_10939,N_9842,N_9015);
and U10940 (N_10940,N_9187,N_9736);
nand U10941 (N_10941,N_9595,N_9403);
nor U10942 (N_10942,N_9123,N_9211);
or U10943 (N_10943,N_9742,N_9682);
nand U10944 (N_10944,N_9579,N_9347);
or U10945 (N_10945,N_9640,N_9912);
xnor U10946 (N_10946,N_9974,N_9360);
or U10947 (N_10947,N_9875,N_9137);
or U10948 (N_10948,N_9285,N_9882);
or U10949 (N_10949,N_9291,N_9347);
or U10950 (N_10950,N_9890,N_9811);
xnor U10951 (N_10951,N_9582,N_9008);
xor U10952 (N_10952,N_9218,N_9834);
and U10953 (N_10953,N_9086,N_9008);
and U10954 (N_10954,N_9912,N_9928);
and U10955 (N_10955,N_9834,N_9029);
nor U10956 (N_10956,N_9752,N_9615);
nor U10957 (N_10957,N_9159,N_9170);
or U10958 (N_10958,N_9404,N_9592);
nand U10959 (N_10959,N_9435,N_9503);
nand U10960 (N_10960,N_9951,N_9822);
nor U10961 (N_10961,N_9828,N_9419);
nor U10962 (N_10962,N_9903,N_9048);
or U10963 (N_10963,N_9670,N_9640);
or U10964 (N_10964,N_9554,N_9527);
xor U10965 (N_10965,N_9963,N_9153);
nand U10966 (N_10966,N_9895,N_9076);
nor U10967 (N_10967,N_9819,N_9211);
nor U10968 (N_10968,N_9382,N_9516);
and U10969 (N_10969,N_9022,N_9450);
xor U10970 (N_10970,N_9740,N_9719);
xor U10971 (N_10971,N_9862,N_9275);
xor U10972 (N_10972,N_9034,N_9783);
xor U10973 (N_10973,N_9308,N_9621);
or U10974 (N_10974,N_9905,N_9167);
or U10975 (N_10975,N_9884,N_9859);
and U10976 (N_10976,N_9500,N_9721);
xnor U10977 (N_10977,N_9926,N_9416);
and U10978 (N_10978,N_9039,N_9057);
xnor U10979 (N_10979,N_9367,N_9015);
xor U10980 (N_10980,N_9544,N_9950);
nor U10981 (N_10981,N_9665,N_9361);
or U10982 (N_10982,N_9011,N_9344);
xor U10983 (N_10983,N_9858,N_9149);
nand U10984 (N_10984,N_9019,N_9741);
xor U10985 (N_10985,N_9759,N_9727);
xor U10986 (N_10986,N_9328,N_9468);
and U10987 (N_10987,N_9311,N_9197);
or U10988 (N_10988,N_9461,N_9222);
and U10989 (N_10989,N_9698,N_9588);
xnor U10990 (N_10990,N_9499,N_9190);
xnor U10991 (N_10991,N_9199,N_9882);
nand U10992 (N_10992,N_9575,N_9253);
and U10993 (N_10993,N_9363,N_9436);
nand U10994 (N_10994,N_9082,N_9890);
nand U10995 (N_10995,N_9777,N_9377);
nand U10996 (N_10996,N_9870,N_9734);
and U10997 (N_10997,N_9605,N_9252);
or U10998 (N_10998,N_9843,N_9342);
nor U10999 (N_10999,N_9780,N_9159);
or U11000 (N_11000,N_10121,N_10859);
and U11001 (N_11001,N_10348,N_10191);
and U11002 (N_11002,N_10056,N_10262);
nor U11003 (N_11003,N_10940,N_10171);
or U11004 (N_11004,N_10016,N_10196);
xor U11005 (N_11005,N_10584,N_10494);
xnor U11006 (N_11006,N_10589,N_10913);
or U11007 (N_11007,N_10547,N_10299);
nand U11008 (N_11008,N_10294,N_10054);
or U11009 (N_11009,N_10004,N_10855);
nor U11010 (N_11010,N_10057,N_10212);
xnor U11011 (N_11011,N_10027,N_10558);
nand U11012 (N_11012,N_10883,N_10879);
nor U11013 (N_11013,N_10190,N_10894);
nor U11014 (N_11014,N_10169,N_10798);
nor U11015 (N_11015,N_10346,N_10587);
xnor U11016 (N_11016,N_10642,N_10469);
xnor U11017 (N_11017,N_10683,N_10555);
nor U11018 (N_11018,N_10439,N_10356);
xnor U11019 (N_11019,N_10824,N_10733);
nand U11020 (N_11020,N_10843,N_10691);
nand U11021 (N_11021,N_10290,N_10833);
and U11022 (N_11022,N_10247,N_10267);
or U11023 (N_11023,N_10856,N_10631);
nor U11024 (N_11024,N_10624,N_10882);
nor U11025 (N_11025,N_10918,N_10523);
nand U11026 (N_11026,N_10662,N_10166);
or U11027 (N_11027,N_10310,N_10285);
nor U11028 (N_11028,N_10092,N_10484);
and U11029 (N_11029,N_10716,N_10134);
xor U11030 (N_11030,N_10556,N_10569);
nand U11031 (N_11031,N_10214,N_10643);
nand U11032 (N_11032,N_10152,N_10229);
or U11033 (N_11033,N_10826,N_10983);
nor U11034 (N_11034,N_10660,N_10493);
nand U11035 (N_11035,N_10546,N_10641);
nand U11036 (N_11036,N_10270,N_10693);
nand U11037 (N_11037,N_10974,N_10891);
xor U11038 (N_11038,N_10761,N_10566);
nor U11039 (N_11039,N_10135,N_10545);
or U11040 (N_11040,N_10963,N_10034);
xor U11041 (N_11041,N_10321,N_10750);
nor U11042 (N_11042,N_10404,N_10551);
or U11043 (N_11043,N_10314,N_10610);
and U11044 (N_11044,N_10123,N_10242);
xor U11045 (N_11045,N_10707,N_10271);
xor U11046 (N_11046,N_10007,N_10260);
and U11047 (N_11047,N_10591,N_10451);
or U11048 (N_11048,N_10769,N_10601);
and U11049 (N_11049,N_10722,N_10064);
and U11050 (N_11050,N_10920,N_10301);
and U11051 (N_11051,N_10175,N_10654);
xnor U11052 (N_11052,N_10470,N_10032);
nand U11053 (N_11053,N_10863,N_10485);
xnor U11054 (N_11054,N_10747,N_10553);
xor U11055 (N_11055,N_10905,N_10185);
and U11056 (N_11056,N_10099,N_10415);
nor U11057 (N_11057,N_10802,N_10880);
nor U11058 (N_11058,N_10120,N_10046);
and U11059 (N_11059,N_10052,N_10808);
xnor U11060 (N_11060,N_10122,N_10237);
xor U11061 (N_11061,N_10816,N_10932);
or U11062 (N_11062,N_10164,N_10038);
and U11063 (N_11063,N_10605,N_10825);
xor U11064 (N_11064,N_10792,N_10499);
xnor U11065 (N_11065,N_10765,N_10162);
nand U11066 (N_11066,N_10414,N_10155);
nor U11067 (N_11067,N_10972,N_10560);
nor U11068 (N_11068,N_10305,N_10534);
or U11069 (N_11069,N_10538,N_10519);
xnor U11070 (N_11070,N_10869,N_10784);
and U11071 (N_11071,N_10465,N_10078);
and U11072 (N_11072,N_10724,N_10363);
nor U11073 (N_11073,N_10364,N_10280);
xor U11074 (N_11074,N_10741,N_10243);
xnor U11075 (N_11075,N_10331,N_10180);
nand U11076 (N_11076,N_10460,N_10987);
nand U11077 (N_11077,N_10089,N_10139);
xnor U11078 (N_11078,N_10150,N_10458);
or U11079 (N_11079,N_10514,N_10115);
nor U11080 (N_11080,N_10725,N_10844);
nand U11081 (N_11081,N_10144,N_10946);
nor U11082 (N_11082,N_10984,N_10791);
and U11083 (N_11083,N_10500,N_10355);
and U11084 (N_11084,N_10788,N_10621);
or U11085 (N_11085,N_10708,N_10885);
xor U11086 (N_11086,N_10362,N_10837);
xor U11087 (N_11087,N_10320,N_10228);
nor U11088 (N_11088,N_10359,N_10506);
nor U11089 (N_11089,N_10933,N_10223);
nor U11090 (N_11090,N_10187,N_10496);
and U11091 (N_11091,N_10440,N_10877);
or U11092 (N_11092,N_10945,N_10737);
xnor U11093 (N_11093,N_10774,N_10955);
nand U11094 (N_11094,N_10995,N_10090);
and U11095 (N_11095,N_10585,N_10073);
nor U11096 (N_11096,N_10559,N_10491);
or U11097 (N_11097,N_10950,N_10338);
nor U11098 (N_11098,N_10618,N_10755);
and U11099 (N_11099,N_10322,N_10518);
and U11100 (N_11100,N_10628,N_10517);
nand U11101 (N_11101,N_10960,N_10680);
nand U11102 (N_11102,N_10537,N_10671);
and U11103 (N_11103,N_10197,N_10463);
and U11104 (N_11104,N_10973,N_10633);
nor U11105 (N_11105,N_10608,N_10350);
nand U11106 (N_11106,N_10498,N_10582);
and U11107 (N_11107,N_10173,N_10893);
nand U11108 (N_11108,N_10847,N_10248);
or U11109 (N_11109,N_10095,N_10809);
nor U11110 (N_11110,N_10873,N_10726);
nand U11111 (N_11111,N_10065,N_10676);
xor U11112 (N_11112,N_10563,N_10783);
and U11113 (N_11113,N_10668,N_10780);
or U11114 (N_11114,N_10813,N_10249);
nor U11115 (N_11115,N_10025,N_10851);
nor U11116 (N_11116,N_10614,N_10335);
or U11117 (N_11117,N_10207,N_10927);
nand U11118 (N_11118,N_10926,N_10282);
xor U11119 (N_11119,N_10764,N_10368);
nand U11120 (N_11120,N_10029,N_10293);
and U11121 (N_11121,N_10533,N_10374);
or U11122 (N_11122,N_10836,N_10705);
nor U11123 (N_11123,N_10107,N_10232);
nand U11124 (N_11124,N_10990,N_10612);
and U11125 (N_11125,N_10970,N_10323);
and U11126 (N_11126,N_10745,N_10377);
xnor U11127 (N_11127,N_10692,N_10637);
or U11128 (N_11128,N_10669,N_10111);
or U11129 (N_11129,N_10014,N_10403);
xnor U11130 (N_11130,N_10428,N_10565);
and U11131 (N_11131,N_10698,N_10209);
nor U11132 (N_11132,N_10200,N_10001);
nor U11133 (N_11133,N_10874,N_10748);
xnor U11134 (N_11134,N_10406,N_10319);
nor U11135 (N_11135,N_10762,N_10831);
or U11136 (N_11136,N_10682,N_10838);
nor U11137 (N_11137,N_10689,N_10898);
nand U11138 (N_11138,N_10245,N_10867);
xnor U11139 (N_11139,N_10807,N_10396);
or U11140 (N_11140,N_10532,N_10444);
or U11141 (N_11141,N_10039,N_10017);
nand U11142 (N_11142,N_10679,N_10806);
and U11143 (N_11143,N_10550,N_10982);
or U11144 (N_11144,N_10609,N_10199);
nand U11145 (N_11145,N_10649,N_10723);
nand U11146 (N_11146,N_10407,N_10220);
xor U11147 (N_11147,N_10467,N_10326);
nor U11148 (N_11148,N_10571,N_10944);
xnor U11149 (N_11149,N_10929,N_10760);
xnor U11150 (N_11150,N_10006,N_10971);
or U11151 (N_11151,N_10210,N_10178);
nand U11152 (N_11152,N_10370,N_10276);
nand U11153 (N_11153,N_10749,N_10481);
nor U11154 (N_11154,N_10670,N_10316);
nor U11155 (N_11155,N_10848,N_10263);
nor U11156 (N_11156,N_10344,N_10184);
nor U11157 (N_11157,N_10174,N_10975);
nor U11158 (N_11158,N_10888,N_10706);
nor U11159 (N_11159,N_10508,N_10098);
and U11160 (N_11160,N_10083,N_10112);
nor U11161 (N_11161,N_10697,N_10858);
nand U11162 (N_11162,N_10509,N_10640);
nor U11163 (N_11163,N_10217,N_10058);
nand U11164 (N_11164,N_10603,N_10731);
or U11165 (N_11165,N_10839,N_10230);
nor U11166 (N_11166,N_10077,N_10024);
or U11167 (N_11167,N_10154,N_10390);
nor U11168 (N_11168,N_10980,N_10163);
nor U11169 (N_11169,N_10158,N_10512);
xor U11170 (N_11170,N_10258,N_10186);
or U11171 (N_11171,N_10810,N_10688);
or U11172 (N_11172,N_10834,N_10992);
xnor U11173 (N_11173,N_10069,N_10629);
and U11174 (N_11174,N_10796,N_10795);
nor U11175 (N_11175,N_10529,N_10264);
and U11176 (N_11176,N_10195,N_10794);
nor U11177 (N_11177,N_10578,N_10181);
or U11178 (N_11178,N_10579,N_10019);
nand U11179 (N_11179,N_10959,N_10372);
or U11180 (N_11180,N_10213,N_10125);
and U11181 (N_11181,N_10653,N_10446);
xor U11182 (N_11182,N_10424,N_10160);
nand U11183 (N_11183,N_10488,N_10543);
and U11184 (N_11184,N_10829,N_10211);
nand U11185 (N_11185,N_10332,N_10906);
nand U11186 (N_11186,N_10567,N_10619);
and U11187 (N_11187,N_10872,N_10703);
nor U11188 (N_11188,N_10473,N_10165);
xor U11189 (N_11189,N_10957,N_10080);
nor U11190 (N_11190,N_10070,N_10744);
or U11191 (N_11191,N_10227,N_10105);
nor U11192 (N_11192,N_10743,N_10457);
nand U11193 (N_11193,N_10934,N_10076);
and U11194 (N_11194,N_10193,N_10352);
xnor U11195 (N_11195,N_10137,N_10239);
nand U11196 (N_11196,N_10079,N_10549);
and U11197 (N_11197,N_10511,N_10763);
nor U11198 (N_11198,N_10395,N_10298);
nand U11199 (N_11199,N_10430,N_10994);
xor U11200 (N_11200,N_10557,N_10900);
nor U11201 (N_11201,N_10988,N_10084);
nor U11202 (N_11202,N_10272,N_10667);
and U11203 (N_11203,N_10754,N_10066);
and U11204 (N_11204,N_10339,N_10379);
nor U11205 (N_11205,N_10235,N_10384);
nand U11206 (N_11206,N_10376,N_10266);
and U11207 (N_11207,N_10148,N_10275);
xor U11208 (N_11208,N_10542,N_10846);
or U11209 (N_11209,N_10766,N_10909);
or U11210 (N_11210,N_10194,N_10255);
and U11211 (N_11211,N_10868,N_10022);
nor U11212 (N_11212,N_10450,N_10206);
nand U11213 (N_11213,N_10313,N_10520);
xnor U11214 (N_11214,N_10562,N_10081);
nand U11215 (N_11215,N_10536,N_10952);
or U11216 (N_11216,N_10059,N_10947);
xnor U11217 (N_11217,N_10307,N_10234);
xor U11218 (N_11218,N_10935,N_10416);
or U11219 (N_11219,N_10840,N_10333);
nor U11220 (N_11220,N_10966,N_10773);
nand U11221 (N_11221,N_10772,N_10422);
or U11222 (N_11222,N_10149,N_10035);
and U11223 (N_11223,N_10969,N_10871);
or U11224 (N_11224,N_10013,N_10759);
or U11225 (N_11225,N_10854,N_10437);
or U11226 (N_11226,N_10675,N_10739);
or U11227 (N_11227,N_10367,N_10596);
and U11228 (N_11228,N_10832,N_10008);
and U11229 (N_11229,N_10903,N_10391);
xnor U11230 (N_11230,N_10189,N_10702);
or U11231 (N_11231,N_10526,N_10231);
nand U11232 (N_11232,N_10811,N_10746);
and U11233 (N_11233,N_10296,N_10658);
xnor U11234 (N_11234,N_10890,N_10131);
nor U11235 (N_11235,N_10548,N_10286);
or U11236 (N_11236,N_10409,N_10274);
nor U11237 (N_11237,N_10283,N_10712);
or U11238 (N_11238,N_10521,N_10928);
or U11239 (N_11239,N_10522,N_10177);
xnor U11240 (N_11240,N_10954,N_10126);
nor U11241 (N_11241,N_10878,N_10815);
or U11242 (N_11242,N_10049,N_10434);
and U11243 (N_11243,N_10828,N_10742);
nor U11244 (N_11244,N_10138,N_10447);
or U11245 (N_11245,N_10435,N_10799);
nand U11246 (N_11246,N_10334,N_10487);
nor U11247 (N_11247,N_10292,N_10208);
nand U11248 (N_11248,N_10156,N_10876);
and U11249 (N_11249,N_10328,N_10136);
or U11250 (N_11250,N_10330,N_10023);
or U11251 (N_11251,N_10480,N_10251);
nand U11252 (N_11252,N_10651,N_10425);
xor U11253 (N_11253,N_10870,N_10393);
or U11254 (N_11254,N_10686,N_10461);
nor U11255 (N_11255,N_10100,N_10622);
nand U11256 (N_11256,N_10524,N_10866);
xor U11257 (N_11257,N_10785,N_10456);
nor U11258 (N_11258,N_10564,N_10398);
nor U11259 (N_11259,N_10597,N_10875);
or U11260 (N_11260,N_10357,N_10613);
xnor U11261 (N_11261,N_10516,N_10454);
and U11262 (N_11262,N_10224,N_10925);
nand U11263 (N_11263,N_10701,N_10340);
and U11264 (N_11264,N_10102,N_10704);
nand U11265 (N_11265,N_10071,N_10110);
nand U11266 (N_11266,N_10586,N_10392);
or U11267 (N_11267,N_10233,N_10647);
nor U11268 (N_11268,N_10418,N_10561);
and U11269 (N_11269,N_10400,N_10273);
or U11270 (N_11270,N_10161,N_10719);
xor U11271 (N_11271,N_10114,N_10221);
xor U11272 (N_11272,N_10599,N_10721);
and U11273 (N_11273,N_10623,N_10575);
nor U11274 (N_11274,N_10801,N_10303);
nor U11275 (N_11275,N_10976,N_10606);
nor U11276 (N_11276,N_10665,N_10044);
or U11277 (N_11277,N_10817,N_10318);
nand U11278 (N_11278,N_10103,N_10779);
nor U11279 (N_11279,N_10311,N_10009);
and U11280 (N_11280,N_10767,N_10188);
and U11281 (N_11281,N_10690,N_10297);
or U11282 (N_11282,N_10617,N_10652);
or U11283 (N_11283,N_10474,N_10709);
and U11284 (N_11284,N_10343,N_10486);
and U11285 (N_11285,N_10087,N_10803);
and U11286 (N_11286,N_10735,N_10075);
nand U11287 (N_11287,N_10253,N_10588);
and U11288 (N_11288,N_10615,N_10300);
or U11289 (N_11289,N_10632,N_10666);
and U11290 (N_11290,N_10345,N_10897);
nor U11291 (N_11291,N_10715,N_10968);
nor U11292 (N_11292,N_10659,N_10892);
nor U11293 (N_11293,N_10673,N_10375);
xor U11294 (N_11294,N_10572,N_10431);
and U11295 (N_11295,N_10937,N_10389);
xor U11296 (N_11296,N_10677,N_10961);
nor U11297 (N_11297,N_10124,N_10861);
or U11298 (N_11298,N_10663,N_10074);
or U11299 (N_11299,N_10886,N_10091);
or U11300 (N_11300,N_10661,N_10590);
or U11301 (N_11301,N_10604,N_10602);
and U11302 (N_11302,N_10192,N_10132);
nor U11303 (N_11303,N_10408,N_10468);
nor U11304 (N_11304,N_10351,N_10449);
xnor U11305 (N_11305,N_10895,N_10205);
and U11306 (N_11306,N_10466,N_10452);
xnor U11307 (N_11307,N_10462,N_10055);
nand U11308 (N_11308,N_10713,N_10655);
or U11309 (N_11309,N_10002,N_10645);
and U11310 (N_11310,N_10315,N_10381);
or U11311 (N_11311,N_10864,N_10353);
nor U11312 (N_11312,N_10684,N_10789);
xnor U11313 (N_11313,N_10770,N_10053);
xnor U11314 (N_11314,N_10953,N_10306);
nor U11315 (N_11315,N_10203,N_10061);
nor U11316 (N_11316,N_10687,N_10729);
and U11317 (N_11317,N_10291,N_10931);
nand U11318 (N_11318,N_10003,N_10246);
nor U11319 (N_11319,N_10845,N_10327);
nand U11320 (N_11320,N_10956,N_10261);
and U11321 (N_11321,N_10777,N_10042);
nand U11322 (N_11322,N_10483,N_10265);
or U11323 (N_11323,N_10085,N_10951);
nor U11324 (N_11324,N_10063,N_10600);
nand U11325 (N_11325,N_10401,N_10495);
xnor U11326 (N_11326,N_10097,N_10753);
and U11327 (N_11327,N_10086,N_10256);
nand U11328 (N_11328,N_10639,N_10540);
nand U11329 (N_11329,N_10453,N_10108);
nand U11330 (N_11330,N_10657,N_10751);
or U11331 (N_11331,N_10930,N_10371);
nor U11332 (N_11332,N_10413,N_10325);
or U11333 (N_11333,N_10051,N_10577);
and U11334 (N_11334,N_10732,N_10923);
xnor U11335 (N_11335,N_10781,N_10917);
or U11336 (N_11336,N_10238,N_10907);
or U11337 (N_11337,N_10436,N_10943);
xor U11338 (N_11338,N_10423,N_10426);
xor U11339 (N_11339,N_10151,N_10530);
or U11340 (N_11340,N_10989,N_10459);
nor U11341 (N_11341,N_10030,N_10922);
and U11342 (N_11342,N_10910,N_10941);
nor U11343 (N_11343,N_10116,N_10268);
xnor U11344 (N_11344,N_10889,N_10887);
nor U11345 (N_11345,N_10373,N_10202);
and U11346 (N_11346,N_10118,N_10849);
nor U11347 (N_11347,N_10996,N_10040);
and U11348 (N_11348,N_10427,N_10443);
nor U11349 (N_11349,N_10634,N_10620);
nor U11350 (N_11350,N_10072,N_10958);
nand U11351 (N_11351,N_10005,N_10757);
and U11352 (N_11352,N_10638,N_10172);
xor U11353 (N_11353,N_10636,N_10860);
nand U11354 (N_11354,N_10841,N_10397);
and U11355 (N_11355,N_10857,N_10096);
nor U11356 (N_11356,N_10936,N_10020);
nor U11357 (N_11357,N_10365,N_10717);
xor U11358 (N_11358,N_10513,N_10576);
nand U11359 (N_11359,N_10573,N_10685);
or U11360 (N_11360,N_10539,N_10380);
xor U11361 (N_11361,N_10093,N_10625);
nor U11362 (N_11362,N_10011,N_10758);
and U11363 (N_11363,N_10349,N_10361);
and U11364 (N_11364,N_10026,N_10244);
nor U11365 (N_11365,N_10101,N_10354);
and U11366 (N_11366,N_10962,N_10616);
nor U11367 (N_11367,N_10018,N_10552);
or U11368 (N_11368,N_10948,N_10800);
nor U11369 (N_11369,N_10583,N_10501);
xnor U11370 (N_11370,N_10050,N_10793);
or U11371 (N_11371,N_10535,N_10015);
nor U11372 (N_11372,N_10225,N_10598);
xor U11373 (N_11373,N_10711,N_10700);
and U11374 (N_11374,N_10412,N_10145);
xnor U11375 (N_11375,N_10835,N_10646);
nor U11376 (N_11376,N_10790,N_10241);
nand U11377 (N_11377,N_10341,N_10916);
nor U11378 (N_11378,N_10921,N_10644);
or U11379 (N_11379,N_10312,N_10896);
xor U11380 (N_11380,N_10419,N_10510);
nand U11381 (N_11381,N_10595,N_10295);
xnor U11382 (N_11382,N_10385,N_10106);
nand U11383 (N_11383,N_10288,N_10525);
nand U11384 (N_11384,N_10257,N_10287);
nor U11385 (N_11385,N_10067,N_10915);
and U11386 (N_11386,N_10279,N_10147);
nand U11387 (N_11387,N_10942,N_10977);
or U11388 (N_11388,N_10738,N_10140);
xnor U11389 (N_11389,N_10218,N_10489);
nand U11390 (N_11390,N_10219,N_10159);
or U11391 (N_11391,N_10281,N_10429);
nor U11392 (N_11392,N_10730,N_10033);
xor U11393 (N_11393,N_10421,N_10455);
xnor U11394 (N_11394,N_10981,N_10047);
nand U11395 (N_11395,N_10236,N_10476);
and U11396 (N_11396,N_10304,N_10507);
and U11397 (N_11397,N_10417,N_10497);
or U11398 (N_11398,N_10531,N_10277);
and U11399 (N_11399,N_10475,N_10527);
xor U11400 (N_11400,N_10490,N_10574);
or U11401 (N_11401,N_10502,N_10993);
nand U11402 (N_11402,N_10949,N_10986);
nor U11403 (N_11403,N_10394,N_10939);
nor U11404 (N_11404,N_10985,N_10329);
xnor U11405 (N_11405,N_10010,N_10317);
nor U11406 (N_11406,N_10179,N_10037);
and U11407 (N_11407,N_10778,N_10648);
nand U11408 (N_11408,N_10768,N_10182);
nand U11409 (N_11409,N_10805,N_10146);
nor U11410 (N_11410,N_10544,N_10541);
nor U11411 (N_11411,N_10388,N_10143);
xor U11412 (N_11412,N_10852,N_10342);
and U11413 (N_11413,N_10133,N_10382);
nor U11414 (N_11414,N_10782,N_10028);
and U11415 (N_11415,N_10911,N_10109);
and U11416 (N_11416,N_10674,N_10471);
nor U11417 (N_11417,N_10853,N_10336);
xnor U11418 (N_11418,N_10804,N_10681);
nor U11419 (N_11419,N_10254,N_10324);
nor U11420 (N_11420,N_10635,N_10611);
xnor U11421 (N_11421,N_10000,N_10360);
or U11422 (N_11422,N_10464,N_10756);
nand U11423 (N_11423,N_10710,N_10119);
and U11424 (N_11424,N_10786,N_10515);
or U11425 (N_11425,N_10998,N_10830);
and U11426 (N_11426,N_10127,N_10978);
and U11427 (N_11427,N_10031,N_10630);
and U11428 (N_11428,N_10420,N_10865);
nand U11429 (N_11429,N_10378,N_10899);
and U11430 (N_11430,N_10167,N_10593);
nand U11431 (N_11431,N_10492,N_10302);
and U11432 (N_11432,N_10201,N_10736);
and U11433 (N_11433,N_10399,N_10337);
and U11434 (N_11434,N_10222,N_10997);
and U11435 (N_11435,N_10062,N_10405);
and U11436 (N_11436,N_10694,N_10820);
and U11437 (N_11437,N_10850,N_10402);
or U11438 (N_11438,N_10358,N_10908);
nand U11439 (N_11439,N_10938,N_10814);
and U11440 (N_11440,N_10226,N_10442);
nand U11441 (N_11441,N_10479,N_10130);
nand U11442 (N_11442,N_10478,N_10818);
nor U11443 (N_11443,N_10088,N_10043);
or U11444 (N_11444,N_10902,N_10819);
nor U11445 (N_11445,N_10664,N_10752);
nor U11446 (N_11446,N_10259,N_10433);
xor U11447 (N_11447,N_10441,N_10884);
and U11448 (N_11448,N_10776,N_10432);
xor U11449 (N_11449,N_10142,N_10965);
nor U11450 (N_11450,N_10472,N_10369);
xnor U11451 (N_11451,N_10964,N_10627);
xor U11452 (N_11452,N_10215,N_10771);
xnor U11453 (N_11453,N_10387,N_10924);
or U11454 (N_11454,N_10672,N_10528);
and U11455 (N_11455,N_10504,N_10157);
nand U11456 (N_11456,N_10117,N_10216);
nor U11457 (N_11457,N_10740,N_10036);
nand U11458 (N_11458,N_10822,N_10082);
or U11459 (N_11459,N_10411,N_10250);
xor U11460 (N_11460,N_10176,N_10198);
or U11461 (N_11461,N_10170,N_10678);
and U11462 (N_11462,N_10594,N_10045);
and U11463 (N_11463,N_10386,N_10581);
nor U11464 (N_11464,N_10570,N_10862);
nand U11465 (N_11465,N_10204,N_10580);
and U11466 (N_11466,N_10812,N_10823);
and U11467 (N_11467,N_10309,N_10068);
nand U11468 (N_11468,N_10503,N_10094);
nand U11469 (N_11469,N_10012,N_10881);
or U11470 (N_11470,N_10048,N_10021);
or U11471 (N_11471,N_10141,N_10289);
xor U11472 (N_11472,N_10797,N_10278);
and U11473 (N_11473,N_10183,N_10104);
xnor U11474 (N_11474,N_10060,N_10477);
xor U11475 (N_11475,N_10728,N_10979);
xnor U11476 (N_11476,N_10448,N_10113);
xnor U11477 (N_11477,N_10699,N_10714);
and U11478 (N_11478,N_10269,N_10718);
xor U11479 (N_11479,N_10967,N_10252);
and U11480 (N_11480,N_10347,N_10383);
nor U11481 (N_11481,N_10650,N_10153);
and U11482 (N_11482,N_10787,N_10240);
xor U11483 (N_11483,N_10129,N_10919);
nand U11484 (N_11484,N_10914,N_10308);
and U11485 (N_11485,N_10991,N_10901);
and U11486 (N_11486,N_10592,N_10482);
or U11487 (N_11487,N_10842,N_10284);
nor U11488 (N_11488,N_10999,N_10438);
nor U11489 (N_11489,N_10727,N_10168);
and U11490 (N_11490,N_10445,N_10626);
nand U11491 (N_11491,N_10912,N_10696);
and U11492 (N_11492,N_10720,N_10041);
nor U11493 (N_11493,N_10827,N_10821);
nand U11494 (N_11494,N_10904,N_10607);
and U11495 (N_11495,N_10695,N_10775);
or U11496 (N_11496,N_10656,N_10366);
xor U11497 (N_11497,N_10568,N_10128);
or U11498 (N_11498,N_10410,N_10554);
xnor U11499 (N_11499,N_10505,N_10734);
nand U11500 (N_11500,N_10134,N_10026);
nor U11501 (N_11501,N_10052,N_10834);
or U11502 (N_11502,N_10608,N_10584);
nand U11503 (N_11503,N_10320,N_10413);
nand U11504 (N_11504,N_10639,N_10201);
nor U11505 (N_11505,N_10727,N_10777);
and U11506 (N_11506,N_10715,N_10230);
nand U11507 (N_11507,N_10903,N_10002);
nor U11508 (N_11508,N_10260,N_10012);
nand U11509 (N_11509,N_10167,N_10140);
and U11510 (N_11510,N_10809,N_10980);
xor U11511 (N_11511,N_10854,N_10783);
and U11512 (N_11512,N_10524,N_10779);
xnor U11513 (N_11513,N_10081,N_10854);
nor U11514 (N_11514,N_10662,N_10598);
nor U11515 (N_11515,N_10757,N_10334);
nand U11516 (N_11516,N_10680,N_10941);
and U11517 (N_11517,N_10371,N_10013);
and U11518 (N_11518,N_10756,N_10660);
or U11519 (N_11519,N_10017,N_10710);
or U11520 (N_11520,N_10639,N_10353);
or U11521 (N_11521,N_10327,N_10822);
or U11522 (N_11522,N_10270,N_10861);
nand U11523 (N_11523,N_10885,N_10335);
or U11524 (N_11524,N_10529,N_10781);
nor U11525 (N_11525,N_10367,N_10024);
and U11526 (N_11526,N_10440,N_10301);
and U11527 (N_11527,N_10322,N_10692);
xor U11528 (N_11528,N_10786,N_10758);
xor U11529 (N_11529,N_10035,N_10503);
xnor U11530 (N_11530,N_10279,N_10910);
nand U11531 (N_11531,N_10230,N_10870);
nand U11532 (N_11532,N_10720,N_10974);
nor U11533 (N_11533,N_10922,N_10977);
nand U11534 (N_11534,N_10313,N_10196);
nand U11535 (N_11535,N_10058,N_10256);
nand U11536 (N_11536,N_10160,N_10757);
nand U11537 (N_11537,N_10148,N_10302);
or U11538 (N_11538,N_10680,N_10041);
nand U11539 (N_11539,N_10475,N_10994);
nor U11540 (N_11540,N_10388,N_10402);
nor U11541 (N_11541,N_10242,N_10158);
xnor U11542 (N_11542,N_10704,N_10028);
xnor U11543 (N_11543,N_10684,N_10662);
nand U11544 (N_11544,N_10111,N_10153);
nor U11545 (N_11545,N_10730,N_10155);
and U11546 (N_11546,N_10046,N_10380);
nand U11547 (N_11547,N_10779,N_10700);
xnor U11548 (N_11548,N_10542,N_10212);
xor U11549 (N_11549,N_10666,N_10261);
and U11550 (N_11550,N_10577,N_10777);
nor U11551 (N_11551,N_10602,N_10757);
and U11552 (N_11552,N_10474,N_10747);
or U11553 (N_11553,N_10787,N_10058);
xnor U11554 (N_11554,N_10059,N_10781);
and U11555 (N_11555,N_10193,N_10332);
or U11556 (N_11556,N_10527,N_10804);
and U11557 (N_11557,N_10365,N_10887);
and U11558 (N_11558,N_10535,N_10455);
and U11559 (N_11559,N_10425,N_10217);
or U11560 (N_11560,N_10227,N_10515);
xor U11561 (N_11561,N_10968,N_10117);
and U11562 (N_11562,N_10252,N_10332);
or U11563 (N_11563,N_10879,N_10473);
nand U11564 (N_11564,N_10425,N_10055);
xnor U11565 (N_11565,N_10245,N_10104);
xor U11566 (N_11566,N_10064,N_10895);
and U11567 (N_11567,N_10578,N_10569);
xnor U11568 (N_11568,N_10185,N_10256);
and U11569 (N_11569,N_10225,N_10505);
xor U11570 (N_11570,N_10430,N_10234);
nand U11571 (N_11571,N_10248,N_10532);
nand U11572 (N_11572,N_10612,N_10188);
and U11573 (N_11573,N_10671,N_10478);
xor U11574 (N_11574,N_10987,N_10891);
or U11575 (N_11575,N_10781,N_10395);
or U11576 (N_11576,N_10233,N_10298);
and U11577 (N_11577,N_10113,N_10201);
xnor U11578 (N_11578,N_10686,N_10533);
or U11579 (N_11579,N_10144,N_10715);
nand U11580 (N_11580,N_10828,N_10055);
xor U11581 (N_11581,N_10118,N_10003);
nand U11582 (N_11582,N_10057,N_10956);
and U11583 (N_11583,N_10011,N_10858);
nand U11584 (N_11584,N_10691,N_10296);
or U11585 (N_11585,N_10822,N_10566);
nor U11586 (N_11586,N_10189,N_10598);
nor U11587 (N_11587,N_10014,N_10152);
and U11588 (N_11588,N_10145,N_10747);
nor U11589 (N_11589,N_10033,N_10014);
nand U11590 (N_11590,N_10974,N_10563);
nor U11591 (N_11591,N_10252,N_10216);
nand U11592 (N_11592,N_10011,N_10310);
or U11593 (N_11593,N_10560,N_10583);
and U11594 (N_11594,N_10317,N_10701);
and U11595 (N_11595,N_10089,N_10558);
nor U11596 (N_11596,N_10798,N_10805);
xor U11597 (N_11597,N_10360,N_10447);
or U11598 (N_11598,N_10423,N_10009);
nand U11599 (N_11599,N_10165,N_10260);
and U11600 (N_11600,N_10619,N_10074);
nor U11601 (N_11601,N_10378,N_10752);
xor U11602 (N_11602,N_10843,N_10526);
nor U11603 (N_11603,N_10744,N_10752);
nor U11604 (N_11604,N_10765,N_10528);
nand U11605 (N_11605,N_10475,N_10124);
or U11606 (N_11606,N_10652,N_10508);
or U11607 (N_11607,N_10324,N_10494);
nor U11608 (N_11608,N_10550,N_10922);
nand U11609 (N_11609,N_10396,N_10570);
xor U11610 (N_11610,N_10848,N_10976);
xnor U11611 (N_11611,N_10647,N_10503);
or U11612 (N_11612,N_10061,N_10262);
nor U11613 (N_11613,N_10681,N_10769);
nand U11614 (N_11614,N_10948,N_10449);
xor U11615 (N_11615,N_10456,N_10339);
xor U11616 (N_11616,N_10145,N_10667);
nand U11617 (N_11617,N_10536,N_10543);
and U11618 (N_11618,N_10315,N_10529);
or U11619 (N_11619,N_10239,N_10761);
nand U11620 (N_11620,N_10797,N_10779);
xnor U11621 (N_11621,N_10469,N_10290);
and U11622 (N_11622,N_10645,N_10710);
nand U11623 (N_11623,N_10551,N_10887);
and U11624 (N_11624,N_10379,N_10632);
or U11625 (N_11625,N_10862,N_10529);
and U11626 (N_11626,N_10056,N_10562);
and U11627 (N_11627,N_10153,N_10529);
and U11628 (N_11628,N_10002,N_10759);
xnor U11629 (N_11629,N_10728,N_10209);
and U11630 (N_11630,N_10174,N_10195);
nand U11631 (N_11631,N_10439,N_10811);
or U11632 (N_11632,N_10884,N_10586);
or U11633 (N_11633,N_10714,N_10402);
nand U11634 (N_11634,N_10035,N_10359);
or U11635 (N_11635,N_10335,N_10254);
nor U11636 (N_11636,N_10254,N_10215);
and U11637 (N_11637,N_10418,N_10449);
nand U11638 (N_11638,N_10702,N_10673);
or U11639 (N_11639,N_10962,N_10403);
xnor U11640 (N_11640,N_10442,N_10219);
nor U11641 (N_11641,N_10349,N_10003);
and U11642 (N_11642,N_10610,N_10085);
nand U11643 (N_11643,N_10697,N_10902);
or U11644 (N_11644,N_10042,N_10818);
xor U11645 (N_11645,N_10608,N_10565);
and U11646 (N_11646,N_10885,N_10971);
or U11647 (N_11647,N_10016,N_10863);
xnor U11648 (N_11648,N_10145,N_10900);
xor U11649 (N_11649,N_10557,N_10737);
nor U11650 (N_11650,N_10731,N_10613);
xnor U11651 (N_11651,N_10889,N_10671);
or U11652 (N_11652,N_10952,N_10310);
xnor U11653 (N_11653,N_10177,N_10902);
or U11654 (N_11654,N_10192,N_10680);
nor U11655 (N_11655,N_10468,N_10828);
nor U11656 (N_11656,N_10652,N_10325);
nand U11657 (N_11657,N_10478,N_10369);
nor U11658 (N_11658,N_10134,N_10807);
nor U11659 (N_11659,N_10078,N_10646);
nand U11660 (N_11660,N_10225,N_10093);
or U11661 (N_11661,N_10884,N_10005);
and U11662 (N_11662,N_10649,N_10185);
nor U11663 (N_11663,N_10341,N_10258);
nand U11664 (N_11664,N_10532,N_10158);
xnor U11665 (N_11665,N_10307,N_10877);
or U11666 (N_11666,N_10104,N_10603);
and U11667 (N_11667,N_10555,N_10102);
and U11668 (N_11668,N_10356,N_10584);
xor U11669 (N_11669,N_10924,N_10260);
nand U11670 (N_11670,N_10205,N_10218);
nand U11671 (N_11671,N_10153,N_10595);
or U11672 (N_11672,N_10857,N_10251);
nand U11673 (N_11673,N_10951,N_10703);
nand U11674 (N_11674,N_10489,N_10569);
or U11675 (N_11675,N_10349,N_10643);
nor U11676 (N_11676,N_10163,N_10199);
or U11677 (N_11677,N_10415,N_10579);
xnor U11678 (N_11678,N_10958,N_10257);
xor U11679 (N_11679,N_10725,N_10342);
nand U11680 (N_11680,N_10802,N_10680);
xnor U11681 (N_11681,N_10072,N_10826);
or U11682 (N_11682,N_10498,N_10422);
nand U11683 (N_11683,N_10934,N_10272);
xnor U11684 (N_11684,N_10877,N_10904);
nor U11685 (N_11685,N_10695,N_10747);
nor U11686 (N_11686,N_10138,N_10946);
nor U11687 (N_11687,N_10063,N_10182);
nand U11688 (N_11688,N_10501,N_10412);
nand U11689 (N_11689,N_10127,N_10566);
nor U11690 (N_11690,N_10704,N_10929);
and U11691 (N_11691,N_10445,N_10636);
nand U11692 (N_11692,N_10572,N_10624);
or U11693 (N_11693,N_10711,N_10550);
and U11694 (N_11694,N_10046,N_10345);
nor U11695 (N_11695,N_10189,N_10768);
xnor U11696 (N_11696,N_10294,N_10715);
nand U11697 (N_11697,N_10750,N_10175);
or U11698 (N_11698,N_10995,N_10804);
nor U11699 (N_11699,N_10177,N_10920);
xnor U11700 (N_11700,N_10183,N_10735);
and U11701 (N_11701,N_10878,N_10966);
nor U11702 (N_11702,N_10984,N_10055);
and U11703 (N_11703,N_10190,N_10163);
xnor U11704 (N_11704,N_10767,N_10446);
xnor U11705 (N_11705,N_10700,N_10786);
and U11706 (N_11706,N_10147,N_10646);
xor U11707 (N_11707,N_10838,N_10591);
xor U11708 (N_11708,N_10243,N_10896);
nand U11709 (N_11709,N_10387,N_10585);
nor U11710 (N_11710,N_10655,N_10180);
nor U11711 (N_11711,N_10729,N_10977);
and U11712 (N_11712,N_10831,N_10694);
and U11713 (N_11713,N_10741,N_10052);
nor U11714 (N_11714,N_10332,N_10427);
and U11715 (N_11715,N_10286,N_10375);
nor U11716 (N_11716,N_10033,N_10126);
nor U11717 (N_11717,N_10137,N_10899);
and U11718 (N_11718,N_10702,N_10640);
nor U11719 (N_11719,N_10062,N_10159);
or U11720 (N_11720,N_10500,N_10705);
and U11721 (N_11721,N_10140,N_10211);
nand U11722 (N_11722,N_10188,N_10337);
nand U11723 (N_11723,N_10862,N_10881);
xor U11724 (N_11724,N_10052,N_10847);
xnor U11725 (N_11725,N_10060,N_10612);
or U11726 (N_11726,N_10030,N_10993);
nor U11727 (N_11727,N_10588,N_10542);
nand U11728 (N_11728,N_10161,N_10083);
nand U11729 (N_11729,N_10819,N_10969);
or U11730 (N_11730,N_10855,N_10341);
nand U11731 (N_11731,N_10812,N_10839);
nand U11732 (N_11732,N_10600,N_10608);
nand U11733 (N_11733,N_10364,N_10687);
nand U11734 (N_11734,N_10376,N_10800);
xor U11735 (N_11735,N_10218,N_10163);
nand U11736 (N_11736,N_10596,N_10709);
nand U11737 (N_11737,N_10659,N_10347);
nor U11738 (N_11738,N_10947,N_10206);
nor U11739 (N_11739,N_10878,N_10419);
or U11740 (N_11740,N_10036,N_10860);
nor U11741 (N_11741,N_10901,N_10115);
and U11742 (N_11742,N_10900,N_10366);
or U11743 (N_11743,N_10595,N_10284);
or U11744 (N_11744,N_10387,N_10284);
and U11745 (N_11745,N_10629,N_10740);
nor U11746 (N_11746,N_10425,N_10913);
and U11747 (N_11747,N_10872,N_10411);
nand U11748 (N_11748,N_10303,N_10824);
or U11749 (N_11749,N_10487,N_10095);
and U11750 (N_11750,N_10049,N_10938);
xnor U11751 (N_11751,N_10336,N_10480);
xnor U11752 (N_11752,N_10914,N_10318);
nand U11753 (N_11753,N_10697,N_10248);
or U11754 (N_11754,N_10809,N_10022);
or U11755 (N_11755,N_10388,N_10629);
nand U11756 (N_11756,N_10310,N_10624);
or U11757 (N_11757,N_10136,N_10607);
and U11758 (N_11758,N_10259,N_10341);
and U11759 (N_11759,N_10332,N_10826);
nor U11760 (N_11760,N_10353,N_10325);
xnor U11761 (N_11761,N_10889,N_10032);
nand U11762 (N_11762,N_10298,N_10139);
and U11763 (N_11763,N_10950,N_10893);
or U11764 (N_11764,N_10507,N_10930);
xnor U11765 (N_11765,N_10365,N_10197);
nand U11766 (N_11766,N_10261,N_10232);
nand U11767 (N_11767,N_10629,N_10009);
xor U11768 (N_11768,N_10638,N_10351);
xor U11769 (N_11769,N_10642,N_10244);
nand U11770 (N_11770,N_10870,N_10515);
or U11771 (N_11771,N_10513,N_10528);
and U11772 (N_11772,N_10787,N_10596);
nor U11773 (N_11773,N_10557,N_10858);
nor U11774 (N_11774,N_10347,N_10656);
nor U11775 (N_11775,N_10235,N_10398);
nor U11776 (N_11776,N_10825,N_10642);
nand U11777 (N_11777,N_10025,N_10196);
xnor U11778 (N_11778,N_10521,N_10021);
and U11779 (N_11779,N_10128,N_10275);
nor U11780 (N_11780,N_10203,N_10917);
xor U11781 (N_11781,N_10564,N_10630);
nor U11782 (N_11782,N_10922,N_10801);
or U11783 (N_11783,N_10071,N_10240);
nand U11784 (N_11784,N_10725,N_10368);
nand U11785 (N_11785,N_10128,N_10004);
and U11786 (N_11786,N_10162,N_10047);
or U11787 (N_11787,N_10887,N_10144);
or U11788 (N_11788,N_10181,N_10673);
nand U11789 (N_11789,N_10077,N_10168);
or U11790 (N_11790,N_10419,N_10995);
or U11791 (N_11791,N_10424,N_10178);
or U11792 (N_11792,N_10552,N_10959);
and U11793 (N_11793,N_10075,N_10842);
and U11794 (N_11794,N_10432,N_10841);
and U11795 (N_11795,N_10395,N_10640);
nor U11796 (N_11796,N_10136,N_10574);
nand U11797 (N_11797,N_10469,N_10574);
nand U11798 (N_11798,N_10679,N_10600);
nand U11799 (N_11799,N_10759,N_10432);
or U11800 (N_11800,N_10493,N_10102);
or U11801 (N_11801,N_10201,N_10095);
and U11802 (N_11802,N_10626,N_10361);
and U11803 (N_11803,N_10876,N_10217);
xor U11804 (N_11804,N_10554,N_10827);
xnor U11805 (N_11805,N_10500,N_10796);
nor U11806 (N_11806,N_10266,N_10772);
nor U11807 (N_11807,N_10010,N_10547);
nand U11808 (N_11808,N_10637,N_10644);
and U11809 (N_11809,N_10866,N_10792);
or U11810 (N_11810,N_10112,N_10730);
or U11811 (N_11811,N_10777,N_10211);
and U11812 (N_11812,N_10226,N_10689);
or U11813 (N_11813,N_10362,N_10380);
xor U11814 (N_11814,N_10912,N_10556);
nand U11815 (N_11815,N_10328,N_10217);
xnor U11816 (N_11816,N_10945,N_10020);
or U11817 (N_11817,N_10283,N_10816);
or U11818 (N_11818,N_10393,N_10958);
and U11819 (N_11819,N_10210,N_10870);
nor U11820 (N_11820,N_10053,N_10574);
nor U11821 (N_11821,N_10327,N_10806);
xnor U11822 (N_11822,N_10378,N_10540);
nand U11823 (N_11823,N_10846,N_10754);
nor U11824 (N_11824,N_10163,N_10287);
or U11825 (N_11825,N_10453,N_10230);
nand U11826 (N_11826,N_10446,N_10824);
nor U11827 (N_11827,N_10242,N_10070);
xnor U11828 (N_11828,N_10403,N_10051);
nand U11829 (N_11829,N_10509,N_10080);
or U11830 (N_11830,N_10744,N_10947);
nor U11831 (N_11831,N_10430,N_10440);
nand U11832 (N_11832,N_10448,N_10687);
xor U11833 (N_11833,N_10679,N_10360);
or U11834 (N_11834,N_10490,N_10822);
or U11835 (N_11835,N_10163,N_10115);
xnor U11836 (N_11836,N_10144,N_10110);
nand U11837 (N_11837,N_10551,N_10117);
xor U11838 (N_11838,N_10219,N_10909);
nand U11839 (N_11839,N_10626,N_10602);
nor U11840 (N_11840,N_10044,N_10510);
and U11841 (N_11841,N_10039,N_10599);
or U11842 (N_11842,N_10991,N_10558);
nand U11843 (N_11843,N_10572,N_10735);
nor U11844 (N_11844,N_10972,N_10326);
or U11845 (N_11845,N_10041,N_10958);
nor U11846 (N_11846,N_10037,N_10098);
and U11847 (N_11847,N_10338,N_10972);
and U11848 (N_11848,N_10910,N_10779);
xnor U11849 (N_11849,N_10488,N_10835);
and U11850 (N_11850,N_10625,N_10945);
nand U11851 (N_11851,N_10602,N_10020);
nand U11852 (N_11852,N_10793,N_10830);
xnor U11853 (N_11853,N_10384,N_10249);
nand U11854 (N_11854,N_10255,N_10591);
nor U11855 (N_11855,N_10039,N_10295);
xnor U11856 (N_11856,N_10922,N_10552);
and U11857 (N_11857,N_10162,N_10493);
and U11858 (N_11858,N_10975,N_10196);
and U11859 (N_11859,N_10993,N_10411);
xor U11860 (N_11860,N_10097,N_10129);
nand U11861 (N_11861,N_10078,N_10086);
nor U11862 (N_11862,N_10010,N_10911);
nor U11863 (N_11863,N_10288,N_10521);
and U11864 (N_11864,N_10360,N_10357);
and U11865 (N_11865,N_10434,N_10251);
xor U11866 (N_11866,N_10204,N_10190);
nand U11867 (N_11867,N_10752,N_10933);
nor U11868 (N_11868,N_10645,N_10694);
xnor U11869 (N_11869,N_10317,N_10064);
nand U11870 (N_11870,N_10982,N_10035);
nand U11871 (N_11871,N_10804,N_10858);
nor U11872 (N_11872,N_10198,N_10474);
nor U11873 (N_11873,N_10127,N_10986);
nor U11874 (N_11874,N_10038,N_10594);
or U11875 (N_11875,N_10204,N_10749);
nand U11876 (N_11876,N_10248,N_10717);
or U11877 (N_11877,N_10030,N_10574);
and U11878 (N_11878,N_10368,N_10161);
and U11879 (N_11879,N_10703,N_10127);
nand U11880 (N_11880,N_10023,N_10742);
or U11881 (N_11881,N_10869,N_10295);
xnor U11882 (N_11882,N_10305,N_10742);
nor U11883 (N_11883,N_10856,N_10762);
nor U11884 (N_11884,N_10698,N_10285);
and U11885 (N_11885,N_10760,N_10415);
nand U11886 (N_11886,N_10382,N_10485);
nand U11887 (N_11887,N_10362,N_10335);
nor U11888 (N_11888,N_10660,N_10160);
and U11889 (N_11889,N_10428,N_10880);
nor U11890 (N_11890,N_10317,N_10406);
or U11891 (N_11891,N_10153,N_10224);
nor U11892 (N_11892,N_10567,N_10380);
and U11893 (N_11893,N_10571,N_10418);
xor U11894 (N_11894,N_10670,N_10366);
nor U11895 (N_11895,N_10223,N_10334);
and U11896 (N_11896,N_10776,N_10950);
or U11897 (N_11897,N_10838,N_10568);
or U11898 (N_11898,N_10978,N_10300);
and U11899 (N_11899,N_10357,N_10269);
xnor U11900 (N_11900,N_10630,N_10986);
xor U11901 (N_11901,N_10866,N_10828);
xor U11902 (N_11902,N_10708,N_10983);
nand U11903 (N_11903,N_10322,N_10556);
or U11904 (N_11904,N_10697,N_10127);
xor U11905 (N_11905,N_10689,N_10527);
and U11906 (N_11906,N_10120,N_10675);
and U11907 (N_11907,N_10723,N_10964);
nand U11908 (N_11908,N_10551,N_10090);
nor U11909 (N_11909,N_10192,N_10930);
or U11910 (N_11910,N_10075,N_10102);
nand U11911 (N_11911,N_10675,N_10262);
xnor U11912 (N_11912,N_10751,N_10862);
and U11913 (N_11913,N_10904,N_10883);
and U11914 (N_11914,N_10632,N_10715);
nor U11915 (N_11915,N_10529,N_10372);
or U11916 (N_11916,N_10553,N_10424);
nor U11917 (N_11917,N_10578,N_10601);
or U11918 (N_11918,N_10669,N_10470);
or U11919 (N_11919,N_10431,N_10954);
and U11920 (N_11920,N_10971,N_10106);
nor U11921 (N_11921,N_10896,N_10819);
and U11922 (N_11922,N_10450,N_10470);
nor U11923 (N_11923,N_10924,N_10148);
nor U11924 (N_11924,N_10939,N_10842);
xnor U11925 (N_11925,N_10575,N_10809);
nor U11926 (N_11926,N_10560,N_10440);
nor U11927 (N_11927,N_10783,N_10482);
xnor U11928 (N_11928,N_10196,N_10985);
nand U11929 (N_11929,N_10547,N_10415);
nor U11930 (N_11930,N_10491,N_10806);
nor U11931 (N_11931,N_10171,N_10652);
xor U11932 (N_11932,N_10698,N_10451);
xnor U11933 (N_11933,N_10283,N_10851);
nand U11934 (N_11934,N_10507,N_10030);
nor U11935 (N_11935,N_10827,N_10422);
or U11936 (N_11936,N_10038,N_10246);
xor U11937 (N_11937,N_10145,N_10314);
and U11938 (N_11938,N_10360,N_10154);
and U11939 (N_11939,N_10360,N_10181);
or U11940 (N_11940,N_10265,N_10478);
nand U11941 (N_11941,N_10738,N_10964);
nand U11942 (N_11942,N_10866,N_10015);
or U11943 (N_11943,N_10543,N_10740);
xor U11944 (N_11944,N_10617,N_10882);
or U11945 (N_11945,N_10816,N_10463);
and U11946 (N_11946,N_10068,N_10095);
or U11947 (N_11947,N_10457,N_10735);
and U11948 (N_11948,N_10722,N_10122);
nor U11949 (N_11949,N_10399,N_10867);
nor U11950 (N_11950,N_10531,N_10956);
and U11951 (N_11951,N_10758,N_10736);
xor U11952 (N_11952,N_10509,N_10798);
nand U11953 (N_11953,N_10768,N_10389);
nand U11954 (N_11954,N_10368,N_10982);
or U11955 (N_11955,N_10344,N_10830);
and U11956 (N_11956,N_10722,N_10890);
nand U11957 (N_11957,N_10802,N_10501);
nor U11958 (N_11958,N_10536,N_10669);
nand U11959 (N_11959,N_10018,N_10746);
xnor U11960 (N_11960,N_10108,N_10244);
and U11961 (N_11961,N_10333,N_10319);
and U11962 (N_11962,N_10538,N_10248);
nand U11963 (N_11963,N_10954,N_10377);
xor U11964 (N_11964,N_10249,N_10255);
nand U11965 (N_11965,N_10806,N_10520);
and U11966 (N_11966,N_10123,N_10790);
or U11967 (N_11967,N_10976,N_10034);
nor U11968 (N_11968,N_10336,N_10083);
nor U11969 (N_11969,N_10504,N_10969);
or U11970 (N_11970,N_10882,N_10130);
or U11971 (N_11971,N_10428,N_10524);
or U11972 (N_11972,N_10392,N_10454);
nand U11973 (N_11973,N_10933,N_10579);
nand U11974 (N_11974,N_10641,N_10353);
or U11975 (N_11975,N_10530,N_10913);
nor U11976 (N_11976,N_10052,N_10176);
nand U11977 (N_11977,N_10869,N_10462);
xnor U11978 (N_11978,N_10588,N_10609);
nand U11979 (N_11979,N_10904,N_10111);
nand U11980 (N_11980,N_10797,N_10446);
nor U11981 (N_11981,N_10463,N_10470);
xnor U11982 (N_11982,N_10763,N_10389);
nor U11983 (N_11983,N_10846,N_10399);
and U11984 (N_11984,N_10289,N_10557);
nand U11985 (N_11985,N_10712,N_10640);
nor U11986 (N_11986,N_10489,N_10834);
or U11987 (N_11987,N_10363,N_10348);
nor U11988 (N_11988,N_10413,N_10029);
or U11989 (N_11989,N_10392,N_10232);
and U11990 (N_11990,N_10390,N_10128);
nor U11991 (N_11991,N_10143,N_10256);
nand U11992 (N_11992,N_10354,N_10956);
nor U11993 (N_11993,N_10790,N_10444);
xnor U11994 (N_11994,N_10426,N_10905);
and U11995 (N_11995,N_10278,N_10108);
and U11996 (N_11996,N_10615,N_10454);
and U11997 (N_11997,N_10386,N_10843);
nor U11998 (N_11998,N_10924,N_10265);
nor U11999 (N_11999,N_10611,N_10616);
and U12000 (N_12000,N_11307,N_11894);
and U12001 (N_12001,N_11407,N_11242);
nand U12002 (N_12002,N_11297,N_11085);
or U12003 (N_12003,N_11926,N_11126);
or U12004 (N_12004,N_11730,N_11445);
nor U12005 (N_12005,N_11501,N_11024);
nand U12006 (N_12006,N_11076,N_11192);
or U12007 (N_12007,N_11149,N_11646);
or U12008 (N_12008,N_11699,N_11986);
and U12009 (N_12009,N_11399,N_11612);
or U12010 (N_12010,N_11892,N_11872);
or U12011 (N_12011,N_11186,N_11613);
nor U12012 (N_12012,N_11084,N_11409);
xor U12013 (N_12013,N_11228,N_11934);
nor U12014 (N_12014,N_11696,N_11584);
nor U12015 (N_12015,N_11095,N_11969);
xnor U12016 (N_12016,N_11680,N_11101);
or U12017 (N_12017,N_11597,N_11248);
and U12018 (N_12018,N_11098,N_11732);
nor U12019 (N_12019,N_11052,N_11321);
nor U12020 (N_12020,N_11203,N_11382);
and U12021 (N_12021,N_11640,N_11289);
nand U12022 (N_12022,N_11863,N_11384);
or U12023 (N_12023,N_11852,N_11470);
xnor U12024 (N_12024,N_11195,N_11756);
nand U12025 (N_12025,N_11386,N_11655);
nand U12026 (N_12026,N_11809,N_11060);
and U12027 (N_12027,N_11104,N_11804);
xnor U12028 (N_12028,N_11325,N_11270);
nor U12029 (N_12029,N_11946,N_11790);
nor U12030 (N_12030,N_11312,N_11155);
nor U12031 (N_12031,N_11212,N_11534);
and U12032 (N_12032,N_11679,N_11835);
nor U12033 (N_12033,N_11274,N_11798);
or U12034 (N_12034,N_11719,N_11910);
or U12035 (N_12035,N_11468,N_11886);
or U12036 (N_12036,N_11308,N_11372);
xor U12037 (N_12037,N_11471,N_11397);
or U12038 (N_12038,N_11654,N_11851);
nor U12039 (N_12039,N_11432,N_11671);
nor U12040 (N_12040,N_11182,N_11704);
xor U12041 (N_12041,N_11258,N_11191);
nand U12042 (N_12042,N_11158,N_11728);
nor U12043 (N_12043,N_11552,N_11209);
and U12044 (N_12044,N_11417,N_11132);
or U12045 (N_12045,N_11588,N_11073);
nand U12046 (N_12046,N_11322,N_11331);
nand U12047 (N_12047,N_11229,N_11766);
nor U12048 (N_12048,N_11023,N_11290);
and U12049 (N_12049,N_11824,N_11473);
nand U12050 (N_12050,N_11941,N_11398);
xor U12051 (N_12051,N_11723,N_11862);
and U12052 (N_12052,N_11772,N_11915);
or U12053 (N_12053,N_11856,N_11278);
or U12054 (N_12054,N_11150,N_11806);
nand U12055 (N_12055,N_11742,N_11648);
nor U12056 (N_12056,N_11922,N_11217);
and U12057 (N_12057,N_11868,N_11357);
nand U12058 (N_12058,N_11879,N_11402);
and U12059 (N_12059,N_11675,N_11998);
xnor U12060 (N_12060,N_11694,N_11000);
xor U12061 (N_12061,N_11722,N_11050);
or U12062 (N_12062,N_11171,N_11649);
xnor U12063 (N_12063,N_11557,N_11829);
or U12064 (N_12064,N_11315,N_11185);
and U12065 (N_12065,N_11611,N_11581);
and U12066 (N_12066,N_11080,N_11446);
nor U12067 (N_12067,N_11013,N_11256);
xnor U12068 (N_12068,N_11583,N_11164);
or U12069 (N_12069,N_11314,N_11461);
nor U12070 (N_12070,N_11647,N_11387);
nand U12071 (N_12071,N_11202,N_11049);
nand U12072 (N_12072,N_11707,N_11978);
nand U12073 (N_12073,N_11606,N_11693);
nand U12074 (N_12074,N_11533,N_11148);
or U12075 (N_12075,N_11792,N_11838);
nor U12076 (N_12076,N_11690,N_11263);
nor U12077 (N_12077,N_11090,N_11210);
nor U12078 (N_12078,N_11528,N_11850);
and U12079 (N_12079,N_11075,N_11960);
and U12080 (N_12080,N_11643,N_11762);
nand U12081 (N_12081,N_11518,N_11444);
and U12082 (N_12082,N_11082,N_11853);
nor U12083 (N_12083,N_11903,N_11069);
and U12084 (N_12084,N_11840,N_11484);
or U12085 (N_12085,N_11036,N_11466);
and U12086 (N_12086,N_11144,N_11428);
or U12087 (N_12087,N_11656,N_11799);
nand U12088 (N_12088,N_11793,N_11423);
nor U12089 (N_12089,N_11535,N_11524);
nor U12090 (N_12090,N_11818,N_11081);
xor U12091 (N_12091,N_11996,N_11854);
xnor U12092 (N_12092,N_11511,N_11939);
xor U12093 (N_12093,N_11598,N_11456);
and U12094 (N_12094,N_11814,N_11162);
or U12095 (N_12095,N_11421,N_11661);
xor U12096 (N_12096,N_11504,N_11875);
nor U12097 (N_12097,N_11190,N_11776);
or U12098 (N_12098,N_11147,N_11514);
xnor U12099 (N_12099,N_11861,N_11108);
nor U12100 (N_12100,N_11898,N_11976);
or U12101 (N_12101,N_11962,N_11356);
nor U12102 (N_12102,N_11682,N_11971);
nand U12103 (N_12103,N_11830,N_11010);
nand U12104 (N_12104,N_11021,N_11726);
and U12105 (N_12105,N_11037,N_11902);
xnor U12106 (N_12106,N_11219,N_11757);
nor U12107 (N_12107,N_11301,N_11179);
nand U12108 (N_12108,N_11542,N_11802);
nor U12109 (N_12109,N_11826,N_11346);
nand U12110 (N_12110,N_11268,N_11053);
and U12111 (N_12111,N_11291,N_11701);
or U12112 (N_12112,N_11751,N_11810);
nor U12113 (N_12113,N_11271,N_11429);
nor U12114 (N_12114,N_11683,N_11235);
or U12115 (N_12115,N_11391,N_11579);
nor U12116 (N_12116,N_11475,N_11687);
xnor U12117 (N_12117,N_11481,N_11296);
or U12118 (N_12118,N_11950,N_11995);
or U12119 (N_12119,N_11964,N_11413);
nand U12120 (N_12120,N_11841,N_11111);
or U12121 (N_12121,N_11717,N_11778);
xor U12122 (N_12122,N_11221,N_11326);
nand U12123 (N_12123,N_11157,N_11561);
xor U12124 (N_12124,N_11645,N_11318);
nand U12125 (N_12125,N_11205,N_11175);
nand U12126 (N_12126,N_11404,N_11593);
and U12127 (N_12127,N_11442,N_11629);
nor U12128 (N_12128,N_11408,N_11727);
and U12129 (N_12129,N_11990,N_11488);
xnor U12130 (N_12130,N_11777,N_11741);
nand U12131 (N_12131,N_11919,N_11497);
or U12132 (N_12132,N_11293,N_11216);
and U12133 (N_12133,N_11364,N_11241);
nand U12134 (N_12134,N_11538,N_11746);
nand U12135 (N_12135,N_11250,N_11617);
nand U12136 (N_12136,N_11887,N_11713);
nand U12137 (N_12137,N_11493,N_11822);
xor U12138 (N_12138,N_11796,N_11869);
and U12139 (N_12139,N_11334,N_11779);
or U12140 (N_12140,N_11540,N_11921);
xnor U12141 (N_12141,N_11254,N_11816);
or U12142 (N_12142,N_11309,N_11449);
xnor U12143 (N_12143,N_11878,N_11945);
nor U12144 (N_12144,N_11403,N_11009);
nand U12145 (N_12145,N_11142,N_11523);
and U12146 (N_12146,N_11393,N_11187);
or U12147 (N_12147,N_11787,N_11341);
nand U12148 (N_12148,N_11441,N_11710);
nand U12149 (N_12149,N_11764,N_11498);
xnor U12150 (N_12150,N_11113,N_11103);
nor U12151 (N_12151,N_11548,N_11238);
and U12152 (N_12152,N_11338,N_11944);
xnor U12153 (N_12153,N_11927,N_11285);
nand U12154 (N_12154,N_11259,N_11530);
or U12155 (N_12155,N_11243,N_11174);
xnor U12156 (N_12156,N_11137,N_11972);
nor U12157 (N_12157,N_11917,N_11345);
and U12158 (N_12158,N_11327,N_11131);
and U12159 (N_12159,N_11156,N_11499);
nand U12160 (N_12160,N_11463,N_11020);
nor U12161 (N_12161,N_11479,N_11625);
or U12162 (N_12162,N_11897,N_11522);
or U12163 (N_12163,N_11980,N_11018);
or U12164 (N_12164,N_11365,N_11328);
xnor U12165 (N_12165,N_11992,N_11952);
nand U12166 (N_12166,N_11070,N_11546);
nand U12167 (N_12167,N_11901,N_11116);
nand U12168 (N_12168,N_11249,N_11665);
nand U12169 (N_12169,N_11916,N_11537);
or U12170 (N_12170,N_11375,N_11725);
nor U12171 (N_12171,N_11477,N_11001);
xnor U12172 (N_12172,N_11230,N_11739);
nand U12173 (N_12173,N_11889,N_11390);
xor U12174 (N_12174,N_11450,N_11666);
nor U12175 (N_12175,N_11770,N_11224);
nor U12176 (N_12176,N_11138,N_11700);
xnor U12177 (N_12177,N_11299,N_11622);
and U12178 (N_12178,N_11983,N_11340);
or U12179 (N_12179,N_11743,N_11607);
and U12180 (N_12180,N_11582,N_11519);
or U12181 (N_12181,N_11933,N_11849);
and U12182 (N_12182,N_11923,N_11025);
and U12183 (N_12183,N_11651,N_11712);
nand U12184 (N_12184,N_11237,N_11760);
or U12185 (N_12185,N_11016,N_11368);
nand U12186 (N_12186,N_11859,N_11339);
xnor U12187 (N_12187,N_11999,N_11545);
and U12188 (N_12188,N_11750,N_11805);
nand U12189 (N_12189,N_11086,N_11797);
and U12190 (N_12190,N_11225,N_11211);
and U12191 (N_12191,N_11685,N_11130);
xor U12192 (N_12192,N_11895,N_11968);
nor U12193 (N_12193,N_11083,N_11536);
nand U12194 (N_12194,N_11636,N_11100);
nand U12195 (N_12195,N_11124,N_11478);
nor U12196 (N_12196,N_11465,N_11193);
or U12197 (N_12197,N_11183,N_11153);
or U12198 (N_12198,N_11317,N_11828);
and U12199 (N_12199,N_11019,N_11286);
nor U12200 (N_12200,N_11206,N_11234);
and U12201 (N_12201,N_11419,N_11748);
nand U12202 (N_12202,N_11168,N_11531);
xor U12203 (N_12203,N_11239,N_11367);
and U12204 (N_12204,N_11691,N_11652);
and U12205 (N_12205,N_11226,N_11269);
nor U12206 (N_12206,N_11508,N_11078);
and U12207 (N_12207,N_11089,N_11152);
nor U12208 (N_12208,N_11698,N_11160);
nand U12209 (N_12209,N_11954,N_11337);
xnor U12210 (N_12210,N_11697,N_11695);
nand U12211 (N_12211,N_11109,N_11426);
nor U12212 (N_12212,N_11821,N_11097);
nand U12213 (N_12213,N_11039,N_11119);
or U12214 (N_12214,N_11997,N_11443);
or U12215 (N_12215,N_11292,N_11008);
nand U12216 (N_12216,N_11352,N_11619);
xnor U12217 (N_12217,N_11015,N_11789);
nor U12218 (N_12218,N_11240,N_11030);
or U12219 (N_12219,N_11313,N_11788);
xnor U12220 (N_12220,N_11931,N_11911);
nand U12221 (N_12221,N_11462,N_11633);
nand U12222 (N_12222,N_11261,N_11763);
nand U12223 (N_12223,N_11918,N_11145);
nand U12224 (N_12224,N_11092,N_11837);
xor U12225 (N_12225,N_11846,N_11663);
nor U12226 (N_12226,N_11855,N_11117);
or U12227 (N_12227,N_11486,N_11414);
nand U12228 (N_12228,N_11987,N_11105);
nor U12229 (N_12229,N_11213,N_11056);
xnor U12230 (N_12230,N_11385,N_11638);
nand U12231 (N_12231,N_11891,N_11112);
xnor U12232 (N_12232,N_11595,N_11961);
xnor U12233 (N_12233,N_11957,N_11882);
and U12234 (N_12234,N_11355,N_11431);
nand U12235 (N_12235,N_11028,N_11173);
nand U12236 (N_12236,N_11564,N_11585);
or U12237 (N_12237,N_11559,N_11106);
nor U12238 (N_12238,N_11689,N_11310);
xnor U12239 (N_12239,N_11295,N_11527);
and U12240 (N_12240,N_11876,N_11420);
or U12241 (N_12241,N_11510,N_11178);
nor U12242 (N_12242,N_11336,N_11383);
nand U12243 (N_12243,N_11159,N_11848);
xor U12244 (N_12244,N_11507,N_11376);
nor U12245 (N_12245,N_11857,N_11121);
nor U12246 (N_12246,N_11379,N_11982);
or U12247 (N_12247,N_11738,N_11642);
or U12248 (N_12248,N_11491,N_11624);
nand U12249 (N_12249,N_11904,N_11556);
or U12250 (N_12250,N_11860,N_11029);
nand U12251 (N_12251,N_11472,N_11304);
nor U12252 (N_12252,N_11204,N_11956);
or U12253 (N_12253,N_11114,N_11517);
and U12254 (N_12254,N_11395,N_11775);
xnor U12255 (N_12255,N_11316,N_11747);
or U12256 (N_12256,N_11394,N_11801);
nor U12257 (N_12257,N_11416,N_11929);
nand U12258 (N_12258,N_11858,N_11664);
xor U12259 (N_12259,N_11731,N_11252);
nand U12260 (N_12260,N_11262,N_11771);
xnor U12261 (N_12261,N_11867,N_11953);
xor U12262 (N_12262,N_11247,N_11184);
and U12263 (N_12263,N_11813,N_11427);
or U12264 (N_12264,N_11963,N_11492);
nor U12265 (N_12265,N_11418,N_11043);
nor U12266 (N_12266,N_11135,N_11733);
and U12267 (N_12267,N_11197,N_11236);
nand U12268 (N_12268,N_11074,N_11288);
and U12269 (N_12269,N_11580,N_11539);
nand U12270 (N_12270,N_11521,N_11358);
nor U12271 (N_12271,N_11866,N_11222);
xnor U12272 (N_12272,N_11893,N_11605);
nor U12273 (N_12273,N_11512,N_11485);
nand U12274 (N_12274,N_11167,N_11094);
xor U12275 (N_12275,N_11373,N_11051);
nand U12276 (N_12276,N_11885,N_11905);
nor U12277 (N_12277,N_11609,N_11761);
nor U12278 (N_12278,N_11396,N_11970);
xnor U12279 (N_12279,N_11574,N_11985);
nor U12280 (N_12280,N_11233,N_11592);
xnor U12281 (N_12281,N_11599,N_11366);
or U12282 (N_12282,N_11565,N_11169);
nand U12283 (N_12283,N_11412,N_11803);
nand U12284 (N_12284,N_11890,N_11012);
nand U12285 (N_12285,N_11631,N_11063);
xor U12286 (N_12286,N_11047,N_11118);
nor U12287 (N_12287,N_11794,N_11305);
and U12288 (N_12288,N_11604,N_11099);
nor U12289 (N_12289,N_11311,N_11811);
and U12290 (N_12290,N_11424,N_11354);
or U12291 (N_12291,N_11332,N_11434);
and U12292 (N_12292,N_11044,N_11096);
or U12293 (N_12293,N_11720,N_11958);
and U12294 (N_12294,N_11637,N_11781);
and U12295 (N_12295,N_11143,N_11758);
nand U12296 (N_12296,N_11287,N_11577);
nor U12297 (N_12297,N_11227,N_11244);
nor U12298 (N_12298,N_11833,N_11672);
or U12299 (N_12299,N_11618,N_11667);
or U12300 (N_12300,N_11549,N_11177);
nand U12301 (N_12301,N_11591,N_11437);
or U12302 (N_12302,N_11260,N_11490);
nand U12303 (N_12303,N_11621,N_11791);
nor U12304 (N_12304,N_11807,N_11973);
or U12305 (N_12305,N_11602,N_11906);
nor U12306 (N_12306,N_11454,N_11808);
and U12307 (N_12307,N_11587,N_11753);
and U12308 (N_12308,N_11482,N_11520);
xnor U12309 (N_12309,N_11275,N_11907);
and U12310 (N_12310,N_11430,N_11207);
nand U12311 (N_12311,N_11626,N_11955);
nor U12312 (N_12312,N_11294,N_11136);
or U12313 (N_12313,N_11842,N_11737);
nand U12314 (N_12314,N_11120,N_11048);
and U12315 (N_12315,N_11817,N_11059);
nand U12316 (N_12316,N_11634,N_11125);
nor U12317 (N_12317,N_11281,N_11688);
xor U12318 (N_12318,N_11087,N_11573);
nor U12319 (N_12319,N_11749,N_11033);
and U12320 (N_12320,N_11388,N_11632);
nand U12321 (N_12321,N_11951,N_11378);
and U12322 (N_12322,N_11107,N_11360);
or U12323 (N_12323,N_11936,N_11977);
xnor U12324 (N_12324,N_11277,N_11067);
nand U12325 (N_12325,N_11920,N_11343);
nand U12326 (N_12326,N_11091,N_11380);
or U12327 (N_12327,N_11401,N_11589);
nor U12328 (N_12328,N_11505,N_11040);
or U12329 (N_12329,N_11134,N_11714);
nor U12330 (N_12330,N_11218,N_11435);
xor U12331 (N_12331,N_11348,N_11610);
and U12332 (N_12332,N_11141,N_11502);
nor U12333 (N_12333,N_11154,N_11513);
and U12334 (N_12334,N_11947,N_11031);
nand U12335 (N_12335,N_11061,N_11034);
nor U12336 (N_12336,N_11272,N_11133);
or U12337 (N_12337,N_11093,N_11864);
nand U12338 (N_12338,N_11452,N_11686);
xnor U12339 (N_12339,N_11754,N_11938);
nor U12340 (N_12340,N_11526,N_11650);
xor U12341 (N_12341,N_11566,N_11670);
nand U12342 (N_12342,N_11344,N_11590);
nor U12343 (N_12343,N_11774,N_11724);
and U12344 (N_12344,N_11433,N_11181);
or U12345 (N_12345,N_11974,N_11991);
and U12346 (N_12346,N_11369,N_11253);
or U12347 (N_12347,N_11653,N_11062);
nor U12348 (N_12348,N_11635,N_11614);
xnor U12349 (N_12349,N_11515,N_11568);
nor U12350 (N_12350,N_11888,N_11320);
and U12351 (N_12351,N_11516,N_11035);
nor U12352 (N_12352,N_11506,N_11881);
nor U12353 (N_12353,N_11659,N_11702);
xnor U12354 (N_12354,N_11601,N_11014);
xnor U12355 (N_12355,N_11457,N_11004);
xor U12356 (N_12356,N_11896,N_11071);
nand U12357 (N_12357,N_11041,N_11800);
nand U12358 (N_12358,N_11752,N_11773);
nand U12359 (N_12359,N_11088,N_11005);
nor U12360 (N_12360,N_11839,N_11425);
or U12361 (N_12361,N_11578,N_11335);
nand U12362 (N_12362,N_11780,N_11819);
nor U12363 (N_12363,N_11989,N_11329);
nand U12364 (N_12364,N_11825,N_11323);
nand U12365 (N_12365,N_11453,N_11669);
nand U12366 (N_12366,N_11381,N_11836);
nor U12367 (N_12367,N_11349,N_11140);
xor U12368 (N_12368,N_11558,N_11003);
and U12369 (N_12369,N_11942,N_11017);
and U12370 (N_12370,N_11608,N_11596);
nand U12371 (N_12371,N_11925,N_11415);
nor U12372 (N_12372,N_11392,N_11827);
or U12373 (N_12373,N_11455,N_11844);
and U12374 (N_12374,N_11820,N_11208);
and U12375 (N_12375,N_11623,N_11966);
xor U12376 (N_12376,N_11735,N_11246);
xnor U12377 (N_12377,N_11055,N_11994);
and U12378 (N_12378,N_11870,N_11706);
nand U12379 (N_12379,N_11146,N_11641);
or U12380 (N_12380,N_11555,N_11439);
and U12381 (N_12381,N_11547,N_11871);
or U12382 (N_12382,N_11660,N_11129);
xnor U12383 (N_12383,N_11509,N_11079);
or U12384 (N_12384,N_11681,N_11543);
xor U12385 (N_12385,N_11845,N_11223);
and U12386 (N_12386,N_11115,N_11438);
xor U12387 (N_12387,N_11967,N_11937);
and U12388 (N_12388,N_11843,N_11949);
nor U12389 (N_12389,N_11302,N_11782);
or U12390 (N_12390,N_11361,N_11544);
nand U12391 (N_12391,N_11324,N_11161);
nor U12392 (N_12392,N_11692,N_11908);
and U12393 (N_12393,N_11189,N_11494);
nor U12394 (N_12394,N_11736,N_11102);
and U12395 (N_12395,N_11716,N_11678);
nand U12396 (N_12396,N_11370,N_11734);
nor U12397 (N_12397,N_11405,N_11077);
nor U12398 (N_12398,N_11460,N_11823);
or U12399 (N_12399,N_11529,N_11628);
nor U12400 (N_12400,N_11884,N_11422);
nand U12401 (N_12401,N_11072,N_11571);
nor U12402 (N_12402,N_11575,N_11279);
xor U12403 (N_12403,N_11483,N_11377);
nand U12404 (N_12404,N_11594,N_11264);
and U12405 (N_12405,N_11058,N_11932);
xor U12406 (N_12406,N_11769,N_11165);
xor U12407 (N_12407,N_11198,N_11899);
xor U12408 (N_12408,N_11795,N_11715);
xor U12409 (N_12409,N_11495,N_11027);
or U12410 (N_12410,N_11616,N_11406);
nor U12411 (N_12411,N_11674,N_11988);
nand U12412 (N_12412,N_11480,N_11708);
xnor U12413 (N_12413,N_11551,N_11487);
nand U12414 (N_12414,N_11064,N_11567);
nor U12415 (N_12415,N_11541,N_11068);
and U12416 (N_12416,N_11451,N_11676);
and U12417 (N_12417,N_11525,N_11353);
and U12418 (N_12418,N_11705,N_11943);
or U12419 (N_12419,N_11847,N_11981);
and U12420 (N_12420,N_11993,N_11576);
or U12421 (N_12421,N_11759,N_11007);
nand U12422 (N_12422,N_11729,N_11300);
and U12423 (N_12423,N_11045,N_11940);
and U12424 (N_12424,N_11603,N_11172);
nor U12425 (N_12425,N_11057,N_11740);
nor U12426 (N_12426,N_11448,N_11002);
nor U12427 (N_12427,N_11054,N_11948);
nor U12428 (N_12428,N_11347,N_11673);
nand U12429 (N_12429,N_11965,N_11280);
or U12430 (N_12430,N_11874,N_11026);
xor U12431 (N_12431,N_11194,N_11880);
xor U12432 (N_12432,N_11066,N_11464);
xnor U12433 (N_12433,N_11127,N_11668);
or U12434 (N_12434,N_11709,N_11215);
or U12435 (N_12435,N_11196,N_11188);
nor U12436 (N_12436,N_11657,N_11658);
nor U12437 (N_12437,N_11459,N_11639);
nor U12438 (N_12438,N_11975,N_11914);
xnor U12439 (N_12439,N_11436,N_11255);
nor U12440 (N_12440,N_11006,N_11042);
nor U12441 (N_12441,N_11935,N_11266);
nor U12442 (N_12442,N_11677,N_11644);
nor U12443 (N_12443,N_11703,N_11038);
nand U12444 (N_12444,N_11267,N_11562);
and U12445 (N_12445,N_11755,N_11815);
xor U12446 (N_12446,N_11333,N_11122);
nand U12447 (N_12447,N_11744,N_11303);
nor U12448 (N_12448,N_11684,N_11011);
xor U12449 (N_12449,N_11718,N_11615);
or U12450 (N_12450,N_11877,N_11912);
nor U12451 (N_12451,N_11572,N_11282);
or U12452 (N_12452,N_11257,N_11458);
xnor U12453 (N_12453,N_11022,N_11831);
and U12454 (N_12454,N_11447,N_11834);
nor U12455 (N_12455,N_11231,N_11476);
nand U12456 (N_12456,N_11768,N_11032);
nor U12457 (N_12457,N_11913,N_11283);
nor U12458 (N_12458,N_11489,N_11553);
or U12459 (N_12459,N_11245,N_11359);
or U12460 (N_12460,N_11812,N_11128);
and U12461 (N_12461,N_11214,N_11959);
nand U12462 (N_12462,N_11350,N_11784);
and U12463 (N_12463,N_11046,N_11469);
xor U12464 (N_12464,N_11832,N_11110);
xnor U12465 (N_12465,N_11273,N_11374);
and U12466 (N_12466,N_11550,N_11474);
and U12467 (N_12467,N_11342,N_11600);
or U12468 (N_12468,N_11200,N_11232);
and U12469 (N_12469,N_11979,N_11865);
xnor U12470 (N_12470,N_11873,N_11276);
and U12471 (N_12471,N_11496,N_11930);
or U12472 (N_12472,N_11123,N_11163);
nand U12473 (N_12473,N_11201,N_11411);
nor U12474 (N_12474,N_11554,N_11176);
or U12475 (N_12475,N_11569,N_11220);
or U12476 (N_12476,N_11319,N_11984);
or U12477 (N_12477,N_11620,N_11251);
and U12478 (N_12478,N_11166,N_11532);
xnor U12479 (N_12479,N_11363,N_11400);
nor U12480 (N_12480,N_11389,N_11767);
nand U12481 (N_12481,N_11170,N_11563);
xor U12482 (N_12482,N_11151,N_11065);
nand U12483 (N_12483,N_11786,N_11180);
xnor U12484 (N_12484,N_11265,N_11586);
and U12485 (N_12485,N_11928,N_11503);
or U12486 (N_12486,N_11721,N_11883);
and U12487 (N_12487,N_11371,N_11924);
or U12488 (N_12488,N_11298,N_11467);
nand U12489 (N_12489,N_11362,N_11909);
nand U12490 (N_12490,N_11351,N_11139);
or U12491 (N_12491,N_11560,N_11199);
nand U12492 (N_12492,N_11783,N_11711);
or U12493 (N_12493,N_11662,N_11570);
nand U12494 (N_12494,N_11500,N_11306);
nor U12495 (N_12495,N_11330,N_11440);
nand U12496 (N_12496,N_11785,N_11630);
and U12497 (N_12497,N_11410,N_11627);
nand U12498 (N_12498,N_11765,N_11284);
xor U12499 (N_12499,N_11900,N_11745);
nand U12500 (N_12500,N_11312,N_11886);
or U12501 (N_12501,N_11801,N_11826);
nor U12502 (N_12502,N_11343,N_11797);
xor U12503 (N_12503,N_11690,N_11667);
and U12504 (N_12504,N_11624,N_11421);
nand U12505 (N_12505,N_11736,N_11193);
nor U12506 (N_12506,N_11677,N_11214);
nand U12507 (N_12507,N_11356,N_11391);
nand U12508 (N_12508,N_11647,N_11171);
and U12509 (N_12509,N_11164,N_11674);
or U12510 (N_12510,N_11519,N_11141);
nand U12511 (N_12511,N_11672,N_11898);
or U12512 (N_12512,N_11780,N_11218);
nand U12513 (N_12513,N_11419,N_11348);
nor U12514 (N_12514,N_11631,N_11094);
xor U12515 (N_12515,N_11813,N_11319);
nor U12516 (N_12516,N_11610,N_11644);
xnor U12517 (N_12517,N_11981,N_11571);
nand U12518 (N_12518,N_11555,N_11975);
and U12519 (N_12519,N_11747,N_11124);
and U12520 (N_12520,N_11842,N_11424);
nand U12521 (N_12521,N_11502,N_11723);
nand U12522 (N_12522,N_11299,N_11200);
or U12523 (N_12523,N_11884,N_11223);
and U12524 (N_12524,N_11656,N_11762);
xnor U12525 (N_12525,N_11073,N_11998);
and U12526 (N_12526,N_11166,N_11056);
nor U12527 (N_12527,N_11497,N_11757);
or U12528 (N_12528,N_11438,N_11777);
and U12529 (N_12529,N_11786,N_11001);
and U12530 (N_12530,N_11856,N_11446);
or U12531 (N_12531,N_11354,N_11089);
and U12532 (N_12532,N_11853,N_11735);
nor U12533 (N_12533,N_11390,N_11100);
xor U12534 (N_12534,N_11970,N_11871);
nand U12535 (N_12535,N_11211,N_11064);
xnor U12536 (N_12536,N_11994,N_11022);
nand U12537 (N_12537,N_11028,N_11744);
or U12538 (N_12538,N_11236,N_11134);
and U12539 (N_12539,N_11583,N_11272);
and U12540 (N_12540,N_11829,N_11335);
or U12541 (N_12541,N_11040,N_11599);
and U12542 (N_12542,N_11564,N_11150);
xor U12543 (N_12543,N_11158,N_11206);
or U12544 (N_12544,N_11044,N_11154);
nand U12545 (N_12545,N_11775,N_11587);
nor U12546 (N_12546,N_11055,N_11786);
or U12547 (N_12547,N_11327,N_11441);
or U12548 (N_12548,N_11244,N_11516);
xor U12549 (N_12549,N_11825,N_11228);
nor U12550 (N_12550,N_11625,N_11462);
nand U12551 (N_12551,N_11425,N_11845);
and U12552 (N_12552,N_11299,N_11338);
xor U12553 (N_12553,N_11325,N_11280);
or U12554 (N_12554,N_11455,N_11341);
or U12555 (N_12555,N_11424,N_11260);
and U12556 (N_12556,N_11845,N_11426);
nand U12557 (N_12557,N_11507,N_11387);
or U12558 (N_12558,N_11147,N_11459);
or U12559 (N_12559,N_11036,N_11112);
nor U12560 (N_12560,N_11316,N_11479);
nand U12561 (N_12561,N_11029,N_11260);
or U12562 (N_12562,N_11571,N_11285);
and U12563 (N_12563,N_11020,N_11936);
nand U12564 (N_12564,N_11951,N_11855);
nand U12565 (N_12565,N_11388,N_11222);
xor U12566 (N_12566,N_11945,N_11770);
nand U12567 (N_12567,N_11397,N_11001);
and U12568 (N_12568,N_11394,N_11553);
nand U12569 (N_12569,N_11125,N_11319);
and U12570 (N_12570,N_11016,N_11906);
or U12571 (N_12571,N_11591,N_11410);
or U12572 (N_12572,N_11135,N_11908);
and U12573 (N_12573,N_11126,N_11495);
nor U12574 (N_12574,N_11235,N_11522);
nand U12575 (N_12575,N_11141,N_11208);
nand U12576 (N_12576,N_11255,N_11145);
and U12577 (N_12577,N_11592,N_11918);
nand U12578 (N_12578,N_11421,N_11385);
nor U12579 (N_12579,N_11034,N_11212);
nand U12580 (N_12580,N_11664,N_11148);
nand U12581 (N_12581,N_11533,N_11578);
nor U12582 (N_12582,N_11098,N_11520);
nor U12583 (N_12583,N_11940,N_11307);
nand U12584 (N_12584,N_11433,N_11239);
nand U12585 (N_12585,N_11048,N_11654);
and U12586 (N_12586,N_11420,N_11509);
and U12587 (N_12587,N_11116,N_11301);
xnor U12588 (N_12588,N_11958,N_11586);
nor U12589 (N_12589,N_11923,N_11617);
nor U12590 (N_12590,N_11055,N_11070);
xnor U12591 (N_12591,N_11246,N_11996);
xor U12592 (N_12592,N_11370,N_11048);
or U12593 (N_12593,N_11919,N_11864);
nor U12594 (N_12594,N_11063,N_11876);
or U12595 (N_12595,N_11051,N_11789);
or U12596 (N_12596,N_11537,N_11509);
and U12597 (N_12597,N_11889,N_11510);
nand U12598 (N_12598,N_11912,N_11327);
nor U12599 (N_12599,N_11443,N_11218);
nor U12600 (N_12600,N_11601,N_11031);
or U12601 (N_12601,N_11608,N_11339);
and U12602 (N_12602,N_11599,N_11246);
xnor U12603 (N_12603,N_11720,N_11009);
and U12604 (N_12604,N_11441,N_11310);
nor U12605 (N_12605,N_11207,N_11845);
nor U12606 (N_12606,N_11000,N_11951);
nor U12607 (N_12607,N_11468,N_11677);
nor U12608 (N_12608,N_11125,N_11240);
and U12609 (N_12609,N_11968,N_11005);
and U12610 (N_12610,N_11619,N_11684);
nand U12611 (N_12611,N_11186,N_11757);
nor U12612 (N_12612,N_11104,N_11659);
xnor U12613 (N_12613,N_11010,N_11925);
nor U12614 (N_12614,N_11136,N_11813);
xnor U12615 (N_12615,N_11802,N_11665);
xor U12616 (N_12616,N_11604,N_11219);
nand U12617 (N_12617,N_11512,N_11802);
and U12618 (N_12618,N_11249,N_11118);
and U12619 (N_12619,N_11236,N_11437);
and U12620 (N_12620,N_11834,N_11113);
nor U12621 (N_12621,N_11700,N_11446);
and U12622 (N_12622,N_11019,N_11102);
or U12623 (N_12623,N_11504,N_11620);
nand U12624 (N_12624,N_11268,N_11766);
or U12625 (N_12625,N_11638,N_11705);
or U12626 (N_12626,N_11537,N_11027);
xnor U12627 (N_12627,N_11243,N_11680);
nand U12628 (N_12628,N_11646,N_11129);
or U12629 (N_12629,N_11537,N_11656);
and U12630 (N_12630,N_11523,N_11149);
nand U12631 (N_12631,N_11219,N_11951);
or U12632 (N_12632,N_11707,N_11643);
or U12633 (N_12633,N_11191,N_11287);
nor U12634 (N_12634,N_11638,N_11237);
xor U12635 (N_12635,N_11095,N_11619);
nand U12636 (N_12636,N_11699,N_11423);
nor U12637 (N_12637,N_11428,N_11814);
and U12638 (N_12638,N_11021,N_11405);
or U12639 (N_12639,N_11993,N_11863);
and U12640 (N_12640,N_11135,N_11483);
nand U12641 (N_12641,N_11716,N_11631);
or U12642 (N_12642,N_11761,N_11300);
nor U12643 (N_12643,N_11429,N_11293);
and U12644 (N_12644,N_11816,N_11113);
and U12645 (N_12645,N_11011,N_11521);
xnor U12646 (N_12646,N_11218,N_11161);
nand U12647 (N_12647,N_11055,N_11421);
and U12648 (N_12648,N_11157,N_11078);
nor U12649 (N_12649,N_11136,N_11888);
and U12650 (N_12650,N_11681,N_11638);
or U12651 (N_12651,N_11806,N_11832);
xnor U12652 (N_12652,N_11382,N_11928);
nor U12653 (N_12653,N_11532,N_11063);
nand U12654 (N_12654,N_11123,N_11572);
or U12655 (N_12655,N_11428,N_11897);
and U12656 (N_12656,N_11169,N_11897);
xor U12657 (N_12657,N_11635,N_11174);
nor U12658 (N_12658,N_11413,N_11113);
xor U12659 (N_12659,N_11808,N_11706);
nor U12660 (N_12660,N_11689,N_11716);
xor U12661 (N_12661,N_11158,N_11269);
and U12662 (N_12662,N_11413,N_11498);
and U12663 (N_12663,N_11889,N_11181);
nor U12664 (N_12664,N_11971,N_11548);
xnor U12665 (N_12665,N_11600,N_11989);
and U12666 (N_12666,N_11222,N_11105);
or U12667 (N_12667,N_11106,N_11560);
xnor U12668 (N_12668,N_11198,N_11521);
nor U12669 (N_12669,N_11047,N_11696);
or U12670 (N_12670,N_11295,N_11094);
or U12671 (N_12671,N_11009,N_11140);
and U12672 (N_12672,N_11463,N_11008);
nor U12673 (N_12673,N_11724,N_11602);
and U12674 (N_12674,N_11141,N_11085);
and U12675 (N_12675,N_11932,N_11545);
nor U12676 (N_12676,N_11738,N_11189);
xor U12677 (N_12677,N_11038,N_11690);
nor U12678 (N_12678,N_11103,N_11692);
xnor U12679 (N_12679,N_11409,N_11185);
nor U12680 (N_12680,N_11858,N_11066);
nor U12681 (N_12681,N_11612,N_11303);
and U12682 (N_12682,N_11872,N_11596);
nor U12683 (N_12683,N_11219,N_11012);
or U12684 (N_12684,N_11759,N_11913);
nand U12685 (N_12685,N_11603,N_11782);
xnor U12686 (N_12686,N_11276,N_11460);
nor U12687 (N_12687,N_11435,N_11475);
and U12688 (N_12688,N_11162,N_11804);
nor U12689 (N_12689,N_11309,N_11458);
and U12690 (N_12690,N_11589,N_11910);
or U12691 (N_12691,N_11623,N_11468);
nor U12692 (N_12692,N_11760,N_11380);
xor U12693 (N_12693,N_11857,N_11894);
xnor U12694 (N_12694,N_11241,N_11795);
nor U12695 (N_12695,N_11106,N_11848);
or U12696 (N_12696,N_11555,N_11721);
xnor U12697 (N_12697,N_11223,N_11256);
xnor U12698 (N_12698,N_11811,N_11701);
and U12699 (N_12699,N_11290,N_11556);
nand U12700 (N_12700,N_11858,N_11300);
nand U12701 (N_12701,N_11325,N_11836);
xor U12702 (N_12702,N_11730,N_11606);
and U12703 (N_12703,N_11526,N_11249);
xor U12704 (N_12704,N_11222,N_11776);
nor U12705 (N_12705,N_11190,N_11089);
nand U12706 (N_12706,N_11347,N_11601);
xor U12707 (N_12707,N_11740,N_11562);
xor U12708 (N_12708,N_11795,N_11004);
nor U12709 (N_12709,N_11505,N_11875);
and U12710 (N_12710,N_11999,N_11042);
and U12711 (N_12711,N_11813,N_11310);
or U12712 (N_12712,N_11505,N_11843);
and U12713 (N_12713,N_11520,N_11802);
nor U12714 (N_12714,N_11583,N_11625);
or U12715 (N_12715,N_11596,N_11954);
xor U12716 (N_12716,N_11631,N_11747);
nand U12717 (N_12717,N_11490,N_11532);
or U12718 (N_12718,N_11473,N_11659);
or U12719 (N_12719,N_11668,N_11782);
nand U12720 (N_12720,N_11739,N_11304);
xnor U12721 (N_12721,N_11771,N_11324);
nand U12722 (N_12722,N_11845,N_11582);
xnor U12723 (N_12723,N_11546,N_11945);
nand U12724 (N_12724,N_11782,N_11905);
xnor U12725 (N_12725,N_11882,N_11538);
nor U12726 (N_12726,N_11161,N_11712);
and U12727 (N_12727,N_11047,N_11775);
xnor U12728 (N_12728,N_11201,N_11330);
or U12729 (N_12729,N_11584,N_11103);
nor U12730 (N_12730,N_11416,N_11186);
xnor U12731 (N_12731,N_11421,N_11379);
xnor U12732 (N_12732,N_11656,N_11776);
nand U12733 (N_12733,N_11238,N_11721);
nand U12734 (N_12734,N_11713,N_11374);
xor U12735 (N_12735,N_11423,N_11493);
or U12736 (N_12736,N_11609,N_11278);
and U12737 (N_12737,N_11769,N_11463);
or U12738 (N_12738,N_11922,N_11723);
nand U12739 (N_12739,N_11235,N_11134);
xnor U12740 (N_12740,N_11847,N_11474);
or U12741 (N_12741,N_11004,N_11078);
xnor U12742 (N_12742,N_11673,N_11853);
or U12743 (N_12743,N_11485,N_11690);
or U12744 (N_12744,N_11944,N_11709);
nor U12745 (N_12745,N_11775,N_11939);
or U12746 (N_12746,N_11770,N_11049);
xor U12747 (N_12747,N_11701,N_11867);
or U12748 (N_12748,N_11158,N_11848);
and U12749 (N_12749,N_11468,N_11316);
or U12750 (N_12750,N_11780,N_11851);
or U12751 (N_12751,N_11552,N_11831);
or U12752 (N_12752,N_11163,N_11510);
xnor U12753 (N_12753,N_11362,N_11641);
nand U12754 (N_12754,N_11986,N_11528);
or U12755 (N_12755,N_11278,N_11822);
nor U12756 (N_12756,N_11660,N_11621);
nand U12757 (N_12757,N_11864,N_11105);
or U12758 (N_12758,N_11943,N_11579);
nand U12759 (N_12759,N_11886,N_11912);
xnor U12760 (N_12760,N_11717,N_11276);
nand U12761 (N_12761,N_11383,N_11645);
xor U12762 (N_12762,N_11533,N_11930);
nor U12763 (N_12763,N_11746,N_11180);
nand U12764 (N_12764,N_11402,N_11973);
nor U12765 (N_12765,N_11402,N_11925);
nor U12766 (N_12766,N_11798,N_11072);
and U12767 (N_12767,N_11423,N_11155);
or U12768 (N_12768,N_11231,N_11675);
nand U12769 (N_12769,N_11130,N_11159);
xor U12770 (N_12770,N_11665,N_11119);
nand U12771 (N_12771,N_11409,N_11139);
xnor U12772 (N_12772,N_11355,N_11804);
nand U12773 (N_12773,N_11689,N_11508);
nand U12774 (N_12774,N_11242,N_11847);
or U12775 (N_12775,N_11463,N_11594);
or U12776 (N_12776,N_11594,N_11975);
nand U12777 (N_12777,N_11745,N_11055);
nor U12778 (N_12778,N_11582,N_11369);
nand U12779 (N_12779,N_11261,N_11615);
or U12780 (N_12780,N_11700,N_11288);
or U12781 (N_12781,N_11601,N_11193);
xor U12782 (N_12782,N_11992,N_11263);
nor U12783 (N_12783,N_11871,N_11056);
xor U12784 (N_12784,N_11899,N_11168);
nand U12785 (N_12785,N_11129,N_11033);
xor U12786 (N_12786,N_11844,N_11353);
xor U12787 (N_12787,N_11695,N_11507);
nand U12788 (N_12788,N_11425,N_11496);
and U12789 (N_12789,N_11887,N_11547);
or U12790 (N_12790,N_11541,N_11973);
nor U12791 (N_12791,N_11837,N_11239);
and U12792 (N_12792,N_11118,N_11273);
nor U12793 (N_12793,N_11141,N_11963);
or U12794 (N_12794,N_11393,N_11528);
nand U12795 (N_12795,N_11966,N_11836);
xor U12796 (N_12796,N_11612,N_11033);
nand U12797 (N_12797,N_11561,N_11781);
xnor U12798 (N_12798,N_11037,N_11307);
nor U12799 (N_12799,N_11114,N_11522);
and U12800 (N_12800,N_11090,N_11642);
and U12801 (N_12801,N_11963,N_11773);
xor U12802 (N_12802,N_11906,N_11069);
and U12803 (N_12803,N_11387,N_11070);
nand U12804 (N_12804,N_11084,N_11332);
and U12805 (N_12805,N_11900,N_11311);
nor U12806 (N_12806,N_11972,N_11901);
nand U12807 (N_12807,N_11355,N_11588);
nand U12808 (N_12808,N_11870,N_11891);
nor U12809 (N_12809,N_11737,N_11456);
xor U12810 (N_12810,N_11292,N_11022);
or U12811 (N_12811,N_11213,N_11595);
and U12812 (N_12812,N_11578,N_11563);
nor U12813 (N_12813,N_11024,N_11667);
nand U12814 (N_12814,N_11516,N_11762);
nor U12815 (N_12815,N_11023,N_11583);
and U12816 (N_12816,N_11571,N_11033);
or U12817 (N_12817,N_11076,N_11985);
nor U12818 (N_12818,N_11356,N_11340);
xor U12819 (N_12819,N_11992,N_11231);
xnor U12820 (N_12820,N_11165,N_11983);
nand U12821 (N_12821,N_11986,N_11299);
nor U12822 (N_12822,N_11428,N_11099);
or U12823 (N_12823,N_11708,N_11291);
nor U12824 (N_12824,N_11577,N_11574);
and U12825 (N_12825,N_11626,N_11291);
or U12826 (N_12826,N_11132,N_11461);
nor U12827 (N_12827,N_11368,N_11758);
and U12828 (N_12828,N_11734,N_11946);
xor U12829 (N_12829,N_11326,N_11556);
and U12830 (N_12830,N_11608,N_11464);
or U12831 (N_12831,N_11874,N_11404);
xnor U12832 (N_12832,N_11705,N_11919);
or U12833 (N_12833,N_11133,N_11849);
nor U12834 (N_12834,N_11330,N_11407);
nand U12835 (N_12835,N_11201,N_11288);
and U12836 (N_12836,N_11492,N_11949);
and U12837 (N_12837,N_11630,N_11178);
and U12838 (N_12838,N_11868,N_11030);
or U12839 (N_12839,N_11390,N_11778);
nand U12840 (N_12840,N_11779,N_11009);
nand U12841 (N_12841,N_11666,N_11702);
and U12842 (N_12842,N_11337,N_11128);
or U12843 (N_12843,N_11180,N_11117);
nor U12844 (N_12844,N_11066,N_11479);
or U12845 (N_12845,N_11137,N_11297);
nand U12846 (N_12846,N_11754,N_11736);
and U12847 (N_12847,N_11664,N_11289);
nor U12848 (N_12848,N_11387,N_11832);
and U12849 (N_12849,N_11116,N_11996);
and U12850 (N_12850,N_11797,N_11050);
nor U12851 (N_12851,N_11905,N_11585);
nand U12852 (N_12852,N_11134,N_11559);
xnor U12853 (N_12853,N_11872,N_11150);
xor U12854 (N_12854,N_11479,N_11190);
or U12855 (N_12855,N_11535,N_11338);
nor U12856 (N_12856,N_11973,N_11558);
nor U12857 (N_12857,N_11483,N_11672);
nor U12858 (N_12858,N_11342,N_11778);
or U12859 (N_12859,N_11251,N_11188);
or U12860 (N_12860,N_11951,N_11102);
and U12861 (N_12861,N_11997,N_11877);
and U12862 (N_12862,N_11301,N_11889);
nor U12863 (N_12863,N_11522,N_11574);
xor U12864 (N_12864,N_11455,N_11648);
nor U12865 (N_12865,N_11621,N_11268);
nor U12866 (N_12866,N_11465,N_11844);
or U12867 (N_12867,N_11922,N_11823);
or U12868 (N_12868,N_11701,N_11760);
nand U12869 (N_12869,N_11235,N_11804);
or U12870 (N_12870,N_11994,N_11518);
xor U12871 (N_12871,N_11346,N_11977);
nor U12872 (N_12872,N_11794,N_11166);
and U12873 (N_12873,N_11733,N_11908);
xnor U12874 (N_12874,N_11549,N_11226);
xnor U12875 (N_12875,N_11778,N_11450);
nor U12876 (N_12876,N_11789,N_11284);
xnor U12877 (N_12877,N_11815,N_11416);
xnor U12878 (N_12878,N_11362,N_11834);
xnor U12879 (N_12879,N_11749,N_11596);
or U12880 (N_12880,N_11574,N_11002);
nor U12881 (N_12881,N_11552,N_11657);
nor U12882 (N_12882,N_11364,N_11471);
xor U12883 (N_12883,N_11692,N_11889);
nand U12884 (N_12884,N_11334,N_11346);
nand U12885 (N_12885,N_11425,N_11125);
nor U12886 (N_12886,N_11396,N_11343);
xor U12887 (N_12887,N_11794,N_11046);
nor U12888 (N_12888,N_11151,N_11937);
or U12889 (N_12889,N_11244,N_11956);
nor U12890 (N_12890,N_11305,N_11147);
and U12891 (N_12891,N_11079,N_11131);
xor U12892 (N_12892,N_11917,N_11735);
nand U12893 (N_12893,N_11536,N_11026);
xnor U12894 (N_12894,N_11489,N_11568);
and U12895 (N_12895,N_11721,N_11278);
and U12896 (N_12896,N_11998,N_11567);
xor U12897 (N_12897,N_11947,N_11227);
xor U12898 (N_12898,N_11122,N_11895);
xor U12899 (N_12899,N_11948,N_11427);
xor U12900 (N_12900,N_11670,N_11545);
xor U12901 (N_12901,N_11312,N_11465);
xor U12902 (N_12902,N_11704,N_11005);
or U12903 (N_12903,N_11565,N_11693);
nor U12904 (N_12904,N_11592,N_11856);
xnor U12905 (N_12905,N_11000,N_11312);
nor U12906 (N_12906,N_11522,N_11327);
and U12907 (N_12907,N_11966,N_11044);
nand U12908 (N_12908,N_11909,N_11198);
or U12909 (N_12909,N_11626,N_11832);
nor U12910 (N_12910,N_11252,N_11245);
and U12911 (N_12911,N_11737,N_11031);
and U12912 (N_12912,N_11022,N_11087);
nor U12913 (N_12913,N_11901,N_11650);
and U12914 (N_12914,N_11886,N_11036);
and U12915 (N_12915,N_11161,N_11099);
and U12916 (N_12916,N_11315,N_11142);
and U12917 (N_12917,N_11948,N_11373);
nand U12918 (N_12918,N_11036,N_11603);
or U12919 (N_12919,N_11920,N_11354);
xor U12920 (N_12920,N_11333,N_11245);
and U12921 (N_12921,N_11175,N_11001);
or U12922 (N_12922,N_11436,N_11382);
nor U12923 (N_12923,N_11197,N_11732);
nor U12924 (N_12924,N_11335,N_11459);
nor U12925 (N_12925,N_11805,N_11255);
or U12926 (N_12926,N_11493,N_11029);
xnor U12927 (N_12927,N_11338,N_11481);
nor U12928 (N_12928,N_11088,N_11734);
nand U12929 (N_12929,N_11108,N_11733);
or U12930 (N_12930,N_11378,N_11275);
nand U12931 (N_12931,N_11666,N_11483);
nor U12932 (N_12932,N_11989,N_11416);
nand U12933 (N_12933,N_11182,N_11338);
and U12934 (N_12934,N_11157,N_11190);
or U12935 (N_12935,N_11063,N_11436);
nand U12936 (N_12936,N_11783,N_11686);
nand U12937 (N_12937,N_11655,N_11722);
nand U12938 (N_12938,N_11882,N_11237);
and U12939 (N_12939,N_11564,N_11204);
or U12940 (N_12940,N_11794,N_11807);
and U12941 (N_12941,N_11334,N_11482);
or U12942 (N_12942,N_11138,N_11370);
and U12943 (N_12943,N_11907,N_11444);
nor U12944 (N_12944,N_11284,N_11640);
or U12945 (N_12945,N_11300,N_11924);
or U12946 (N_12946,N_11130,N_11528);
xor U12947 (N_12947,N_11396,N_11692);
nor U12948 (N_12948,N_11752,N_11572);
or U12949 (N_12949,N_11998,N_11927);
nor U12950 (N_12950,N_11866,N_11078);
nand U12951 (N_12951,N_11876,N_11628);
or U12952 (N_12952,N_11419,N_11841);
xor U12953 (N_12953,N_11650,N_11094);
and U12954 (N_12954,N_11671,N_11088);
and U12955 (N_12955,N_11639,N_11819);
and U12956 (N_12956,N_11698,N_11380);
or U12957 (N_12957,N_11713,N_11207);
or U12958 (N_12958,N_11712,N_11134);
nand U12959 (N_12959,N_11842,N_11574);
and U12960 (N_12960,N_11347,N_11279);
and U12961 (N_12961,N_11443,N_11688);
nor U12962 (N_12962,N_11728,N_11525);
xnor U12963 (N_12963,N_11838,N_11227);
and U12964 (N_12964,N_11620,N_11877);
nand U12965 (N_12965,N_11550,N_11744);
xnor U12966 (N_12966,N_11477,N_11588);
and U12967 (N_12967,N_11497,N_11554);
nor U12968 (N_12968,N_11868,N_11653);
and U12969 (N_12969,N_11060,N_11709);
xor U12970 (N_12970,N_11257,N_11465);
xor U12971 (N_12971,N_11435,N_11681);
or U12972 (N_12972,N_11801,N_11299);
nor U12973 (N_12973,N_11534,N_11187);
nand U12974 (N_12974,N_11196,N_11279);
nor U12975 (N_12975,N_11693,N_11311);
nor U12976 (N_12976,N_11094,N_11949);
xnor U12977 (N_12977,N_11230,N_11733);
nand U12978 (N_12978,N_11888,N_11865);
nor U12979 (N_12979,N_11442,N_11435);
nor U12980 (N_12980,N_11328,N_11629);
xor U12981 (N_12981,N_11567,N_11685);
nand U12982 (N_12982,N_11298,N_11203);
or U12983 (N_12983,N_11138,N_11083);
nor U12984 (N_12984,N_11601,N_11322);
nor U12985 (N_12985,N_11934,N_11049);
nor U12986 (N_12986,N_11889,N_11756);
xor U12987 (N_12987,N_11899,N_11572);
or U12988 (N_12988,N_11976,N_11299);
nor U12989 (N_12989,N_11059,N_11223);
nor U12990 (N_12990,N_11210,N_11108);
nor U12991 (N_12991,N_11392,N_11996);
or U12992 (N_12992,N_11946,N_11159);
nor U12993 (N_12993,N_11449,N_11418);
nor U12994 (N_12994,N_11904,N_11711);
nor U12995 (N_12995,N_11935,N_11987);
nor U12996 (N_12996,N_11550,N_11917);
and U12997 (N_12997,N_11431,N_11665);
xnor U12998 (N_12998,N_11467,N_11925);
or U12999 (N_12999,N_11657,N_11754);
and U13000 (N_13000,N_12317,N_12556);
xnor U13001 (N_13001,N_12587,N_12925);
or U13002 (N_13002,N_12467,N_12130);
or U13003 (N_13003,N_12448,N_12847);
xor U13004 (N_13004,N_12204,N_12672);
xor U13005 (N_13005,N_12215,N_12503);
xor U13006 (N_13006,N_12733,N_12165);
or U13007 (N_13007,N_12606,N_12398);
xor U13008 (N_13008,N_12299,N_12761);
nand U13009 (N_13009,N_12133,N_12937);
or U13010 (N_13010,N_12458,N_12452);
and U13011 (N_13011,N_12703,N_12167);
and U13012 (N_13012,N_12978,N_12891);
or U13013 (N_13013,N_12478,N_12386);
nor U13014 (N_13014,N_12298,N_12081);
nand U13015 (N_13015,N_12617,N_12673);
and U13016 (N_13016,N_12479,N_12849);
and U13017 (N_13017,N_12786,N_12820);
nand U13018 (N_13018,N_12529,N_12087);
nand U13019 (N_13019,N_12865,N_12358);
nor U13020 (N_13020,N_12561,N_12474);
nor U13021 (N_13021,N_12676,N_12366);
nor U13022 (N_13022,N_12486,N_12570);
or U13023 (N_13023,N_12579,N_12297);
nand U13024 (N_13024,N_12367,N_12116);
xor U13025 (N_13025,N_12435,N_12287);
xor U13026 (N_13026,N_12874,N_12641);
or U13027 (N_13027,N_12235,N_12692);
nor U13028 (N_13028,N_12150,N_12686);
or U13029 (N_13029,N_12885,N_12162);
xor U13030 (N_13030,N_12019,N_12433);
and U13031 (N_13031,N_12875,N_12163);
and U13032 (N_13032,N_12645,N_12110);
and U13033 (N_13033,N_12039,N_12611);
and U13034 (N_13034,N_12376,N_12113);
nor U13035 (N_13035,N_12199,N_12091);
or U13036 (N_13036,N_12315,N_12043);
xor U13037 (N_13037,N_12040,N_12950);
and U13038 (N_13038,N_12339,N_12998);
nor U13039 (N_13039,N_12881,N_12258);
xor U13040 (N_13040,N_12807,N_12890);
and U13041 (N_13041,N_12249,N_12330);
xnor U13042 (N_13042,N_12603,N_12077);
and U13043 (N_13043,N_12922,N_12500);
xor U13044 (N_13044,N_12403,N_12082);
or U13045 (N_13045,N_12661,N_12624);
and U13046 (N_13046,N_12353,N_12909);
and U13047 (N_13047,N_12089,N_12418);
xor U13048 (N_13048,N_12602,N_12827);
nand U13049 (N_13049,N_12651,N_12101);
nand U13050 (N_13050,N_12578,N_12908);
xor U13051 (N_13051,N_12273,N_12001);
nand U13052 (N_13052,N_12805,N_12658);
xor U13053 (N_13053,N_12528,N_12377);
and U13054 (N_13054,N_12427,N_12128);
xnor U13055 (N_13055,N_12970,N_12341);
or U13056 (N_13056,N_12011,N_12973);
xnor U13057 (N_13057,N_12322,N_12927);
xnor U13058 (N_13058,N_12473,N_12111);
nor U13059 (N_13059,N_12234,N_12489);
or U13060 (N_13060,N_12835,N_12302);
xor U13061 (N_13061,N_12421,N_12904);
nor U13062 (N_13062,N_12949,N_12387);
nor U13063 (N_13063,N_12018,N_12092);
nor U13064 (N_13064,N_12769,N_12394);
xnor U13065 (N_13065,N_12056,N_12153);
xnor U13066 (N_13066,N_12717,N_12682);
xor U13067 (N_13067,N_12806,N_12269);
and U13068 (N_13068,N_12918,N_12044);
nor U13069 (N_13069,N_12935,N_12510);
nand U13070 (N_13070,N_12469,N_12090);
nor U13071 (N_13071,N_12329,N_12375);
nand U13072 (N_13072,N_12758,N_12751);
and U13073 (N_13073,N_12824,N_12552);
xnor U13074 (N_13074,N_12272,N_12408);
nor U13075 (N_13075,N_12047,N_12161);
nand U13076 (N_13076,N_12430,N_12357);
and U13077 (N_13077,N_12100,N_12932);
and U13078 (N_13078,N_12213,N_12714);
nand U13079 (N_13079,N_12581,N_12863);
and U13080 (N_13080,N_12356,N_12680);
nor U13081 (N_13081,N_12247,N_12037);
nor U13082 (N_13082,N_12837,N_12476);
nor U13083 (N_13083,N_12811,N_12447);
nor U13084 (N_13084,N_12814,N_12822);
and U13085 (N_13085,N_12248,N_12880);
and U13086 (N_13086,N_12777,N_12347);
nand U13087 (N_13087,N_12054,N_12208);
nand U13088 (N_13088,N_12886,N_12194);
xnor U13089 (N_13089,N_12156,N_12482);
nor U13090 (N_13090,N_12210,N_12472);
nand U13091 (N_13091,N_12862,N_12960);
or U13092 (N_13092,N_12228,N_12283);
nand U13093 (N_13093,N_12220,N_12155);
or U13094 (N_13094,N_12568,N_12064);
nand U13095 (N_13095,N_12866,N_12559);
nor U13096 (N_13096,N_12939,N_12662);
nand U13097 (N_13097,N_12523,N_12059);
and U13098 (N_13098,N_12031,N_12384);
xor U13099 (N_13099,N_12691,N_12744);
and U13100 (N_13100,N_12237,N_12615);
nand U13101 (N_13101,N_12493,N_12346);
and U13102 (N_13102,N_12506,N_12522);
nor U13103 (N_13103,N_12170,N_12901);
nand U13104 (N_13104,N_12225,N_12352);
nor U13105 (N_13105,N_12631,N_12738);
nor U13106 (N_13106,N_12134,N_12505);
and U13107 (N_13107,N_12660,N_12069);
and U13108 (N_13108,N_12079,N_12099);
xnor U13109 (N_13109,N_12028,N_12034);
xnor U13110 (N_13110,N_12223,N_12819);
nand U13111 (N_13111,N_12203,N_12311);
or U13112 (N_13112,N_12067,N_12701);
nor U13113 (N_13113,N_12218,N_12548);
nand U13114 (N_13114,N_12294,N_12838);
xnor U13115 (N_13115,N_12928,N_12956);
and U13116 (N_13116,N_12191,N_12335);
xor U13117 (N_13117,N_12931,N_12852);
nand U13118 (N_13118,N_12279,N_12491);
or U13119 (N_13119,N_12321,N_12245);
or U13120 (N_13120,N_12251,N_12065);
or U13121 (N_13121,N_12966,N_12685);
nor U13122 (N_13122,N_12817,N_12823);
nand U13123 (N_13123,N_12541,N_12834);
nand U13124 (N_13124,N_12816,N_12916);
and U13125 (N_13125,N_12637,N_12792);
nor U13126 (N_13126,N_12010,N_12072);
nand U13127 (N_13127,N_12889,N_12566);
nor U13128 (N_13128,N_12504,N_12319);
nand U13129 (N_13129,N_12549,N_12695);
nand U13130 (N_13130,N_12118,N_12564);
and U13131 (N_13131,N_12576,N_12991);
or U13132 (N_13132,N_12976,N_12182);
and U13133 (N_13133,N_12188,N_12732);
and U13134 (N_13134,N_12005,N_12129);
nor U13135 (N_13135,N_12774,N_12597);
and U13136 (N_13136,N_12871,N_12303);
nand U13137 (N_13137,N_12396,N_12078);
xnor U13138 (N_13138,N_12798,N_12599);
or U13139 (N_13139,N_12052,N_12584);
nor U13140 (N_13140,N_12892,N_12953);
xnor U13141 (N_13141,N_12519,N_12093);
xor U13142 (N_13142,N_12135,N_12669);
xnor U13143 (N_13143,N_12230,N_12944);
nand U13144 (N_13144,N_12759,N_12531);
or U13145 (N_13145,N_12270,N_12754);
nor U13146 (N_13146,N_12259,N_12829);
xnor U13147 (N_13147,N_12562,N_12762);
or U13148 (N_13148,N_12923,N_12502);
nand U13149 (N_13149,N_12912,N_12670);
and U13150 (N_13150,N_12383,N_12989);
and U13151 (N_13151,N_12217,N_12640);
xnor U13152 (N_13152,N_12420,N_12105);
or U13153 (N_13153,N_12103,N_12859);
xor U13154 (N_13154,N_12511,N_12098);
xor U13155 (N_13155,N_12285,N_12626);
xnor U13156 (N_13156,N_12343,N_12195);
or U13157 (N_13157,N_12015,N_12715);
xnor U13158 (N_13158,N_12961,N_12588);
xor U13159 (N_13159,N_12119,N_12924);
nor U13160 (N_13160,N_12955,N_12021);
and U13161 (N_13161,N_12483,N_12362);
or U13162 (N_13162,N_12630,N_12437);
xor U13163 (N_13163,N_12485,N_12409);
nor U13164 (N_13164,N_12340,N_12397);
and U13165 (N_13165,N_12982,N_12905);
and U13166 (N_13166,N_12184,N_12494);
or U13167 (N_13167,N_12591,N_12075);
xor U13168 (N_13168,N_12898,N_12202);
nand U13169 (N_13169,N_12550,N_12694);
xnor U13170 (N_13170,N_12333,N_12414);
and U13171 (N_13171,N_12328,N_12567);
xor U13172 (N_13172,N_12913,N_12756);
nand U13173 (N_13173,N_12013,N_12232);
nor U13174 (N_13174,N_12413,N_12757);
and U13175 (N_13175,N_12041,N_12618);
xor U13176 (N_13176,N_12647,N_12058);
and U13177 (N_13177,N_12836,N_12320);
xnor U13178 (N_13178,N_12154,N_12546);
nor U13179 (N_13179,N_12117,N_12716);
nand U13180 (N_13180,N_12266,N_12454);
or U13181 (N_13181,N_12586,N_12623);
xnor U13182 (N_13182,N_12760,N_12293);
nand U13183 (N_13183,N_12492,N_12276);
nor U13184 (N_13184,N_12309,N_12793);
and U13185 (N_13185,N_12697,N_12974);
nand U13186 (N_13186,N_12867,N_12709);
nand U13187 (N_13187,N_12783,N_12943);
and U13188 (N_13188,N_12080,N_12284);
and U13189 (N_13189,N_12419,N_12780);
nand U13190 (N_13190,N_12390,N_12027);
nand U13191 (N_13191,N_12126,N_12681);
nand U13192 (N_13192,N_12903,N_12629);
nor U13193 (N_13193,N_12209,N_12667);
xnor U13194 (N_13194,N_12710,N_12085);
nor U13195 (N_13195,N_12378,N_12896);
nand U13196 (N_13196,N_12766,N_12275);
nor U13197 (N_13197,N_12149,N_12304);
or U13198 (N_13198,N_12845,N_12261);
xnor U13199 (N_13199,N_12712,N_12456);
or U13200 (N_13200,N_12198,N_12380);
or U13201 (N_13201,N_12742,N_12288);
or U13202 (N_13202,N_12665,N_12609);
or U13203 (N_13203,N_12003,N_12241);
or U13204 (N_13204,N_12365,N_12997);
nand U13205 (N_13205,N_12264,N_12590);
and U13206 (N_13206,N_12171,N_12671);
and U13207 (N_13207,N_12410,N_12625);
and U13208 (N_13208,N_12547,N_12515);
xnor U13209 (N_13209,N_12812,N_12291);
and U13210 (N_13210,N_12239,N_12879);
and U13211 (N_13211,N_12533,N_12233);
and U13212 (N_13212,N_12652,N_12152);
nor U13213 (N_13213,N_12364,N_12371);
nand U13214 (N_13214,N_12514,N_12443);
nand U13215 (N_13215,N_12577,N_12596);
or U13216 (N_13216,N_12450,N_12363);
and U13217 (N_13217,N_12109,N_12628);
nand U13218 (N_13218,N_12844,N_12051);
xnor U13219 (N_13219,N_12265,N_12422);
xnor U13220 (N_13220,N_12172,N_12643);
nor U13221 (N_13221,N_12538,N_12983);
xor U13222 (N_13222,N_12157,N_12164);
and U13223 (N_13223,N_12555,N_12839);
or U13224 (N_13224,N_12663,N_12438);
and U13225 (N_13225,N_12023,N_12608);
and U13226 (N_13226,N_12726,N_12114);
and U13227 (N_13227,N_12711,N_12342);
xor U13228 (N_13228,N_12029,N_12799);
nand U13229 (N_13229,N_12179,N_12132);
or U13230 (N_13230,N_12992,N_12038);
nand U13231 (N_13231,N_12461,N_12959);
nand U13232 (N_13232,N_12169,N_12719);
and U13233 (N_13233,N_12189,N_12668);
xnor U13234 (N_13234,N_12996,N_12930);
and U13235 (N_13235,N_12086,N_12281);
or U13236 (N_13236,N_12873,N_12739);
and U13237 (N_13237,N_12292,N_12148);
xor U13238 (N_13238,N_12355,N_12583);
or U13239 (N_13239,N_12470,N_12369);
xor U13240 (N_13240,N_12988,N_12395);
or U13241 (N_13241,N_12030,N_12296);
nand U13242 (N_13242,N_12706,N_12635);
or U13243 (N_13243,N_12776,N_12809);
xor U13244 (N_13244,N_12735,N_12573);
or U13245 (N_13245,N_12620,N_12929);
xor U13246 (N_13246,N_12053,N_12429);
xor U13247 (N_13247,N_12804,N_12004);
and U13248 (N_13248,N_12687,N_12083);
xor U13249 (N_13249,N_12700,N_12379);
nor U13250 (N_13250,N_12604,N_12073);
xnor U13251 (N_13251,N_12723,N_12752);
nand U13252 (N_13252,N_12071,N_12894);
and U13253 (N_13253,N_12477,N_12778);
and U13254 (N_13254,N_12813,N_12840);
or U13255 (N_13255,N_12598,N_12971);
and U13256 (N_13256,N_12858,N_12061);
xor U13257 (N_13257,N_12571,N_12619);
or U13258 (N_13258,N_12183,N_12785);
xnor U13259 (N_13259,N_12545,N_12987);
and U13260 (N_13260,N_12775,N_12747);
nand U13261 (N_13261,N_12144,N_12262);
nor U13262 (N_13262,N_12893,N_12428);
or U13263 (N_13263,N_12440,N_12490);
and U13264 (N_13264,N_12451,N_12818);
xor U13265 (N_13265,N_12475,N_12301);
or U13266 (N_13266,N_12076,N_12108);
and U13267 (N_13267,N_12354,N_12800);
xor U13268 (N_13268,N_12095,N_12808);
nor U13269 (N_13269,N_12593,N_12316);
xnor U13270 (N_13270,N_12666,N_12802);
nor U13271 (N_13271,N_12268,N_12853);
and U13272 (N_13272,N_12878,N_12979);
nand U13273 (N_13273,N_12012,N_12260);
and U13274 (N_13274,N_12190,N_12951);
or U13275 (N_13275,N_12580,N_12734);
xor U13276 (N_13276,N_12883,N_12627);
xnor U13277 (N_13277,N_12737,N_12002);
nor U13278 (N_13278,N_12977,N_12934);
xnor U13279 (N_13279,N_12045,N_12096);
nor U13280 (N_13280,N_12147,N_12324);
xnor U13281 (N_13281,N_12240,N_12351);
nor U13282 (N_13282,N_12280,N_12825);
and U13283 (N_13283,N_12677,N_12787);
nand U13284 (N_13284,N_12389,N_12142);
or U13285 (N_13285,N_12035,N_12212);
nor U13286 (N_13286,N_12616,N_12050);
nand U13287 (N_13287,N_12911,N_12753);
nor U13288 (N_13288,N_12193,N_12882);
or U13289 (N_13289,N_12139,N_12516);
nor U13290 (N_13290,N_12917,N_12244);
nor U13291 (N_13291,N_12958,N_12632);
nor U13292 (N_13292,N_12622,N_12789);
xnor U13293 (N_13293,N_12993,N_12196);
xor U13294 (N_13294,N_12967,N_12143);
nor U13295 (N_13295,N_12984,N_12674);
nor U13296 (N_13296,N_12690,N_12860);
and U13297 (N_13297,N_12205,N_12401);
nand U13298 (N_13298,N_12382,N_12920);
nand U13299 (N_13299,N_12595,N_12610);
and U13300 (N_13300,N_12138,N_12256);
nand U13301 (N_13301,N_12543,N_12495);
nor U13302 (N_13302,N_12306,N_12068);
or U13303 (N_13303,N_12381,N_12634);
and U13304 (N_13304,N_12392,N_12323);
or U13305 (N_13305,N_12400,N_12286);
and U13306 (N_13306,N_12565,N_12066);
nand U13307 (N_13307,N_12036,N_12530);
nand U13308 (N_13308,N_12872,N_12963);
nor U13309 (N_13309,N_12417,N_12919);
and U13310 (N_13310,N_12185,N_12946);
and U13311 (N_13311,N_12063,N_12947);
nand U13312 (N_13312,N_12763,N_12981);
nor U13313 (N_13313,N_12022,N_12411);
xor U13314 (N_13314,N_12954,N_12334);
or U13315 (N_13315,N_12795,N_12915);
nor U13316 (N_13316,N_12062,N_12102);
xnor U13317 (N_13317,N_12656,N_12704);
nor U13318 (N_13318,N_12601,N_12277);
xor U13319 (N_13319,N_12553,N_12788);
xor U13320 (N_13320,N_12459,N_12254);
or U13321 (N_13321,N_12646,N_12856);
xor U13322 (N_13322,N_12746,N_12537);
xnor U13323 (N_13323,N_12696,N_12074);
nand U13324 (N_13324,N_12655,N_12024);
and U13325 (N_13325,N_12159,N_12846);
nand U13326 (N_13326,N_12173,N_12527);
and U13327 (N_13327,N_12621,N_12832);
xor U13328 (N_13328,N_12471,N_12263);
nor U13329 (N_13329,N_12166,N_12344);
and U13330 (N_13330,N_12693,N_12921);
and U13331 (N_13331,N_12563,N_12532);
nand U13332 (N_13332,N_12325,N_12684);
and U13333 (N_13333,N_12121,N_12509);
and U13334 (N_13334,N_12941,N_12033);
or U13335 (N_13335,N_12999,N_12048);
and U13336 (N_13336,N_12679,N_12815);
xor U13337 (N_13337,N_12942,N_12592);
xor U13338 (N_13338,N_12453,N_12614);
or U13339 (N_13339,N_12952,N_12252);
nand U13340 (N_13340,N_12174,N_12388);
and U13341 (N_13341,N_12231,N_12736);
and U13342 (N_13342,N_12508,N_12902);
and U13343 (N_13343,N_12442,N_12446);
xor U13344 (N_13344,N_12675,N_12463);
xnor U13345 (N_13345,N_12131,N_12897);
and U13346 (N_13346,N_12855,N_12006);
and U13347 (N_13347,N_12496,N_12748);
or U13348 (N_13348,N_12243,N_12227);
nand U13349 (N_13349,N_12585,N_12698);
nor U13350 (N_13350,N_12124,N_12416);
and U13351 (N_13351,N_12107,N_12965);
or U13352 (N_13352,N_12187,N_12370);
nor U13353 (N_13353,N_12449,N_12644);
nand U13354 (N_13354,N_12542,N_12127);
xnor U13355 (N_13355,N_12851,N_12554);
nor U13356 (N_13356,N_12801,N_12831);
or U13357 (N_13357,N_12141,N_12192);
xor U13358 (N_13358,N_12841,N_12600);
nand U13359 (N_13359,N_12740,N_12374);
xor U13360 (N_13360,N_12525,N_12638);
and U13361 (N_13361,N_12308,N_12899);
or U13362 (N_13362,N_12009,N_12368);
or U13363 (N_13363,N_12995,N_12331);
nor U13364 (N_13364,N_12750,N_12488);
xor U13365 (N_13365,N_12558,N_12854);
and U13366 (N_13366,N_12499,N_12313);
nor U13367 (N_13367,N_12178,N_12391);
xor U13368 (N_13368,N_12794,N_12796);
nor U13369 (N_13369,N_12907,N_12683);
xor U13370 (N_13370,N_12295,N_12821);
nand U13371 (N_13371,N_12426,N_12791);
xor U13372 (N_13372,N_12945,N_12664);
xnor U13373 (N_13373,N_12481,N_12876);
nand U13374 (N_13374,N_12016,N_12201);
or U13375 (N_13375,N_12415,N_12106);
nand U13376 (N_13376,N_12372,N_12200);
xor U13377 (N_13377,N_12968,N_12221);
nand U13378 (N_13378,N_12137,N_12650);
and U13379 (N_13379,N_12526,N_12219);
nand U13380 (N_13380,N_12521,N_12713);
nor U13381 (N_13381,N_12699,N_12432);
and U13382 (N_13382,N_12348,N_12112);
xnor U13383 (N_13383,N_12517,N_12910);
nor U13384 (N_13384,N_12975,N_12326);
and U13385 (N_13385,N_12678,N_12764);
xor U13386 (N_13386,N_12688,N_12868);
nand U13387 (N_13387,N_12255,N_12743);
nand U13388 (N_13388,N_12345,N_12007);
and U13389 (N_13389,N_12642,N_12771);
nor U13390 (N_13390,N_12933,N_12373);
xor U13391 (N_13391,N_12540,N_12175);
nor U13392 (N_13392,N_12722,N_12008);
and U13393 (N_13393,N_12507,N_12441);
or U13394 (N_13394,N_12468,N_12307);
xnor U13395 (N_13395,N_12487,N_12431);
xnor U13396 (N_13396,N_12745,N_12572);
and U13397 (N_13397,N_12749,N_12728);
nand U13398 (N_13398,N_12768,N_12123);
nor U13399 (N_13399,N_12501,N_12861);
nor U13400 (N_13400,N_12790,N_12659);
xor U13401 (N_13401,N_12057,N_12779);
xor U13402 (N_13402,N_12569,N_12186);
and U13403 (N_13403,N_12848,N_12434);
nand U13404 (N_13404,N_12639,N_12484);
xnor U13405 (N_13405,N_12551,N_12936);
xnor U13406 (N_13406,N_12151,N_12407);
xor U13407 (N_13407,N_12177,N_12765);
xor U13408 (N_13408,N_12888,N_12842);
nor U13409 (N_13409,N_12857,N_12594);
xnor U13410 (N_13410,N_12120,N_12636);
nor U13411 (N_13411,N_12877,N_12439);
xnor U13412 (N_13412,N_12870,N_12084);
nor U13413 (N_13413,N_12957,N_12654);
or U13414 (N_13414,N_12513,N_12246);
xor U13415 (N_13415,N_12168,N_12136);
xor U13416 (N_13416,N_12055,N_12257);
or U13417 (N_13417,N_12406,N_12338);
and U13418 (N_13418,N_12725,N_12094);
and U13419 (N_13419,N_12361,N_12727);
and U13420 (N_13420,N_12560,N_12582);
nor U13421 (N_13421,N_12480,N_12990);
nand U13422 (N_13422,N_12702,N_12412);
and U13423 (N_13423,N_12557,N_12349);
or U13424 (N_13424,N_12884,N_12803);
or U13425 (N_13425,N_12327,N_12336);
xnor U13426 (N_13426,N_12176,N_12300);
nor U13427 (N_13427,N_12305,N_12088);
and U13428 (N_13428,N_12657,N_12278);
xnor U13429 (N_13429,N_12207,N_12964);
and U13430 (N_13430,N_12773,N_12539);
xor U13431 (N_13431,N_12574,N_12310);
and U13432 (N_13432,N_12536,N_12402);
or U13433 (N_13433,N_12140,N_12000);
nand U13434 (N_13434,N_12181,N_12455);
nand U13435 (N_13435,N_12843,N_12986);
and U13436 (N_13436,N_12466,N_12026);
nand U13437 (N_13437,N_12914,N_12464);
and U13438 (N_13438,N_12253,N_12014);
xnor U13439 (N_13439,N_12158,N_12980);
nor U13440 (N_13440,N_12830,N_12948);
nand U13441 (N_13441,N_12332,N_12512);
nor U13442 (N_13442,N_12236,N_12544);
nand U13443 (N_13443,N_12046,N_12613);
nor U13444 (N_13444,N_12767,N_12729);
xnor U13445 (N_13445,N_12360,N_12926);
nand U13446 (N_13446,N_12520,N_12720);
nand U13447 (N_13447,N_12070,N_12274);
or U13448 (N_13448,N_12772,N_12985);
nor U13449 (N_13449,N_12457,N_12906);
or U13450 (N_13450,N_12810,N_12589);
xor U13451 (N_13451,N_12730,N_12721);
or U13452 (N_13452,N_12180,N_12900);
nand U13453 (N_13453,N_12689,N_12850);
xor U13454 (N_13454,N_12049,N_12424);
nor U13455 (N_13455,N_12969,N_12755);
and U13456 (N_13456,N_12146,N_12648);
xnor U13457 (N_13457,N_12828,N_12032);
and U13458 (N_13458,N_12497,N_12797);
nor U13459 (N_13459,N_12115,N_12020);
and U13460 (N_13460,N_12518,N_12607);
and U13461 (N_13461,N_12781,N_12226);
or U13462 (N_13462,N_12887,N_12465);
nor U13463 (N_13463,N_12864,N_12318);
nor U13464 (N_13464,N_12229,N_12612);
and U13465 (N_13465,N_12122,N_12826);
nand U13466 (N_13466,N_12242,N_12404);
or U13467 (N_13467,N_12962,N_12312);
xor U13468 (N_13468,N_12206,N_12605);
xor U13469 (N_13469,N_12445,N_12423);
and U13470 (N_13470,N_12160,N_12104);
nand U13471 (N_13471,N_12940,N_12633);
nor U13472 (N_13472,N_12267,N_12385);
xnor U13473 (N_13473,N_12216,N_12708);
nor U13474 (N_13474,N_12718,N_12994);
xor U13475 (N_13475,N_12833,N_12425);
and U13476 (N_13476,N_12271,N_12222);
nor U13477 (N_13477,N_12337,N_12314);
or U13478 (N_13478,N_12224,N_12741);
xor U13479 (N_13479,N_12462,N_12350);
or U13480 (N_13480,N_12869,N_12705);
nand U13481 (N_13481,N_12653,N_12972);
or U13482 (N_13482,N_12444,N_12405);
nor U13483 (N_13483,N_12290,N_12782);
nor U13484 (N_13484,N_12197,N_12707);
xnor U13485 (N_13485,N_12289,N_12524);
and U13486 (N_13486,N_12724,N_12731);
nor U13487 (N_13487,N_12393,N_12784);
xnor U13488 (N_13488,N_12498,N_12895);
or U13489 (N_13489,N_12534,N_12025);
nand U13490 (N_13490,N_12535,N_12282);
nand U13491 (N_13491,N_12359,N_12399);
nor U13492 (N_13492,N_12017,N_12145);
or U13493 (N_13493,N_12214,N_12250);
and U13494 (N_13494,N_12125,N_12042);
nand U13495 (N_13495,N_12211,N_12649);
xnor U13496 (N_13496,N_12770,N_12060);
or U13497 (N_13497,N_12097,N_12575);
and U13498 (N_13498,N_12460,N_12938);
and U13499 (N_13499,N_12238,N_12436);
nand U13500 (N_13500,N_12055,N_12866);
nor U13501 (N_13501,N_12883,N_12571);
nor U13502 (N_13502,N_12855,N_12749);
and U13503 (N_13503,N_12484,N_12420);
and U13504 (N_13504,N_12481,N_12087);
nor U13505 (N_13505,N_12002,N_12828);
xor U13506 (N_13506,N_12893,N_12483);
xor U13507 (N_13507,N_12849,N_12854);
or U13508 (N_13508,N_12747,N_12594);
nand U13509 (N_13509,N_12043,N_12505);
nand U13510 (N_13510,N_12822,N_12881);
nand U13511 (N_13511,N_12000,N_12453);
nand U13512 (N_13512,N_12261,N_12796);
nor U13513 (N_13513,N_12319,N_12490);
and U13514 (N_13514,N_12879,N_12657);
and U13515 (N_13515,N_12015,N_12975);
nor U13516 (N_13516,N_12182,N_12974);
nand U13517 (N_13517,N_12768,N_12677);
or U13518 (N_13518,N_12130,N_12147);
xnor U13519 (N_13519,N_12845,N_12309);
xor U13520 (N_13520,N_12263,N_12547);
or U13521 (N_13521,N_12049,N_12055);
nor U13522 (N_13522,N_12447,N_12367);
xor U13523 (N_13523,N_12771,N_12098);
or U13524 (N_13524,N_12501,N_12085);
nand U13525 (N_13525,N_12311,N_12610);
nand U13526 (N_13526,N_12781,N_12299);
and U13527 (N_13527,N_12173,N_12828);
nor U13528 (N_13528,N_12016,N_12234);
and U13529 (N_13529,N_12953,N_12121);
xor U13530 (N_13530,N_12121,N_12817);
and U13531 (N_13531,N_12648,N_12687);
and U13532 (N_13532,N_12480,N_12779);
xor U13533 (N_13533,N_12375,N_12801);
and U13534 (N_13534,N_12372,N_12554);
and U13535 (N_13535,N_12460,N_12794);
and U13536 (N_13536,N_12853,N_12761);
nand U13537 (N_13537,N_12838,N_12471);
nor U13538 (N_13538,N_12380,N_12017);
xor U13539 (N_13539,N_12071,N_12006);
nor U13540 (N_13540,N_12757,N_12848);
nor U13541 (N_13541,N_12080,N_12470);
xor U13542 (N_13542,N_12741,N_12937);
xor U13543 (N_13543,N_12905,N_12367);
nor U13544 (N_13544,N_12550,N_12281);
nand U13545 (N_13545,N_12991,N_12141);
and U13546 (N_13546,N_12247,N_12113);
or U13547 (N_13547,N_12266,N_12554);
and U13548 (N_13548,N_12077,N_12395);
xnor U13549 (N_13549,N_12454,N_12838);
nand U13550 (N_13550,N_12255,N_12267);
and U13551 (N_13551,N_12228,N_12999);
nor U13552 (N_13552,N_12197,N_12990);
and U13553 (N_13553,N_12945,N_12292);
xnor U13554 (N_13554,N_12249,N_12849);
nor U13555 (N_13555,N_12793,N_12924);
and U13556 (N_13556,N_12714,N_12007);
xor U13557 (N_13557,N_12605,N_12786);
nand U13558 (N_13558,N_12443,N_12587);
nor U13559 (N_13559,N_12666,N_12882);
nor U13560 (N_13560,N_12645,N_12528);
and U13561 (N_13561,N_12086,N_12835);
nand U13562 (N_13562,N_12362,N_12635);
nor U13563 (N_13563,N_12846,N_12037);
xnor U13564 (N_13564,N_12087,N_12674);
and U13565 (N_13565,N_12857,N_12366);
and U13566 (N_13566,N_12110,N_12056);
nand U13567 (N_13567,N_12058,N_12914);
nand U13568 (N_13568,N_12171,N_12706);
or U13569 (N_13569,N_12407,N_12815);
nor U13570 (N_13570,N_12918,N_12406);
and U13571 (N_13571,N_12294,N_12848);
nand U13572 (N_13572,N_12622,N_12800);
nor U13573 (N_13573,N_12161,N_12948);
or U13574 (N_13574,N_12747,N_12936);
nor U13575 (N_13575,N_12074,N_12976);
and U13576 (N_13576,N_12976,N_12736);
nand U13577 (N_13577,N_12983,N_12671);
nor U13578 (N_13578,N_12934,N_12917);
nand U13579 (N_13579,N_12565,N_12651);
or U13580 (N_13580,N_12057,N_12036);
or U13581 (N_13581,N_12867,N_12972);
and U13582 (N_13582,N_12196,N_12937);
nand U13583 (N_13583,N_12498,N_12084);
nor U13584 (N_13584,N_12157,N_12504);
xor U13585 (N_13585,N_12555,N_12393);
xor U13586 (N_13586,N_12650,N_12236);
nor U13587 (N_13587,N_12395,N_12782);
or U13588 (N_13588,N_12729,N_12673);
xor U13589 (N_13589,N_12624,N_12216);
or U13590 (N_13590,N_12474,N_12118);
nand U13591 (N_13591,N_12600,N_12788);
and U13592 (N_13592,N_12027,N_12958);
nand U13593 (N_13593,N_12114,N_12492);
and U13594 (N_13594,N_12221,N_12456);
or U13595 (N_13595,N_12990,N_12937);
nor U13596 (N_13596,N_12954,N_12870);
xnor U13597 (N_13597,N_12815,N_12915);
nand U13598 (N_13598,N_12092,N_12430);
nand U13599 (N_13599,N_12699,N_12132);
nand U13600 (N_13600,N_12112,N_12370);
nand U13601 (N_13601,N_12138,N_12022);
xnor U13602 (N_13602,N_12864,N_12690);
or U13603 (N_13603,N_12012,N_12305);
xnor U13604 (N_13604,N_12373,N_12004);
and U13605 (N_13605,N_12232,N_12086);
and U13606 (N_13606,N_12044,N_12448);
xnor U13607 (N_13607,N_12894,N_12916);
and U13608 (N_13608,N_12937,N_12284);
nor U13609 (N_13609,N_12126,N_12233);
nor U13610 (N_13610,N_12882,N_12581);
and U13611 (N_13611,N_12871,N_12849);
or U13612 (N_13612,N_12607,N_12313);
nand U13613 (N_13613,N_12955,N_12957);
or U13614 (N_13614,N_12858,N_12087);
xor U13615 (N_13615,N_12142,N_12301);
nand U13616 (N_13616,N_12392,N_12705);
or U13617 (N_13617,N_12784,N_12375);
nand U13618 (N_13618,N_12924,N_12084);
xor U13619 (N_13619,N_12243,N_12076);
nand U13620 (N_13620,N_12340,N_12574);
xnor U13621 (N_13621,N_12811,N_12820);
and U13622 (N_13622,N_12044,N_12912);
and U13623 (N_13623,N_12636,N_12656);
or U13624 (N_13624,N_12861,N_12202);
nand U13625 (N_13625,N_12140,N_12696);
xnor U13626 (N_13626,N_12889,N_12488);
nand U13627 (N_13627,N_12189,N_12403);
or U13628 (N_13628,N_12450,N_12188);
or U13629 (N_13629,N_12433,N_12441);
and U13630 (N_13630,N_12451,N_12312);
nand U13631 (N_13631,N_12871,N_12542);
and U13632 (N_13632,N_12508,N_12874);
or U13633 (N_13633,N_12180,N_12979);
xor U13634 (N_13634,N_12651,N_12033);
or U13635 (N_13635,N_12692,N_12707);
xnor U13636 (N_13636,N_12870,N_12381);
nand U13637 (N_13637,N_12119,N_12611);
and U13638 (N_13638,N_12192,N_12056);
nand U13639 (N_13639,N_12063,N_12720);
nand U13640 (N_13640,N_12182,N_12229);
or U13641 (N_13641,N_12007,N_12238);
nor U13642 (N_13642,N_12826,N_12531);
or U13643 (N_13643,N_12896,N_12977);
or U13644 (N_13644,N_12496,N_12907);
and U13645 (N_13645,N_12999,N_12459);
xor U13646 (N_13646,N_12273,N_12492);
xnor U13647 (N_13647,N_12380,N_12747);
nor U13648 (N_13648,N_12197,N_12100);
and U13649 (N_13649,N_12988,N_12002);
and U13650 (N_13650,N_12546,N_12620);
nand U13651 (N_13651,N_12782,N_12026);
xnor U13652 (N_13652,N_12911,N_12797);
xor U13653 (N_13653,N_12367,N_12564);
xnor U13654 (N_13654,N_12463,N_12829);
xor U13655 (N_13655,N_12191,N_12823);
and U13656 (N_13656,N_12420,N_12792);
and U13657 (N_13657,N_12934,N_12371);
and U13658 (N_13658,N_12525,N_12457);
and U13659 (N_13659,N_12169,N_12277);
nand U13660 (N_13660,N_12189,N_12920);
and U13661 (N_13661,N_12179,N_12131);
or U13662 (N_13662,N_12189,N_12022);
and U13663 (N_13663,N_12935,N_12833);
xor U13664 (N_13664,N_12716,N_12414);
xor U13665 (N_13665,N_12480,N_12900);
and U13666 (N_13666,N_12461,N_12692);
xnor U13667 (N_13667,N_12413,N_12485);
nand U13668 (N_13668,N_12012,N_12516);
and U13669 (N_13669,N_12572,N_12246);
nand U13670 (N_13670,N_12477,N_12417);
nand U13671 (N_13671,N_12513,N_12278);
or U13672 (N_13672,N_12975,N_12640);
and U13673 (N_13673,N_12379,N_12555);
nor U13674 (N_13674,N_12380,N_12718);
or U13675 (N_13675,N_12732,N_12740);
and U13676 (N_13676,N_12632,N_12308);
nand U13677 (N_13677,N_12409,N_12120);
and U13678 (N_13678,N_12376,N_12098);
nor U13679 (N_13679,N_12835,N_12190);
or U13680 (N_13680,N_12623,N_12426);
and U13681 (N_13681,N_12384,N_12693);
or U13682 (N_13682,N_12132,N_12162);
and U13683 (N_13683,N_12387,N_12689);
or U13684 (N_13684,N_12964,N_12429);
or U13685 (N_13685,N_12713,N_12028);
or U13686 (N_13686,N_12444,N_12809);
xnor U13687 (N_13687,N_12498,N_12205);
xnor U13688 (N_13688,N_12411,N_12240);
nor U13689 (N_13689,N_12204,N_12906);
nor U13690 (N_13690,N_12279,N_12929);
xnor U13691 (N_13691,N_12446,N_12677);
xor U13692 (N_13692,N_12634,N_12649);
nand U13693 (N_13693,N_12223,N_12678);
xor U13694 (N_13694,N_12029,N_12635);
and U13695 (N_13695,N_12439,N_12548);
nor U13696 (N_13696,N_12949,N_12003);
nor U13697 (N_13697,N_12267,N_12280);
or U13698 (N_13698,N_12755,N_12688);
xor U13699 (N_13699,N_12160,N_12704);
xnor U13700 (N_13700,N_12570,N_12827);
nand U13701 (N_13701,N_12289,N_12190);
and U13702 (N_13702,N_12797,N_12146);
nor U13703 (N_13703,N_12500,N_12520);
nor U13704 (N_13704,N_12544,N_12377);
or U13705 (N_13705,N_12466,N_12438);
or U13706 (N_13706,N_12872,N_12100);
or U13707 (N_13707,N_12785,N_12361);
nand U13708 (N_13708,N_12179,N_12219);
or U13709 (N_13709,N_12434,N_12466);
xor U13710 (N_13710,N_12329,N_12679);
and U13711 (N_13711,N_12522,N_12977);
or U13712 (N_13712,N_12733,N_12565);
xnor U13713 (N_13713,N_12743,N_12077);
or U13714 (N_13714,N_12171,N_12379);
xnor U13715 (N_13715,N_12131,N_12004);
and U13716 (N_13716,N_12797,N_12734);
nand U13717 (N_13717,N_12059,N_12571);
and U13718 (N_13718,N_12554,N_12501);
nor U13719 (N_13719,N_12022,N_12960);
xor U13720 (N_13720,N_12887,N_12827);
or U13721 (N_13721,N_12195,N_12245);
or U13722 (N_13722,N_12213,N_12401);
nor U13723 (N_13723,N_12840,N_12938);
or U13724 (N_13724,N_12174,N_12474);
or U13725 (N_13725,N_12381,N_12519);
and U13726 (N_13726,N_12409,N_12823);
nand U13727 (N_13727,N_12572,N_12501);
nand U13728 (N_13728,N_12350,N_12876);
or U13729 (N_13729,N_12771,N_12858);
and U13730 (N_13730,N_12805,N_12076);
or U13731 (N_13731,N_12628,N_12572);
and U13732 (N_13732,N_12338,N_12483);
xor U13733 (N_13733,N_12206,N_12038);
or U13734 (N_13734,N_12723,N_12046);
and U13735 (N_13735,N_12861,N_12289);
nand U13736 (N_13736,N_12253,N_12363);
nor U13737 (N_13737,N_12933,N_12708);
or U13738 (N_13738,N_12928,N_12631);
nor U13739 (N_13739,N_12047,N_12789);
nor U13740 (N_13740,N_12888,N_12284);
and U13741 (N_13741,N_12949,N_12690);
and U13742 (N_13742,N_12509,N_12911);
and U13743 (N_13743,N_12174,N_12663);
nand U13744 (N_13744,N_12711,N_12736);
and U13745 (N_13745,N_12256,N_12243);
or U13746 (N_13746,N_12950,N_12601);
or U13747 (N_13747,N_12108,N_12613);
nor U13748 (N_13748,N_12827,N_12820);
or U13749 (N_13749,N_12896,N_12850);
or U13750 (N_13750,N_12066,N_12224);
xor U13751 (N_13751,N_12941,N_12362);
nand U13752 (N_13752,N_12880,N_12268);
or U13753 (N_13753,N_12806,N_12228);
and U13754 (N_13754,N_12167,N_12025);
nor U13755 (N_13755,N_12646,N_12983);
and U13756 (N_13756,N_12672,N_12996);
and U13757 (N_13757,N_12721,N_12399);
or U13758 (N_13758,N_12016,N_12453);
nand U13759 (N_13759,N_12004,N_12081);
and U13760 (N_13760,N_12662,N_12289);
xnor U13761 (N_13761,N_12097,N_12822);
nor U13762 (N_13762,N_12276,N_12336);
nand U13763 (N_13763,N_12045,N_12892);
or U13764 (N_13764,N_12082,N_12819);
nor U13765 (N_13765,N_12352,N_12350);
or U13766 (N_13766,N_12925,N_12283);
nor U13767 (N_13767,N_12359,N_12430);
nand U13768 (N_13768,N_12139,N_12736);
xnor U13769 (N_13769,N_12964,N_12998);
nand U13770 (N_13770,N_12668,N_12751);
or U13771 (N_13771,N_12184,N_12199);
nor U13772 (N_13772,N_12125,N_12380);
nor U13773 (N_13773,N_12262,N_12196);
xnor U13774 (N_13774,N_12247,N_12449);
or U13775 (N_13775,N_12755,N_12527);
nor U13776 (N_13776,N_12945,N_12179);
nor U13777 (N_13777,N_12594,N_12746);
and U13778 (N_13778,N_12731,N_12832);
and U13779 (N_13779,N_12978,N_12584);
xor U13780 (N_13780,N_12256,N_12494);
nor U13781 (N_13781,N_12159,N_12756);
or U13782 (N_13782,N_12561,N_12825);
nand U13783 (N_13783,N_12195,N_12941);
or U13784 (N_13784,N_12037,N_12396);
or U13785 (N_13785,N_12512,N_12392);
nor U13786 (N_13786,N_12941,N_12271);
and U13787 (N_13787,N_12470,N_12296);
or U13788 (N_13788,N_12287,N_12733);
xor U13789 (N_13789,N_12581,N_12735);
nand U13790 (N_13790,N_12160,N_12931);
and U13791 (N_13791,N_12364,N_12683);
and U13792 (N_13792,N_12689,N_12475);
and U13793 (N_13793,N_12710,N_12884);
and U13794 (N_13794,N_12859,N_12560);
nand U13795 (N_13795,N_12634,N_12832);
or U13796 (N_13796,N_12817,N_12166);
nor U13797 (N_13797,N_12497,N_12312);
and U13798 (N_13798,N_12186,N_12078);
nor U13799 (N_13799,N_12950,N_12165);
and U13800 (N_13800,N_12584,N_12576);
xor U13801 (N_13801,N_12306,N_12233);
nor U13802 (N_13802,N_12954,N_12004);
nor U13803 (N_13803,N_12604,N_12587);
and U13804 (N_13804,N_12840,N_12581);
xor U13805 (N_13805,N_12606,N_12266);
xor U13806 (N_13806,N_12746,N_12140);
and U13807 (N_13807,N_12690,N_12032);
nand U13808 (N_13808,N_12930,N_12828);
xnor U13809 (N_13809,N_12406,N_12491);
and U13810 (N_13810,N_12729,N_12012);
and U13811 (N_13811,N_12023,N_12905);
xor U13812 (N_13812,N_12977,N_12280);
nor U13813 (N_13813,N_12422,N_12685);
and U13814 (N_13814,N_12542,N_12261);
or U13815 (N_13815,N_12694,N_12498);
or U13816 (N_13816,N_12423,N_12191);
or U13817 (N_13817,N_12526,N_12694);
and U13818 (N_13818,N_12734,N_12352);
xor U13819 (N_13819,N_12453,N_12841);
xnor U13820 (N_13820,N_12735,N_12781);
xnor U13821 (N_13821,N_12375,N_12341);
and U13822 (N_13822,N_12858,N_12249);
nand U13823 (N_13823,N_12974,N_12083);
or U13824 (N_13824,N_12923,N_12944);
and U13825 (N_13825,N_12227,N_12630);
nand U13826 (N_13826,N_12085,N_12193);
xnor U13827 (N_13827,N_12048,N_12403);
and U13828 (N_13828,N_12722,N_12173);
nand U13829 (N_13829,N_12690,N_12511);
nor U13830 (N_13830,N_12995,N_12961);
xnor U13831 (N_13831,N_12747,N_12005);
nand U13832 (N_13832,N_12281,N_12329);
nand U13833 (N_13833,N_12324,N_12198);
or U13834 (N_13834,N_12957,N_12243);
nor U13835 (N_13835,N_12399,N_12162);
and U13836 (N_13836,N_12657,N_12135);
or U13837 (N_13837,N_12565,N_12520);
nand U13838 (N_13838,N_12263,N_12464);
xnor U13839 (N_13839,N_12568,N_12119);
nand U13840 (N_13840,N_12447,N_12878);
nand U13841 (N_13841,N_12008,N_12844);
nand U13842 (N_13842,N_12853,N_12640);
or U13843 (N_13843,N_12430,N_12526);
xnor U13844 (N_13844,N_12254,N_12763);
nor U13845 (N_13845,N_12546,N_12290);
nor U13846 (N_13846,N_12887,N_12405);
xor U13847 (N_13847,N_12093,N_12558);
xor U13848 (N_13848,N_12715,N_12775);
nor U13849 (N_13849,N_12528,N_12631);
nor U13850 (N_13850,N_12665,N_12980);
and U13851 (N_13851,N_12843,N_12110);
nor U13852 (N_13852,N_12867,N_12988);
or U13853 (N_13853,N_12765,N_12220);
and U13854 (N_13854,N_12305,N_12299);
xor U13855 (N_13855,N_12549,N_12440);
nor U13856 (N_13856,N_12207,N_12963);
nor U13857 (N_13857,N_12050,N_12250);
nor U13858 (N_13858,N_12798,N_12984);
nor U13859 (N_13859,N_12289,N_12371);
or U13860 (N_13860,N_12897,N_12379);
and U13861 (N_13861,N_12941,N_12269);
and U13862 (N_13862,N_12869,N_12601);
and U13863 (N_13863,N_12854,N_12770);
nand U13864 (N_13864,N_12965,N_12036);
and U13865 (N_13865,N_12144,N_12967);
nand U13866 (N_13866,N_12371,N_12844);
nand U13867 (N_13867,N_12594,N_12044);
nand U13868 (N_13868,N_12296,N_12152);
nor U13869 (N_13869,N_12540,N_12664);
xor U13870 (N_13870,N_12719,N_12679);
xnor U13871 (N_13871,N_12269,N_12599);
xnor U13872 (N_13872,N_12184,N_12822);
or U13873 (N_13873,N_12370,N_12979);
nand U13874 (N_13874,N_12313,N_12167);
xor U13875 (N_13875,N_12883,N_12358);
nand U13876 (N_13876,N_12764,N_12354);
and U13877 (N_13877,N_12415,N_12594);
and U13878 (N_13878,N_12771,N_12502);
nand U13879 (N_13879,N_12499,N_12157);
nand U13880 (N_13880,N_12841,N_12260);
xor U13881 (N_13881,N_12903,N_12291);
nor U13882 (N_13882,N_12333,N_12382);
xor U13883 (N_13883,N_12964,N_12577);
nand U13884 (N_13884,N_12248,N_12116);
nor U13885 (N_13885,N_12054,N_12455);
and U13886 (N_13886,N_12756,N_12048);
and U13887 (N_13887,N_12688,N_12105);
and U13888 (N_13888,N_12552,N_12610);
xor U13889 (N_13889,N_12635,N_12567);
and U13890 (N_13890,N_12214,N_12933);
or U13891 (N_13891,N_12483,N_12360);
and U13892 (N_13892,N_12564,N_12314);
nor U13893 (N_13893,N_12682,N_12714);
nor U13894 (N_13894,N_12054,N_12557);
nor U13895 (N_13895,N_12875,N_12698);
nor U13896 (N_13896,N_12871,N_12838);
nand U13897 (N_13897,N_12624,N_12981);
xnor U13898 (N_13898,N_12730,N_12406);
xnor U13899 (N_13899,N_12509,N_12902);
nand U13900 (N_13900,N_12503,N_12811);
and U13901 (N_13901,N_12791,N_12797);
xor U13902 (N_13902,N_12150,N_12373);
nand U13903 (N_13903,N_12736,N_12544);
and U13904 (N_13904,N_12553,N_12365);
or U13905 (N_13905,N_12247,N_12252);
nor U13906 (N_13906,N_12862,N_12389);
nor U13907 (N_13907,N_12916,N_12891);
xnor U13908 (N_13908,N_12149,N_12937);
and U13909 (N_13909,N_12660,N_12699);
or U13910 (N_13910,N_12486,N_12037);
xor U13911 (N_13911,N_12846,N_12623);
nand U13912 (N_13912,N_12948,N_12603);
nor U13913 (N_13913,N_12657,N_12875);
and U13914 (N_13914,N_12509,N_12992);
nor U13915 (N_13915,N_12783,N_12028);
nand U13916 (N_13916,N_12399,N_12655);
nor U13917 (N_13917,N_12339,N_12280);
and U13918 (N_13918,N_12803,N_12296);
and U13919 (N_13919,N_12968,N_12028);
and U13920 (N_13920,N_12503,N_12339);
nor U13921 (N_13921,N_12885,N_12267);
nor U13922 (N_13922,N_12133,N_12086);
nand U13923 (N_13923,N_12028,N_12544);
and U13924 (N_13924,N_12466,N_12117);
xor U13925 (N_13925,N_12936,N_12501);
nand U13926 (N_13926,N_12273,N_12910);
nand U13927 (N_13927,N_12255,N_12757);
and U13928 (N_13928,N_12507,N_12545);
or U13929 (N_13929,N_12197,N_12241);
nor U13930 (N_13930,N_12662,N_12445);
or U13931 (N_13931,N_12550,N_12595);
xnor U13932 (N_13932,N_12657,N_12039);
and U13933 (N_13933,N_12042,N_12327);
xor U13934 (N_13934,N_12466,N_12632);
nor U13935 (N_13935,N_12772,N_12580);
and U13936 (N_13936,N_12637,N_12866);
nand U13937 (N_13937,N_12829,N_12489);
nand U13938 (N_13938,N_12823,N_12412);
nand U13939 (N_13939,N_12531,N_12709);
nor U13940 (N_13940,N_12480,N_12765);
nor U13941 (N_13941,N_12897,N_12187);
or U13942 (N_13942,N_12177,N_12449);
and U13943 (N_13943,N_12601,N_12434);
xnor U13944 (N_13944,N_12124,N_12099);
and U13945 (N_13945,N_12138,N_12429);
xnor U13946 (N_13946,N_12786,N_12885);
or U13947 (N_13947,N_12043,N_12024);
or U13948 (N_13948,N_12879,N_12359);
or U13949 (N_13949,N_12128,N_12379);
nor U13950 (N_13950,N_12483,N_12883);
and U13951 (N_13951,N_12669,N_12050);
or U13952 (N_13952,N_12694,N_12341);
xnor U13953 (N_13953,N_12438,N_12083);
and U13954 (N_13954,N_12110,N_12355);
nor U13955 (N_13955,N_12875,N_12109);
nor U13956 (N_13956,N_12507,N_12250);
nor U13957 (N_13957,N_12831,N_12854);
or U13958 (N_13958,N_12740,N_12245);
nand U13959 (N_13959,N_12716,N_12513);
or U13960 (N_13960,N_12678,N_12135);
nand U13961 (N_13961,N_12099,N_12524);
or U13962 (N_13962,N_12113,N_12390);
and U13963 (N_13963,N_12847,N_12269);
nand U13964 (N_13964,N_12179,N_12659);
and U13965 (N_13965,N_12758,N_12321);
xor U13966 (N_13966,N_12290,N_12666);
and U13967 (N_13967,N_12975,N_12999);
or U13968 (N_13968,N_12259,N_12283);
nand U13969 (N_13969,N_12928,N_12067);
or U13970 (N_13970,N_12024,N_12701);
nor U13971 (N_13971,N_12401,N_12803);
nor U13972 (N_13972,N_12892,N_12283);
or U13973 (N_13973,N_12117,N_12311);
and U13974 (N_13974,N_12205,N_12701);
and U13975 (N_13975,N_12291,N_12189);
or U13976 (N_13976,N_12011,N_12536);
nand U13977 (N_13977,N_12641,N_12698);
nand U13978 (N_13978,N_12801,N_12018);
and U13979 (N_13979,N_12503,N_12424);
xor U13980 (N_13980,N_12600,N_12032);
nor U13981 (N_13981,N_12145,N_12380);
and U13982 (N_13982,N_12227,N_12253);
and U13983 (N_13983,N_12183,N_12844);
nor U13984 (N_13984,N_12742,N_12293);
and U13985 (N_13985,N_12590,N_12142);
nand U13986 (N_13986,N_12484,N_12762);
xor U13987 (N_13987,N_12723,N_12089);
xnor U13988 (N_13988,N_12439,N_12486);
and U13989 (N_13989,N_12968,N_12507);
and U13990 (N_13990,N_12446,N_12899);
and U13991 (N_13991,N_12888,N_12578);
nand U13992 (N_13992,N_12024,N_12275);
xor U13993 (N_13993,N_12771,N_12294);
or U13994 (N_13994,N_12377,N_12280);
xor U13995 (N_13995,N_12995,N_12645);
nor U13996 (N_13996,N_12400,N_12084);
or U13997 (N_13997,N_12787,N_12199);
or U13998 (N_13998,N_12565,N_12244);
and U13999 (N_13999,N_12187,N_12538);
nor U14000 (N_14000,N_13024,N_13136);
or U14001 (N_14001,N_13298,N_13500);
and U14002 (N_14002,N_13846,N_13595);
or U14003 (N_14003,N_13008,N_13634);
xnor U14004 (N_14004,N_13711,N_13625);
or U14005 (N_14005,N_13991,N_13566);
nand U14006 (N_14006,N_13454,N_13170);
xnor U14007 (N_14007,N_13231,N_13320);
nand U14008 (N_14008,N_13134,N_13153);
and U14009 (N_14009,N_13203,N_13986);
or U14010 (N_14010,N_13564,N_13234);
nand U14011 (N_14011,N_13310,N_13013);
and U14012 (N_14012,N_13823,N_13764);
nor U14013 (N_14013,N_13061,N_13580);
nor U14014 (N_14014,N_13861,N_13867);
nor U14015 (N_14015,N_13257,N_13720);
nor U14016 (N_14016,N_13446,N_13302);
nand U14017 (N_14017,N_13238,N_13987);
nor U14018 (N_14018,N_13078,N_13596);
and U14019 (N_14019,N_13043,N_13751);
nand U14020 (N_14020,N_13871,N_13841);
xnor U14021 (N_14021,N_13091,N_13392);
xnor U14022 (N_14022,N_13103,N_13311);
or U14023 (N_14023,N_13723,N_13358);
and U14024 (N_14024,N_13090,N_13479);
and U14025 (N_14025,N_13958,N_13968);
nor U14026 (N_14026,N_13156,N_13756);
nand U14027 (N_14027,N_13424,N_13609);
xnor U14028 (N_14028,N_13931,N_13220);
xor U14029 (N_14029,N_13264,N_13330);
and U14030 (N_14030,N_13184,N_13662);
nor U14031 (N_14031,N_13534,N_13222);
and U14032 (N_14032,N_13438,N_13807);
nor U14033 (N_14033,N_13005,N_13747);
and U14034 (N_14034,N_13100,N_13567);
and U14035 (N_14035,N_13197,N_13201);
or U14036 (N_14036,N_13229,N_13526);
and U14037 (N_14037,N_13622,N_13762);
and U14038 (N_14038,N_13389,N_13906);
nor U14039 (N_14039,N_13810,N_13832);
and U14040 (N_14040,N_13189,N_13195);
or U14041 (N_14041,N_13670,N_13521);
or U14042 (N_14042,N_13668,N_13959);
nor U14043 (N_14043,N_13323,N_13243);
nor U14044 (N_14044,N_13887,N_13890);
and U14045 (N_14045,N_13192,N_13929);
nor U14046 (N_14046,N_13822,N_13317);
nand U14047 (N_14047,N_13633,N_13465);
nor U14048 (N_14048,N_13087,N_13441);
and U14049 (N_14049,N_13047,N_13672);
or U14050 (N_14050,N_13088,N_13857);
xnor U14051 (N_14051,N_13737,N_13181);
or U14052 (N_14052,N_13436,N_13554);
or U14053 (N_14053,N_13806,N_13833);
or U14054 (N_14054,N_13313,N_13150);
or U14055 (N_14055,N_13666,N_13419);
or U14056 (N_14056,N_13434,N_13749);
or U14057 (N_14057,N_13387,N_13196);
and U14058 (N_14058,N_13880,N_13485);
and U14059 (N_14059,N_13159,N_13287);
or U14060 (N_14060,N_13054,N_13831);
or U14061 (N_14061,N_13910,N_13135);
nand U14062 (N_14062,N_13004,N_13464);
or U14063 (N_14063,N_13328,N_13585);
xnor U14064 (N_14064,N_13027,N_13506);
nor U14065 (N_14065,N_13350,N_13586);
and U14066 (N_14066,N_13916,N_13025);
or U14067 (N_14067,N_13525,N_13496);
and U14068 (N_14068,N_13045,N_13778);
nand U14069 (N_14069,N_13845,N_13267);
or U14070 (N_14070,N_13453,N_13932);
and U14071 (N_14071,N_13028,N_13112);
xnor U14072 (N_14072,N_13902,N_13707);
and U14073 (N_14073,N_13793,N_13637);
nand U14074 (N_14074,N_13335,N_13759);
nand U14075 (N_14075,N_13117,N_13780);
xor U14076 (N_14076,N_13029,N_13381);
and U14077 (N_14077,N_13509,N_13937);
nor U14078 (N_14078,N_13966,N_13581);
xnor U14079 (N_14079,N_13856,N_13085);
or U14080 (N_14080,N_13621,N_13239);
nor U14081 (N_14081,N_13213,N_13256);
nand U14082 (N_14082,N_13305,N_13770);
and U14083 (N_14083,N_13699,N_13225);
and U14084 (N_14084,N_13133,N_13086);
nor U14085 (N_14085,N_13615,N_13038);
or U14086 (N_14086,N_13131,N_13891);
nand U14087 (N_14087,N_13276,N_13011);
and U14088 (N_14088,N_13002,N_13605);
xor U14089 (N_14089,N_13970,N_13640);
and U14090 (N_14090,N_13370,N_13221);
nor U14091 (N_14091,N_13975,N_13855);
or U14092 (N_14092,N_13836,N_13817);
nor U14093 (N_14093,N_13894,N_13990);
and U14094 (N_14094,N_13097,N_13944);
nand U14095 (N_14095,N_13226,N_13486);
nand U14096 (N_14096,N_13205,N_13934);
nand U14097 (N_14097,N_13563,N_13076);
xor U14098 (N_14098,N_13108,N_13685);
nor U14099 (N_14099,N_13223,N_13623);
xnor U14100 (N_14100,N_13557,N_13726);
xor U14101 (N_14101,N_13800,N_13157);
nor U14102 (N_14102,N_13340,N_13361);
nand U14103 (N_14103,N_13366,N_13251);
nand U14104 (N_14104,N_13187,N_13882);
or U14105 (N_14105,N_13468,N_13332);
xor U14106 (N_14106,N_13068,N_13303);
and U14107 (N_14107,N_13655,N_13368);
or U14108 (N_14108,N_13808,N_13379);
nand U14109 (N_14109,N_13618,N_13113);
nor U14110 (N_14110,N_13235,N_13653);
xor U14111 (N_14111,N_13344,N_13035);
nor U14112 (N_14112,N_13907,N_13612);
or U14113 (N_14113,N_13040,N_13847);
xor U14114 (N_14114,N_13296,N_13953);
or U14115 (N_14115,N_13216,N_13292);
and U14116 (N_14116,N_13401,N_13299);
nand U14117 (N_14117,N_13702,N_13347);
nand U14118 (N_14118,N_13752,N_13760);
or U14119 (N_14119,N_13741,N_13865);
xor U14120 (N_14120,N_13673,N_13104);
nand U14121 (N_14121,N_13917,N_13830);
or U14122 (N_14122,N_13400,N_13481);
nor U14123 (N_14123,N_13694,N_13301);
or U14124 (N_14124,N_13761,N_13771);
xor U14125 (N_14125,N_13367,N_13147);
and U14126 (N_14126,N_13385,N_13407);
nor U14127 (N_14127,N_13674,N_13343);
nand U14128 (N_14128,N_13409,N_13306);
nor U14129 (N_14129,N_13740,N_13642);
nand U14130 (N_14130,N_13565,N_13217);
nand U14131 (N_14131,N_13981,N_13241);
xor U14132 (N_14132,N_13881,N_13448);
xor U14133 (N_14133,N_13530,N_13675);
nor U14134 (N_14134,N_13875,N_13152);
xnor U14135 (N_14135,N_13792,N_13208);
or U14136 (N_14136,N_13173,N_13322);
xor U14137 (N_14137,N_13645,N_13594);
xnor U14138 (N_14138,N_13911,N_13519);
and U14139 (N_14139,N_13177,N_13092);
xnor U14140 (N_14140,N_13592,N_13656);
or U14141 (N_14141,N_13692,N_13919);
or U14142 (N_14142,N_13731,N_13065);
nor U14143 (N_14143,N_13562,N_13456);
or U14144 (N_14144,N_13601,N_13466);
xor U14145 (N_14145,N_13155,N_13491);
nor U14146 (N_14146,N_13098,N_13297);
and U14147 (N_14147,N_13360,N_13651);
or U14148 (N_14148,N_13540,N_13717);
nor U14149 (N_14149,N_13888,N_13433);
and U14150 (N_14150,N_13574,N_13023);
and U14151 (N_14151,N_13275,N_13105);
nand U14152 (N_14152,N_13458,N_13872);
xor U14153 (N_14153,N_13682,N_13815);
or U14154 (N_14154,N_13009,N_13044);
and U14155 (N_14155,N_13034,N_13460);
nand U14156 (N_14156,N_13254,N_13404);
and U14157 (N_14157,N_13643,N_13026);
nor U14158 (N_14158,N_13750,N_13753);
nor U14159 (N_14159,N_13073,N_13200);
or U14160 (N_14160,N_13265,N_13403);
or U14161 (N_14161,N_13449,N_13420);
or U14162 (N_14162,N_13021,N_13654);
or U14163 (N_14163,N_13947,N_13704);
nor U14164 (N_14164,N_13118,N_13743);
xor U14165 (N_14165,N_13001,N_13638);
and U14166 (N_14166,N_13619,N_13825);
and U14167 (N_14167,N_13333,N_13051);
xnor U14168 (N_14168,N_13139,N_13160);
and U14169 (N_14169,N_13459,N_13163);
and U14170 (N_14170,N_13669,N_13397);
and U14171 (N_14171,N_13308,N_13179);
and U14172 (N_14172,N_13019,N_13678);
nand U14173 (N_14173,N_13383,N_13336);
nor U14174 (N_14174,N_13489,N_13188);
nor U14175 (N_14175,N_13236,N_13372);
xnor U14176 (N_14176,N_13998,N_13733);
xnor U14177 (N_14177,N_13979,N_13543);
or U14178 (N_14178,N_13079,N_13356);
xor U14179 (N_14179,N_13194,N_13253);
or U14180 (N_14180,N_13327,N_13329);
nand U14181 (N_14181,N_13735,N_13375);
or U14182 (N_14182,N_13274,N_13337);
or U14183 (N_14183,N_13266,N_13897);
nand U14184 (N_14184,N_13925,N_13262);
and U14185 (N_14185,N_13948,N_13659);
nor U14186 (N_14186,N_13868,N_13785);
nand U14187 (N_14187,N_13537,N_13923);
xor U14188 (N_14188,N_13973,N_13570);
and U14189 (N_14189,N_13539,N_13960);
nand U14190 (N_14190,N_13081,N_13721);
and U14191 (N_14191,N_13757,N_13119);
xor U14192 (N_14192,N_13165,N_13627);
nand U14193 (N_14193,N_13149,N_13282);
and U14194 (N_14194,N_13819,N_13850);
and U14195 (N_14195,N_13763,N_13942);
nand U14196 (N_14196,N_13729,N_13176);
xor U14197 (N_14197,N_13550,N_13121);
or U14198 (N_14198,N_13652,N_13607);
and U14199 (N_14199,N_13950,N_13742);
xnor U14200 (N_14200,N_13736,N_13909);
nor U14201 (N_14201,N_13781,N_13204);
nand U14202 (N_14202,N_13395,N_13072);
nand U14203 (N_14203,N_13983,N_13210);
nor U14204 (N_14204,N_13422,N_13854);
xor U14205 (N_14205,N_13590,N_13148);
nor U14206 (N_14206,N_13237,N_13671);
nand U14207 (N_14207,N_13342,N_13351);
nand U14208 (N_14208,N_13289,N_13561);
and U14209 (N_14209,N_13687,N_13089);
or U14210 (N_14210,N_13202,N_13151);
nand U14211 (N_14211,N_13132,N_13690);
nor U14212 (N_14212,N_13144,N_13374);
and U14213 (N_14213,N_13473,N_13965);
nor U14214 (N_14214,N_13175,N_13697);
nor U14215 (N_14215,N_13031,N_13487);
or U14216 (N_14216,N_13660,N_13876);
nand U14217 (N_14217,N_13745,N_13066);
nand U14218 (N_14218,N_13432,N_13258);
nand U14219 (N_14219,N_13837,N_13576);
nand U14220 (N_14220,N_13193,N_13591);
nand U14221 (N_14221,N_13143,N_13558);
nand U14222 (N_14222,N_13007,N_13405);
nand U14223 (N_14223,N_13614,N_13190);
nor U14224 (N_14224,N_13844,N_13548);
xnor U14225 (N_14225,N_13994,N_13504);
xor U14226 (N_14226,N_13315,N_13616);
and U14227 (N_14227,N_13325,N_13501);
or U14228 (N_14228,N_13610,N_13507);
xnor U14229 (N_14229,N_13014,N_13584);
and U14230 (N_14230,N_13982,N_13138);
and U14231 (N_14231,N_13688,N_13233);
nor U14232 (N_14232,N_13198,N_13748);
and U14233 (N_14233,N_13095,N_13644);
nor U14234 (N_14234,N_13346,N_13706);
nor U14235 (N_14235,N_13712,N_13255);
nor U14236 (N_14236,N_13452,N_13331);
or U14237 (N_14237,N_13630,N_13545);
or U14238 (N_14238,N_13490,N_13495);
nand U14239 (N_14239,N_13814,N_13765);
nor U14240 (N_14240,N_13898,N_13773);
nand U14241 (N_14241,N_13345,N_13939);
and U14242 (N_14242,N_13511,N_13715);
or U14243 (N_14243,N_13058,N_13394);
nand U14244 (N_14244,N_13037,N_13971);
xor U14245 (N_14245,N_13278,N_13956);
nand U14246 (N_14246,N_13538,N_13447);
or U14247 (N_14247,N_13532,N_13709);
or U14248 (N_14248,N_13294,N_13316);
xnor U14249 (N_14249,N_13877,N_13041);
nor U14250 (N_14250,N_13398,N_13547);
xor U14251 (N_14251,N_13862,N_13658);
or U14252 (N_14252,N_13996,N_13722);
and U14253 (N_14253,N_13437,N_13186);
and U14254 (N_14254,N_13377,N_13146);
xor U14255 (N_14255,N_13869,N_13701);
nor U14256 (N_14256,N_13636,N_13813);
nand U14257 (N_14257,N_13474,N_13805);
and U14258 (N_14258,N_13484,N_13922);
nand U14259 (N_14259,N_13866,N_13206);
or U14260 (N_14260,N_13641,N_13246);
nor U14261 (N_14261,N_13006,N_13639);
nor U14262 (N_14262,N_13293,N_13488);
nand U14263 (N_14263,N_13291,N_13502);
xnor U14264 (N_14264,N_13102,N_13363);
nand U14265 (N_14265,N_13228,N_13602);
or U14266 (N_14266,N_13508,N_13099);
or U14267 (N_14267,N_13141,N_13457);
xor U14268 (N_14268,N_13126,N_13801);
nand U14269 (N_14269,N_13626,N_13517);
or U14270 (N_14270,N_13499,N_13069);
nand U14271 (N_14271,N_13914,N_13578);
and U14272 (N_14272,N_13926,N_13732);
and U14273 (N_14273,N_13124,N_13107);
xor U14274 (N_14274,N_13480,N_13211);
nor U14275 (N_14275,N_13110,N_13199);
and U14276 (N_14276,N_13492,N_13154);
nand U14277 (N_14277,N_13999,N_13111);
or U14278 (N_14278,N_13541,N_13811);
and U14279 (N_14279,N_13598,N_13840);
and U14280 (N_14280,N_13946,N_13046);
xor U14281 (N_14281,N_13518,N_13874);
nor U14282 (N_14282,N_13744,N_13560);
or U14283 (N_14283,N_13787,N_13522);
nand U14284 (N_14284,N_13443,N_13664);
xnor U14285 (N_14285,N_13018,N_13657);
xnor U14286 (N_14286,N_13349,N_13588);
xor U14287 (N_14287,N_13758,N_13467);
and U14288 (N_14288,N_13738,N_13632);
nor U14289 (N_14289,N_13573,N_13290);
nand U14290 (N_14290,N_13476,N_13984);
nand U14291 (N_14291,N_13421,N_13362);
nor U14292 (N_14292,N_13774,N_13804);
xnor U14293 (N_14293,N_13597,N_13191);
nor U14294 (N_14294,N_13042,N_13020);
and U14295 (N_14295,N_13772,N_13714);
nor U14296 (N_14296,N_13365,N_13988);
nor U14297 (N_14297,N_13312,N_13075);
and U14298 (N_14298,N_13661,N_13679);
xnor U14299 (N_14299,N_13798,N_13551);
xnor U14300 (N_14300,N_13512,N_13995);
and U14301 (N_14301,N_13039,N_13497);
nor U14302 (N_14302,N_13912,N_13728);
and U14303 (N_14303,N_13273,N_13430);
xnor U14304 (N_14304,N_13413,N_13915);
and U14305 (N_14305,N_13777,N_13553);
or U14306 (N_14306,N_13171,N_13782);
or U14307 (N_14307,N_13992,N_13408);
nor U14308 (N_14308,N_13314,N_13535);
nand U14309 (N_14309,N_13015,N_13396);
nor U14310 (N_14310,N_13884,N_13427);
or U14311 (N_14311,N_13858,N_13938);
xnor U14312 (N_14312,N_13477,N_13769);
nand U14313 (N_14313,N_13895,N_13247);
xnor U14314 (N_14314,N_13883,N_13224);
or U14315 (N_14315,N_13482,N_13663);
nand U14316 (N_14316,N_13790,N_13440);
or U14317 (N_14317,N_13429,N_13724);
xnor U14318 (N_14318,N_13901,N_13283);
nor U14319 (N_14319,N_13978,N_13423);
and U14320 (N_14320,N_13326,N_13277);
and U14321 (N_14321,N_13167,N_13261);
nand U14322 (N_14322,N_13727,N_13084);
nor U14323 (N_14323,N_13339,N_13941);
or U14324 (N_14324,N_13710,N_13353);
nand U14325 (N_14325,N_13794,N_13628);
xnor U14326 (N_14326,N_13617,N_13680);
and U14327 (N_14327,N_13120,N_13166);
xor U14328 (N_14328,N_13129,N_13271);
or U14329 (N_14329,N_13713,N_13583);
nor U14330 (N_14330,N_13493,N_13544);
nand U14331 (N_14331,N_13571,N_13376);
nand U14332 (N_14332,N_13402,N_13913);
or U14333 (N_14333,N_13060,N_13052);
nor U14334 (N_14334,N_13848,N_13796);
and U14335 (N_14335,N_13268,N_13359);
and U14336 (N_14336,N_13527,N_13520);
or U14337 (N_14337,N_13354,N_13603);
xor U14338 (N_14338,N_13700,N_13852);
nor U14339 (N_14339,N_13215,N_13516);
nor U14340 (N_14340,N_13838,N_13803);
xnor U14341 (N_14341,N_13444,N_13693);
or U14342 (N_14342,N_13115,N_13304);
nand U14343 (N_14343,N_13083,N_13599);
and U14344 (N_14344,N_13260,N_13892);
and U14345 (N_14345,N_13263,N_13945);
and U14346 (N_14346,N_13786,N_13927);
nor U14347 (N_14347,N_13049,N_13352);
and U14348 (N_14348,N_13093,N_13012);
nand U14349 (N_14349,N_13435,N_13835);
and U14350 (N_14350,N_13373,N_13940);
nand U14351 (N_14351,N_13684,N_13218);
or U14352 (N_14352,N_13364,N_13016);
nor U14353 (N_14353,N_13579,N_13463);
or U14354 (N_14354,N_13439,N_13033);
xor U14355 (N_14355,N_13022,N_13647);
nor U14356 (N_14356,N_13784,N_13300);
xnor U14357 (N_14357,N_13936,N_13935);
and U14358 (N_14358,N_13905,N_13426);
nand U14359 (N_14359,N_13168,N_13380);
xnor U14360 (N_14360,N_13878,N_13559);
or U14361 (N_14361,N_13677,N_13829);
nand U14362 (N_14362,N_13067,N_13318);
or U14363 (N_14363,N_13050,N_13789);
nor U14364 (N_14364,N_13431,N_13207);
nand U14365 (N_14365,N_13142,N_13248);
or U14366 (N_14366,N_13860,N_13334);
or U14367 (N_14367,N_13414,N_13130);
nand U14368 (N_14368,N_13886,N_13106);
and U14369 (N_14369,N_13783,N_13478);
nor U14370 (N_14370,N_13161,N_13498);
and U14371 (N_14371,N_13471,N_13080);
and U14372 (N_14372,N_13272,N_13140);
xnor U14373 (N_14373,N_13980,N_13445);
nand U14374 (N_14374,N_13624,N_13734);
nor U14375 (N_14375,N_13900,N_13003);
nor U14376 (N_14376,N_13920,N_13828);
and U14377 (N_14377,N_13952,N_13809);
and U14378 (N_14378,N_13219,N_13169);
xor U14379 (N_14379,N_13415,N_13698);
xnor U14380 (N_14380,N_13820,N_13776);
or U14381 (N_14381,N_13589,N_13338);
nor U14382 (N_14382,N_13577,N_13017);
nor U14383 (N_14383,N_13470,N_13321);
or U14384 (N_14384,N_13077,N_13649);
or U14385 (N_14385,N_13683,N_13635);
or U14386 (N_14386,N_13214,N_13851);
nand U14387 (N_14387,N_13137,N_13826);
or U14388 (N_14388,N_13555,N_13716);
nor U14389 (N_14389,N_13949,N_13357);
xor U14390 (N_14390,N_13178,N_13839);
and U14391 (N_14391,N_13842,N_13057);
or U14392 (N_14392,N_13324,N_13469);
xor U14393 (N_14393,N_13442,N_13245);
and U14394 (N_14394,N_13125,N_13410);
and U14395 (N_14395,N_13053,N_13288);
nor U14396 (N_14396,N_13962,N_13921);
nor U14397 (N_14397,N_13284,N_13523);
xnor U14398 (N_14398,N_13494,N_13483);
or U14399 (N_14399,N_13094,N_13587);
and U14400 (N_14400,N_13873,N_13388);
xor U14401 (N_14401,N_13209,N_13812);
nor U14402 (N_14402,N_13821,N_13754);
and U14403 (N_14403,N_13230,N_13843);
nor U14404 (N_14404,N_13768,N_13341);
or U14405 (N_14405,N_13182,N_13977);
nor U14406 (N_14406,N_13064,N_13957);
and U14407 (N_14407,N_13172,N_13425);
or U14408 (N_14408,N_13696,N_13604);
xor U14409 (N_14409,N_13461,N_13739);
nor U14410 (N_14410,N_13390,N_13667);
or U14411 (N_14411,N_13533,N_13549);
nor U14412 (N_14412,N_13412,N_13648);
and U14413 (N_14413,N_13164,N_13386);
nor U14414 (N_14414,N_13063,N_13885);
nor U14415 (N_14415,N_13295,N_13791);
nand U14416 (N_14416,N_13930,N_13528);
or U14417 (N_14417,N_13062,N_13145);
and U14418 (N_14418,N_13967,N_13279);
or U14419 (N_14419,N_13122,N_13568);
or U14420 (N_14420,N_13070,N_13719);
or U14421 (N_14421,N_13455,N_13055);
nand U14422 (N_14422,N_13893,N_13391);
and U14423 (N_14423,N_13746,N_13378);
xnor U14424 (N_14424,N_13162,N_13393);
and U14425 (N_14425,N_13505,N_13795);
or U14426 (N_14426,N_13000,N_13799);
nor U14427 (N_14427,N_13542,N_13127);
and U14428 (N_14428,N_13082,N_13827);
nor U14429 (N_14429,N_13879,N_13280);
nand U14430 (N_14430,N_13056,N_13689);
xnor U14431 (N_14431,N_13240,N_13174);
or U14432 (N_14432,N_13569,N_13406);
or U14433 (N_14433,N_13955,N_13766);
and U14434 (N_14434,N_13416,N_13514);
nand U14435 (N_14435,N_13114,N_13059);
and U14436 (N_14436,N_13116,N_13032);
nand U14437 (N_14437,N_13676,N_13963);
or U14438 (N_14438,N_13646,N_13109);
and U14439 (N_14439,N_13227,N_13681);
nor U14440 (N_14440,N_13384,N_13524);
xnor U14441 (N_14441,N_13101,N_13924);
nor U14442 (N_14442,N_13954,N_13834);
xor U14443 (N_14443,N_13259,N_13918);
xnor U14444 (N_14444,N_13158,N_13185);
and U14445 (N_14445,N_13472,N_13348);
nand U14446 (N_14446,N_13575,N_13411);
or U14447 (N_14447,N_13036,N_13515);
and U14448 (N_14448,N_13613,N_13450);
xnor U14449 (N_14449,N_13418,N_13943);
nand U14450 (N_14450,N_13546,N_13629);
and U14451 (N_14451,N_13128,N_13428);
or U14452 (N_14452,N_13903,N_13725);
nand U14453 (N_14453,N_13307,N_13933);
xor U14454 (N_14454,N_13928,N_13849);
and U14455 (N_14455,N_13475,N_13969);
and U14456 (N_14456,N_13775,N_13285);
nor U14457 (N_14457,N_13048,N_13961);
xor U14458 (N_14458,N_13212,N_13870);
or U14459 (N_14459,N_13985,N_13997);
xnor U14460 (N_14460,N_13853,N_13816);
nand U14461 (N_14461,N_13964,N_13382);
and U14462 (N_14462,N_13863,N_13703);
or U14463 (N_14463,N_13270,N_13989);
nor U14464 (N_14464,N_13510,N_13650);
xnor U14465 (N_14465,N_13572,N_13993);
nor U14466 (N_14466,N_13797,N_13531);
nand U14467 (N_14467,N_13755,N_13889);
xnor U14468 (N_14468,N_13695,N_13859);
nand U14469 (N_14469,N_13582,N_13974);
nor U14470 (N_14470,N_13552,N_13123);
and U14471 (N_14471,N_13269,N_13818);
xnor U14472 (N_14472,N_13250,N_13691);
nor U14473 (N_14473,N_13686,N_13462);
nor U14474 (N_14474,N_13232,N_13071);
nand U14475 (N_14475,N_13665,N_13183);
nor U14476 (N_14476,N_13824,N_13399);
nand U14477 (N_14477,N_13730,N_13536);
xnor U14478 (N_14478,N_13503,N_13556);
nor U14479 (N_14479,N_13451,N_13319);
nand U14480 (N_14480,N_13767,N_13600);
and U14481 (N_14481,N_13631,N_13779);
nor U14482 (N_14482,N_13802,N_13608);
and U14483 (N_14483,N_13864,N_13529);
nand U14484 (N_14484,N_13951,N_13242);
or U14485 (N_14485,N_13369,N_13611);
nand U14486 (N_14486,N_13252,N_13074);
nand U14487 (N_14487,N_13371,N_13606);
nor U14488 (N_14488,N_13096,N_13593);
xnor U14489 (N_14489,N_13899,N_13620);
nand U14490 (N_14490,N_13896,N_13718);
or U14491 (N_14491,N_13513,N_13972);
nand U14492 (N_14492,N_13417,N_13708);
xnor U14493 (N_14493,N_13976,N_13010);
nor U14494 (N_14494,N_13309,N_13705);
nand U14495 (N_14495,N_13244,N_13908);
nor U14496 (N_14496,N_13180,N_13904);
and U14497 (N_14497,N_13355,N_13281);
and U14498 (N_14498,N_13030,N_13286);
and U14499 (N_14499,N_13788,N_13249);
and U14500 (N_14500,N_13902,N_13771);
or U14501 (N_14501,N_13153,N_13729);
and U14502 (N_14502,N_13264,N_13738);
nand U14503 (N_14503,N_13543,N_13064);
xor U14504 (N_14504,N_13141,N_13719);
nor U14505 (N_14505,N_13924,N_13847);
and U14506 (N_14506,N_13167,N_13722);
or U14507 (N_14507,N_13407,N_13696);
xnor U14508 (N_14508,N_13510,N_13124);
and U14509 (N_14509,N_13095,N_13298);
xnor U14510 (N_14510,N_13050,N_13348);
nor U14511 (N_14511,N_13411,N_13443);
nor U14512 (N_14512,N_13933,N_13236);
nor U14513 (N_14513,N_13147,N_13810);
and U14514 (N_14514,N_13849,N_13635);
nand U14515 (N_14515,N_13048,N_13749);
and U14516 (N_14516,N_13431,N_13448);
nand U14517 (N_14517,N_13684,N_13777);
or U14518 (N_14518,N_13080,N_13348);
or U14519 (N_14519,N_13871,N_13445);
xnor U14520 (N_14520,N_13978,N_13557);
nor U14521 (N_14521,N_13343,N_13167);
and U14522 (N_14522,N_13885,N_13345);
nor U14523 (N_14523,N_13577,N_13663);
or U14524 (N_14524,N_13485,N_13851);
nor U14525 (N_14525,N_13435,N_13069);
xnor U14526 (N_14526,N_13092,N_13482);
or U14527 (N_14527,N_13587,N_13837);
nand U14528 (N_14528,N_13560,N_13660);
and U14529 (N_14529,N_13220,N_13606);
and U14530 (N_14530,N_13466,N_13341);
xor U14531 (N_14531,N_13484,N_13514);
or U14532 (N_14532,N_13402,N_13309);
nor U14533 (N_14533,N_13356,N_13404);
and U14534 (N_14534,N_13112,N_13327);
xnor U14535 (N_14535,N_13463,N_13291);
and U14536 (N_14536,N_13868,N_13264);
xnor U14537 (N_14537,N_13250,N_13922);
xor U14538 (N_14538,N_13436,N_13874);
xor U14539 (N_14539,N_13643,N_13970);
or U14540 (N_14540,N_13417,N_13820);
or U14541 (N_14541,N_13578,N_13497);
nor U14542 (N_14542,N_13427,N_13855);
nand U14543 (N_14543,N_13952,N_13063);
nor U14544 (N_14544,N_13361,N_13518);
nor U14545 (N_14545,N_13709,N_13761);
nand U14546 (N_14546,N_13908,N_13874);
and U14547 (N_14547,N_13487,N_13993);
and U14548 (N_14548,N_13033,N_13399);
or U14549 (N_14549,N_13066,N_13736);
xor U14550 (N_14550,N_13126,N_13259);
and U14551 (N_14551,N_13786,N_13917);
nor U14552 (N_14552,N_13854,N_13701);
or U14553 (N_14553,N_13775,N_13338);
nand U14554 (N_14554,N_13076,N_13021);
xor U14555 (N_14555,N_13323,N_13422);
or U14556 (N_14556,N_13051,N_13887);
nand U14557 (N_14557,N_13625,N_13966);
nor U14558 (N_14558,N_13327,N_13903);
and U14559 (N_14559,N_13032,N_13706);
and U14560 (N_14560,N_13033,N_13250);
nor U14561 (N_14561,N_13492,N_13727);
xnor U14562 (N_14562,N_13273,N_13554);
nor U14563 (N_14563,N_13583,N_13128);
and U14564 (N_14564,N_13708,N_13059);
xor U14565 (N_14565,N_13227,N_13056);
and U14566 (N_14566,N_13024,N_13962);
xor U14567 (N_14567,N_13209,N_13656);
nor U14568 (N_14568,N_13692,N_13111);
or U14569 (N_14569,N_13336,N_13785);
and U14570 (N_14570,N_13296,N_13016);
nand U14571 (N_14571,N_13392,N_13306);
or U14572 (N_14572,N_13416,N_13989);
xor U14573 (N_14573,N_13360,N_13314);
nand U14574 (N_14574,N_13370,N_13169);
and U14575 (N_14575,N_13142,N_13323);
and U14576 (N_14576,N_13873,N_13505);
or U14577 (N_14577,N_13534,N_13296);
xnor U14578 (N_14578,N_13993,N_13025);
nand U14579 (N_14579,N_13217,N_13591);
or U14580 (N_14580,N_13118,N_13141);
or U14581 (N_14581,N_13503,N_13801);
nor U14582 (N_14582,N_13134,N_13532);
nand U14583 (N_14583,N_13717,N_13570);
or U14584 (N_14584,N_13799,N_13815);
nand U14585 (N_14585,N_13770,N_13599);
and U14586 (N_14586,N_13171,N_13836);
or U14587 (N_14587,N_13110,N_13604);
or U14588 (N_14588,N_13942,N_13677);
nand U14589 (N_14589,N_13630,N_13911);
nor U14590 (N_14590,N_13601,N_13854);
nor U14591 (N_14591,N_13206,N_13941);
or U14592 (N_14592,N_13633,N_13293);
and U14593 (N_14593,N_13234,N_13175);
or U14594 (N_14594,N_13892,N_13803);
or U14595 (N_14595,N_13053,N_13163);
nor U14596 (N_14596,N_13890,N_13028);
nor U14597 (N_14597,N_13235,N_13759);
nand U14598 (N_14598,N_13454,N_13615);
and U14599 (N_14599,N_13695,N_13036);
or U14600 (N_14600,N_13660,N_13782);
xor U14601 (N_14601,N_13263,N_13220);
and U14602 (N_14602,N_13855,N_13251);
or U14603 (N_14603,N_13201,N_13934);
nor U14604 (N_14604,N_13877,N_13551);
or U14605 (N_14605,N_13737,N_13344);
and U14606 (N_14606,N_13255,N_13821);
xnor U14607 (N_14607,N_13940,N_13643);
nand U14608 (N_14608,N_13152,N_13198);
and U14609 (N_14609,N_13647,N_13050);
xor U14610 (N_14610,N_13649,N_13901);
or U14611 (N_14611,N_13605,N_13550);
or U14612 (N_14612,N_13048,N_13920);
and U14613 (N_14613,N_13515,N_13060);
nand U14614 (N_14614,N_13536,N_13981);
xnor U14615 (N_14615,N_13957,N_13019);
nand U14616 (N_14616,N_13252,N_13183);
xor U14617 (N_14617,N_13303,N_13204);
nor U14618 (N_14618,N_13629,N_13683);
and U14619 (N_14619,N_13385,N_13017);
or U14620 (N_14620,N_13282,N_13917);
xnor U14621 (N_14621,N_13769,N_13910);
xor U14622 (N_14622,N_13949,N_13324);
or U14623 (N_14623,N_13047,N_13172);
and U14624 (N_14624,N_13702,N_13353);
and U14625 (N_14625,N_13787,N_13680);
and U14626 (N_14626,N_13607,N_13004);
or U14627 (N_14627,N_13401,N_13208);
and U14628 (N_14628,N_13713,N_13166);
nand U14629 (N_14629,N_13745,N_13573);
nor U14630 (N_14630,N_13760,N_13157);
xor U14631 (N_14631,N_13917,N_13284);
or U14632 (N_14632,N_13827,N_13968);
nor U14633 (N_14633,N_13625,N_13898);
or U14634 (N_14634,N_13088,N_13453);
or U14635 (N_14635,N_13733,N_13671);
nand U14636 (N_14636,N_13631,N_13282);
nand U14637 (N_14637,N_13119,N_13649);
nor U14638 (N_14638,N_13501,N_13664);
nand U14639 (N_14639,N_13385,N_13313);
xor U14640 (N_14640,N_13070,N_13914);
xnor U14641 (N_14641,N_13365,N_13843);
nand U14642 (N_14642,N_13765,N_13918);
nand U14643 (N_14643,N_13006,N_13770);
or U14644 (N_14644,N_13700,N_13448);
and U14645 (N_14645,N_13917,N_13870);
nor U14646 (N_14646,N_13132,N_13214);
nor U14647 (N_14647,N_13001,N_13678);
or U14648 (N_14648,N_13269,N_13404);
nor U14649 (N_14649,N_13732,N_13416);
nand U14650 (N_14650,N_13423,N_13804);
or U14651 (N_14651,N_13299,N_13008);
nand U14652 (N_14652,N_13162,N_13546);
nor U14653 (N_14653,N_13328,N_13558);
nor U14654 (N_14654,N_13790,N_13794);
nor U14655 (N_14655,N_13481,N_13854);
or U14656 (N_14656,N_13745,N_13194);
or U14657 (N_14657,N_13097,N_13764);
xnor U14658 (N_14658,N_13486,N_13468);
nand U14659 (N_14659,N_13463,N_13263);
or U14660 (N_14660,N_13032,N_13494);
and U14661 (N_14661,N_13142,N_13847);
or U14662 (N_14662,N_13478,N_13179);
xnor U14663 (N_14663,N_13951,N_13421);
or U14664 (N_14664,N_13020,N_13931);
xor U14665 (N_14665,N_13461,N_13407);
and U14666 (N_14666,N_13296,N_13102);
xor U14667 (N_14667,N_13744,N_13584);
and U14668 (N_14668,N_13242,N_13800);
and U14669 (N_14669,N_13293,N_13330);
nand U14670 (N_14670,N_13607,N_13716);
nand U14671 (N_14671,N_13933,N_13848);
or U14672 (N_14672,N_13813,N_13756);
and U14673 (N_14673,N_13384,N_13082);
nor U14674 (N_14674,N_13482,N_13735);
or U14675 (N_14675,N_13432,N_13680);
xnor U14676 (N_14676,N_13286,N_13242);
xnor U14677 (N_14677,N_13927,N_13964);
and U14678 (N_14678,N_13607,N_13149);
and U14679 (N_14679,N_13262,N_13797);
xnor U14680 (N_14680,N_13818,N_13391);
xor U14681 (N_14681,N_13646,N_13948);
nor U14682 (N_14682,N_13102,N_13981);
nor U14683 (N_14683,N_13344,N_13841);
and U14684 (N_14684,N_13844,N_13979);
nand U14685 (N_14685,N_13169,N_13588);
or U14686 (N_14686,N_13501,N_13960);
nand U14687 (N_14687,N_13443,N_13104);
and U14688 (N_14688,N_13860,N_13385);
and U14689 (N_14689,N_13784,N_13499);
or U14690 (N_14690,N_13846,N_13868);
nor U14691 (N_14691,N_13044,N_13718);
nand U14692 (N_14692,N_13004,N_13468);
nand U14693 (N_14693,N_13986,N_13829);
and U14694 (N_14694,N_13441,N_13543);
or U14695 (N_14695,N_13623,N_13684);
nand U14696 (N_14696,N_13405,N_13212);
xnor U14697 (N_14697,N_13043,N_13056);
and U14698 (N_14698,N_13603,N_13053);
and U14699 (N_14699,N_13589,N_13056);
or U14700 (N_14700,N_13091,N_13291);
or U14701 (N_14701,N_13878,N_13055);
or U14702 (N_14702,N_13006,N_13502);
nor U14703 (N_14703,N_13967,N_13618);
and U14704 (N_14704,N_13473,N_13133);
xnor U14705 (N_14705,N_13121,N_13984);
xor U14706 (N_14706,N_13786,N_13402);
nor U14707 (N_14707,N_13024,N_13618);
or U14708 (N_14708,N_13727,N_13574);
xnor U14709 (N_14709,N_13353,N_13751);
nor U14710 (N_14710,N_13034,N_13326);
nor U14711 (N_14711,N_13093,N_13363);
or U14712 (N_14712,N_13622,N_13890);
xor U14713 (N_14713,N_13980,N_13854);
nor U14714 (N_14714,N_13038,N_13026);
and U14715 (N_14715,N_13227,N_13087);
nor U14716 (N_14716,N_13303,N_13893);
nor U14717 (N_14717,N_13389,N_13913);
xor U14718 (N_14718,N_13524,N_13986);
nor U14719 (N_14719,N_13304,N_13009);
and U14720 (N_14720,N_13147,N_13006);
nor U14721 (N_14721,N_13526,N_13345);
nor U14722 (N_14722,N_13819,N_13444);
and U14723 (N_14723,N_13117,N_13792);
nand U14724 (N_14724,N_13779,N_13005);
and U14725 (N_14725,N_13951,N_13211);
or U14726 (N_14726,N_13698,N_13212);
nand U14727 (N_14727,N_13880,N_13707);
or U14728 (N_14728,N_13263,N_13843);
nand U14729 (N_14729,N_13590,N_13233);
nand U14730 (N_14730,N_13004,N_13475);
nor U14731 (N_14731,N_13289,N_13929);
nand U14732 (N_14732,N_13106,N_13202);
nand U14733 (N_14733,N_13708,N_13996);
or U14734 (N_14734,N_13981,N_13967);
and U14735 (N_14735,N_13886,N_13311);
nor U14736 (N_14736,N_13094,N_13979);
nand U14737 (N_14737,N_13251,N_13588);
xor U14738 (N_14738,N_13975,N_13670);
and U14739 (N_14739,N_13771,N_13603);
and U14740 (N_14740,N_13178,N_13270);
xnor U14741 (N_14741,N_13773,N_13887);
or U14742 (N_14742,N_13635,N_13620);
and U14743 (N_14743,N_13681,N_13980);
and U14744 (N_14744,N_13947,N_13564);
and U14745 (N_14745,N_13357,N_13728);
and U14746 (N_14746,N_13009,N_13337);
and U14747 (N_14747,N_13359,N_13074);
and U14748 (N_14748,N_13889,N_13385);
and U14749 (N_14749,N_13005,N_13920);
xor U14750 (N_14750,N_13101,N_13457);
nor U14751 (N_14751,N_13661,N_13824);
and U14752 (N_14752,N_13061,N_13415);
nor U14753 (N_14753,N_13960,N_13145);
or U14754 (N_14754,N_13622,N_13111);
or U14755 (N_14755,N_13268,N_13394);
xnor U14756 (N_14756,N_13129,N_13815);
xor U14757 (N_14757,N_13134,N_13641);
nor U14758 (N_14758,N_13684,N_13388);
nor U14759 (N_14759,N_13398,N_13773);
nand U14760 (N_14760,N_13007,N_13186);
nand U14761 (N_14761,N_13525,N_13004);
and U14762 (N_14762,N_13490,N_13675);
nor U14763 (N_14763,N_13515,N_13907);
nor U14764 (N_14764,N_13225,N_13437);
nand U14765 (N_14765,N_13762,N_13367);
or U14766 (N_14766,N_13197,N_13570);
nor U14767 (N_14767,N_13075,N_13563);
or U14768 (N_14768,N_13140,N_13835);
nor U14769 (N_14769,N_13163,N_13927);
xnor U14770 (N_14770,N_13864,N_13527);
nand U14771 (N_14771,N_13347,N_13740);
or U14772 (N_14772,N_13315,N_13204);
or U14773 (N_14773,N_13370,N_13760);
nand U14774 (N_14774,N_13656,N_13776);
xor U14775 (N_14775,N_13939,N_13338);
or U14776 (N_14776,N_13697,N_13107);
nand U14777 (N_14777,N_13341,N_13110);
xnor U14778 (N_14778,N_13367,N_13012);
xor U14779 (N_14779,N_13259,N_13606);
or U14780 (N_14780,N_13048,N_13146);
and U14781 (N_14781,N_13628,N_13927);
nor U14782 (N_14782,N_13607,N_13166);
xor U14783 (N_14783,N_13897,N_13039);
or U14784 (N_14784,N_13937,N_13964);
or U14785 (N_14785,N_13076,N_13705);
or U14786 (N_14786,N_13760,N_13081);
or U14787 (N_14787,N_13618,N_13268);
nand U14788 (N_14788,N_13257,N_13816);
or U14789 (N_14789,N_13548,N_13445);
xor U14790 (N_14790,N_13076,N_13507);
xnor U14791 (N_14791,N_13634,N_13976);
and U14792 (N_14792,N_13255,N_13494);
or U14793 (N_14793,N_13620,N_13607);
or U14794 (N_14794,N_13758,N_13683);
nand U14795 (N_14795,N_13041,N_13973);
or U14796 (N_14796,N_13705,N_13103);
xor U14797 (N_14797,N_13245,N_13342);
or U14798 (N_14798,N_13444,N_13682);
or U14799 (N_14799,N_13887,N_13077);
nor U14800 (N_14800,N_13681,N_13120);
or U14801 (N_14801,N_13752,N_13140);
xor U14802 (N_14802,N_13703,N_13443);
xnor U14803 (N_14803,N_13468,N_13983);
nor U14804 (N_14804,N_13831,N_13228);
and U14805 (N_14805,N_13741,N_13807);
or U14806 (N_14806,N_13666,N_13143);
xor U14807 (N_14807,N_13032,N_13487);
xnor U14808 (N_14808,N_13148,N_13283);
nor U14809 (N_14809,N_13075,N_13283);
xor U14810 (N_14810,N_13803,N_13257);
xnor U14811 (N_14811,N_13688,N_13782);
or U14812 (N_14812,N_13694,N_13532);
and U14813 (N_14813,N_13991,N_13358);
xor U14814 (N_14814,N_13745,N_13455);
xnor U14815 (N_14815,N_13121,N_13129);
or U14816 (N_14816,N_13739,N_13217);
or U14817 (N_14817,N_13918,N_13847);
or U14818 (N_14818,N_13001,N_13761);
xnor U14819 (N_14819,N_13665,N_13605);
and U14820 (N_14820,N_13664,N_13709);
or U14821 (N_14821,N_13777,N_13143);
nor U14822 (N_14822,N_13511,N_13609);
nand U14823 (N_14823,N_13703,N_13893);
xnor U14824 (N_14824,N_13808,N_13435);
and U14825 (N_14825,N_13024,N_13315);
nand U14826 (N_14826,N_13504,N_13820);
and U14827 (N_14827,N_13874,N_13894);
nor U14828 (N_14828,N_13097,N_13665);
and U14829 (N_14829,N_13755,N_13395);
and U14830 (N_14830,N_13447,N_13816);
and U14831 (N_14831,N_13573,N_13177);
xor U14832 (N_14832,N_13832,N_13879);
nand U14833 (N_14833,N_13873,N_13243);
nand U14834 (N_14834,N_13941,N_13647);
and U14835 (N_14835,N_13026,N_13448);
or U14836 (N_14836,N_13240,N_13108);
and U14837 (N_14837,N_13672,N_13805);
nand U14838 (N_14838,N_13933,N_13991);
or U14839 (N_14839,N_13915,N_13559);
or U14840 (N_14840,N_13886,N_13676);
nand U14841 (N_14841,N_13036,N_13576);
nand U14842 (N_14842,N_13803,N_13827);
xor U14843 (N_14843,N_13120,N_13997);
and U14844 (N_14844,N_13010,N_13059);
xnor U14845 (N_14845,N_13849,N_13643);
and U14846 (N_14846,N_13879,N_13710);
nand U14847 (N_14847,N_13267,N_13637);
nand U14848 (N_14848,N_13745,N_13324);
nor U14849 (N_14849,N_13852,N_13548);
xnor U14850 (N_14850,N_13115,N_13870);
and U14851 (N_14851,N_13671,N_13341);
and U14852 (N_14852,N_13671,N_13594);
nor U14853 (N_14853,N_13728,N_13914);
nand U14854 (N_14854,N_13055,N_13931);
or U14855 (N_14855,N_13374,N_13525);
nand U14856 (N_14856,N_13876,N_13931);
nor U14857 (N_14857,N_13358,N_13666);
nor U14858 (N_14858,N_13363,N_13995);
xnor U14859 (N_14859,N_13811,N_13489);
and U14860 (N_14860,N_13404,N_13616);
xnor U14861 (N_14861,N_13799,N_13617);
and U14862 (N_14862,N_13928,N_13329);
nand U14863 (N_14863,N_13008,N_13219);
nand U14864 (N_14864,N_13026,N_13634);
and U14865 (N_14865,N_13792,N_13342);
or U14866 (N_14866,N_13146,N_13233);
and U14867 (N_14867,N_13695,N_13170);
and U14868 (N_14868,N_13384,N_13260);
or U14869 (N_14869,N_13009,N_13467);
nand U14870 (N_14870,N_13611,N_13799);
and U14871 (N_14871,N_13267,N_13471);
nand U14872 (N_14872,N_13642,N_13341);
and U14873 (N_14873,N_13287,N_13466);
or U14874 (N_14874,N_13386,N_13481);
and U14875 (N_14875,N_13049,N_13496);
nand U14876 (N_14876,N_13463,N_13217);
nand U14877 (N_14877,N_13006,N_13108);
xnor U14878 (N_14878,N_13159,N_13338);
and U14879 (N_14879,N_13446,N_13344);
and U14880 (N_14880,N_13190,N_13430);
xnor U14881 (N_14881,N_13633,N_13497);
or U14882 (N_14882,N_13770,N_13442);
nand U14883 (N_14883,N_13185,N_13807);
or U14884 (N_14884,N_13062,N_13240);
xor U14885 (N_14885,N_13139,N_13740);
nand U14886 (N_14886,N_13657,N_13775);
nand U14887 (N_14887,N_13373,N_13029);
or U14888 (N_14888,N_13570,N_13779);
xnor U14889 (N_14889,N_13587,N_13098);
and U14890 (N_14890,N_13710,N_13872);
nor U14891 (N_14891,N_13108,N_13755);
and U14892 (N_14892,N_13223,N_13960);
xnor U14893 (N_14893,N_13608,N_13654);
and U14894 (N_14894,N_13435,N_13339);
nand U14895 (N_14895,N_13810,N_13255);
xor U14896 (N_14896,N_13385,N_13201);
nor U14897 (N_14897,N_13501,N_13072);
or U14898 (N_14898,N_13910,N_13809);
xor U14899 (N_14899,N_13803,N_13668);
or U14900 (N_14900,N_13908,N_13754);
xor U14901 (N_14901,N_13461,N_13001);
nor U14902 (N_14902,N_13360,N_13030);
and U14903 (N_14903,N_13321,N_13512);
xnor U14904 (N_14904,N_13584,N_13353);
xnor U14905 (N_14905,N_13658,N_13653);
nand U14906 (N_14906,N_13769,N_13407);
xor U14907 (N_14907,N_13231,N_13772);
nand U14908 (N_14908,N_13853,N_13088);
nor U14909 (N_14909,N_13785,N_13952);
nand U14910 (N_14910,N_13597,N_13895);
nand U14911 (N_14911,N_13897,N_13184);
xor U14912 (N_14912,N_13975,N_13598);
and U14913 (N_14913,N_13547,N_13199);
nand U14914 (N_14914,N_13265,N_13887);
xor U14915 (N_14915,N_13353,N_13934);
nand U14916 (N_14916,N_13493,N_13114);
and U14917 (N_14917,N_13125,N_13748);
nand U14918 (N_14918,N_13801,N_13156);
or U14919 (N_14919,N_13909,N_13211);
nor U14920 (N_14920,N_13758,N_13580);
nand U14921 (N_14921,N_13423,N_13684);
xor U14922 (N_14922,N_13951,N_13853);
or U14923 (N_14923,N_13777,N_13720);
nand U14924 (N_14924,N_13418,N_13577);
xnor U14925 (N_14925,N_13560,N_13374);
xor U14926 (N_14926,N_13734,N_13127);
nand U14927 (N_14927,N_13465,N_13850);
xnor U14928 (N_14928,N_13245,N_13905);
nand U14929 (N_14929,N_13175,N_13286);
or U14930 (N_14930,N_13810,N_13753);
xor U14931 (N_14931,N_13278,N_13653);
and U14932 (N_14932,N_13227,N_13909);
xnor U14933 (N_14933,N_13159,N_13947);
xor U14934 (N_14934,N_13403,N_13728);
and U14935 (N_14935,N_13473,N_13717);
xor U14936 (N_14936,N_13571,N_13616);
or U14937 (N_14937,N_13975,N_13804);
or U14938 (N_14938,N_13677,N_13174);
nand U14939 (N_14939,N_13833,N_13667);
nand U14940 (N_14940,N_13647,N_13955);
or U14941 (N_14941,N_13485,N_13897);
nor U14942 (N_14942,N_13783,N_13581);
nand U14943 (N_14943,N_13981,N_13042);
or U14944 (N_14944,N_13266,N_13032);
or U14945 (N_14945,N_13141,N_13423);
xnor U14946 (N_14946,N_13616,N_13882);
xor U14947 (N_14947,N_13801,N_13464);
nand U14948 (N_14948,N_13029,N_13654);
nand U14949 (N_14949,N_13044,N_13571);
or U14950 (N_14950,N_13019,N_13170);
xor U14951 (N_14951,N_13400,N_13420);
xor U14952 (N_14952,N_13777,N_13953);
nor U14953 (N_14953,N_13088,N_13195);
or U14954 (N_14954,N_13389,N_13641);
nand U14955 (N_14955,N_13728,N_13188);
nand U14956 (N_14956,N_13250,N_13975);
xor U14957 (N_14957,N_13153,N_13757);
nand U14958 (N_14958,N_13647,N_13926);
nor U14959 (N_14959,N_13745,N_13125);
nand U14960 (N_14960,N_13020,N_13416);
or U14961 (N_14961,N_13671,N_13124);
nand U14962 (N_14962,N_13401,N_13079);
and U14963 (N_14963,N_13720,N_13332);
and U14964 (N_14964,N_13440,N_13073);
and U14965 (N_14965,N_13305,N_13062);
nand U14966 (N_14966,N_13889,N_13845);
and U14967 (N_14967,N_13650,N_13757);
nand U14968 (N_14968,N_13733,N_13625);
or U14969 (N_14969,N_13471,N_13078);
nor U14970 (N_14970,N_13447,N_13327);
nor U14971 (N_14971,N_13167,N_13804);
nand U14972 (N_14972,N_13689,N_13841);
xnor U14973 (N_14973,N_13324,N_13901);
or U14974 (N_14974,N_13234,N_13141);
nand U14975 (N_14975,N_13647,N_13563);
nor U14976 (N_14976,N_13980,N_13145);
or U14977 (N_14977,N_13170,N_13767);
or U14978 (N_14978,N_13699,N_13688);
xor U14979 (N_14979,N_13310,N_13911);
nand U14980 (N_14980,N_13577,N_13429);
xnor U14981 (N_14981,N_13481,N_13266);
nand U14982 (N_14982,N_13572,N_13222);
xnor U14983 (N_14983,N_13181,N_13862);
nor U14984 (N_14984,N_13403,N_13493);
xnor U14985 (N_14985,N_13590,N_13901);
and U14986 (N_14986,N_13264,N_13429);
nand U14987 (N_14987,N_13953,N_13248);
or U14988 (N_14988,N_13623,N_13558);
and U14989 (N_14989,N_13600,N_13273);
or U14990 (N_14990,N_13042,N_13149);
or U14991 (N_14991,N_13998,N_13416);
nor U14992 (N_14992,N_13813,N_13518);
or U14993 (N_14993,N_13931,N_13968);
nand U14994 (N_14994,N_13066,N_13232);
and U14995 (N_14995,N_13094,N_13584);
or U14996 (N_14996,N_13690,N_13663);
and U14997 (N_14997,N_13799,N_13407);
nand U14998 (N_14998,N_13378,N_13861);
or U14999 (N_14999,N_13318,N_13079);
xnor UO_0 (O_0,N_14912,N_14334);
xor UO_1 (O_1,N_14482,N_14389);
nand UO_2 (O_2,N_14790,N_14857);
and UO_3 (O_3,N_14698,N_14124);
nor UO_4 (O_4,N_14766,N_14425);
nor UO_5 (O_5,N_14304,N_14097);
or UO_6 (O_6,N_14629,N_14803);
and UO_7 (O_7,N_14974,N_14746);
or UO_8 (O_8,N_14264,N_14432);
xor UO_9 (O_9,N_14694,N_14494);
and UO_10 (O_10,N_14162,N_14599);
xnor UO_11 (O_11,N_14420,N_14214);
xor UO_12 (O_12,N_14937,N_14479);
or UO_13 (O_13,N_14869,N_14745);
nand UO_14 (O_14,N_14961,N_14696);
and UO_15 (O_15,N_14598,N_14801);
and UO_16 (O_16,N_14738,N_14414);
xnor UO_17 (O_17,N_14680,N_14895);
nor UO_18 (O_18,N_14426,N_14915);
and UO_19 (O_19,N_14095,N_14930);
or UO_20 (O_20,N_14554,N_14679);
xor UO_21 (O_21,N_14613,N_14837);
xnor UO_22 (O_22,N_14643,N_14972);
and UO_23 (O_23,N_14617,N_14717);
nor UO_24 (O_24,N_14932,N_14891);
and UO_25 (O_25,N_14569,N_14834);
nand UO_26 (O_26,N_14605,N_14678);
or UO_27 (O_27,N_14435,N_14486);
and UO_28 (O_28,N_14656,N_14688);
or UO_29 (O_29,N_14503,N_14245);
or UO_30 (O_30,N_14959,N_14773);
and UO_31 (O_31,N_14042,N_14589);
and UO_32 (O_32,N_14765,N_14517);
nor UO_33 (O_33,N_14362,N_14971);
xor UO_34 (O_34,N_14390,N_14787);
nand UO_35 (O_35,N_14507,N_14575);
and UO_36 (O_36,N_14951,N_14906);
and UO_37 (O_37,N_14229,N_14927);
nand UO_38 (O_38,N_14037,N_14129);
xor UO_39 (O_39,N_14113,N_14463);
nor UO_40 (O_40,N_14004,N_14422);
nor UO_41 (O_41,N_14860,N_14441);
or UO_42 (O_42,N_14614,N_14813);
or UO_43 (O_43,N_14317,N_14371);
and UO_44 (O_44,N_14563,N_14898);
xnor UO_45 (O_45,N_14257,N_14663);
and UO_46 (O_46,N_14763,N_14006);
nand UO_47 (O_47,N_14594,N_14017);
nand UO_48 (O_48,N_14111,N_14190);
and UO_49 (O_49,N_14373,N_14865);
and UO_50 (O_50,N_14612,N_14168);
nor UO_51 (O_51,N_14883,N_14026);
nor UO_52 (O_52,N_14847,N_14743);
nand UO_53 (O_53,N_14173,N_14641);
and UO_54 (O_54,N_14545,N_14965);
nor UO_55 (O_55,N_14565,N_14789);
or UO_56 (O_56,N_14988,N_14704);
nor UO_57 (O_57,N_14293,N_14091);
nor UO_58 (O_58,N_14196,N_14066);
xnor UO_59 (O_59,N_14332,N_14513);
and UO_60 (O_60,N_14272,N_14300);
nand UO_61 (O_61,N_14203,N_14938);
or UO_62 (O_62,N_14606,N_14966);
xor UO_63 (O_63,N_14917,N_14438);
or UO_64 (O_64,N_14265,N_14281);
and UO_65 (O_65,N_14417,N_14537);
nor UO_66 (O_66,N_14053,N_14364);
or UO_67 (O_67,N_14924,N_14387);
and UO_68 (O_68,N_14327,N_14902);
nand UO_69 (O_69,N_14046,N_14237);
xor UO_70 (O_70,N_14261,N_14123);
nor UO_71 (O_71,N_14899,N_14716);
and UO_72 (O_72,N_14199,N_14761);
or UO_73 (O_73,N_14475,N_14511);
or UO_74 (O_74,N_14023,N_14114);
nand UO_75 (O_75,N_14806,N_14419);
nand UO_76 (O_76,N_14805,N_14268);
xor UO_77 (O_77,N_14999,N_14071);
nor UO_78 (O_78,N_14025,N_14952);
nor UO_79 (O_79,N_14838,N_14897);
and UO_80 (O_80,N_14050,N_14049);
or UO_81 (O_81,N_14205,N_14980);
and UO_82 (O_82,N_14428,N_14630);
nand UO_83 (O_83,N_14526,N_14666);
nor UO_84 (O_84,N_14263,N_14028);
and UO_85 (O_85,N_14771,N_14008);
and UO_86 (O_86,N_14351,N_14206);
xnor UO_87 (O_87,N_14607,N_14379);
nand UO_88 (O_88,N_14107,N_14142);
and UO_89 (O_89,N_14177,N_14741);
nand UO_90 (O_90,N_14442,N_14520);
nand UO_91 (O_91,N_14054,N_14730);
xor UO_92 (O_92,N_14885,N_14677);
xor UO_93 (O_93,N_14154,N_14892);
and UO_94 (O_94,N_14359,N_14833);
nand UO_95 (O_95,N_14143,N_14636);
or UO_96 (O_96,N_14628,N_14845);
nor UO_97 (O_97,N_14238,N_14207);
or UO_98 (O_98,N_14233,N_14112);
nor UO_99 (O_99,N_14712,N_14609);
and UO_100 (O_100,N_14243,N_14276);
xnor UO_101 (O_101,N_14910,N_14474);
xnor UO_102 (O_102,N_14780,N_14015);
nor UO_103 (O_103,N_14926,N_14187);
nor UO_104 (O_104,N_14156,N_14699);
nand UO_105 (O_105,N_14323,N_14374);
nor UO_106 (O_106,N_14828,N_14181);
or UO_107 (O_107,N_14434,N_14278);
nand UO_108 (O_108,N_14076,N_14559);
nor UO_109 (O_109,N_14752,N_14189);
nand UO_110 (O_110,N_14027,N_14361);
nand UO_111 (O_111,N_14851,N_14856);
or UO_112 (O_112,N_14476,N_14724);
nand UO_113 (O_113,N_14160,N_14218);
xnor UO_114 (O_114,N_14370,N_14638);
and UO_115 (O_115,N_14401,N_14574);
or UO_116 (O_116,N_14673,N_14500);
xnor UO_117 (O_117,N_14939,N_14600);
and UO_118 (O_118,N_14247,N_14282);
or UO_119 (O_119,N_14088,N_14991);
xnor UO_120 (O_120,N_14204,N_14538);
or UO_121 (O_121,N_14796,N_14943);
or UO_122 (O_122,N_14179,N_14650);
and UO_123 (O_123,N_14504,N_14175);
nor UO_124 (O_124,N_14848,N_14288);
or UO_125 (O_125,N_14251,N_14172);
and UO_126 (O_126,N_14769,N_14477);
and UO_127 (O_127,N_14552,N_14620);
nand UO_128 (O_128,N_14778,N_14530);
nand UO_129 (O_129,N_14038,N_14051);
and UO_130 (O_130,N_14239,N_14702);
or UO_131 (O_131,N_14692,N_14903);
nand UO_132 (O_132,N_14956,N_14874);
nor UO_133 (O_133,N_14399,N_14940);
nand UO_134 (O_134,N_14349,N_14336);
nand UO_135 (O_135,N_14515,N_14000);
nand UO_136 (O_136,N_14819,N_14485);
and UO_137 (O_137,N_14198,N_14985);
nor UO_138 (O_138,N_14918,N_14242);
nor UO_139 (O_139,N_14667,N_14708);
and UO_140 (O_140,N_14352,N_14764);
and UO_141 (O_141,N_14793,N_14122);
and UO_142 (O_142,N_14843,N_14270);
or UO_143 (O_143,N_14138,N_14627);
and UO_144 (O_144,N_14126,N_14659);
or UO_145 (O_145,N_14832,N_14465);
and UO_146 (O_146,N_14063,N_14292);
and UO_147 (O_147,N_14208,N_14227);
or UO_148 (O_148,N_14171,N_14383);
and UO_149 (O_149,N_14505,N_14445);
xnor UO_150 (O_150,N_14460,N_14496);
nand UO_151 (O_151,N_14608,N_14186);
and UO_152 (O_152,N_14169,N_14130);
or UO_153 (O_153,N_14751,N_14416);
xnor UO_154 (O_154,N_14909,N_14841);
and UO_155 (O_155,N_14089,N_14020);
nand UO_156 (O_156,N_14424,N_14521);
or UO_157 (O_157,N_14522,N_14307);
and UO_158 (O_158,N_14928,N_14984);
nand UO_159 (O_159,N_14150,N_14532);
nor UO_160 (O_160,N_14735,N_14954);
nor UO_161 (O_161,N_14440,N_14676);
nand UO_162 (O_162,N_14873,N_14774);
xor UO_163 (O_163,N_14758,N_14061);
or UO_164 (O_164,N_14427,N_14802);
nand UO_165 (O_165,N_14115,N_14753);
nor UO_166 (O_166,N_14092,N_14375);
nand UO_167 (O_167,N_14703,N_14945);
nand UO_168 (O_168,N_14710,N_14035);
or UO_169 (O_169,N_14353,N_14669);
and UO_170 (O_170,N_14622,N_14473);
xnor UO_171 (O_171,N_14674,N_14378);
nand UO_172 (O_172,N_14635,N_14280);
or UO_173 (O_173,N_14498,N_14182);
nand UO_174 (O_174,N_14534,N_14615);
nand UO_175 (O_175,N_14396,N_14106);
xnor UO_176 (O_176,N_14262,N_14525);
or UO_177 (O_177,N_14583,N_14623);
xnor UO_178 (O_178,N_14978,N_14550);
nor UO_179 (O_179,N_14369,N_14007);
nand UO_180 (O_180,N_14573,N_14217);
xnor UO_181 (O_181,N_14977,N_14893);
or UO_182 (O_182,N_14604,N_14029);
nand UO_183 (O_183,N_14081,N_14877);
and UO_184 (O_184,N_14824,N_14570);
or UO_185 (O_185,N_14448,N_14625);
xnor UO_186 (O_186,N_14481,N_14592);
and UO_187 (O_187,N_14571,N_14328);
or UO_188 (O_188,N_14256,N_14785);
nand UO_189 (O_189,N_14603,N_14754);
nor UO_190 (O_190,N_14222,N_14982);
and UO_191 (O_191,N_14810,N_14742);
or UO_192 (O_192,N_14315,N_14979);
xnor UO_193 (O_193,N_14346,N_14193);
nor UO_194 (O_194,N_14493,N_14719);
xor UO_195 (O_195,N_14707,N_14421);
or UO_196 (O_196,N_14737,N_14531);
and UO_197 (O_197,N_14639,N_14291);
nand UO_198 (O_198,N_14901,N_14911);
or UO_199 (O_199,N_14986,N_14516);
nor UO_200 (O_200,N_14104,N_14510);
xnor UO_201 (O_201,N_14544,N_14941);
nand UO_202 (O_202,N_14273,N_14740);
or UO_203 (O_203,N_14045,N_14040);
nand UO_204 (O_204,N_14458,N_14086);
xor UO_205 (O_205,N_14826,N_14788);
xor UO_206 (O_206,N_14944,N_14842);
nand UO_207 (O_207,N_14284,N_14644);
nand UO_208 (O_208,N_14632,N_14983);
or UO_209 (O_209,N_14110,N_14128);
or UO_210 (O_210,N_14118,N_14823);
nand UO_211 (O_211,N_14240,N_14070);
nand UO_212 (O_212,N_14394,N_14365);
and UO_213 (O_213,N_14827,N_14997);
xnor UO_214 (O_214,N_14957,N_14878);
xor UO_215 (O_215,N_14393,N_14726);
xor UO_216 (O_216,N_14800,N_14502);
or UO_217 (O_217,N_14541,N_14508);
nor UO_218 (O_218,N_14149,N_14593);
xor UO_219 (O_219,N_14405,N_14850);
xor UO_220 (O_220,N_14320,N_14555);
xnor UO_221 (O_221,N_14557,N_14277);
xnor UO_222 (O_222,N_14354,N_14407);
xnor UO_223 (O_223,N_14561,N_14167);
xnor UO_224 (O_224,N_14791,N_14658);
or UO_225 (O_225,N_14558,N_14335);
nand UO_226 (O_226,N_14949,N_14528);
and UO_227 (O_227,N_14385,N_14331);
xor UO_228 (O_228,N_14921,N_14372);
or UO_229 (O_229,N_14781,N_14451);
nor UO_230 (O_230,N_14109,N_14672);
xnor UO_231 (O_231,N_14194,N_14226);
nand UO_232 (O_232,N_14241,N_14514);
xnor UO_233 (O_233,N_14811,N_14572);
xnor UO_234 (O_234,N_14855,N_14818);
nor UO_235 (O_235,N_14079,N_14055);
and UO_236 (O_236,N_14152,N_14798);
nand UO_237 (O_237,N_14990,N_14144);
nand UO_238 (O_238,N_14799,N_14881);
nor UO_239 (O_239,N_14854,N_14147);
xor UO_240 (O_240,N_14436,N_14030);
nor UO_241 (O_241,N_14085,N_14987);
nor UO_242 (O_242,N_14914,N_14074);
xnor UO_243 (O_243,N_14931,N_14408);
xnor UO_244 (O_244,N_14259,N_14543);
nand UO_245 (O_245,N_14311,N_14859);
or UO_246 (O_246,N_14119,N_14887);
nor UO_247 (O_247,N_14995,N_14302);
and UO_248 (O_248,N_14595,N_14964);
nor UO_249 (O_249,N_14464,N_14794);
nor UO_250 (O_250,N_14760,N_14621);
and UO_251 (O_251,N_14453,N_14069);
xor UO_252 (O_252,N_14862,N_14922);
nand UO_253 (O_253,N_14768,N_14064);
nor UO_254 (O_254,N_14388,N_14861);
or UO_255 (O_255,N_14989,N_14718);
and UO_256 (O_256,N_14402,N_14014);
or UO_257 (O_257,N_14755,N_14398);
or UO_258 (O_258,N_14449,N_14670);
and UO_259 (O_259,N_14671,N_14096);
nor UO_260 (O_260,N_14444,N_14197);
nor UO_261 (O_261,N_14524,N_14624);
nor UO_262 (O_262,N_14312,N_14447);
nor UO_263 (O_263,N_14047,N_14337);
and UO_264 (O_264,N_14231,N_14568);
nand UO_265 (O_265,N_14835,N_14645);
and UO_266 (O_266,N_14075,N_14059);
or UO_267 (O_267,N_14715,N_14660);
or UO_268 (O_268,N_14219,N_14258);
or UO_269 (O_269,N_14133,N_14863);
nor UO_270 (O_270,N_14105,N_14936);
nor UO_271 (O_271,N_14299,N_14021);
and UO_272 (O_272,N_14184,N_14981);
nor UO_273 (O_273,N_14341,N_14750);
xnor UO_274 (O_274,N_14216,N_14736);
and UO_275 (O_275,N_14080,N_14062);
and UO_276 (O_276,N_14466,N_14546);
nor UO_277 (O_277,N_14722,N_14308);
or UO_278 (O_278,N_14876,N_14587);
or UO_279 (O_279,N_14711,N_14461);
nor UO_280 (O_280,N_14326,N_14094);
xnor UO_281 (O_281,N_14779,N_14815);
and UO_282 (O_282,N_14963,N_14333);
or UO_283 (O_283,N_14478,N_14343);
nand UO_284 (O_284,N_14749,N_14471);
xor UO_285 (O_285,N_14301,N_14356);
and UO_286 (O_286,N_14437,N_14597);
xor UO_287 (O_287,N_14536,N_14136);
nand UO_288 (O_288,N_14099,N_14489);
xnor UO_289 (O_289,N_14290,N_14303);
nor UO_290 (O_290,N_14720,N_14324);
nor UO_291 (O_291,N_14888,N_14005);
and UO_292 (O_292,N_14610,N_14784);
xnor UO_293 (O_293,N_14697,N_14423);
or UO_294 (O_294,N_14232,N_14358);
xor UO_295 (O_295,N_14675,N_14920);
or UO_296 (O_296,N_14322,N_14446);
and UO_297 (O_297,N_14034,N_14866);
or UO_298 (O_298,N_14889,N_14579);
and UO_299 (O_299,N_14215,N_14691);
or UO_300 (O_300,N_14433,N_14289);
nor UO_301 (O_301,N_14491,N_14221);
and UO_302 (O_302,N_14919,N_14795);
or UO_303 (O_303,N_14732,N_14844);
and UO_304 (O_304,N_14487,N_14868);
or UO_305 (O_305,N_14705,N_14117);
nand UO_306 (O_306,N_14472,N_14266);
or UO_307 (O_307,N_14533,N_14973);
xnor UO_308 (O_308,N_14413,N_14905);
nand UO_309 (O_309,N_14542,N_14586);
or UO_310 (O_310,N_14211,N_14392);
nand UO_311 (O_311,N_14596,N_14872);
nand UO_312 (O_312,N_14611,N_14452);
xnor UO_313 (O_313,N_14223,N_14495);
nand UO_314 (O_314,N_14016,N_14041);
and UO_315 (O_315,N_14523,N_14512);
or UO_316 (O_316,N_14376,N_14996);
nand UO_317 (O_317,N_14907,N_14654);
and UO_318 (O_318,N_14871,N_14830);
nor UO_319 (O_319,N_14849,N_14430);
or UO_320 (O_320,N_14509,N_14879);
and UO_321 (O_321,N_14825,N_14633);
nand UO_322 (O_322,N_14224,N_14900);
nor UO_323 (O_323,N_14338,N_14455);
xor UO_324 (O_324,N_14381,N_14640);
nand UO_325 (O_325,N_14244,N_14391);
nor UO_326 (O_326,N_14116,N_14649);
xnor UO_327 (O_327,N_14431,N_14072);
and UO_328 (O_328,N_14342,N_14101);
or UO_329 (O_329,N_14068,N_14191);
or UO_330 (O_330,N_14220,N_14783);
xor UO_331 (O_331,N_14816,N_14011);
and UO_332 (O_332,N_14748,N_14867);
nor UO_333 (O_333,N_14141,N_14032);
nor UO_334 (O_334,N_14652,N_14411);
and UO_335 (O_335,N_14295,N_14706);
or UO_336 (O_336,N_14180,N_14298);
xnor UO_337 (O_337,N_14321,N_14083);
or UO_338 (O_338,N_14044,N_14807);
and UO_339 (O_339,N_14585,N_14368);
nand UO_340 (O_340,N_14274,N_14934);
nor UO_341 (O_341,N_14693,N_14131);
nand UO_342 (O_342,N_14882,N_14916);
and UO_343 (O_343,N_14875,N_14820);
and UO_344 (O_344,N_14657,N_14057);
nand UO_345 (O_345,N_14384,N_14084);
nor UO_346 (O_346,N_14454,N_14380);
and UO_347 (O_347,N_14056,N_14287);
xor UO_348 (O_348,N_14929,N_14584);
nor UO_349 (O_349,N_14969,N_14013);
xnor UO_350 (O_350,N_14817,N_14252);
and UO_351 (O_351,N_14024,N_14852);
and UO_352 (O_352,N_14499,N_14976);
nand UO_353 (O_353,N_14450,N_14003);
and UO_354 (O_354,N_14950,N_14067);
or UO_355 (O_355,N_14560,N_14782);
nor UO_356 (O_356,N_14562,N_14853);
xor UO_357 (O_357,N_14551,N_14357);
nor UO_358 (O_358,N_14134,N_14188);
xor UO_359 (O_359,N_14733,N_14022);
or UO_360 (O_360,N_14812,N_14283);
xnor UO_361 (O_361,N_14060,N_14683);
nor UO_362 (O_362,N_14567,N_14043);
nand UO_363 (O_363,N_14468,N_14155);
nand UO_364 (O_364,N_14582,N_14153);
nor UO_365 (O_365,N_14814,N_14344);
or UO_366 (O_366,N_14870,N_14310);
xnor UO_367 (O_367,N_14200,N_14403);
xnor UO_368 (O_368,N_14686,N_14935);
and UO_369 (O_369,N_14962,N_14662);
nor UO_370 (O_370,N_14618,N_14925);
xor UO_371 (O_371,N_14137,N_14121);
nand UO_372 (O_372,N_14540,N_14098);
nor UO_373 (O_373,N_14340,N_14684);
nor UO_374 (O_374,N_14165,N_14090);
nand UO_375 (O_375,N_14201,N_14183);
or UO_376 (O_376,N_14619,N_14174);
xor UO_377 (O_377,N_14125,N_14386);
or UO_378 (O_378,N_14588,N_14576);
xor UO_379 (O_379,N_14178,N_14467);
or UO_380 (O_380,N_14564,N_14260);
nand UO_381 (O_381,N_14234,N_14469);
or UO_382 (O_382,N_14923,N_14527);
nor UO_383 (O_383,N_14580,N_14230);
and UO_384 (O_384,N_14484,N_14501);
nand UO_385 (O_385,N_14958,N_14553);
and UO_386 (O_386,N_14689,N_14626);
nand UO_387 (O_387,N_14347,N_14809);
and UO_388 (O_388,N_14225,N_14884);
nand UO_389 (O_389,N_14202,N_14255);
nand UO_390 (O_390,N_14739,N_14100);
or UO_391 (O_391,N_14661,N_14547);
and UO_392 (O_392,N_14457,N_14195);
or UO_393 (O_393,N_14470,N_14729);
or UO_394 (O_394,N_14313,N_14363);
xor UO_395 (O_395,N_14590,N_14395);
xnor UO_396 (O_396,N_14329,N_14170);
xnor UO_397 (O_397,N_14767,N_14176);
nor UO_398 (O_398,N_14968,N_14275);
and UO_399 (O_399,N_14157,N_14139);
and UO_400 (O_400,N_14151,N_14960);
nand UO_401 (O_401,N_14776,N_14490);
nand UO_402 (O_402,N_14325,N_14880);
or UO_403 (O_403,N_14992,N_14757);
and UO_404 (O_404,N_14518,N_14886);
and UO_405 (O_405,N_14808,N_14655);
nor UO_406 (O_406,N_14161,N_14286);
and UO_407 (O_407,N_14734,N_14459);
or UO_408 (O_408,N_14519,N_14836);
xor UO_409 (O_409,N_14946,N_14839);
and UO_410 (O_410,N_14665,N_14690);
and UO_411 (O_411,N_14078,N_14093);
or UO_412 (O_412,N_14132,N_14001);
xnor UO_413 (O_413,N_14591,N_14355);
nand UO_414 (O_414,N_14728,N_14314);
nor UO_415 (O_415,N_14019,N_14249);
xnor UO_416 (O_416,N_14727,N_14581);
nor UO_417 (O_417,N_14148,N_14488);
xor UO_418 (O_418,N_14831,N_14804);
xnor UO_419 (O_419,N_14345,N_14942);
nor UO_420 (O_420,N_14998,N_14566);
or UO_421 (O_421,N_14506,N_14330);
or UO_422 (O_422,N_14339,N_14412);
nor UO_423 (O_423,N_14382,N_14777);
nand UO_424 (O_424,N_14377,N_14653);
and UO_425 (O_425,N_14770,N_14246);
xor UO_426 (O_426,N_14319,N_14350);
xor UO_427 (O_427,N_14140,N_14146);
nor UO_428 (O_428,N_14822,N_14577);
and UO_429 (O_429,N_14406,N_14253);
xnor UO_430 (O_430,N_14668,N_14158);
nor UO_431 (O_431,N_14418,N_14642);
and UO_432 (O_432,N_14462,N_14185);
and UO_433 (O_433,N_14695,N_14556);
and UO_434 (O_434,N_14012,N_14018);
or UO_435 (O_435,N_14975,N_14967);
xor UO_436 (O_436,N_14549,N_14775);
or UO_437 (O_437,N_14756,N_14052);
xnor UO_438 (O_438,N_14723,N_14772);
and UO_439 (O_439,N_14058,N_14637);
or UO_440 (O_440,N_14166,N_14073);
nor UO_441 (O_441,N_14578,N_14483);
xnor UO_442 (O_442,N_14908,N_14953);
and UO_443 (O_443,N_14647,N_14439);
xnor UO_444 (O_444,N_14294,N_14309);
nor UO_445 (O_445,N_14318,N_14039);
or UO_446 (O_446,N_14682,N_14360);
xnor UO_447 (O_447,N_14009,N_14700);
xnor UO_448 (O_448,N_14002,N_14415);
or UO_449 (O_449,N_14648,N_14108);
xnor UO_450 (O_450,N_14762,N_14994);
nand UO_451 (O_451,N_14145,N_14316);
nand UO_452 (O_452,N_14948,N_14236);
or UO_453 (O_453,N_14497,N_14228);
and UO_454 (O_454,N_14993,N_14970);
nand UO_455 (O_455,N_14159,N_14048);
and UO_456 (O_456,N_14456,N_14404);
or UO_457 (O_457,N_14367,N_14306);
nand UO_458 (O_458,N_14731,N_14209);
and UO_459 (O_459,N_14409,N_14548);
nor UO_460 (O_460,N_14858,N_14297);
nor UO_461 (O_461,N_14864,N_14120);
xnor UO_462 (O_462,N_14492,N_14759);
and UO_463 (O_463,N_14933,N_14267);
nand UO_464 (O_464,N_14010,N_14601);
xor UO_465 (O_465,N_14033,N_14947);
xor UO_466 (O_466,N_14792,N_14210);
xnor UO_467 (O_467,N_14087,N_14721);
nand UO_468 (O_468,N_14631,N_14480);
or UO_469 (O_469,N_14366,N_14685);
nand UO_470 (O_470,N_14602,N_14429);
nand UO_471 (O_471,N_14077,N_14410);
or UO_472 (O_472,N_14913,N_14285);
or UO_473 (O_473,N_14248,N_14713);
or UO_474 (O_474,N_14955,N_14701);
nand UO_475 (O_475,N_14646,N_14296);
nor UO_476 (O_476,N_14192,N_14539);
or UO_477 (O_477,N_14269,N_14786);
nor UO_478 (O_478,N_14254,N_14127);
nand UO_479 (O_479,N_14031,N_14535);
and UO_480 (O_480,N_14102,N_14135);
nand UO_481 (O_481,N_14687,N_14797);
nor UO_482 (O_482,N_14894,N_14747);
nand UO_483 (O_483,N_14829,N_14714);
or UO_484 (O_484,N_14036,N_14279);
nand UO_485 (O_485,N_14212,N_14271);
and UO_486 (O_486,N_14305,N_14681);
nor UO_487 (O_487,N_14213,N_14400);
and UO_488 (O_488,N_14821,N_14348);
xor UO_489 (O_489,N_14065,N_14725);
and UO_490 (O_490,N_14529,N_14103);
nor UO_491 (O_491,N_14664,N_14744);
nand UO_492 (O_492,N_14651,N_14616);
or UO_493 (O_493,N_14163,N_14890);
nand UO_494 (O_494,N_14896,N_14164);
xor UO_495 (O_495,N_14235,N_14634);
xor UO_496 (O_496,N_14443,N_14840);
xnor UO_497 (O_497,N_14082,N_14250);
nand UO_498 (O_498,N_14846,N_14709);
xor UO_499 (O_499,N_14904,N_14397);
nor UO_500 (O_500,N_14050,N_14512);
or UO_501 (O_501,N_14132,N_14930);
and UO_502 (O_502,N_14872,N_14542);
xor UO_503 (O_503,N_14761,N_14489);
nand UO_504 (O_504,N_14985,N_14766);
or UO_505 (O_505,N_14426,N_14118);
and UO_506 (O_506,N_14939,N_14903);
and UO_507 (O_507,N_14648,N_14969);
xor UO_508 (O_508,N_14001,N_14445);
nor UO_509 (O_509,N_14135,N_14913);
nor UO_510 (O_510,N_14958,N_14642);
nand UO_511 (O_511,N_14175,N_14593);
or UO_512 (O_512,N_14639,N_14205);
and UO_513 (O_513,N_14073,N_14114);
and UO_514 (O_514,N_14119,N_14638);
and UO_515 (O_515,N_14255,N_14340);
xnor UO_516 (O_516,N_14854,N_14455);
nand UO_517 (O_517,N_14565,N_14024);
or UO_518 (O_518,N_14254,N_14465);
nand UO_519 (O_519,N_14511,N_14946);
or UO_520 (O_520,N_14850,N_14201);
or UO_521 (O_521,N_14870,N_14788);
and UO_522 (O_522,N_14030,N_14750);
or UO_523 (O_523,N_14897,N_14537);
and UO_524 (O_524,N_14365,N_14793);
nor UO_525 (O_525,N_14092,N_14419);
and UO_526 (O_526,N_14186,N_14831);
or UO_527 (O_527,N_14020,N_14877);
nand UO_528 (O_528,N_14663,N_14486);
and UO_529 (O_529,N_14480,N_14753);
nor UO_530 (O_530,N_14077,N_14225);
and UO_531 (O_531,N_14896,N_14105);
nand UO_532 (O_532,N_14403,N_14173);
nand UO_533 (O_533,N_14667,N_14219);
nor UO_534 (O_534,N_14627,N_14454);
xor UO_535 (O_535,N_14602,N_14204);
and UO_536 (O_536,N_14665,N_14151);
nand UO_537 (O_537,N_14624,N_14733);
nand UO_538 (O_538,N_14057,N_14546);
or UO_539 (O_539,N_14730,N_14356);
xor UO_540 (O_540,N_14719,N_14635);
or UO_541 (O_541,N_14619,N_14491);
xnor UO_542 (O_542,N_14673,N_14060);
or UO_543 (O_543,N_14046,N_14605);
or UO_544 (O_544,N_14203,N_14589);
nor UO_545 (O_545,N_14342,N_14112);
or UO_546 (O_546,N_14801,N_14466);
xor UO_547 (O_547,N_14767,N_14975);
or UO_548 (O_548,N_14131,N_14595);
nor UO_549 (O_549,N_14321,N_14810);
nor UO_550 (O_550,N_14947,N_14828);
and UO_551 (O_551,N_14785,N_14481);
xnor UO_552 (O_552,N_14614,N_14840);
nor UO_553 (O_553,N_14790,N_14166);
xnor UO_554 (O_554,N_14675,N_14012);
nand UO_555 (O_555,N_14693,N_14383);
nand UO_556 (O_556,N_14132,N_14981);
and UO_557 (O_557,N_14381,N_14937);
and UO_558 (O_558,N_14355,N_14634);
and UO_559 (O_559,N_14059,N_14006);
and UO_560 (O_560,N_14797,N_14547);
or UO_561 (O_561,N_14378,N_14368);
or UO_562 (O_562,N_14464,N_14161);
and UO_563 (O_563,N_14375,N_14119);
and UO_564 (O_564,N_14216,N_14375);
nor UO_565 (O_565,N_14312,N_14701);
nand UO_566 (O_566,N_14211,N_14894);
and UO_567 (O_567,N_14509,N_14626);
nand UO_568 (O_568,N_14903,N_14286);
and UO_569 (O_569,N_14883,N_14744);
or UO_570 (O_570,N_14842,N_14656);
nand UO_571 (O_571,N_14486,N_14969);
nor UO_572 (O_572,N_14491,N_14286);
and UO_573 (O_573,N_14433,N_14036);
xor UO_574 (O_574,N_14805,N_14400);
or UO_575 (O_575,N_14000,N_14390);
nand UO_576 (O_576,N_14308,N_14046);
or UO_577 (O_577,N_14571,N_14188);
and UO_578 (O_578,N_14208,N_14822);
nand UO_579 (O_579,N_14194,N_14611);
xnor UO_580 (O_580,N_14816,N_14935);
nor UO_581 (O_581,N_14009,N_14816);
or UO_582 (O_582,N_14545,N_14417);
xor UO_583 (O_583,N_14446,N_14147);
and UO_584 (O_584,N_14771,N_14813);
nand UO_585 (O_585,N_14495,N_14924);
xnor UO_586 (O_586,N_14049,N_14798);
and UO_587 (O_587,N_14407,N_14623);
nand UO_588 (O_588,N_14770,N_14789);
nor UO_589 (O_589,N_14773,N_14297);
and UO_590 (O_590,N_14284,N_14172);
nor UO_591 (O_591,N_14991,N_14370);
nand UO_592 (O_592,N_14737,N_14911);
or UO_593 (O_593,N_14651,N_14173);
nand UO_594 (O_594,N_14769,N_14674);
and UO_595 (O_595,N_14365,N_14254);
nor UO_596 (O_596,N_14796,N_14039);
nand UO_597 (O_597,N_14066,N_14639);
and UO_598 (O_598,N_14199,N_14247);
or UO_599 (O_599,N_14139,N_14879);
and UO_600 (O_600,N_14422,N_14444);
or UO_601 (O_601,N_14267,N_14490);
or UO_602 (O_602,N_14260,N_14230);
nor UO_603 (O_603,N_14082,N_14550);
nor UO_604 (O_604,N_14576,N_14803);
or UO_605 (O_605,N_14718,N_14660);
or UO_606 (O_606,N_14417,N_14880);
xnor UO_607 (O_607,N_14419,N_14794);
or UO_608 (O_608,N_14468,N_14658);
nor UO_609 (O_609,N_14424,N_14282);
nand UO_610 (O_610,N_14031,N_14582);
nand UO_611 (O_611,N_14391,N_14826);
nand UO_612 (O_612,N_14971,N_14430);
and UO_613 (O_613,N_14621,N_14601);
nand UO_614 (O_614,N_14213,N_14694);
nand UO_615 (O_615,N_14822,N_14617);
xnor UO_616 (O_616,N_14068,N_14010);
and UO_617 (O_617,N_14405,N_14727);
xor UO_618 (O_618,N_14299,N_14884);
xor UO_619 (O_619,N_14244,N_14760);
nand UO_620 (O_620,N_14555,N_14027);
nand UO_621 (O_621,N_14201,N_14179);
nor UO_622 (O_622,N_14856,N_14340);
xor UO_623 (O_623,N_14458,N_14028);
and UO_624 (O_624,N_14337,N_14683);
or UO_625 (O_625,N_14099,N_14705);
and UO_626 (O_626,N_14129,N_14785);
or UO_627 (O_627,N_14745,N_14137);
nor UO_628 (O_628,N_14495,N_14020);
xnor UO_629 (O_629,N_14900,N_14036);
xor UO_630 (O_630,N_14455,N_14063);
nand UO_631 (O_631,N_14138,N_14076);
nor UO_632 (O_632,N_14878,N_14762);
nor UO_633 (O_633,N_14342,N_14749);
nor UO_634 (O_634,N_14218,N_14782);
nor UO_635 (O_635,N_14887,N_14144);
nand UO_636 (O_636,N_14939,N_14132);
or UO_637 (O_637,N_14622,N_14321);
nand UO_638 (O_638,N_14810,N_14248);
xor UO_639 (O_639,N_14371,N_14491);
and UO_640 (O_640,N_14157,N_14083);
or UO_641 (O_641,N_14559,N_14498);
xnor UO_642 (O_642,N_14309,N_14048);
xor UO_643 (O_643,N_14832,N_14837);
nor UO_644 (O_644,N_14078,N_14343);
nor UO_645 (O_645,N_14525,N_14825);
xor UO_646 (O_646,N_14782,N_14008);
xor UO_647 (O_647,N_14486,N_14130);
xnor UO_648 (O_648,N_14302,N_14988);
and UO_649 (O_649,N_14766,N_14322);
nor UO_650 (O_650,N_14175,N_14800);
nand UO_651 (O_651,N_14501,N_14777);
nor UO_652 (O_652,N_14287,N_14327);
or UO_653 (O_653,N_14110,N_14108);
nor UO_654 (O_654,N_14756,N_14616);
nor UO_655 (O_655,N_14958,N_14718);
nand UO_656 (O_656,N_14437,N_14222);
nand UO_657 (O_657,N_14249,N_14935);
and UO_658 (O_658,N_14735,N_14139);
nor UO_659 (O_659,N_14270,N_14408);
nor UO_660 (O_660,N_14232,N_14979);
and UO_661 (O_661,N_14975,N_14955);
nor UO_662 (O_662,N_14613,N_14638);
and UO_663 (O_663,N_14754,N_14141);
xor UO_664 (O_664,N_14989,N_14990);
nor UO_665 (O_665,N_14997,N_14479);
and UO_666 (O_666,N_14206,N_14599);
and UO_667 (O_667,N_14217,N_14829);
nand UO_668 (O_668,N_14032,N_14356);
nor UO_669 (O_669,N_14735,N_14322);
nor UO_670 (O_670,N_14986,N_14419);
or UO_671 (O_671,N_14302,N_14905);
nand UO_672 (O_672,N_14894,N_14165);
nand UO_673 (O_673,N_14843,N_14765);
nand UO_674 (O_674,N_14121,N_14261);
or UO_675 (O_675,N_14831,N_14023);
and UO_676 (O_676,N_14911,N_14342);
xor UO_677 (O_677,N_14675,N_14633);
nor UO_678 (O_678,N_14888,N_14955);
or UO_679 (O_679,N_14485,N_14573);
nand UO_680 (O_680,N_14987,N_14238);
and UO_681 (O_681,N_14505,N_14640);
xor UO_682 (O_682,N_14795,N_14102);
xnor UO_683 (O_683,N_14642,N_14145);
nor UO_684 (O_684,N_14812,N_14881);
and UO_685 (O_685,N_14879,N_14946);
and UO_686 (O_686,N_14018,N_14859);
or UO_687 (O_687,N_14624,N_14513);
nand UO_688 (O_688,N_14774,N_14507);
or UO_689 (O_689,N_14031,N_14061);
and UO_690 (O_690,N_14532,N_14842);
xnor UO_691 (O_691,N_14971,N_14133);
or UO_692 (O_692,N_14160,N_14455);
and UO_693 (O_693,N_14384,N_14223);
nand UO_694 (O_694,N_14796,N_14224);
or UO_695 (O_695,N_14328,N_14685);
and UO_696 (O_696,N_14085,N_14058);
or UO_697 (O_697,N_14313,N_14389);
and UO_698 (O_698,N_14061,N_14057);
and UO_699 (O_699,N_14189,N_14923);
nor UO_700 (O_700,N_14411,N_14993);
xor UO_701 (O_701,N_14477,N_14040);
and UO_702 (O_702,N_14867,N_14455);
nand UO_703 (O_703,N_14113,N_14771);
or UO_704 (O_704,N_14644,N_14236);
and UO_705 (O_705,N_14967,N_14350);
and UO_706 (O_706,N_14553,N_14783);
nor UO_707 (O_707,N_14405,N_14800);
nand UO_708 (O_708,N_14113,N_14593);
and UO_709 (O_709,N_14623,N_14895);
or UO_710 (O_710,N_14650,N_14889);
or UO_711 (O_711,N_14425,N_14751);
nand UO_712 (O_712,N_14028,N_14772);
nand UO_713 (O_713,N_14629,N_14925);
nand UO_714 (O_714,N_14469,N_14360);
nor UO_715 (O_715,N_14468,N_14234);
or UO_716 (O_716,N_14092,N_14387);
nand UO_717 (O_717,N_14565,N_14165);
nor UO_718 (O_718,N_14379,N_14706);
and UO_719 (O_719,N_14937,N_14150);
nand UO_720 (O_720,N_14411,N_14034);
nand UO_721 (O_721,N_14020,N_14326);
and UO_722 (O_722,N_14152,N_14795);
nor UO_723 (O_723,N_14843,N_14051);
or UO_724 (O_724,N_14890,N_14433);
xor UO_725 (O_725,N_14102,N_14670);
and UO_726 (O_726,N_14843,N_14746);
nor UO_727 (O_727,N_14284,N_14731);
or UO_728 (O_728,N_14812,N_14239);
or UO_729 (O_729,N_14968,N_14001);
or UO_730 (O_730,N_14357,N_14884);
and UO_731 (O_731,N_14500,N_14615);
or UO_732 (O_732,N_14995,N_14619);
nor UO_733 (O_733,N_14858,N_14583);
or UO_734 (O_734,N_14328,N_14393);
xor UO_735 (O_735,N_14293,N_14905);
nand UO_736 (O_736,N_14634,N_14386);
and UO_737 (O_737,N_14944,N_14830);
xnor UO_738 (O_738,N_14137,N_14977);
xnor UO_739 (O_739,N_14324,N_14044);
and UO_740 (O_740,N_14075,N_14177);
xnor UO_741 (O_741,N_14508,N_14817);
nand UO_742 (O_742,N_14303,N_14782);
nand UO_743 (O_743,N_14964,N_14539);
or UO_744 (O_744,N_14873,N_14469);
and UO_745 (O_745,N_14933,N_14175);
nand UO_746 (O_746,N_14703,N_14510);
nand UO_747 (O_747,N_14401,N_14413);
nand UO_748 (O_748,N_14752,N_14762);
nor UO_749 (O_749,N_14660,N_14301);
and UO_750 (O_750,N_14216,N_14448);
nand UO_751 (O_751,N_14432,N_14454);
nor UO_752 (O_752,N_14190,N_14648);
or UO_753 (O_753,N_14354,N_14135);
or UO_754 (O_754,N_14760,N_14136);
and UO_755 (O_755,N_14359,N_14617);
nor UO_756 (O_756,N_14721,N_14559);
or UO_757 (O_757,N_14345,N_14045);
or UO_758 (O_758,N_14866,N_14988);
or UO_759 (O_759,N_14023,N_14310);
nand UO_760 (O_760,N_14980,N_14105);
xor UO_761 (O_761,N_14360,N_14906);
xor UO_762 (O_762,N_14250,N_14123);
xor UO_763 (O_763,N_14292,N_14821);
xnor UO_764 (O_764,N_14871,N_14509);
nand UO_765 (O_765,N_14152,N_14345);
nor UO_766 (O_766,N_14225,N_14906);
nor UO_767 (O_767,N_14270,N_14189);
xor UO_768 (O_768,N_14368,N_14800);
or UO_769 (O_769,N_14032,N_14574);
or UO_770 (O_770,N_14181,N_14535);
nor UO_771 (O_771,N_14481,N_14997);
xnor UO_772 (O_772,N_14776,N_14619);
xnor UO_773 (O_773,N_14951,N_14202);
nand UO_774 (O_774,N_14988,N_14870);
nand UO_775 (O_775,N_14036,N_14679);
and UO_776 (O_776,N_14652,N_14837);
xor UO_777 (O_777,N_14141,N_14158);
nor UO_778 (O_778,N_14373,N_14649);
xor UO_779 (O_779,N_14156,N_14851);
nor UO_780 (O_780,N_14993,N_14663);
nor UO_781 (O_781,N_14304,N_14206);
nand UO_782 (O_782,N_14578,N_14273);
xnor UO_783 (O_783,N_14327,N_14354);
and UO_784 (O_784,N_14657,N_14654);
nor UO_785 (O_785,N_14078,N_14641);
xor UO_786 (O_786,N_14864,N_14769);
or UO_787 (O_787,N_14072,N_14595);
nor UO_788 (O_788,N_14469,N_14133);
xor UO_789 (O_789,N_14478,N_14139);
or UO_790 (O_790,N_14204,N_14217);
or UO_791 (O_791,N_14689,N_14812);
or UO_792 (O_792,N_14601,N_14741);
xnor UO_793 (O_793,N_14317,N_14926);
nor UO_794 (O_794,N_14112,N_14715);
nand UO_795 (O_795,N_14264,N_14780);
and UO_796 (O_796,N_14458,N_14608);
or UO_797 (O_797,N_14573,N_14951);
or UO_798 (O_798,N_14521,N_14597);
xnor UO_799 (O_799,N_14392,N_14432);
nand UO_800 (O_800,N_14729,N_14082);
nor UO_801 (O_801,N_14975,N_14926);
and UO_802 (O_802,N_14517,N_14838);
or UO_803 (O_803,N_14935,N_14123);
and UO_804 (O_804,N_14536,N_14637);
xnor UO_805 (O_805,N_14540,N_14096);
nand UO_806 (O_806,N_14141,N_14765);
or UO_807 (O_807,N_14060,N_14214);
nor UO_808 (O_808,N_14209,N_14001);
or UO_809 (O_809,N_14446,N_14999);
and UO_810 (O_810,N_14265,N_14939);
xnor UO_811 (O_811,N_14319,N_14615);
and UO_812 (O_812,N_14385,N_14620);
xnor UO_813 (O_813,N_14541,N_14491);
xor UO_814 (O_814,N_14462,N_14274);
and UO_815 (O_815,N_14011,N_14396);
nand UO_816 (O_816,N_14168,N_14009);
xnor UO_817 (O_817,N_14209,N_14348);
or UO_818 (O_818,N_14767,N_14661);
nand UO_819 (O_819,N_14647,N_14247);
xor UO_820 (O_820,N_14815,N_14047);
nor UO_821 (O_821,N_14813,N_14630);
nor UO_822 (O_822,N_14669,N_14303);
nand UO_823 (O_823,N_14770,N_14098);
or UO_824 (O_824,N_14456,N_14839);
or UO_825 (O_825,N_14246,N_14970);
and UO_826 (O_826,N_14033,N_14915);
xnor UO_827 (O_827,N_14351,N_14504);
nand UO_828 (O_828,N_14823,N_14778);
nor UO_829 (O_829,N_14274,N_14611);
xnor UO_830 (O_830,N_14309,N_14177);
or UO_831 (O_831,N_14922,N_14887);
or UO_832 (O_832,N_14391,N_14726);
and UO_833 (O_833,N_14605,N_14377);
xor UO_834 (O_834,N_14497,N_14706);
nor UO_835 (O_835,N_14041,N_14538);
or UO_836 (O_836,N_14268,N_14327);
or UO_837 (O_837,N_14867,N_14127);
and UO_838 (O_838,N_14776,N_14621);
nor UO_839 (O_839,N_14153,N_14141);
and UO_840 (O_840,N_14430,N_14677);
and UO_841 (O_841,N_14690,N_14628);
or UO_842 (O_842,N_14979,N_14701);
and UO_843 (O_843,N_14492,N_14584);
nand UO_844 (O_844,N_14356,N_14051);
nand UO_845 (O_845,N_14962,N_14399);
nand UO_846 (O_846,N_14665,N_14317);
xor UO_847 (O_847,N_14097,N_14456);
xnor UO_848 (O_848,N_14778,N_14827);
nor UO_849 (O_849,N_14228,N_14601);
nor UO_850 (O_850,N_14428,N_14607);
xor UO_851 (O_851,N_14309,N_14299);
and UO_852 (O_852,N_14603,N_14325);
or UO_853 (O_853,N_14468,N_14380);
nor UO_854 (O_854,N_14339,N_14168);
and UO_855 (O_855,N_14817,N_14006);
nand UO_856 (O_856,N_14911,N_14113);
nand UO_857 (O_857,N_14705,N_14516);
xnor UO_858 (O_858,N_14286,N_14870);
and UO_859 (O_859,N_14960,N_14810);
xor UO_860 (O_860,N_14598,N_14392);
and UO_861 (O_861,N_14336,N_14816);
xor UO_862 (O_862,N_14224,N_14411);
or UO_863 (O_863,N_14082,N_14587);
nand UO_864 (O_864,N_14490,N_14695);
nand UO_865 (O_865,N_14674,N_14533);
nor UO_866 (O_866,N_14459,N_14143);
nand UO_867 (O_867,N_14370,N_14601);
and UO_868 (O_868,N_14084,N_14154);
nand UO_869 (O_869,N_14101,N_14220);
nand UO_870 (O_870,N_14153,N_14937);
nor UO_871 (O_871,N_14147,N_14219);
or UO_872 (O_872,N_14644,N_14315);
and UO_873 (O_873,N_14228,N_14608);
or UO_874 (O_874,N_14335,N_14572);
and UO_875 (O_875,N_14279,N_14246);
and UO_876 (O_876,N_14389,N_14933);
nand UO_877 (O_877,N_14357,N_14245);
nor UO_878 (O_878,N_14109,N_14852);
xor UO_879 (O_879,N_14303,N_14023);
or UO_880 (O_880,N_14024,N_14475);
xor UO_881 (O_881,N_14906,N_14352);
or UO_882 (O_882,N_14677,N_14035);
nand UO_883 (O_883,N_14669,N_14054);
nand UO_884 (O_884,N_14430,N_14762);
xor UO_885 (O_885,N_14865,N_14070);
nor UO_886 (O_886,N_14627,N_14540);
or UO_887 (O_887,N_14864,N_14138);
and UO_888 (O_888,N_14678,N_14430);
xnor UO_889 (O_889,N_14938,N_14476);
xor UO_890 (O_890,N_14177,N_14745);
and UO_891 (O_891,N_14313,N_14298);
nand UO_892 (O_892,N_14640,N_14652);
nor UO_893 (O_893,N_14553,N_14735);
nor UO_894 (O_894,N_14721,N_14806);
or UO_895 (O_895,N_14335,N_14993);
and UO_896 (O_896,N_14201,N_14917);
xor UO_897 (O_897,N_14713,N_14702);
nand UO_898 (O_898,N_14990,N_14405);
xnor UO_899 (O_899,N_14881,N_14188);
and UO_900 (O_900,N_14817,N_14078);
or UO_901 (O_901,N_14915,N_14863);
and UO_902 (O_902,N_14960,N_14549);
or UO_903 (O_903,N_14455,N_14007);
nand UO_904 (O_904,N_14370,N_14471);
nor UO_905 (O_905,N_14917,N_14003);
xor UO_906 (O_906,N_14034,N_14150);
nand UO_907 (O_907,N_14302,N_14232);
or UO_908 (O_908,N_14474,N_14384);
nand UO_909 (O_909,N_14109,N_14068);
or UO_910 (O_910,N_14383,N_14053);
and UO_911 (O_911,N_14190,N_14857);
or UO_912 (O_912,N_14584,N_14549);
and UO_913 (O_913,N_14363,N_14898);
or UO_914 (O_914,N_14533,N_14477);
xor UO_915 (O_915,N_14936,N_14829);
nand UO_916 (O_916,N_14167,N_14756);
or UO_917 (O_917,N_14348,N_14936);
and UO_918 (O_918,N_14124,N_14452);
nor UO_919 (O_919,N_14482,N_14511);
nor UO_920 (O_920,N_14644,N_14475);
xor UO_921 (O_921,N_14797,N_14714);
nand UO_922 (O_922,N_14830,N_14784);
nor UO_923 (O_923,N_14230,N_14072);
nand UO_924 (O_924,N_14952,N_14611);
and UO_925 (O_925,N_14306,N_14578);
xor UO_926 (O_926,N_14678,N_14523);
and UO_927 (O_927,N_14901,N_14272);
and UO_928 (O_928,N_14519,N_14887);
nand UO_929 (O_929,N_14814,N_14158);
nand UO_930 (O_930,N_14387,N_14135);
or UO_931 (O_931,N_14386,N_14451);
nand UO_932 (O_932,N_14282,N_14996);
or UO_933 (O_933,N_14015,N_14896);
nand UO_934 (O_934,N_14701,N_14522);
or UO_935 (O_935,N_14222,N_14568);
and UO_936 (O_936,N_14831,N_14151);
xnor UO_937 (O_937,N_14187,N_14533);
xnor UO_938 (O_938,N_14794,N_14890);
and UO_939 (O_939,N_14811,N_14840);
nand UO_940 (O_940,N_14927,N_14218);
or UO_941 (O_941,N_14721,N_14757);
nor UO_942 (O_942,N_14884,N_14591);
and UO_943 (O_943,N_14231,N_14873);
or UO_944 (O_944,N_14887,N_14330);
nand UO_945 (O_945,N_14389,N_14289);
or UO_946 (O_946,N_14507,N_14047);
and UO_947 (O_947,N_14347,N_14632);
nand UO_948 (O_948,N_14300,N_14632);
or UO_949 (O_949,N_14795,N_14783);
nand UO_950 (O_950,N_14592,N_14805);
and UO_951 (O_951,N_14503,N_14681);
nand UO_952 (O_952,N_14070,N_14820);
xnor UO_953 (O_953,N_14030,N_14638);
nand UO_954 (O_954,N_14600,N_14412);
xor UO_955 (O_955,N_14629,N_14927);
nor UO_956 (O_956,N_14772,N_14709);
and UO_957 (O_957,N_14993,N_14346);
or UO_958 (O_958,N_14278,N_14237);
and UO_959 (O_959,N_14653,N_14866);
and UO_960 (O_960,N_14437,N_14294);
nand UO_961 (O_961,N_14907,N_14646);
nor UO_962 (O_962,N_14223,N_14111);
nor UO_963 (O_963,N_14834,N_14815);
and UO_964 (O_964,N_14600,N_14250);
or UO_965 (O_965,N_14202,N_14614);
or UO_966 (O_966,N_14227,N_14108);
and UO_967 (O_967,N_14722,N_14700);
or UO_968 (O_968,N_14120,N_14593);
nor UO_969 (O_969,N_14035,N_14747);
nand UO_970 (O_970,N_14566,N_14921);
or UO_971 (O_971,N_14351,N_14667);
or UO_972 (O_972,N_14408,N_14990);
and UO_973 (O_973,N_14263,N_14265);
nand UO_974 (O_974,N_14931,N_14558);
or UO_975 (O_975,N_14033,N_14392);
and UO_976 (O_976,N_14844,N_14782);
xor UO_977 (O_977,N_14892,N_14769);
or UO_978 (O_978,N_14939,N_14246);
or UO_979 (O_979,N_14202,N_14785);
nor UO_980 (O_980,N_14956,N_14150);
or UO_981 (O_981,N_14488,N_14652);
nor UO_982 (O_982,N_14193,N_14843);
xor UO_983 (O_983,N_14918,N_14593);
nor UO_984 (O_984,N_14446,N_14611);
and UO_985 (O_985,N_14134,N_14459);
nor UO_986 (O_986,N_14602,N_14455);
or UO_987 (O_987,N_14395,N_14968);
nand UO_988 (O_988,N_14043,N_14040);
or UO_989 (O_989,N_14688,N_14298);
nor UO_990 (O_990,N_14658,N_14698);
nor UO_991 (O_991,N_14535,N_14113);
nand UO_992 (O_992,N_14663,N_14151);
xnor UO_993 (O_993,N_14487,N_14414);
xor UO_994 (O_994,N_14225,N_14669);
or UO_995 (O_995,N_14645,N_14346);
or UO_996 (O_996,N_14222,N_14052);
xor UO_997 (O_997,N_14456,N_14163);
xnor UO_998 (O_998,N_14425,N_14314);
nor UO_999 (O_999,N_14991,N_14296);
xor UO_1000 (O_1000,N_14490,N_14478);
nor UO_1001 (O_1001,N_14605,N_14584);
nor UO_1002 (O_1002,N_14832,N_14057);
xnor UO_1003 (O_1003,N_14805,N_14818);
nand UO_1004 (O_1004,N_14605,N_14910);
or UO_1005 (O_1005,N_14625,N_14143);
nand UO_1006 (O_1006,N_14227,N_14583);
or UO_1007 (O_1007,N_14249,N_14963);
xnor UO_1008 (O_1008,N_14492,N_14813);
nor UO_1009 (O_1009,N_14703,N_14050);
nor UO_1010 (O_1010,N_14380,N_14929);
xnor UO_1011 (O_1011,N_14878,N_14066);
nand UO_1012 (O_1012,N_14290,N_14133);
and UO_1013 (O_1013,N_14622,N_14246);
or UO_1014 (O_1014,N_14619,N_14630);
xnor UO_1015 (O_1015,N_14025,N_14384);
nand UO_1016 (O_1016,N_14508,N_14724);
xnor UO_1017 (O_1017,N_14308,N_14442);
xor UO_1018 (O_1018,N_14143,N_14038);
and UO_1019 (O_1019,N_14060,N_14254);
nand UO_1020 (O_1020,N_14824,N_14082);
or UO_1021 (O_1021,N_14319,N_14283);
nand UO_1022 (O_1022,N_14264,N_14267);
nor UO_1023 (O_1023,N_14234,N_14096);
xor UO_1024 (O_1024,N_14279,N_14967);
nand UO_1025 (O_1025,N_14412,N_14944);
and UO_1026 (O_1026,N_14445,N_14428);
or UO_1027 (O_1027,N_14063,N_14236);
xnor UO_1028 (O_1028,N_14514,N_14269);
or UO_1029 (O_1029,N_14494,N_14386);
or UO_1030 (O_1030,N_14268,N_14393);
or UO_1031 (O_1031,N_14235,N_14838);
nor UO_1032 (O_1032,N_14874,N_14072);
and UO_1033 (O_1033,N_14155,N_14439);
and UO_1034 (O_1034,N_14533,N_14621);
or UO_1035 (O_1035,N_14607,N_14710);
and UO_1036 (O_1036,N_14686,N_14889);
nor UO_1037 (O_1037,N_14404,N_14928);
nand UO_1038 (O_1038,N_14304,N_14818);
nor UO_1039 (O_1039,N_14681,N_14424);
nand UO_1040 (O_1040,N_14064,N_14268);
and UO_1041 (O_1041,N_14298,N_14824);
nor UO_1042 (O_1042,N_14525,N_14433);
or UO_1043 (O_1043,N_14636,N_14411);
and UO_1044 (O_1044,N_14371,N_14361);
nor UO_1045 (O_1045,N_14665,N_14515);
xor UO_1046 (O_1046,N_14387,N_14125);
nor UO_1047 (O_1047,N_14918,N_14518);
and UO_1048 (O_1048,N_14926,N_14516);
xnor UO_1049 (O_1049,N_14079,N_14338);
or UO_1050 (O_1050,N_14062,N_14686);
and UO_1051 (O_1051,N_14628,N_14905);
nand UO_1052 (O_1052,N_14988,N_14960);
and UO_1053 (O_1053,N_14230,N_14351);
xor UO_1054 (O_1054,N_14681,N_14266);
nand UO_1055 (O_1055,N_14709,N_14435);
xor UO_1056 (O_1056,N_14463,N_14137);
nand UO_1057 (O_1057,N_14942,N_14420);
or UO_1058 (O_1058,N_14525,N_14830);
nor UO_1059 (O_1059,N_14931,N_14487);
xnor UO_1060 (O_1060,N_14738,N_14444);
and UO_1061 (O_1061,N_14950,N_14579);
nand UO_1062 (O_1062,N_14939,N_14985);
nand UO_1063 (O_1063,N_14100,N_14420);
and UO_1064 (O_1064,N_14362,N_14656);
and UO_1065 (O_1065,N_14745,N_14294);
or UO_1066 (O_1066,N_14359,N_14851);
and UO_1067 (O_1067,N_14320,N_14645);
nor UO_1068 (O_1068,N_14821,N_14531);
xnor UO_1069 (O_1069,N_14588,N_14721);
nand UO_1070 (O_1070,N_14984,N_14489);
and UO_1071 (O_1071,N_14519,N_14358);
xnor UO_1072 (O_1072,N_14815,N_14007);
and UO_1073 (O_1073,N_14285,N_14041);
or UO_1074 (O_1074,N_14542,N_14407);
and UO_1075 (O_1075,N_14019,N_14623);
nor UO_1076 (O_1076,N_14473,N_14898);
nor UO_1077 (O_1077,N_14160,N_14708);
nor UO_1078 (O_1078,N_14564,N_14240);
and UO_1079 (O_1079,N_14863,N_14129);
or UO_1080 (O_1080,N_14000,N_14723);
xor UO_1081 (O_1081,N_14722,N_14467);
nand UO_1082 (O_1082,N_14133,N_14618);
xor UO_1083 (O_1083,N_14607,N_14291);
and UO_1084 (O_1084,N_14622,N_14680);
nor UO_1085 (O_1085,N_14001,N_14281);
or UO_1086 (O_1086,N_14107,N_14857);
nor UO_1087 (O_1087,N_14911,N_14325);
nor UO_1088 (O_1088,N_14764,N_14265);
nand UO_1089 (O_1089,N_14703,N_14406);
nand UO_1090 (O_1090,N_14490,N_14768);
nand UO_1091 (O_1091,N_14303,N_14999);
nor UO_1092 (O_1092,N_14116,N_14794);
nand UO_1093 (O_1093,N_14354,N_14431);
xor UO_1094 (O_1094,N_14041,N_14826);
nor UO_1095 (O_1095,N_14202,N_14011);
nand UO_1096 (O_1096,N_14921,N_14297);
nand UO_1097 (O_1097,N_14488,N_14566);
nor UO_1098 (O_1098,N_14742,N_14100);
or UO_1099 (O_1099,N_14247,N_14676);
and UO_1100 (O_1100,N_14493,N_14445);
and UO_1101 (O_1101,N_14796,N_14259);
xnor UO_1102 (O_1102,N_14929,N_14053);
and UO_1103 (O_1103,N_14756,N_14223);
nand UO_1104 (O_1104,N_14355,N_14913);
and UO_1105 (O_1105,N_14852,N_14660);
and UO_1106 (O_1106,N_14444,N_14815);
nand UO_1107 (O_1107,N_14788,N_14089);
xor UO_1108 (O_1108,N_14932,N_14565);
nor UO_1109 (O_1109,N_14990,N_14717);
nor UO_1110 (O_1110,N_14155,N_14138);
nand UO_1111 (O_1111,N_14960,N_14742);
or UO_1112 (O_1112,N_14992,N_14952);
nand UO_1113 (O_1113,N_14486,N_14915);
xor UO_1114 (O_1114,N_14720,N_14386);
nor UO_1115 (O_1115,N_14763,N_14315);
xor UO_1116 (O_1116,N_14582,N_14721);
xor UO_1117 (O_1117,N_14235,N_14553);
nor UO_1118 (O_1118,N_14465,N_14862);
xnor UO_1119 (O_1119,N_14686,N_14176);
nor UO_1120 (O_1120,N_14921,N_14825);
xor UO_1121 (O_1121,N_14194,N_14917);
and UO_1122 (O_1122,N_14138,N_14964);
or UO_1123 (O_1123,N_14836,N_14842);
and UO_1124 (O_1124,N_14881,N_14755);
or UO_1125 (O_1125,N_14003,N_14527);
nand UO_1126 (O_1126,N_14939,N_14823);
or UO_1127 (O_1127,N_14821,N_14067);
nand UO_1128 (O_1128,N_14811,N_14587);
xnor UO_1129 (O_1129,N_14694,N_14906);
nand UO_1130 (O_1130,N_14124,N_14931);
and UO_1131 (O_1131,N_14990,N_14388);
or UO_1132 (O_1132,N_14540,N_14101);
nor UO_1133 (O_1133,N_14908,N_14408);
and UO_1134 (O_1134,N_14231,N_14266);
nor UO_1135 (O_1135,N_14882,N_14267);
or UO_1136 (O_1136,N_14243,N_14418);
xor UO_1137 (O_1137,N_14810,N_14755);
xnor UO_1138 (O_1138,N_14195,N_14943);
xor UO_1139 (O_1139,N_14195,N_14928);
nand UO_1140 (O_1140,N_14143,N_14830);
or UO_1141 (O_1141,N_14415,N_14426);
and UO_1142 (O_1142,N_14227,N_14497);
nor UO_1143 (O_1143,N_14665,N_14813);
nand UO_1144 (O_1144,N_14384,N_14715);
or UO_1145 (O_1145,N_14041,N_14913);
nor UO_1146 (O_1146,N_14543,N_14782);
and UO_1147 (O_1147,N_14960,N_14843);
xor UO_1148 (O_1148,N_14620,N_14074);
and UO_1149 (O_1149,N_14719,N_14055);
or UO_1150 (O_1150,N_14556,N_14902);
nor UO_1151 (O_1151,N_14656,N_14910);
nand UO_1152 (O_1152,N_14039,N_14080);
and UO_1153 (O_1153,N_14419,N_14187);
and UO_1154 (O_1154,N_14852,N_14183);
xor UO_1155 (O_1155,N_14906,N_14484);
nand UO_1156 (O_1156,N_14390,N_14756);
nor UO_1157 (O_1157,N_14232,N_14356);
nand UO_1158 (O_1158,N_14628,N_14124);
nor UO_1159 (O_1159,N_14217,N_14704);
nand UO_1160 (O_1160,N_14628,N_14862);
xnor UO_1161 (O_1161,N_14884,N_14955);
and UO_1162 (O_1162,N_14959,N_14528);
nor UO_1163 (O_1163,N_14365,N_14478);
and UO_1164 (O_1164,N_14614,N_14531);
and UO_1165 (O_1165,N_14259,N_14539);
nand UO_1166 (O_1166,N_14377,N_14457);
nor UO_1167 (O_1167,N_14663,N_14493);
and UO_1168 (O_1168,N_14113,N_14863);
nor UO_1169 (O_1169,N_14531,N_14526);
nand UO_1170 (O_1170,N_14003,N_14370);
and UO_1171 (O_1171,N_14445,N_14491);
nor UO_1172 (O_1172,N_14966,N_14882);
xor UO_1173 (O_1173,N_14414,N_14592);
or UO_1174 (O_1174,N_14192,N_14147);
xor UO_1175 (O_1175,N_14260,N_14309);
or UO_1176 (O_1176,N_14655,N_14730);
nand UO_1177 (O_1177,N_14734,N_14473);
xnor UO_1178 (O_1178,N_14960,N_14974);
and UO_1179 (O_1179,N_14495,N_14661);
nand UO_1180 (O_1180,N_14838,N_14632);
nand UO_1181 (O_1181,N_14429,N_14336);
nor UO_1182 (O_1182,N_14396,N_14791);
nand UO_1183 (O_1183,N_14315,N_14629);
nand UO_1184 (O_1184,N_14570,N_14883);
and UO_1185 (O_1185,N_14662,N_14821);
nand UO_1186 (O_1186,N_14814,N_14134);
xnor UO_1187 (O_1187,N_14143,N_14631);
nor UO_1188 (O_1188,N_14808,N_14467);
nor UO_1189 (O_1189,N_14786,N_14930);
nand UO_1190 (O_1190,N_14320,N_14964);
nand UO_1191 (O_1191,N_14910,N_14564);
xor UO_1192 (O_1192,N_14652,N_14154);
or UO_1193 (O_1193,N_14475,N_14972);
nor UO_1194 (O_1194,N_14315,N_14612);
nor UO_1195 (O_1195,N_14987,N_14708);
or UO_1196 (O_1196,N_14286,N_14851);
and UO_1197 (O_1197,N_14385,N_14095);
and UO_1198 (O_1198,N_14296,N_14200);
nor UO_1199 (O_1199,N_14334,N_14830);
and UO_1200 (O_1200,N_14486,N_14224);
nand UO_1201 (O_1201,N_14691,N_14121);
or UO_1202 (O_1202,N_14921,N_14685);
nand UO_1203 (O_1203,N_14543,N_14652);
and UO_1204 (O_1204,N_14479,N_14793);
and UO_1205 (O_1205,N_14222,N_14413);
xor UO_1206 (O_1206,N_14324,N_14802);
xor UO_1207 (O_1207,N_14204,N_14799);
and UO_1208 (O_1208,N_14752,N_14026);
xnor UO_1209 (O_1209,N_14332,N_14772);
xnor UO_1210 (O_1210,N_14475,N_14649);
or UO_1211 (O_1211,N_14360,N_14230);
nor UO_1212 (O_1212,N_14547,N_14287);
or UO_1213 (O_1213,N_14382,N_14789);
xor UO_1214 (O_1214,N_14766,N_14268);
or UO_1215 (O_1215,N_14104,N_14968);
nand UO_1216 (O_1216,N_14541,N_14516);
and UO_1217 (O_1217,N_14834,N_14654);
or UO_1218 (O_1218,N_14814,N_14100);
nand UO_1219 (O_1219,N_14879,N_14024);
or UO_1220 (O_1220,N_14149,N_14468);
nor UO_1221 (O_1221,N_14299,N_14035);
or UO_1222 (O_1222,N_14815,N_14405);
and UO_1223 (O_1223,N_14969,N_14868);
nand UO_1224 (O_1224,N_14321,N_14268);
xnor UO_1225 (O_1225,N_14137,N_14640);
nor UO_1226 (O_1226,N_14797,N_14383);
nor UO_1227 (O_1227,N_14188,N_14032);
xor UO_1228 (O_1228,N_14809,N_14689);
xor UO_1229 (O_1229,N_14573,N_14713);
xnor UO_1230 (O_1230,N_14043,N_14583);
or UO_1231 (O_1231,N_14051,N_14585);
nor UO_1232 (O_1232,N_14469,N_14765);
nor UO_1233 (O_1233,N_14893,N_14334);
and UO_1234 (O_1234,N_14266,N_14161);
nand UO_1235 (O_1235,N_14723,N_14625);
nor UO_1236 (O_1236,N_14740,N_14214);
and UO_1237 (O_1237,N_14152,N_14111);
xnor UO_1238 (O_1238,N_14765,N_14680);
and UO_1239 (O_1239,N_14380,N_14675);
nand UO_1240 (O_1240,N_14062,N_14497);
xor UO_1241 (O_1241,N_14601,N_14964);
and UO_1242 (O_1242,N_14821,N_14920);
nor UO_1243 (O_1243,N_14237,N_14972);
nand UO_1244 (O_1244,N_14095,N_14809);
and UO_1245 (O_1245,N_14651,N_14592);
or UO_1246 (O_1246,N_14422,N_14574);
nor UO_1247 (O_1247,N_14232,N_14517);
and UO_1248 (O_1248,N_14066,N_14204);
nor UO_1249 (O_1249,N_14239,N_14401);
or UO_1250 (O_1250,N_14336,N_14937);
nand UO_1251 (O_1251,N_14314,N_14828);
xnor UO_1252 (O_1252,N_14558,N_14408);
or UO_1253 (O_1253,N_14849,N_14464);
xor UO_1254 (O_1254,N_14717,N_14450);
and UO_1255 (O_1255,N_14844,N_14152);
or UO_1256 (O_1256,N_14409,N_14876);
or UO_1257 (O_1257,N_14812,N_14622);
nand UO_1258 (O_1258,N_14529,N_14955);
nand UO_1259 (O_1259,N_14996,N_14032);
or UO_1260 (O_1260,N_14735,N_14768);
or UO_1261 (O_1261,N_14902,N_14154);
xor UO_1262 (O_1262,N_14748,N_14181);
or UO_1263 (O_1263,N_14461,N_14636);
nor UO_1264 (O_1264,N_14958,N_14076);
nor UO_1265 (O_1265,N_14161,N_14281);
nor UO_1266 (O_1266,N_14250,N_14341);
nand UO_1267 (O_1267,N_14760,N_14736);
or UO_1268 (O_1268,N_14618,N_14066);
nand UO_1269 (O_1269,N_14804,N_14838);
nor UO_1270 (O_1270,N_14011,N_14504);
nand UO_1271 (O_1271,N_14890,N_14668);
xor UO_1272 (O_1272,N_14489,N_14351);
nor UO_1273 (O_1273,N_14551,N_14238);
nand UO_1274 (O_1274,N_14374,N_14994);
and UO_1275 (O_1275,N_14729,N_14228);
xor UO_1276 (O_1276,N_14025,N_14104);
xnor UO_1277 (O_1277,N_14574,N_14083);
xor UO_1278 (O_1278,N_14314,N_14871);
nand UO_1279 (O_1279,N_14286,N_14332);
nor UO_1280 (O_1280,N_14317,N_14741);
nand UO_1281 (O_1281,N_14277,N_14000);
nand UO_1282 (O_1282,N_14977,N_14696);
nand UO_1283 (O_1283,N_14768,N_14744);
and UO_1284 (O_1284,N_14721,N_14832);
and UO_1285 (O_1285,N_14568,N_14705);
xnor UO_1286 (O_1286,N_14712,N_14264);
xnor UO_1287 (O_1287,N_14748,N_14962);
and UO_1288 (O_1288,N_14388,N_14732);
and UO_1289 (O_1289,N_14269,N_14781);
nand UO_1290 (O_1290,N_14410,N_14666);
and UO_1291 (O_1291,N_14959,N_14925);
and UO_1292 (O_1292,N_14443,N_14848);
nor UO_1293 (O_1293,N_14094,N_14979);
and UO_1294 (O_1294,N_14815,N_14732);
or UO_1295 (O_1295,N_14388,N_14702);
or UO_1296 (O_1296,N_14361,N_14909);
nand UO_1297 (O_1297,N_14208,N_14892);
xor UO_1298 (O_1298,N_14905,N_14493);
and UO_1299 (O_1299,N_14616,N_14145);
and UO_1300 (O_1300,N_14076,N_14354);
xnor UO_1301 (O_1301,N_14479,N_14911);
or UO_1302 (O_1302,N_14122,N_14248);
nand UO_1303 (O_1303,N_14204,N_14187);
nand UO_1304 (O_1304,N_14103,N_14210);
and UO_1305 (O_1305,N_14986,N_14914);
or UO_1306 (O_1306,N_14752,N_14819);
or UO_1307 (O_1307,N_14356,N_14434);
and UO_1308 (O_1308,N_14003,N_14020);
nor UO_1309 (O_1309,N_14988,N_14156);
or UO_1310 (O_1310,N_14345,N_14027);
xnor UO_1311 (O_1311,N_14406,N_14552);
nand UO_1312 (O_1312,N_14115,N_14065);
nand UO_1313 (O_1313,N_14596,N_14654);
and UO_1314 (O_1314,N_14750,N_14167);
nor UO_1315 (O_1315,N_14958,N_14862);
xor UO_1316 (O_1316,N_14263,N_14849);
xor UO_1317 (O_1317,N_14338,N_14145);
xnor UO_1318 (O_1318,N_14699,N_14385);
xor UO_1319 (O_1319,N_14551,N_14575);
nand UO_1320 (O_1320,N_14862,N_14449);
and UO_1321 (O_1321,N_14700,N_14046);
or UO_1322 (O_1322,N_14892,N_14653);
nand UO_1323 (O_1323,N_14378,N_14635);
nand UO_1324 (O_1324,N_14171,N_14481);
xnor UO_1325 (O_1325,N_14065,N_14108);
nand UO_1326 (O_1326,N_14536,N_14703);
nand UO_1327 (O_1327,N_14598,N_14320);
xnor UO_1328 (O_1328,N_14266,N_14041);
xnor UO_1329 (O_1329,N_14123,N_14638);
and UO_1330 (O_1330,N_14345,N_14223);
and UO_1331 (O_1331,N_14813,N_14823);
or UO_1332 (O_1332,N_14224,N_14918);
xor UO_1333 (O_1333,N_14794,N_14166);
nor UO_1334 (O_1334,N_14126,N_14048);
nand UO_1335 (O_1335,N_14743,N_14889);
or UO_1336 (O_1336,N_14089,N_14910);
nor UO_1337 (O_1337,N_14533,N_14769);
nand UO_1338 (O_1338,N_14768,N_14310);
and UO_1339 (O_1339,N_14844,N_14879);
nor UO_1340 (O_1340,N_14961,N_14587);
nand UO_1341 (O_1341,N_14432,N_14947);
nand UO_1342 (O_1342,N_14031,N_14293);
or UO_1343 (O_1343,N_14333,N_14340);
nor UO_1344 (O_1344,N_14844,N_14768);
or UO_1345 (O_1345,N_14564,N_14920);
nand UO_1346 (O_1346,N_14488,N_14989);
or UO_1347 (O_1347,N_14642,N_14949);
xnor UO_1348 (O_1348,N_14148,N_14362);
xor UO_1349 (O_1349,N_14964,N_14532);
xnor UO_1350 (O_1350,N_14639,N_14260);
or UO_1351 (O_1351,N_14410,N_14356);
nand UO_1352 (O_1352,N_14386,N_14752);
and UO_1353 (O_1353,N_14100,N_14407);
xor UO_1354 (O_1354,N_14569,N_14197);
nor UO_1355 (O_1355,N_14977,N_14883);
or UO_1356 (O_1356,N_14387,N_14472);
xnor UO_1357 (O_1357,N_14584,N_14887);
nor UO_1358 (O_1358,N_14893,N_14756);
and UO_1359 (O_1359,N_14314,N_14030);
nand UO_1360 (O_1360,N_14113,N_14345);
xor UO_1361 (O_1361,N_14250,N_14657);
nor UO_1362 (O_1362,N_14279,N_14356);
and UO_1363 (O_1363,N_14942,N_14341);
and UO_1364 (O_1364,N_14812,N_14594);
xor UO_1365 (O_1365,N_14544,N_14506);
and UO_1366 (O_1366,N_14897,N_14997);
and UO_1367 (O_1367,N_14243,N_14901);
and UO_1368 (O_1368,N_14093,N_14455);
nand UO_1369 (O_1369,N_14855,N_14930);
nor UO_1370 (O_1370,N_14245,N_14241);
nand UO_1371 (O_1371,N_14298,N_14862);
and UO_1372 (O_1372,N_14698,N_14517);
xnor UO_1373 (O_1373,N_14693,N_14678);
nor UO_1374 (O_1374,N_14709,N_14246);
nand UO_1375 (O_1375,N_14060,N_14858);
nor UO_1376 (O_1376,N_14593,N_14533);
nor UO_1377 (O_1377,N_14777,N_14779);
nor UO_1378 (O_1378,N_14858,N_14116);
or UO_1379 (O_1379,N_14982,N_14179);
or UO_1380 (O_1380,N_14673,N_14691);
nor UO_1381 (O_1381,N_14760,N_14065);
nor UO_1382 (O_1382,N_14666,N_14951);
or UO_1383 (O_1383,N_14375,N_14607);
nor UO_1384 (O_1384,N_14143,N_14412);
nor UO_1385 (O_1385,N_14166,N_14694);
or UO_1386 (O_1386,N_14861,N_14614);
xnor UO_1387 (O_1387,N_14377,N_14236);
and UO_1388 (O_1388,N_14780,N_14539);
nand UO_1389 (O_1389,N_14597,N_14419);
nand UO_1390 (O_1390,N_14869,N_14710);
nor UO_1391 (O_1391,N_14396,N_14501);
nand UO_1392 (O_1392,N_14063,N_14755);
nor UO_1393 (O_1393,N_14825,N_14401);
nand UO_1394 (O_1394,N_14263,N_14315);
and UO_1395 (O_1395,N_14526,N_14923);
nor UO_1396 (O_1396,N_14999,N_14809);
or UO_1397 (O_1397,N_14919,N_14131);
nand UO_1398 (O_1398,N_14521,N_14390);
nor UO_1399 (O_1399,N_14452,N_14278);
and UO_1400 (O_1400,N_14756,N_14178);
nand UO_1401 (O_1401,N_14976,N_14546);
xor UO_1402 (O_1402,N_14782,N_14713);
nand UO_1403 (O_1403,N_14146,N_14974);
and UO_1404 (O_1404,N_14126,N_14222);
xor UO_1405 (O_1405,N_14736,N_14085);
nand UO_1406 (O_1406,N_14901,N_14779);
or UO_1407 (O_1407,N_14997,N_14330);
nor UO_1408 (O_1408,N_14286,N_14092);
nor UO_1409 (O_1409,N_14069,N_14595);
nor UO_1410 (O_1410,N_14068,N_14755);
nand UO_1411 (O_1411,N_14943,N_14664);
nor UO_1412 (O_1412,N_14472,N_14881);
nand UO_1413 (O_1413,N_14300,N_14502);
nor UO_1414 (O_1414,N_14283,N_14703);
xor UO_1415 (O_1415,N_14343,N_14566);
or UO_1416 (O_1416,N_14550,N_14392);
or UO_1417 (O_1417,N_14400,N_14349);
nor UO_1418 (O_1418,N_14735,N_14140);
nand UO_1419 (O_1419,N_14044,N_14486);
and UO_1420 (O_1420,N_14659,N_14183);
xor UO_1421 (O_1421,N_14629,N_14044);
nor UO_1422 (O_1422,N_14226,N_14570);
nor UO_1423 (O_1423,N_14348,N_14447);
xor UO_1424 (O_1424,N_14042,N_14238);
or UO_1425 (O_1425,N_14955,N_14252);
nand UO_1426 (O_1426,N_14128,N_14036);
xor UO_1427 (O_1427,N_14434,N_14404);
nor UO_1428 (O_1428,N_14240,N_14650);
nor UO_1429 (O_1429,N_14524,N_14560);
nor UO_1430 (O_1430,N_14690,N_14475);
xnor UO_1431 (O_1431,N_14031,N_14795);
and UO_1432 (O_1432,N_14759,N_14765);
nand UO_1433 (O_1433,N_14247,N_14275);
nor UO_1434 (O_1434,N_14952,N_14318);
nand UO_1435 (O_1435,N_14316,N_14364);
nor UO_1436 (O_1436,N_14275,N_14308);
xor UO_1437 (O_1437,N_14251,N_14592);
nand UO_1438 (O_1438,N_14042,N_14793);
nand UO_1439 (O_1439,N_14867,N_14939);
xnor UO_1440 (O_1440,N_14867,N_14234);
or UO_1441 (O_1441,N_14036,N_14972);
or UO_1442 (O_1442,N_14414,N_14434);
or UO_1443 (O_1443,N_14173,N_14833);
nor UO_1444 (O_1444,N_14423,N_14673);
nand UO_1445 (O_1445,N_14842,N_14528);
nor UO_1446 (O_1446,N_14518,N_14013);
nor UO_1447 (O_1447,N_14155,N_14010);
nor UO_1448 (O_1448,N_14228,N_14689);
and UO_1449 (O_1449,N_14880,N_14834);
and UO_1450 (O_1450,N_14812,N_14741);
or UO_1451 (O_1451,N_14051,N_14974);
and UO_1452 (O_1452,N_14967,N_14260);
nand UO_1453 (O_1453,N_14607,N_14406);
xor UO_1454 (O_1454,N_14617,N_14771);
xnor UO_1455 (O_1455,N_14641,N_14924);
and UO_1456 (O_1456,N_14077,N_14202);
nor UO_1457 (O_1457,N_14759,N_14928);
nand UO_1458 (O_1458,N_14167,N_14718);
xnor UO_1459 (O_1459,N_14341,N_14100);
nor UO_1460 (O_1460,N_14863,N_14258);
and UO_1461 (O_1461,N_14143,N_14951);
nor UO_1462 (O_1462,N_14536,N_14521);
xnor UO_1463 (O_1463,N_14153,N_14711);
nand UO_1464 (O_1464,N_14526,N_14387);
nor UO_1465 (O_1465,N_14026,N_14015);
and UO_1466 (O_1466,N_14578,N_14823);
nor UO_1467 (O_1467,N_14290,N_14245);
xnor UO_1468 (O_1468,N_14931,N_14726);
xnor UO_1469 (O_1469,N_14461,N_14964);
or UO_1470 (O_1470,N_14494,N_14447);
or UO_1471 (O_1471,N_14505,N_14999);
or UO_1472 (O_1472,N_14279,N_14595);
nand UO_1473 (O_1473,N_14352,N_14270);
xnor UO_1474 (O_1474,N_14852,N_14879);
nor UO_1475 (O_1475,N_14296,N_14695);
and UO_1476 (O_1476,N_14302,N_14725);
nor UO_1477 (O_1477,N_14715,N_14999);
and UO_1478 (O_1478,N_14211,N_14131);
nand UO_1479 (O_1479,N_14999,N_14883);
nor UO_1480 (O_1480,N_14689,N_14433);
and UO_1481 (O_1481,N_14557,N_14500);
and UO_1482 (O_1482,N_14061,N_14711);
xnor UO_1483 (O_1483,N_14048,N_14762);
or UO_1484 (O_1484,N_14998,N_14899);
and UO_1485 (O_1485,N_14863,N_14204);
nor UO_1486 (O_1486,N_14112,N_14007);
and UO_1487 (O_1487,N_14911,N_14319);
and UO_1488 (O_1488,N_14297,N_14049);
nand UO_1489 (O_1489,N_14335,N_14578);
nor UO_1490 (O_1490,N_14103,N_14955);
and UO_1491 (O_1491,N_14208,N_14145);
nand UO_1492 (O_1492,N_14433,N_14415);
nand UO_1493 (O_1493,N_14481,N_14104);
or UO_1494 (O_1494,N_14572,N_14552);
nand UO_1495 (O_1495,N_14850,N_14360);
or UO_1496 (O_1496,N_14574,N_14240);
nand UO_1497 (O_1497,N_14660,N_14721);
and UO_1498 (O_1498,N_14894,N_14081);
nand UO_1499 (O_1499,N_14138,N_14340);
or UO_1500 (O_1500,N_14730,N_14524);
or UO_1501 (O_1501,N_14823,N_14222);
nand UO_1502 (O_1502,N_14599,N_14079);
nand UO_1503 (O_1503,N_14815,N_14546);
or UO_1504 (O_1504,N_14424,N_14257);
nand UO_1505 (O_1505,N_14103,N_14741);
xnor UO_1506 (O_1506,N_14951,N_14207);
xnor UO_1507 (O_1507,N_14213,N_14580);
nand UO_1508 (O_1508,N_14640,N_14317);
and UO_1509 (O_1509,N_14871,N_14219);
and UO_1510 (O_1510,N_14232,N_14348);
xor UO_1511 (O_1511,N_14677,N_14580);
nand UO_1512 (O_1512,N_14967,N_14492);
or UO_1513 (O_1513,N_14570,N_14154);
nand UO_1514 (O_1514,N_14140,N_14657);
nand UO_1515 (O_1515,N_14842,N_14953);
xnor UO_1516 (O_1516,N_14734,N_14002);
or UO_1517 (O_1517,N_14358,N_14720);
nand UO_1518 (O_1518,N_14051,N_14003);
nand UO_1519 (O_1519,N_14522,N_14975);
or UO_1520 (O_1520,N_14605,N_14176);
and UO_1521 (O_1521,N_14858,N_14134);
nand UO_1522 (O_1522,N_14785,N_14773);
nand UO_1523 (O_1523,N_14617,N_14211);
nand UO_1524 (O_1524,N_14051,N_14423);
xor UO_1525 (O_1525,N_14000,N_14309);
xor UO_1526 (O_1526,N_14190,N_14421);
and UO_1527 (O_1527,N_14371,N_14761);
or UO_1528 (O_1528,N_14149,N_14647);
nand UO_1529 (O_1529,N_14861,N_14180);
nand UO_1530 (O_1530,N_14652,N_14776);
nand UO_1531 (O_1531,N_14137,N_14832);
and UO_1532 (O_1532,N_14955,N_14473);
or UO_1533 (O_1533,N_14864,N_14560);
nand UO_1534 (O_1534,N_14177,N_14655);
nand UO_1535 (O_1535,N_14503,N_14963);
nor UO_1536 (O_1536,N_14318,N_14649);
nand UO_1537 (O_1537,N_14203,N_14506);
and UO_1538 (O_1538,N_14254,N_14556);
or UO_1539 (O_1539,N_14236,N_14093);
xor UO_1540 (O_1540,N_14086,N_14540);
and UO_1541 (O_1541,N_14872,N_14809);
xnor UO_1542 (O_1542,N_14348,N_14592);
xnor UO_1543 (O_1543,N_14398,N_14051);
or UO_1544 (O_1544,N_14423,N_14311);
nand UO_1545 (O_1545,N_14847,N_14248);
and UO_1546 (O_1546,N_14132,N_14564);
or UO_1547 (O_1547,N_14592,N_14032);
or UO_1548 (O_1548,N_14693,N_14559);
or UO_1549 (O_1549,N_14229,N_14814);
xor UO_1550 (O_1550,N_14924,N_14129);
xnor UO_1551 (O_1551,N_14715,N_14149);
xor UO_1552 (O_1552,N_14857,N_14202);
nand UO_1553 (O_1553,N_14492,N_14809);
nor UO_1554 (O_1554,N_14170,N_14014);
or UO_1555 (O_1555,N_14278,N_14315);
nor UO_1556 (O_1556,N_14538,N_14882);
nor UO_1557 (O_1557,N_14243,N_14344);
nor UO_1558 (O_1558,N_14773,N_14481);
and UO_1559 (O_1559,N_14334,N_14624);
nand UO_1560 (O_1560,N_14986,N_14465);
or UO_1561 (O_1561,N_14049,N_14376);
and UO_1562 (O_1562,N_14803,N_14328);
and UO_1563 (O_1563,N_14515,N_14593);
xnor UO_1564 (O_1564,N_14191,N_14849);
and UO_1565 (O_1565,N_14067,N_14338);
and UO_1566 (O_1566,N_14185,N_14175);
or UO_1567 (O_1567,N_14655,N_14749);
nor UO_1568 (O_1568,N_14058,N_14936);
nor UO_1569 (O_1569,N_14355,N_14912);
and UO_1570 (O_1570,N_14554,N_14484);
or UO_1571 (O_1571,N_14877,N_14289);
or UO_1572 (O_1572,N_14715,N_14702);
nand UO_1573 (O_1573,N_14504,N_14646);
or UO_1574 (O_1574,N_14963,N_14953);
nand UO_1575 (O_1575,N_14556,N_14299);
nand UO_1576 (O_1576,N_14587,N_14160);
nor UO_1577 (O_1577,N_14977,N_14329);
and UO_1578 (O_1578,N_14809,N_14232);
nor UO_1579 (O_1579,N_14909,N_14563);
nor UO_1580 (O_1580,N_14399,N_14572);
nor UO_1581 (O_1581,N_14851,N_14123);
nor UO_1582 (O_1582,N_14770,N_14178);
nand UO_1583 (O_1583,N_14015,N_14992);
nor UO_1584 (O_1584,N_14877,N_14119);
nor UO_1585 (O_1585,N_14315,N_14054);
and UO_1586 (O_1586,N_14143,N_14334);
nor UO_1587 (O_1587,N_14137,N_14278);
or UO_1588 (O_1588,N_14527,N_14484);
nor UO_1589 (O_1589,N_14089,N_14964);
and UO_1590 (O_1590,N_14288,N_14521);
nor UO_1591 (O_1591,N_14277,N_14076);
nor UO_1592 (O_1592,N_14062,N_14483);
or UO_1593 (O_1593,N_14183,N_14843);
nand UO_1594 (O_1594,N_14020,N_14213);
xnor UO_1595 (O_1595,N_14798,N_14821);
nand UO_1596 (O_1596,N_14379,N_14458);
nor UO_1597 (O_1597,N_14978,N_14273);
or UO_1598 (O_1598,N_14772,N_14724);
xnor UO_1599 (O_1599,N_14295,N_14533);
or UO_1600 (O_1600,N_14038,N_14906);
or UO_1601 (O_1601,N_14963,N_14295);
nor UO_1602 (O_1602,N_14295,N_14892);
nor UO_1603 (O_1603,N_14104,N_14558);
nor UO_1604 (O_1604,N_14019,N_14047);
nor UO_1605 (O_1605,N_14495,N_14902);
and UO_1606 (O_1606,N_14419,N_14732);
and UO_1607 (O_1607,N_14842,N_14219);
or UO_1608 (O_1608,N_14622,N_14112);
or UO_1609 (O_1609,N_14496,N_14308);
xor UO_1610 (O_1610,N_14700,N_14882);
or UO_1611 (O_1611,N_14108,N_14641);
and UO_1612 (O_1612,N_14792,N_14271);
and UO_1613 (O_1613,N_14313,N_14417);
or UO_1614 (O_1614,N_14633,N_14567);
nor UO_1615 (O_1615,N_14950,N_14972);
xnor UO_1616 (O_1616,N_14066,N_14666);
and UO_1617 (O_1617,N_14404,N_14570);
nor UO_1618 (O_1618,N_14566,N_14163);
nand UO_1619 (O_1619,N_14312,N_14932);
or UO_1620 (O_1620,N_14757,N_14801);
nor UO_1621 (O_1621,N_14492,N_14346);
or UO_1622 (O_1622,N_14535,N_14041);
and UO_1623 (O_1623,N_14205,N_14905);
or UO_1624 (O_1624,N_14036,N_14378);
nor UO_1625 (O_1625,N_14583,N_14474);
nor UO_1626 (O_1626,N_14434,N_14797);
or UO_1627 (O_1627,N_14390,N_14356);
and UO_1628 (O_1628,N_14342,N_14458);
xnor UO_1629 (O_1629,N_14530,N_14731);
or UO_1630 (O_1630,N_14695,N_14674);
xnor UO_1631 (O_1631,N_14033,N_14068);
nor UO_1632 (O_1632,N_14036,N_14376);
or UO_1633 (O_1633,N_14720,N_14182);
xnor UO_1634 (O_1634,N_14337,N_14490);
xnor UO_1635 (O_1635,N_14870,N_14003);
nand UO_1636 (O_1636,N_14752,N_14231);
or UO_1637 (O_1637,N_14292,N_14310);
xor UO_1638 (O_1638,N_14967,N_14555);
xnor UO_1639 (O_1639,N_14285,N_14512);
or UO_1640 (O_1640,N_14356,N_14732);
nand UO_1641 (O_1641,N_14314,N_14034);
nand UO_1642 (O_1642,N_14607,N_14717);
or UO_1643 (O_1643,N_14438,N_14782);
nand UO_1644 (O_1644,N_14348,N_14524);
nor UO_1645 (O_1645,N_14894,N_14171);
or UO_1646 (O_1646,N_14578,N_14395);
nand UO_1647 (O_1647,N_14511,N_14942);
nand UO_1648 (O_1648,N_14434,N_14660);
nor UO_1649 (O_1649,N_14374,N_14937);
nor UO_1650 (O_1650,N_14960,N_14700);
nor UO_1651 (O_1651,N_14776,N_14274);
xnor UO_1652 (O_1652,N_14110,N_14635);
nor UO_1653 (O_1653,N_14216,N_14782);
nor UO_1654 (O_1654,N_14656,N_14206);
or UO_1655 (O_1655,N_14703,N_14594);
nand UO_1656 (O_1656,N_14195,N_14499);
nor UO_1657 (O_1657,N_14384,N_14939);
and UO_1658 (O_1658,N_14427,N_14262);
nor UO_1659 (O_1659,N_14998,N_14116);
or UO_1660 (O_1660,N_14552,N_14429);
nor UO_1661 (O_1661,N_14418,N_14401);
nor UO_1662 (O_1662,N_14054,N_14767);
xor UO_1663 (O_1663,N_14974,N_14847);
xnor UO_1664 (O_1664,N_14296,N_14230);
or UO_1665 (O_1665,N_14495,N_14950);
xnor UO_1666 (O_1666,N_14215,N_14331);
xor UO_1667 (O_1667,N_14628,N_14804);
nor UO_1668 (O_1668,N_14779,N_14538);
and UO_1669 (O_1669,N_14478,N_14831);
nand UO_1670 (O_1670,N_14251,N_14503);
or UO_1671 (O_1671,N_14388,N_14798);
and UO_1672 (O_1672,N_14335,N_14857);
nand UO_1673 (O_1673,N_14883,N_14598);
xor UO_1674 (O_1674,N_14897,N_14726);
nand UO_1675 (O_1675,N_14859,N_14865);
xor UO_1676 (O_1676,N_14168,N_14708);
and UO_1677 (O_1677,N_14293,N_14185);
nand UO_1678 (O_1678,N_14891,N_14213);
and UO_1679 (O_1679,N_14925,N_14559);
and UO_1680 (O_1680,N_14257,N_14898);
and UO_1681 (O_1681,N_14920,N_14859);
nor UO_1682 (O_1682,N_14060,N_14083);
or UO_1683 (O_1683,N_14582,N_14294);
and UO_1684 (O_1684,N_14792,N_14807);
or UO_1685 (O_1685,N_14535,N_14204);
or UO_1686 (O_1686,N_14545,N_14884);
nor UO_1687 (O_1687,N_14523,N_14969);
or UO_1688 (O_1688,N_14796,N_14517);
and UO_1689 (O_1689,N_14680,N_14595);
nor UO_1690 (O_1690,N_14908,N_14189);
nor UO_1691 (O_1691,N_14211,N_14679);
nand UO_1692 (O_1692,N_14589,N_14860);
xor UO_1693 (O_1693,N_14782,N_14382);
xor UO_1694 (O_1694,N_14203,N_14488);
or UO_1695 (O_1695,N_14089,N_14997);
nand UO_1696 (O_1696,N_14301,N_14726);
nor UO_1697 (O_1697,N_14205,N_14146);
xnor UO_1698 (O_1698,N_14231,N_14317);
and UO_1699 (O_1699,N_14832,N_14541);
nor UO_1700 (O_1700,N_14224,N_14346);
nand UO_1701 (O_1701,N_14737,N_14170);
nand UO_1702 (O_1702,N_14213,N_14354);
xor UO_1703 (O_1703,N_14296,N_14585);
nor UO_1704 (O_1704,N_14662,N_14650);
nor UO_1705 (O_1705,N_14626,N_14643);
nand UO_1706 (O_1706,N_14807,N_14361);
nand UO_1707 (O_1707,N_14535,N_14328);
and UO_1708 (O_1708,N_14165,N_14968);
or UO_1709 (O_1709,N_14465,N_14728);
nand UO_1710 (O_1710,N_14433,N_14245);
xor UO_1711 (O_1711,N_14577,N_14570);
or UO_1712 (O_1712,N_14530,N_14428);
or UO_1713 (O_1713,N_14766,N_14044);
xor UO_1714 (O_1714,N_14716,N_14483);
or UO_1715 (O_1715,N_14129,N_14039);
nor UO_1716 (O_1716,N_14357,N_14773);
nand UO_1717 (O_1717,N_14706,N_14849);
and UO_1718 (O_1718,N_14060,N_14194);
or UO_1719 (O_1719,N_14327,N_14868);
nand UO_1720 (O_1720,N_14282,N_14352);
nand UO_1721 (O_1721,N_14391,N_14415);
and UO_1722 (O_1722,N_14591,N_14066);
nor UO_1723 (O_1723,N_14717,N_14428);
nor UO_1724 (O_1724,N_14820,N_14434);
nand UO_1725 (O_1725,N_14457,N_14313);
or UO_1726 (O_1726,N_14432,N_14228);
nor UO_1727 (O_1727,N_14778,N_14610);
or UO_1728 (O_1728,N_14128,N_14834);
or UO_1729 (O_1729,N_14750,N_14169);
or UO_1730 (O_1730,N_14174,N_14834);
nand UO_1731 (O_1731,N_14245,N_14282);
nand UO_1732 (O_1732,N_14453,N_14147);
nand UO_1733 (O_1733,N_14912,N_14007);
nand UO_1734 (O_1734,N_14959,N_14768);
xnor UO_1735 (O_1735,N_14350,N_14841);
nor UO_1736 (O_1736,N_14730,N_14653);
or UO_1737 (O_1737,N_14913,N_14356);
nor UO_1738 (O_1738,N_14220,N_14929);
nand UO_1739 (O_1739,N_14820,N_14702);
or UO_1740 (O_1740,N_14371,N_14820);
xnor UO_1741 (O_1741,N_14155,N_14054);
xor UO_1742 (O_1742,N_14040,N_14227);
and UO_1743 (O_1743,N_14288,N_14320);
or UO_1744 (O_1744,N_14988,N_14662);
and UO_1745 (O_1745,N_14741,N_14557);
nor UO_1746 (O_1746,N_14647,N_14134);
nor UO_1747 (O_1747,N_14538,N_14076);
xor UO_1748 (O_1748,N_14828,N_14320);
or UO_1749 (O_1749,N_14655,N_14502);
nand UO_1750 (O_1750,N_14300,N_14561);
xor UO_1751 (O_1751,N_14164,N_14256);
or UO_1752 (O_1752,N_14289,N_14809);
nand UO_1753 (O_1753,N_14691,N_14649);
xnor UO_1754 (O_1754,N_14086,N_14745);
or UO_1755 (O_1755,N_14332,N_14011);
xnor UO_1756 (O_1756,N_14850,N_14344);
and UO_1757 (O_1757,N_14876,N_14100);
xor UO_1758 (O_1758,N_14114,N_14369);
and UO_1759 (O_1759,N_14617,N_14166);
or UO_1760 (O_1760,N_14583,N_14141);
nor UO_1761 (O_1761,N_14186,N_14573);
nor UO_1762 (O_1762,N_14588,N_14341);
xor UO_1763 (O_1763,N_14536,N_14149);
nand UO_1764 (O_1764,N_14723,N_14039);
nor UO_1765 (O_1765,N_14138,N_14322);
or UO_1766 (O_1766,N_14638,N_14509);
and UO_1767 (O_1767,N_14592,N_14542);
and UO_1768 (O_1768,N_14484,N_14303);
nand UO_1769 (O_1769,N_14998,N_14065);
or UO_1770 (O_1770,N_14719,N_14664);
and UO_1771 (O_1771,N_14336,N_14913);
or UO_1772 (O_1772,N_14829,N_14977);
nor UO_1773 (O_1773,N_14324,N_14304);
nor UO_1774 (O_1774,N_14196,N_14727);
and UO_1775 (O_1775,N_14555,N_14601);
xor UO_1776 (O_1776,N_14313,N_14548);
and UO_1777 (O_1777,N_14048,N_14037);
and UO_1778 (O_1778,N_14045,N_14552);
nand UO_1779 (O_1779,N_14403,N_14338);
nor UO_1780 (O_1780,N_14848,N_14397);
nand UO_1781 (O_1781,N_14804,N_14826);
nor UO_1782 (O_1782,N_14991,N_14236);
or UO_1783 (O_1783,N_14667,N_14952);
nand UO_1784 (O_1784,N_14989,N_14102);
and UO_1785 (O_1785,N_14786,N_14116);
and UO_1786 (O_1786,N_14741,N_14087);
nand UO_1787 (O_1787,N_14744,N_14540);
or UO_1788 (O_1788,N_14165,N_14706);
or UO_1789 (O_1789,N_14912,N_14356);
or UO_1790 (O_1790,N_14804,N_14395);
nand UO_1791 (O_1791,N_14870,N_14993);
and UO_1792 (O_1792,N_14213,N_14156);
and UO_1793 (O_1793,N_14218,N_14134);
or UO_1794 (O_1794,N_14702,N_14682);
xnor UO_1795 (O_1795,N_14243,N_14765);
or UO_1796 (O_1796,N_14833,N_14491);
nor UO_1797 (O_1797,N_14951,N_14838);
and UO_1798 (O_1798,N_14207,N_14682);
or UO_1799 (O_1799,N_14852,N_14120);
nand UO_1800 (O_1800,N_14213,N_14847);
xor UO_1801 (O_1801,N_14206,N_14353);
xor UO_1802 (O_1802,N_14476,N_14905);
or UO_1803 (O_1803,N_14750,N_14621);
or UO_1804 (O_1804,N_14020,N_14248);
nand UO_1805 (O_1805,N_14142,N_14614);
nor UO_1806 (O_1806,N_14528,N_14467);
or UO_1807 (O_1807,N_14415,N_14564);
and UO_1808 (O_1808,N_14449,N_14837);
and UO_1809 (O_1809,N_14904,N_14091);
nor UO_1810 (O_1810,N_14185,N_14648);
and UO_1811 (O_1811,N_14381,N_14633);
or UO_1812 (O_1812,N_14995,N_14162);
nand UO_1813 (O_1813,N_14391,N_14797);
nand UO_1814 (O_1814,N_14522,N_14144);
nand UO_1815 (O_1815,N_14848,N_14922);
nand UO_1816 (O_1816,N_14261,N_14419);
xor UO_1817 (O_1817,N_14508,N_14244);
xnor UO_1818 (O_1818,N_14242,N_14343);
and UO_1819 (O_1819,N_14559,N_14263);
and UO_1820 (O_1820,N_14482,N_14870);
nand UO_1821 (O_1821,N_14222,N_14361);
nor UO_1822 (O_1822,N_14170,N_14142);
xnor UO_1823 (O_1823,N_14999,N_14176);
and UO_1824 (O_1824,N_14596,N_14234);
nand UO_1825 (O_1825,N_14708,N_14592);
nand UO_1826 (O_1826,N_14529,N_14457);
or UO_1827 (O_1827,N_14672,N_14478);
or UO_1828 (O_1828,N_14541,N_14161);
nor UO_1829 (O_1829,N_14699,N_14234);
nand UO_1830 (O_1830,N_14075,N_14881);
and UO_1831 (O_1831,N_14608,N_14359);
nor UO_1832 (O_1832,N_14960,N_14266);
and UO_1833 (O_1833,N_14406,N_14614);
nand UO_1834 (O_1834,N_14996,N_14456);
or UO_1835 (O_1835,N_14298,N_14152);
nor UO_1836 (O_1836,N_14480,N_14277);
or UO_1837 (O_1837,N_14578,N_14141);
or UO_1838 (O_1838,N_14094,N_14237);
and UO_1839 (O_1839,N_14752,N_14090);
nor UO_1840 (O_1840,N_14133,N_14952);
and UO_1841 (O_1841,N_14076,N_14917);
or UO_1842 (O_1842,N_14021,N_14029);
nor UO_1843 (O_1843,N_14913,N_14923);
xor UO_1844 (O_1844,N_14171,N_14407);
nand UO_1845 (O_1845,N_14097,N_14318);
nand UO_1846 (O_1846,N_14089,N_14454);
nor UO_1847 (O_1847,N_14049,N_14895);
xnor UO_1848 (O_1848,N_14608,N_14387);
and UO_1849 (O_1849,N_14706,N_14762);
or UO_1850 (O_1850,N_14717,N_14514);
nor UO_1851 (O_1851,N_14307,N_14389);
and UO_1852 (O_1852,N_14364,N_14564);
and UO_1853 (O_1853,N_14742,N_14322);
nand UO_1854 (O_1854,N_14548,N_14054);
nor UO_1855 (O_1855,N_14587,N_14179);
or UO_1856 (O_1856,N_14102,N_14965);
nand UO_1857 (O_1857,N_14346,N_14170);
or UO_1858 (O_1858,N_14529,N_14675);
or UO_1859 (O_1859,N_14799,N_14074);
nor UO_1860 (O_1860,N_14075,N_14239);
nor UO_1861 (O_1861,N_14348,N_14152);
and UO_1862 (O_1862,N_14812,N_14962);
or UO_1863 (O_1863,N_14195,N_14142);
nand UO_1864 (O_1864,N_14103,N_14775);
xor UO_1865 (O_1865,N_14726,N_14093);
nand UO_1866 (O_1866,N_14761,N_14743);
or UO_1867 (O_1867,N_14776,N_14376);
nor UO_1868 (O_1868,N_14792,N_14934);
nand UO_1869 (O_1869,N_14565,N_14360);
or UO_1870 (O_1870,N_14776,N_14056);
or UO_1871 (O_1871,N_14516,N_14894);
nor UO_1872 (O_1872,N_14151,N_14217);
xor UO_1873 (O_1873,N_14325,N_14770);
or UO_1874 (O_1874,N_14322,N_14770);
nand UO_1875 (O_1875,N_14031,N_14334);
and UO_1876 (O_1876,N_14711,N_14620);
or UO_1877 (O_1877,N_14332,N_14257);
xnor UO_1878 (O_1878,N_14509,N_14068);
and UO_1879 (O_1879,N_14981,N_14540);
xor UO_1880 (O_1880,N_14671,N_14347);
or UO_1881 (O_1881,N_14161,N_14289);
and UO_1882 (O_1882,N_14653,N_14798);
nand UO_1883 (O_1883,N_14329,N_14839);
xor UO_1884 (O_1884,N_14730,N_14027);
or UO_1885 (O_1885,N_14875,N_14476);
nand UO_1886 (O_1886,N_14642,N_14989);
or UO_1887 (O_1887,N_14756,N_14755);
and UO_1888 (O_1888,N_14453,N_14481);
nor UO_1889 (O_1889,N_14093,N_14645);
nor UO_1890 (O_1890,N_14641,N_14041);
or UO_1891 (O_1891,N_14041,N_14719);
nand UO_1892 (O_1892,N_14024,N_14408);
nand UO_1893 (O_1893,N_14246,N_14426);
nor UO_1894 (O_1894,N_14145,N_14650);
xnor UO_1895 (O_1895,N_14097,N_14316);
and UO_1896 (O_1896,N_14524,N_14397);
nand UO_1897 (O_1897,N_14990,N_14092);
nand UO_1898 (O_1898,N_14555,N_14128);
or UO_1899 (O_1899,N_14781,N_14190);
or UO_1900 (O_1900,N_14698,N_14841);
nor UO_1901 (O_1901,N_14363,N_14040);
and UO_1902 (O_1902,N_14186,N_14750);
xnor UO_1903 (O_1903,N_14325,N_14412);
nor UO_1904 (O_1904,N_14223,N_14865);
nor UO_1905 (O_1905,N_14202,N_14588);
or UO_1906 (O_1906,N_14607,N_14669);
xnor UO_1907 (O_1907,N_14161,N_14287);
nor UO_1908 (O_1908,N_14290,N_14948);
nor UO_1909 (O_1909,N_14413,N_14887);
xor UO_1910 (O_1910,N_14780,N_14360);
nand UO_1911 (O_1911,N_14523,N_14088);
xor UO_1912 (O_1912,N_14594,N_14857);
or UO_1913 (O_1913,N_14672,N_14325);
or UO_1914 (O_1914,N_14736,N_14224);
xor UO_1915 (O_1915,N_14183,N_14853);
nand UO_1916 (O_1916,N_14652,N_14467);
and UO_1917 (O_1917,N_14818,N_14420);
or UO_1918 (O_1918,N_14805,N_14995);
and UO_1919 (O_1919,N_14084,N_14565);
xor UO_1920 (O_1920,N_14384,N_14661);
or UO_1921 (O_1921,N_14847,N_14177);
nand UO_1922 (O_1922,N_14459,N_14239);
nor UO_1923 (O_1923,N_14959,N_14431);
xnor UO_1924 (O_1924,N_14933,N_14758);
and UO_1925 (O_1925,N_14631,N_14810);
nand UO_1926 (O_1926,N_14982,N_14860);
xor UO_1927 (O_1927,N_14754,N_14836);
nor UO_1928 (O_1928,N_14864,N_14129);
nor UO_1929 (O_1929,N_14656,N_14923);
nor UO_1930 (O_1930,N_14154,N_14048);
or UO_1931 (O_1931,N_14088,N_14684);
or UO_1932 (O_1932,N_14592,N_14914);
and UO_1933 (O_1933,N_14459,N_14219);
nand UO_1934 (O_1934,N_14628,N_14314);
nor UO_1935 (O_1935,N_14920,N_14620);
and UO_1936 (O_1936,N_14532,N_14884);
or UO_1937 (O_1937,N_14876,N_14898);
nor UO_1938 (O_1938,N_14029,N_14965);
and UO_1939 (O_1939,N_14469,N_14588);
or UO_1940 (O_1940,N_14751,N_14733);
nor UO_1941 (O_1941,N_14347,N_14007);
nand UO_1942 (O_1942,N_14265,N_14948);
or UO_1943 (O_1943,N_14098,N_14413);
or UO_1944 (O_1944,N_14649,N_14881);
and UO_1945 (O_1945,N_14089,N_14019);
xor UO_1946 (O_1946,N_14517,N_14983);
nand UO_1947 (O_1947,N_14301,N_14200);
and UO_1948 (O_1948,N_14231,N_14430);
nand UO_1949 (O_1949,N_14720,N_14638);
xor UO_1950 (O_1950,N_14638,N_14800);
nor UO_1951 (O_1951,N_14670,N_14188);
xnor UO_1952 (O_1952,N_14107,N_14131);
xnor UO_1953 (O_1953,N_14739,N_14908);
and UO_1954 (O_1954,N_14064,N_14682);
nand UO_1955 (O_1955,N_14508,N_14950);
and UO_1956 (O_1956,N_14090,N_14704);
xor UO_1957 (O_1957,N_14476,N_14167);
nor UO_1958 (O_1958,N_14044,N_14460);
and UO_1959 (O_1959,N_14231,N_14821);
and UO_1960 (O_1960,N_14936,N_14990);
and UO_1961 (O_1961,N_14263,N_14470);
nor UO_1962 (O_1962,N_14242,N_14240);
nand UO_1963 (O_1963,N_14042,N_14176);
and UO_1964 (O_1964,N_14241,N_14718);
nor UO_1965 (O_1965,N_14476,N_14828);
nand UO_1966 (O_1966,N_14130,N_14444);
nor UO_1967 (O_1967,N_14717,N_14096);
and UO_1968 (O_1968,N_14398,N_14710);
nor UO_1969 (O_1969,N_14898,N_14715);
nor UO_1970 (O_1970,N_14060,N_14961);
nand UO_1971 (O_1971,N_14497,N_14231);
nor UO_1972 (O_1972,N_14731,N_14640);
or UO_1973 (O_1973,N_14487,N_14605);
or UO_1974 (O_1974,N_14998,N_14458);
and UO_1975 (O_1975,N_14283,N_14082);
nand UO_1976 (O_1976,N_14267,N_14713);
xnor UO_1977 (O_1977,N_14877,N_14924);
xor UO_1978 (O_1978,N_14068,N_14759);
xor UO_1979 (O_1979,N_14075,N_14968);
nand UO_1980 (O_1980,N_14421,N_14628);
and UO_1981 (O_1981,N_14924,N_14428);
or UO_1982 (O_1982,N_14140,N_14169);
xnor UO_1983 (O_1983,N_14858,N_14430);
nor UO_1984 (O_1984,N_14390,N_14863);
and UO_1985 (O_1985,N_14987,N_14535);
and UO_1986 (O_1986,N_14181,N_14062);
xnor UO_1987 (O_1987,N_14019,N_14964);
and UO_1988 (O_1988,N_14703,N_14214);
xnor UO_1989 (O_1989,N_14687,N_14319);
nand UO_1990 (O_1990,N_14087,N_14334);
or UO_1991 (O_1991,N_14382,N_14590);
and UO_1992 (O_1992,N_14445,N_14378);
and UO_1993 (O_1993,N_14090,N_14619);
nor UO_1994 (O_1994,N_14621,N_14231);
and UO_1995 (O_1995,N_14478,N_14090);
or UO_1996 (O_1996,N_14452,N_14072);
nor UO_1997 (O_1997,N_14773,N_14487);
and UO_1998 (O_1998,N_14379,N_14900);
or UO_1999 (O_1999,N_14985,N_14727);
endmodule