module basic_1000_10000_1500_100_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_533,In_121);
nor U1 (N_1,In_979,In_725);
and U2 (N_2,In_21,In_126);
nor U3 (N_3,In_704,In_931);
nor U4 (N_4,In_230,In_404);
nor U5 (N_5,In_60,In_705);
and U6 (N_6,In_500,In_922);
nor U7 (N_7,In_496,In_640);
nor U8 (N_8,In_795,In_754);
or U9 (N_9,In_497,In_880);
xnor U10 (N_10,In_962,In_84);
nor U11 (N_11,In_732,In_133);
or U12 (N_12,In_251,In_426);
nand U13 (N_13,In_364,In_183);
or U14 (N_14,In_680,In_332);
nand U15 (N_15,In_787,In_843);
nor U16 (N_16,In_434,In_446);
or U17 (N_17,In_585,In_886);
nand U18 (N_18,In_637,In_663);
or U19 (N_19,In_806,In_878);
or U20 (N_20,In_98,In_653);
or U21 (N_21,In_944,In_214);
and U22 (N_22,In_905,In_847);
nor U23 (N_23,In_887,In_210);
nand U24 (N_24,In_4,In_372);
or U25 (N_25,In_515,In_852);
and U26 (N_26,In_552,In_863);
nand U27 (N_27,In_453,In_297);
and U28 (N_28,In_14,In_984);
xor U29 (N_29,In_18,In_826);
nor U30 (N_30,In_987,In_667);
xnor U31 (N_31,In_716,In_238);
and U32 (N_32,In_975,In_553);
and U33 (N_33,In_528,In_478);
and U34 (N_34,In_738,In_36);
and U35 (N_35,In_235,In_571);
or U36 (N_36,In_417,In_392);
nor U37 (N_37,In_956,In_236);
nor U38 (N_38,In_408,In_110);
nand U39 (N_39,In_591,In_714);
or U40 (N_40,In_699,In_662);
xnor U41 (N_41,In_567,In_914);
and U42 (N_42,In_520,In_947);
xor U43 (N_43,In_815,In_598);
and U44 (N_44,In_796,In_17);
nor U45 (N_45,In_678,In_652);
nand U46 (N_46,In_656,In_940);
nand U47 (N_47,In_93,In_470);
or U48 (N_48,In_835,In_248);
nand U49 (N_49,In_649,In_522);
nor U50 (N_50,In_829,In_564);
nand U51 (N_51,In_285,In_724);
and U52 (N_52,In_237,In_576);
nand U53 (N_53,In_658,In_872);
nand U54 (N_54,In_926,In_969);
nor U55 (N_55,In_390,In_643);
or U56 (N_56,In_952,In_566);
nor U57 (N_57,In_890,In_124);
nor U58 (N_58,In_70,In_81);
or U59 (N_59,In_486,In_211);
and U60 (N_60,In_166,In_68);
nor U61 (N_61,In_170,In_180);
and U62 (N_62,In_540,In_734);
or U63 (N_63,In_212,In_433);
nand U64 (N_64,In_774,In_701);
and U65 (N_65,In_670,In_273);
and U66 (N_66,In_537,In_411);
and U67 (N_67,In_785,In_672);
nor U68 (N_68,In_839,In_336);
and U69 (N_69,In_638,In_61);
and U70 (N_70,In_594,In_90);
or U71 (N_71,In_57,In_582);
nand U72 (N_72,In_554,In_673);
xor U73 (N_73,In_59,In_335);
nand U74 (N_74,In_513,In_963);
and U75 (N_75,In_47,In_740);
nor U76 (N_76,In_423,In_458);
and U77 (N_77,In_903,In_213);
and U78 (N_78,In_250,In_25);
nor U79 (N_79,In_810,In_267);
and U80 (N_80,In_971,In_937);
or U81 (N_81,In_460,In_832);
xor U82 (N_82,In_702,In_33);
nor U83 (N_83,In_174,In_642);
nor U84 (N_84,In_197,In_836);
and U85 (N_85,In_960,In_595);
or U86 (N_86,In_599,In_659);
and U87 (N_87,In_337,In_402);
and U88 (N_88,In_116,In_964);
or U89 (N_89,In_312,In_946);
or U90 (N_90,In_179,In_243);
xnor U91 (N_91,In_572,In_748);
or U92 (N_92,In_601,In_505);
nand U93 (N_93,In_583,In_651);
nand U94 (N_94,In_375,In_590);
or U95 (N_95,In_930,In_921);
or U96 (N_96,In_193,In_902);
or U97 (N_97,In_646,In_783);
or U98 (N_98,In_233,In_64);
or U99 (N_99,In_563,In_586);
xnor U100 (N_100,In_481,In_950);
or U101 (N_101,In_524,In_153);
xor U102 (N_102,In_827,In_442);
or U103 (N_103,In_295,In_252);
nor U104 (N_104,In_492,In_519);
nor U105 (N_105,In_209,N_85);
nand U106 (N_106,In_62,In_789);
nand U107 (N_107,In_727,In_321);
or U108 (N_108,In_39,In_41);
and U109 (N_109,In_397,In_574);
nand U110 (N_110,In_866,In_750);
nand U111 (N_111,In_915,In_53);
xor U112 (N_112,In_362,In_88);
and U113 (N_113,In_148,In_227);
nor U114 (N_114,In_924,In_284);
or U115 (N_115,In_634,In_874);
or U116 (N_116,In_526,In_52);
nor U117 (N_117,In_228,In_896);
nand U118 (N_118,In_360,In_244);
and U119 (N_119,In_483,In_198);
nand U120 (N_120,In_812,In_269);
nor U121 (N_121,In_281,In_293);
and U122 (N_122,N_68,In_387);
xor U123 (N_123,In_809,In_468);
and U124 (N_124,In_970,In_927);
nand U125 (N_125,In_428,In_710);
nand U126 (N_126,In_79,In_986);
or U127 (N_127,In_814,In_339);
and U128 (N_128,In_194,In_311);
or U129 (N_129,In_942,In_418);
and U130 (N_130,In_983,In_104);
and U131 (N_131,In_684,In_461);
xor U132 (N_132,In_438,In_908);
and U133 (N_133,In_331,In_232);
nor U134 (N_134,In_441,In_780);
nand U135 (N_135,In_884,In_629);
xnor U136 (N_136,In_76,In_650);
nand U137 (N_137,In_118,In_163);
or U138 (N_138,In_491,In_117);
nand U139 (N_139,In_633,N_15);
nand U140 (N_140,In_420,In_995);
nor U141 (N_141,In_488,In_393);
nand U142 (N_142,In_484,In_317);
nand U143 (N_143,In_42,In_287);
xor U144 (N_144,In_388,In_407);
nand U145 (N_145,In_135,In_838);
or U146 (N_146,In_561,In_772);
nand U147 (N_147,In_114,In_792);
nor U148 (N_148,In_55,In_63);
and U149 (N_149,In_607,In_181);
nor U150 (N_150,N_26,In_192);
nor U151 (N_151,In_344,In_669);
and U152 (N_152,In_152,In_741);
and U153 (N_153,In_119,In_432);
nor U154 (N_154,In_389,In_26);
nor U155 (N_155,In_38,In_203);
nor U156 (N_156,In_425,In_266);
xor U157 (N_157,In_534,In_377);
and U158 (N_158,In_419,In_802);
nand U159 (N_159,In_630,In_208);
and U160 (N_160,N_95,In_20);
or U161 (N_161,In_588,N_25);
xor U162 (N_162,In_749,In_304);
nand U163 (N_163,In_489,In_562);
nand U164 (N_164,In_856,In_800);
and U165 (N_165,In_6,In_318);
nand U166 (N_166,In_240,In_790);
or U167 (N_167,N_0,In_200);
or U168 (N_168,In_910,In_906);
or U169 (N_169,In_395,In_289);
nand U170 (N_170,In_2,In_99);
nand U171 (N_171,In_988,N_35);
nor U172 (N_172,In_215,In_415);
xnor U173 (N_173,In_525,In_165);
or U174 (N_174,N_88,In_11);
or U175 (N_175,In_794,In_568);
or U176 (N_176,N_96,N_92);
or U177 (N_177,In_167,In_406);
or U178 (N_178,In_299,In_265);
or U179 (N_179,In_711,In_542);
or U180 (N_180,In_693,In_306);
or U181 (N_181,In_222,In_282);
nor U182 (N_182,In_31,In_19);
nor U183 (N_183,In_862,In_833);
nand U184 (N_184,N_22,In_29);
nor U185 (N_185,In_363,In_159);
nand U186 (N_186,In_674,N_9);
or U187 (N_187,In_686,In_218);
nand U188 (N_188,In_398,N_1);
xor U189 (N_189,In_523,In_142);
nand U190 (N_190,In_474,In_147);
and U191 (N_191,In_189,In_918);
nor U192 (N_192,In_898,In_7);
and U193 (N_193,In_647,In_369);
or U194 (N_194,In_349,In_195);
or U195 (N_195,In_108,In_909);
and U196 (N_196,In_512,In_288);
and U197 (N_197,N_78,In_535);
or U198 (N_198,N_67,In_329);
and U199 (N_199,In_756,In_224);
and U200 (N_200,In_690,In_394);
nand U201 (N_201,In_703,In_254);
or U202 (N_202,In_365,N_31);
nand U203 (N_203,N_38,N_133);
and U204 (N_204,N_150,In_296);
or U205 (N_205,N_58,In_187);
or U206 (N_206,In_531,In_615);
or U207 (N_207,In_958,In_378);
nand U208 (N_208,N_168,In_323);
xnor U209 (N_209,In_80,In_616);
nand U210 (N_210,In_16,N_36);
nand U211 (N_211,In_801,In_463);
or U212 (N_212,In_793,In_846);
or U213 (N_213,N_93,N_164);
nor U214 (N_214,In_275,In_454);
and U215 (N_215,In_412,In_28);
and U216 (N_216,In_954,In_824);
and U217 (N_217,In_72,In_632);
nand U218 (N_218,In_13,N_17);
nand U219 (N_219,In_345,In_767);
or U220 (N_220,N_198,N_129);
and U221 (N_221,In_437,In_82);
nand U222 (N_222,In_391,In_246);
nor U223 (N_223,In_457,In_851);
nor U224 (N_224,In_145,In_443);
nand U225 (N_225,N_176,In_9);
nor U226 (N_226,N_24,In_469);
or U227 (N_227,In_837,In_682);
and U228 (N_228,In_894,In_155);
nand U229 (N_229,In_308,N_39);
nand U230 (N_230,N_66,In_511);
nor U231 (N_231,In_459,In_596);
and U232 (N_232,In_374,In_544);
or U233 (N_233,In_804,In_757);
and U234 (N_234,In_171,In_507);
nand U235 (N_235,N_196,In_712);
or U236 (N_236,In_817,In_216);
nor U237 (N_237,In_482,N_184);
nand U238 (N_238,In_593,In_292);
nor U239 (N_239,In_74,In_990);
nand U240 (N_240,In_998,In_831);
nor U241 (N_241,In_695,In_22);
or U242 (N_242,In_277,In_580);
or U243 (N_243,In_66,In_993);
xnor U244 (N_244,In_328,In_786);
nor U245 (N_245,In_48,In_361);
nor U246 (N_246,In_421,N_11);
nand U247 (N_247,In_938,In_521);
nor U248 (N_248,In_888,In_69);
and U249 (N_249,In_405,In_92);
and U250 (N_250,In_45,In_161);
and U251 (N_251,In_530,N_77);
and U252 (N_252,In_150,In_50);
nand U253 (N_253,N_84,N_172);
nor U254 (N_254,In_300,In_123);
or U255 (N_255,In_310,In_177);
or U256 (N_256,In_901,In_353);
nand U257 (N_257,In_334,N_56);
nor U258 (N_258,In_822,In_840);
nand U259 (N_259,In_536,In_911);
nand U260 (N_260,In_134,In_700);
nand U261 (N_261,In_627,In_154);
or U262 (N_262,N_152,In_396);
xor U263 (N_263,In_0,N_19);
xnor U264 (N_264,N_43,In_448);
nand U265 (N_265,N_30,In_413);
or U266 (N_266,In_980,In_113);
xor U267 (N_267,N_158,In_436);
and U268 (N_268,In_268,In_717);
nor U269 (N_269,In_139,In_858);
nand U270 (N_270,In_737,In_845);
or U271 (N_271,In_422,In_314);
xnor U272 (N_272,In_538,In_913);
xnor U273 (N_273,In_263,N_60);
nand U274 (N_274,In_307,In_270);
and U275 (N_275,N_120,In_225);
or U276 (N_276,N_147,In_753);
nand U277 (N_277,N_145,In_925);
and U278 (N_278,N_4,In_782);
nor U279 (N_279,In_494,In_623);
xor U280 (N_280,In_560,In_955);
nand U281 (N_281,In_342,In_357);
and U282 (N_282,In_264,N_143);
or U283 (N_283,In_755,In_132);
or U284 (N_284,In_450,N_179);
xnor U285 (N_285,In_828,In_15);
nor U286 (N_286,In_529,N_157);
nand U287 (N_287,In_294,N_122);
and U288 (N_288,In_234,In_91);
or U289 (N_289,N_76,In_477);
or U290 (N_290,In_621,N_55);
nand U291 (N_291,In_302,In_726);
nor U292 (N_292,In_626,In_67);
nor U293 (N_293,In_414,In_784);
nand U294 (N_294,N_100,N_14);
or U295 (N_295,In_698,In_645);
and U296 (N_296,In_834,In_451);
or U297 (N_297,N_101,In_473);
nand U298 (N_298,In_602,In_614);
nor U299 (N_299,In_777,In_445);
nor U300 (N_300,N_247,In_985);
nand U301 (N_301,N_221,In_859);
and U302 (N_302,In_510,In_509);
or U303 (N_303,In_948,In_694);
nor U304 (N_304,N_50,N_117);
nor U305 (N_305,In_668,In_427);
nor U306 (N_306,N_255,In_639);
or U307 (N_307,In_733,In_881);
or U308 (N_308,N_284,In_532);
nand U309 (N_309,In_464,N_274);
or U310 (N_310,N_218,In_162);
and U311 (N_311,In_897,N_131);
nor U312 (N_312,In_356,In_661);
nand U313 (N_313,In_128,In_981);
nand U314 (N_314,N_108,In_850);
or U315 (N_315,In_578,N_259);
or U316 (N_316,In_729,N_249);
nor U317 (N_317,In_348,In_697);
or U318 (N_318,N_182,In_860);
nand U319 (N_319,In_107,In_373);
and U320 (N_320,In_498,N_267);
xnor U321 (N_321,N_23,In_957);
nor U322 (N_322,N_70,N_252);
nand U323 (N_323,In_3,In_770);
or U324 (N_324,N_275,In_429);
nand U325 (N_325,In_713,In_876);
and U326 (N_326,N_175,N_87);
or U327 (N_327,N_113,N_174);
and U328 (N_328,In_49,In_327);
or U329 (N_329,In_386,N_228);
nand U330 (N_330,In_548,N_73);
nand U331 (N_331,In_291,In_143);
nand U332 (N_332,N_52,N_266);
nand U333 (N_333,N_211,In_403);
or U334 (N_334,In_354,In_959);
nor U335 (N_335,N_295,In_821);
and U336 (N_336,In_410,In_358);
nor U337 (N_337,In_849,In_625);
and U338 (N_338,In_655,N_7);
nand U339 (N_339,In_176,N_127);
and U340 (N_340,In_366,In_779);
or U341 (N_341,In_719,In_557);
or U342 (N_342,In_720,N_167);
and U343 (N_343,N_98,In_56);
xor U344 (N_344,N_21,N_233);
nor U345 (N_345,In_487,N_187);
and U346 (N_346,N_289,N_239);
or U347 (N_347,In_751,N_299);
nand U348 (N_348,In_112,In_503);
nor U349 (N_349,In_272,N_273);
nor U350 (N_350,N_162,In_604);
nand U351 (N_351,In_589,N_107);
and U352 (N_352,N_149,In_343);
or U353 (N_353,In_274,In_797);
nand U354 (N_354,N_90,In_325);
and U355 (N_355,In_696,In_592);
xor U356 (N_356,In_83,In_929);
and U357 (N_357,N_154,In_359);
xor U358 (N_358,In_660,N_34);
or U359 (N_359,In_199,N_64);
nand U360 (N_360,N_10,In_506);
nor U361 (N_361,In_207,In_555);
xnor U362 (N_362,In_675,In_46);
nand U363 (N_363,In_330,In_764);
and U364 (N_364,In_584,In_654);
nand U365 (N_365,N_69,In_943);
nand U366 (N_366,N_219,In_204);
nand U367 (N_367,In_636,In_577);
xnor U368 (N_368,In_517,In_706);
xor U369 (N_369,N_204,In_175);
xnor U370 (N_370,In_895,In_781);
xnor U371 (N_371,N_200,In_945);
nand U372 (N_372,In_617,In_788);
nor U373 (N_373,In_539,In_977);
nor U374 (N_374,In_350,N_238);
or U375 (N_375,In_260,In_644);
or U376 (N_376,In_994,In_864);
nor U377 (N_377,In_115,In_932);
nor U378 (N_378,N_136,In_624);
and U379 (N_379,In_516,N_271);
nand U380 (N_380,In_191,In_182);
nand U381 (N_381,In_941,In_504);
or U382 (N_382,N_135,In_467);
nand U383 (N_383,In_605,In_613);
nand U384 (N_384,In_514,N_232);
and U385 (N_385,In_742,In_923);
and U386 (N_386,In_160,In_346);
nor U387 (N_387,In_168,In_889);
nor U388 (N_388,N_45,In_805);
and U389 (N_389,N_111,In_844);
xnor U390 (N_390,In_976,In_401);
nor U391 (N_391,In_186,N_207);
and U392 (N_392,In_255,In_309);
and U393 (N_393,In_384,N_75);
nor U394 (N_394,In_111,N_216);
nand U395 (N_395,In_628,In_620);
xnor U396 (N_396,N_62,In_982);
nor U397 (N_397,In_44,In_127);
nor U398 (N_398,N_291,In_303);
nor U399 (N_399,N_37,N_159);
and U400 (N_400,In_820,N_302);
nand U401 (N_401,In_131,N_188);
xnor U402 (N_402,N_140,In_546);
nand U403 (N_403,N_306,In_570);
and U404 (N_404,N_310,In_495);
nand U405 (N_405,N_33,N_372);
nand U406 (N_406,N_178,N_390);
and U407 (N_407,N_396,N_296);
and U408 (N_408,In_664,In_919);
nand U409 (N_409,In_608,N_340);
nor U410 (N_410,In_324,N_276);
or U411 (N_411,N_327,In_35);
nand U412 (N_412,N_321,In_631);
and U413 (N_413,N_210,N_380);
nand U414 (N_414,In_169,N_304);
nor U415 (N_415,In_619,N_116);
or U416 (N_416,N_74,N_91);
or U417 (N_417,In_258,N_280);
nor U418 (N_418,In_543,In_871);
or U419 (N_419,In_424,N_209);
nand U420 (N_420,In_996,In_89);
and U421 (N_421,N_298,In_231);
nor U422 (N_422,In_676,N_386);
or U423 (N_423,In_745,N_54);
nor U424 (N_424,In_769,In_379);
nand U425 (N_425,In_305,In_456);
or U426 (N_426,In_877,In_808);
or U427 (N_427,N_2,N_370);
and U428 (N_428,In_773,N_364);
and U429 (N_429,N_119,N_338);
nor U430 (N_430,In_791,N_236);
nor U431 (N_431,In_476,In_689);
or U432 (N_432,In_261,N_13);
nor U433 (N_433,In_550,In_799);
or U434 (N_434,In_870,N_20);
and U435 (N_435,In_140,In_239);
xor U436 (N_436,In_935,In_765);
and U437 (N_437,In_439,N_253);
or U438 (N_438,In_811,In_989);
and U439 (N_439,In_761,In_257);
or U440 (N_440,N_375,In_103);
nand U441 (N_441,N_303,N_367);
or U442 (N_442,In_965,In_367);
and U443 (N_443,In_666,In_768);
and U444 (N_444,N_205,In_692);
nand U445 (N_445,N_345,In_137);
xor U446 (N_446,In_333,In_485);
or U447 (N_447,In_992,In_618);
or U448 (N_448,In_400,In_149);
nand U449 (N_449,In_435,N_155);
nand U450 (N_450,In_766,In_721);
and U451 (N_451,In_579,In_867);
nand U452 (N_452,In_253,In_184);
nand U453 (N_453,In_735,N_318);
nand U454 (N_454,N_389,N_248);
or U455 (N_455,In_276,N_123);
nor U456 (N_456,N_86,N_378);
and U457 (N_457,In_885,N_348);
and U458 (N_458,In_606,N_217);
xnor U459 (N_459,N_201,In_762);
xnor U460 (N_460,In_54,In_280);
nor U461 (N_461,In_313,In_597);
nand U462 (N_462,In_928,N_137);
xnor U463 (N_463,N_300,In_472);
nand U464 (N_464,In_156,N_257);
nand U465 (N_465,In_97,N_242);
and U466 (N_466,N_360,N_260);
nand U467 (N_467,N_351,N_124);
or U468 (N_468,In_541,N_244);
and U469 (N_469,N_132,N_48);
nand U470 (N_470,N_379,N_118);
and U471 (N_471,In_728,In_933);
xnor U472 (N_472,N_330,In_722);
and U473 (N_473,N_112,In_823);
or U474 (N_474,In_892,N_171);
nand U475 (N_475,N_5,N_341);
xnor U476 (N_476,In_743,In_816);
xnor U477 (N_477,N_82,In_78);
or U478 (N_478,N_397,N_393);
and U479 (N_479,In_245,In_259);
or U480 (N_480,N_334,In_818);
nand U481 (N_481,In_279,In_290);
and U482 (N_482,In_688,In_196);
nand U483 (N_483,N_16,N_72);
nor U484 (N_484,In_206,N_241);
or U485 (N_485,N_18,In_462);
and U486 (N_486,In_452,N_227);
nand U487 (N_487,In_775,In_351);
nor U488 (N_488,N_192,In_853);
nor U489 (N_489,N_350,In_912);
nor U490 (N_490,N_349,N_278);
xnor U491 (N_491,In_249,N_134);
and U492 (N_492,In_974,N_191);
nand U493 (N_493,In_43,N_28);
or U494 (N_494,In_444,N_353);
or U495 (N_495,In_229,In_157);
nand U496 (N_496,N_254,In_77);
or U497 (N_497,In_622,N_317);
nand U498 (N_498,N_246,In_609);
and U499 (N_499,In_219,In_376);
nand U500 (N_500,N_347,In_144);
or U501 (N_501,In_278,N_286);
nor U502 (N_502,N_400,In_549);
nor U503 (N_503,N_47,N_440);
nor U504 (N_504,N_153,N_438);
and U505 (N_505,N_424,N_53);
nand U506 (N_506,In_776,N_427);
and U507 (N_507,N_105,N_439);
and U508 (N_508,In_449,N_442);
nor U509 (N_509,In_803,N_466);
nor U510 (N_510,N_166,In_164);
xnor U511 (N_511,N_437,N_388);
nand U512 (N_512,N_165,N_308);
and U513 (N_513,In_893,N_336);
xnor U514 (N_514,N_464,N_316);
nand U515 (N_515,N_434,In_869);
and U516 (N_516,N_477,N_250);
or U517 (N_517,In_527,N_177);
nor U518 (N_518,N_475,N_27);
and U519 (N_519,In_466,In_430);
and U520 (N_520,N_382,N_495);
nand U521 (N_521,N_368,N_224);
nor U522 (N_522,N_362,In_848);
xor U523 (N_523,N_343,In_315);
or U524 (N_524,N_494,N_229);
nor U525 (N_525,In_556,N_463);
nand U526 (N_526,In_600,N_468);
nor U527 (N_527,In_547,In_86);
and U528 (N_528,In_138,N_366);
nand U529 (N_529,In_899,In_648);
nand U530 (N_530,N_309,N_376);
nor U531 (N_531,In_879,N_194);
nor U532 (N_532,In_657,In_934);
nand U533 (N_533,N_139,N_496);
and U534 (N_534,N_208,In_746);
or U535 (N_535,N_456,N_40);
xor U536 (N_536,In_27,N_130);
and U537 (N_537,N_417,N_264);
nand U538 (N_538,In_301,In_545);
nor U539 (N_539,In_807,N_8);
xor U540 (N_540,N_344,N_425);
nor U541 (N_541,In_286,In_771);
or U542 (N_542,N_80,In_747);
xor U543 (N_543,N_81,In_247);
nor U544 (N_544,N_335,In_271);
nor U545 (N_545,N_311,N_346);
nor U546 (N_546,N_461,In_34);
nor U547 (N_547,N_315,N_474);
nor U548 (N_548,In_94,In_883);
nor U549 (N_549,N_290,In_217);
nor U550 (N_550,N_281,N_395);
or U551 (N_551,N_265,In_861);
and U552 (N_552,N_333,N_183);
nor U553 (N_553,N_231,In_875);
and U554 (N_554,In_322,In_475);
nand U555 (N_555,N_381,N_89);
nor U556 (N_556,N_460,N_206);
or U557 (N_557,In_731,In_978);
and U558 (N_558,N_287,N_471);
nor U559 (N_559,In_635,In_409);
xor U560 (N_560,N_447,N_180);
xnor U561 (N_561,N_436,N_214);
and U562 (N_562,In_677,In_569);
nand U563 (N_563,N_237,In_739);
or U564 (N_564,In_106,In_96);
xnor U565 (N_565,In_71,In_102);
nand U566 (N_566,N_384,In_185);
xor U567 (N_567,N_355,In_151);
and U568 (N_568,N_408,In_380);
nor U569 (N_569,N_41,N_251);
or U570 (N_570,In_968,N_498);
nor U571 (N_571,N_458,N_288);
or U572 (N_572,N_487,N_65);
nor U573 (N_573,N_450,N_385);
xnor U574 (N_574,In_709,N_313);
nor U575 (N_575,In_900,N_220);
nor U576 (N_576,N_245,In_87);
nor U577 (N_577,N_59,N_444);
nand U578 (N_578,In_141,N_469);
nor U579 (N_579,N_240,N_32);
and U580 (N_580,In_122,In_37);
nor U581 (N_581,In_715,N_126);
nor U582 (N_582,N_223,In_671);
xnor U583 (N_583,In_573,N_476);
nor U584 (N_584,In_370,N_369);
or U585 (N_585,In_825,N_186);
nor U586 (N_586,N_359,N_419);
nand U587 (N_587,N_181,N_446);
and U588 (N_588,In_502,N_314);
or U589 (N_589,N_230,In_758);
xor U590 (N_590,In_158,In_223);
nand U591 (N_591,In_707,In_8);
and U592 (N_592,N_449,N_323);
nand U593 (N_593,N_151,N_103);
or U594 (N_594,In_5,In_221);
or U595 (N_595,N_322,In_340);
or U596 (N_596,N_320,In_40);
and U597 (N_597,In_907,N_337);
nand U598 (N_598,In_65,N_409);
nand U599 (N_599,N_269,N_146);
nor U600 (N_600,In_917,N_465);
nand U601 (N_601,N_109,N_587);
or U602 (N_602,N_71,N_537);
nand U603 (N_603,N_292,N_564);
nand U604 (N_604,In_873,In_882);
nand U605 (N_605,N_410,N_156);
or U606 (N_606,N_594,N_391);
nand U607 (N_607,N_392,N_63);
nor U608 (N_608,N_582,In_508);
and U609 (N_609,N_524,N_560);
or U610 (N_610,N_416,In_100);
xnor U611 (N_611,N_554,N_510);
nand U612 (N_612,N_312,N_258);
nand U613 (N_613,N_462,N_285);
nor U614 (N_614,N_421,N_459);
or U615 (N_615,N_467,N_199);
and U616 (N_616,N_521,N_377);
and U617 (N_617,In_1,N_42);
and U618 (N_618,N_319,In_972);
nor U619 (N_619,N_552,N_520);
nor U620 (N_620,In_501,N_544);
or U621 (N_621,N_581,In_146);
nand U622 (N_622,In_58,N_558);
xnor U623 (N_623,N_339,In_480);
or U624 (N_624,N_293,N_301);
or U625 (N_625,N_574,In_830);
xor U626 (N_626,N_297,N_557);
or U627 (N_627,N_202,N_529);
nor U628 (N_628,N_542,In_51);
and U629 (N_629,In_610,N_546);
or U630 (N_630,N_550,N_441);
nor U631 (N_631,N_383,N_361);
or U632 (N_632,In_383,N_428);
nand U633 (N_633,N_457,In_973);
and U634 (N_634,N_595,In_226);
nand U635 (N_635,In_904,N_279);
nand U636 (N_636,In_551,In_691);
and U637 (N_637,N_549,In_416);
nand U638 (N_638,N_115,N_527);
nor U639 (N_639,In_685,In_752);
nand U640 (N_640,N_226,In_868);
nand U641 (N_641,N_448,In_961);
nor U642 (N_642,N_512,N_332);
or U643 (N_643,N_583,N_79);
nor U644 (N_644,In_813,N_481);
nor U645 (N_645,N_530,N_485);
or U646 (N_646,N_282,In_368);
nor U647 (N_647,In_10,N_144);
or U648 (N_648,N_516,N_517);
nand U649 (N_649,N_189,N_6);
and U650 (N_650,N_403,N_420);
and U651 (N_651,In_798,In_347);
or U652 (N_652,In_842,N_329);
and U653 (N_653,N_535,In_744);
nor U654 (N_654,N_110,N_586);
and U655 (N_655,N_94,In_316);
or U656 (N_656,N_592,N_114);
nor U657 (N_657,N_499,N_102);
or U658 (N_658,N_185,In_202);
nor U659 (N_659,N_591,N_536);
nor U660 (N_660,In_854,N_526);
nor U661 (N_661,N_553,N_331);
and U662 (N_662,N_484,In_936);
nor U663 (N_663,N_422,N_328);
and U664 (N_664,In_730,N_454);
nand U665 (N_665,In_683,N_193);
or U666 (N_666,In_763,In_355);
nor U667 (N_667,N_324,N_169);
and U668 (N_668,N_443,In_338);
or U669 (N_669,In_920,In_493);
nor U670 (N_670,N_596,N_402);
and U671 (N_671,In_178,In_603);
nand U672 (N_672,In_687,In_381);
nand U673 (N_673,In_129,N_399);
and U674 (N_674,In_201,N_429);
nand U675 (N_675,In_172,N_234);
nand U676 (N_676,N_215,In_399);
nand U677 (N_677,N_500,N_545);
nor U678 (N_678,N_561,In_951);
and U679 (N_679,N_472,N_431);
nand U680 (N_680,N_261,N_426);
nand U681 (N_681,In_455,In_109);
or U682 (N_682,N_508,N_480);
and U683 (N_683,N_365,N_504);
or U684 (N_684,In_612,In_465);
nand U685 (N_685,In_136,In_256);
nand U686 (N_686,N_593,In_125);
nor U687 (N_687,N_262,N_489);
nor U688 (N_688,In_855,N_543);
and U689 (N_689,N_578,N_541);
and U690 (N_690,In_857,N_555);
nor U691 (N_691,N_212,In_723);
or U692 (N_692,N_492,N_413);
xnor U693 (N_693,N_435,N_570);
nand U694 (N_694,N_551,In_75);
or U695 (N_695,N_599,N_562);
or U696 (N_696,N_490,N_473);
or U697 (N_697,N_46,N_29);
or U698 (N_698,N_161,N_514);
or U699 (N_699,N_356,N_407);
xnor U700 (N_700,N_432,N_651);
nand U701 (N_701,N_470,In_220);
or U702 (N_702,N_679,N_525);
or U703 (N_703,N_699,In_708);
or U704 (N_704,N_479,N_577);
nor U705 (N_705,In_967,N_575);
nor U706 (N_706,N_677,N_121);
or U707 (N_707,N_608,In_431);
or U708 (N_708,N_579,In_759);
or U709 (N_709,N_654,N_641);
nand U710 (N_710,N_452,N_610);
nor U711 (N_711,N_695,N_672);
or U712 (N_712,N_61,N_628);
nor U713 (N_713,N_405,N_373);
xor U714 (N_714,In_447,In_499);
nor U715 (N_715,N_686,N_358);
nor U716 (N_716,N_502,N_671);
xnor U717 (N_717,N_566,N_488);
nor U718 (N_718,N_268,N_615);
nor U719 (N_719,N_631,N_411);
nand U720 (N_720,N_572,N_160);
nor U721 (N_721,In_479,In_371);
or U722 (N_722,In_558,N_141);
or U723 (N_723,N_190,N_605);
xor U724 (N_724,In_95,N_616);
nand U725 (N_725,N_646,N_128);
nand U726 (N_726,In_352,N_270);
and U727 (N_727,In_73,N_676);
or U728 (N_728,N_600,N_604);
xnor U729 (N_729,In_241,N_614);
nand U730 (N_730,N_538,In_382);
or U731 (N_731,N_513,N_401);
nand U732 (N_732,In_997,In_939);
and U733 (N_733,N_106,N_57);
and U734 (N_734,N_272,In_565);
nand U735 (N_735,N_540,N_352);
and U736 (N_736,N_478,In_575);
nor U737 (N_737,N_283,N_580);
nand U738 (N_738,N_612,N_12);
nor U739 (N_739,N_173,N_698);
or U740 (N_740,In_190,N_637);
nand U741 (N_741,N_573,N_644);
nand U742 (N_742,N_415,N_569);
nand U743 (N_743,In_262,N_648);
xor U744 (N_744,N_406,N_305);
and U745 (N_745,N_626,N_618);
and U746 (N_746,N_639,N_433);
or U747 (N_747,N_606,N_613);
xnor U748 (N_748,N_506,N_621);
nor U749 (N_749,N_547,N_451);
nor U750 (N_750,In_23,N_325);
and U751 (N_751,N_568,In_320);
nor U752 (N_752,N_622,N_624);
nand U753 (N_753,In_736,N_197);
nor U754 (N_754,N_418,N_49);
nand U755 (N_755,N_342,N_138);
and U756 (N_756,N_455,In_953);
nor U757 (N_757,N_680,N_104);
and U758 (N_758,N_507,N_497);
and U759 (N_759,In_679,N_486);
nor U760 (N_760,N_681,N_354);
xnor U761 (N_761,N_657,N_515);
nor U762 (N_762,In_966,N_664);
xor U763 (N_763,N_493,N_633);
or U764 (N_764,N_256,N_656);
nor U765 (N_765,In_30,N_584);
and U766 (N_766,In_440,N_630);
or U767 (N_767,N_678,N_453);
and U768 (N_768,N_326,N_585);
nand U769 (N_769,N_83,In_188);
or U770 (N_770,N_51,In_32);
and U771 (N_771,N_692,N_689);
or U772 (N_772,In_819,In_173);
or U773 (N_773,N_632,N_598);
nand U774 (N_774,N_539,In_85);
nor U775 (N_775,N_99,N_696);
or U776 (N_776,N_590,N_412);
or U777 (N_777,N_263,N_667);
or U778 (N_778,In_490,N_669);
nand U779 (N_779,N_142,N_636);
nor U780 (N_780,N_645,N_394);
or U781 (N_781,N_522,N_195);
nor U782 (N_782,In_12,N_668);
nor U783 (N_783,N_482,In_341);
or U784 (N_784,In_283,N_661);
and U785 (N_785,N_567,N_653);
xnor U786 (N_786,In_298,N_602);
nor U787 (N_787,N_652,N_635);
or U788 (N_788,In_559,In_681);
xnor U789 (N_789,N_503,In_665);
or U790 (N_790,N_647,In_319);
or U791 (N_791,N_404,N_532);
xnor U792 (N_792,N_222,N_509);
and U793 (N_793,N_690,N_533);
and U794 (N_794,N_629,N_277);
and U795 (N_795,In_205,N_663);
nand U796 (N_796,In_518,N_148);
or U797 (N_797,N_374,N_518);
or U798 (N_798,N_642,N_97);
nand U799 (N_799,In_999,N_627);
or U800 (N_800,In_587,N_658);
and U801 (N_801,N_740,N_728);
nor U802 (N_802,N_620,N_747);
and U803 (N_803,N_721,N_523);
nor U804 (N_804,N_719,N_748);
nand U805 (N_805,N_125,N_609);
nor U806 (N_806,N_768,N_718);
nor U807 (N_807,N_794,N_640);
xor U808 (N_808,N_733,N_727);
xnor U809 (N_809,N_662,In_581);
nor U810 (N_810,In_385,N_773);
nor U811 (N_811,N_704,In_778);
or U812 (N_812,In_611,N_203);
and U813 (N_813,N_44,N_398);
nor U814 (N_814,N_701,N_709);
nor U815 (N_815,N_737,N_722);
and U816 (N_816,N_738,N_655);
nand U817 (N_817,N_674,N_548);
xor U818 (N_818,N_682,N_225);
and U819 (N_819,N_714,In_991);
nor U820 (N_820,N_734,N_746);
nand U821 (N_821,N_625,N_743);
nand U822 (N_822,N_729,N_753);
or U823 (N_823,N_731,N_707);
or U824 (N_824,N_163,N_796);
nor U825 (N_825,N_708,N_491);
and U826 (N_826,N_756,N_673);
and U827 (N_827,N_732,N_213);
and U828 (N_828,N_601,N_736);
and U829 (N_829,N_589,N_775);
nand U830 (N_830,N_769,N_713);
nand U831 (N_831,N_776,N_534);
and U832 (N_832,N_638,N_665);
nand U833 (N_833,N_650,N_643);
nand U834 (N_834,In_242,N_795);
or U835 (N_835,N_559,N_725);
and U836 (N_836,N_623,In_760);
nor U837 (N_837,N_783,N_685);
nor U838 (N_838,N_697,N_706);
or U839 (N_839,N_483,N_790);
or U840 (N_840,N_576,In_130);
and U841 (N_841,N_691,N_754);
nor U842 (N_842,N_563,N_675);
nor U843 (N_843,N_797,N_742);
and U844 (N_844,N_597,N_774);
nor U845 (N_845,In_891,N_371);
nand U846 (N_846,N_588,N_715);
nand U847 (N_847,N_779,In_718);
nand U848 (N_848,N_785,N_741);
or U849 (N_849,N_666,N_784);
nand U850 (N_850,N_3,N_720);
or U851 (N_851,N_703,N_724);
xor U852 (N_852,N_751,N_735);
or U853 (N_853,N_781,In_841);
nor U854 (N_854,In_120,N_670);
nor U855 (N_855,In_24,N_792);
and U856 (N_856,N_767,In_101);
or U857 (N_857,N_235,N_780);
or U858 (N_858,N_387,N_565);
or U859 (N_859,N_634,N_649);
or U860 (N_860,N_617,N_750);
nor U861 (N_861,N_798,N_705);
nor U862 (N_862,N_771,N_726);
or U863 (N_863,N_430,N_762);
and U864 (N_864,N_752,In_641);
xor U865 (N_865,In_949,In_105);
nor U866 (N_866,N_772,N_716);
and U867 (N_867,N_745,N_723);
and U868 (N_868,N_744,N_683);
and U869 (N_869,N_659,N_793);
nor U870 (N_870,N_757,N_764);
nand U871 (N_871,N_717,N_414);
nand U872 (N_872,N_505,N_519);
nand U873 (N_873,N_749,In_916);
or U874 (N_874,N_766,N_556);
and U875 (N_875,N_739,N_357);
xnor U876 (N_876,N_694,N_511);
nand U877 (N_877,N_761,In_471);
nand U878 (N_878,N_787,N_730);
xnor U879 (N_879,N_758,N_712);
nand U880 (N_880,In_326,In_865);
or U881 (N_881,N_501,N_759);
or U882 (N_882,N_755,N_799);
or U883 (N_883,N_363,N_170);
nand U884 (N_884,N_660,N_763);
nor U885 (N_885,N_531,N_791);
and U886 (N_886,N_760,N_711);
and U887 (N_887,N_777,N_619);
nor U888 (N_888,N_782,N_710);
nand U889 (N_889,N_770,N_702);
nand U890 (N_890,N_778,N_788);
or U891 (N_891,N_684,N_445);
nand U892 (N_892,N_603,N_294);
and U893 (N_893,N_607,N_789);
or U894 (N_894,N_693,N_700);
or U895 (N_895,N_243,N_687);
nand U896 (N_896,N_786,N_423);
or U897 (N_897,N_611,N_765);
nand U898 (N_898,N_528,N_688);
xnor U899 (N_899,N_571,N_307);
and U900 (N_900,N_871,N_895);
nand U901 (N_901,N_834,N_827);
nand U902 (N_902,N_868,N_858);
and U903 (N_903,N_887,N_814);
xor U904 (N_904,N_864,N_846);
and U905 (N_905,N_855,N_844);
or U906 (N_906,N_815,N_883);
nor U907 (N_907,N_802,N_831);
nand U908 (N_908,N_836,N_841);
or U909 (N_909,N_897,N_892);
and U910 (N_910,N_854,N_866);
nand U911 (N_911,N_879,N_817);
and U912 (N_912,N_851,N_804);
xor U913 (N_913,N_820,N_806);
or U914 (N_914,N_852,N_878);
and U915 (N_915,N_899,N_875);
nor U916 (N_916,N_853,N_889);
or U917 (N_917,N_888,N_821);
nand U918 (N_918,N_850,N_891);
or U919 (N_919,N_828,N_819);
nand U920 (N_920,N_863,N_812);
and U921 (N_921,N_876,N_823);
and U922 (N_922,N_893,N_825);
nor U923 (N_923,N_898,N_816);
nor U924 (N_924,N_837,N_881);
or U925 (N_925,N_890,N_860);
or U926 (N_926,N_809,N_859);
nor U927 (N_927,N_873,N_849);
and U928 (N_928,N_877,N_856);
nand U929 (N_929,N_848,N_861);
and U930 (N_930,N_896,N_808);
and U931 (N_931,N_839,N_800);
or U932 (N_932,N_880,N_805);
or U933 (N_933,N_832,N_838);
and U934 (N_934,N_865,N_840);
nor U935 (N_935,N_835,N_842);
nand U936 (N_936,N_826,N_807);
and U937 (N_937,N_885,N_829);
nor U938 (N_938,N_886,N_872);
nor U939 (N_939,N_894,N_884);
and U940 (N_940,N_869,N_870);
or U941 (N_941,N_843,N_824);
or U942 (N_942,N_833,N_811);
nor U943 (N_943,N_803,N_830);
xor U944 (N_944,N_862,N_857);
or U945 (N_945,N_847,N_810);
nand U946 (N_946,N_867,N_882);
xnor U947 (N_947,N_801,N_813);
nor U948 (N_948,N_845,N_874);
nor U949 (N_949,N_818,N_822);
xor U950 (N_950,N_895,N_843);
nor U951 (N_951,N_875,N_879);
or U952 (N_952,N_897,N_818);
or U953 (N_953,N_836,N_879);
or U954 (N_954,N_853,N_856);
or U955 (N_955,N_815,N_840);
xor U956 (N_956,N_853,N_804);
nand U957 (N_957,N_880,N_827);
and U958 (N_958,N_885,N_825);
or U959 (N_959,N_811,N_844);
and U960 (N_960,N_831,N_896);
nand U961 (N_961,N_839,N_870);
and U962 (N_962,N_882,N_849);
xnor U963 (N_963,N_864,N_810);
or U964 (N_964,N_884,N_864);
or U965 (N_965,N_876,N_812);
nand U966 (N_966,N_840,N_898);
nor U967 (N_967,N_869,N_816);
and U968 (N_968,N_864,N_866);
nor U969 (N_969,N_879,N_891);
nor U970 (N_970,N_835,N_860);
nand U971 (N_971,N_876,N_818);
nor U972 (N_972,N_806,N_866);
and U973 (N_973,N_870,N_885);
nor U974 (N_974,N_819,N_868);
nor U975 (N_975,N_870,N_891);
nand U976 (N_976,N_806,N_886);
nor U977 (N_977,N_828,N_897);
nor U978 (N_978,N_818,N_815);
and U979 (N_979,N_847,N_886);
nand U980 (N_980,N_836,N_814);
nand U981 (N_981,N_883,N_800);
or U982 (N_982,N_832,N_853);
nand U983 (N_983,N_810,N_870);
nor U984 (N_984,N_873,N_822);
nor U985 (N_985,N_873,N_883);
nor U986 (N_986,N_809,N_862);
xnor U987 (N_987,N_852,N_853);
and U988 (N_988,N_821,N_839);
xnor U989 (N_989,N_891,N_877);
and U990 (N_990,N_813,N_857);
nand U991 (N_991,N_815,N_889);
nand U992 (N_992,N_825,N_827);
xor U993 (N_993,N_872,N_834);
nand U994 (N_994,N_832,N_855);
and U995 (N_995,N_810,N_807);
nor U996 (N_996,N_874,N_829);
or U997 (N_997,N_832,N_860);
xnor U998 (N_998,N_898,N_804);
and U999 (N_999,N_810,N_884);
or U1000 (N_1000,N_903,N_994);
nand U1001 (N_1001,N_968,N_999);
and U1002 (N_1002,N_938,N_974);
and U1003 (N_1003,N_904,N_939);
xnor U1004 (N_1004,N_911,N_922);
or U1005 (N_1005,N_998,N_929);
or U1006 (N_1006,N_918,N_983);
nand U1007 (N_1007,N_957,N_991);
or U1008 (N_1008,N_978,N_937);
or U1009 (N_1009,N_934,N_984);
nand U1010 (N_1010,N_928,N_945);
or U1011 (N_1011,N_956,N_959);
nor U1012 (N_1012,N_988,N_990);
nor U1013 (N_1013,N_950,N_920);
or U1014 (N_1014,N_917,N_923);
xnor U1015 (N_1015,N_931,N_935);
nand U1016 (N_1016,N_985,N_912);
nor U1017 (N_1017,N_947,N_952);
and U1018 (N_1018,N_976,N_973);
or U1019 (N_1019,N_986,N_961);
or U1020 (N_1020,N_967,N_936);
and U1021 (N_1021,N_906,N_948);
nand U1022 (N_1022,N_966,N_942);
and U1023 (N_1023,N_930,N_979);
and U1024 (N_1024,N_981,N_971);
nor U1025 (N_1025,N_989,N_905);
and U1026 (N_1026,N_946,N_995);
nand U1027 (N_1027,N_970,N_933);
xor U1028 (N_1028,N_982,N_914);
and U1029 (N_1029,N_907,N_975);
nor U1030 (N_1030,N_943,N_964);
or U1031 (N_1031,N_962,N_915);
and U1032 (N_1032,N_908,N_963);
and U1033 (N_1033,N_954,N_924);
nor U1034 (N_1034,N_926,N_960);
and U1035 (N_1035,N_900,N_941);
and U1036 (N_1036,N_965,N_972);
nand U1037 (N_1037,N_913,N_901);
or U1038 (N_1038,N_902,N_916);
xnor U1039 (N_1039,N_925,N_909);
nand U1040 (N_1040,N_949,N_940);
nor U1041 (N_1041,N_969,N_993);
and U1042 (N_1042,N_944,N_977);
nand U1043 (N_1043,N_919,N_996);
or U1044 (N_1044,N_921,N_992);
nand U1045 (N_1045,N_958,N_927);
and U1046 (N_1046,N_987,N_953);
nand U1047 (N_1047,N_951,N_955);
nand U1048 (N_1048,N_932,N_910);
or U1049 (N_1049,N_980,N_997);
nor U1050 (N_1050,N_993,N_912);
and U1051 (N_1051,N_926,N_971);
and U1052 (N_1052,N_986,N_927);
and U1053 (N_1053,N_917,N_938);
and U1054 (N_1054,N_928,N_919);
or U1055 (N_1055,N_911,N_994);
or U1056 (N_1056,N_928,N_938);
nand U1057 (N_1057,N_900,N_989);
or U1058 (N_1058,N_975,N_912);
and U1059 (N_1059,N_986,N_985);
and U1060 (N_1060,N_955,N_972);
nor U1061 (N_1061,N_947,N_961);
and U1062 (N_1062,N_908,N_902);
or U1063 (N_1063,N_907,N_935);
and U1064 (N_1064,N_937,N_910);
or U1065 (N_1065,N_952,N_974);
or U1066 (N_1066,N_940,N_995);
or U1067 (N_1067,N_904,N_968);
xor U1068 (N_1068,N_927,N_976);
xor U1069 (N_1069,N_934,N_948);
and U1070 (N_1070,N_968,N_952);
nor U1071 (N_1071,N_914,N_918);
or U1072 (N_1072,N_904,N_910);
nor U1073 (N_1073,N_994,N_906);
nand U1074 (N_1074,N_951,N_953);
and U1075 (N_1075,N_972,N_995);
xor U1076 (N_1076,N_982,N_953);
and U1077 (N_1077,N_937,N_932);
or U1078 (N_1078,N_952,N_950);
nand U1079 (N_1079,N_950,N_978);
nand U1080 (N_1080,N_905,N_954);
nand U1081 (N_1081,N_979,N_907);
nor U1082 (N_1082,N_950,N_979);
xnor U1083 (N_1083,N_958,N_955);
or U1084 (N_1084,N_944,N_916);
nand U1085 (N_1085,N_979,N_928);
and U1086 (N_1086,N_993,N_979);
nand U1087 (N_1087,N_964,N_976);
and U1088 (N_1088,N_900,N_916);
and U1089 (N_1089,N_931,N_978);
or U1090 (N_1090,N_968,N_953);
and U1091 (N_1091,N_954,N_994);
and U1092 (N_1092,N_910,N_940);
nor U1093 (N_1093,N_922,N_983);
or U1094 (N_1094,N_973,N_912);
or U1095 (N_1095,N_980,N_910);
or U1096 (N_1096,N_944,N_929);
and U1097 (N_1097,N_904,N_957);
nand U1098 (N_1098,N_985,N_929);
and U1099 (N_1099,N_992,N_987);
nand U1100 (N_1100,N_1083,N_1037);
nand U1101 (N_1101,N_1097,N_1098);
nand U1102 (N_1102,N_1054,N_1024);
nand U1103 (N_1103,N_1022,N_1034);
or U1104 (N_1104,N_1011,N_1018);
and U1105 (N_1105,N_1073,N_1081);
nand U1106 (N_1106,N_1046,N_1093);
nand U1107 (N_1107,N_1056,N_1033);
nand U1108 (N_1108,N_1091,N_1087);
nand U1109 (N_1109,N_1031,N_1029);
nand U1110 (N_1110,N_1021,N_1064);
or U1111 (N_1111,N_1045,N_1027);
or U1112 (N_1112,N_1025,N_1089);
or U1113 (N_1113,N_1012,N_1032);
xor U1114 (N_1114,N_1006,N_1069);
and U1115 (N_1115,N_1079,N_1071);
xnor U1116 (N_1116,N_1058,N_1043);
and U1117 (N_1117,N_1020,N_1044);
nand U1118 (N_1118,N_1062,N_1059);
nand U1119 (N_1119,N_1035,N_1070);
nor U1120 (N_1120,N_1092,N_1082);
and U1121 (N_1121,N_1023,N_1036);
and U1122 (N_1122,N_1026,N_1077);
and U1123 (N_1123,N_1051,N_1055);
nand U1124 (N_1124,N_1075,N_1017);
nand U1125 (N_1125,N_1090,N_1001);
xnor U1126 (N_1126,N_1039,N_1084);
and U1127 (N_1127,N_1004,N_1067);
and U1128 (N_1128,N_1072,N_1050);
and U1129 (N_1129,N_1040,N_1053);
nand U1130 (N_1130,N_1038,N_1048);
nand U1131 (N_1131,N_1085,N_1009);
nand U1132 (N_1132,N_1003,N_1095);
nor U1133 (N_1133,N_1099,N_1010);
nand U1134 (N_1134,N_1000,N_1014);
nand U1135 (N_1135,N_1008,N_1078);
or U1136 (N_1136,N_1063,N_1065);
xnor U1137 (N_1137,N_1061,N_1088);
xnor U1138 (N_1138,N_1066,N_1002);
and U1139 (N_1139,N_1019,N_1076);
xnor U1140 (N_1140,N_1086,N_1060);
or U1141 (N_1141,N_1068,N_1052);
nand U1142 (N_1142,N_1015,N_1049);
xnor U1143 (N_1143,N_1057,N_1007);
nor U1144 (N_1144,N_1094,N_1042);
nand U1145 (N_1145,N_1074,N_1028);
nor U1146 (N_1146,N_1005,N_1096);
or U1147 (N_1147,N_1047,N_1030);
or U1148 (N_1148,N_1080,N_1041);
nor U1149 (N_1149,N_1013,N_1016);
and U1150 (N_1150,N_1005,N_1089);
and U1151 (N_1151,N_1063,N_1015);
or U1152 (N_1152,N_1086,N_1044);
nor U1153 (N_1153,N_1070,N_1044);
and U1154 (N_1154,N_1057,N_1051);
nor U1155 (N_1155,N_1062,N_1037);
nor U1156 (N_1156,N_1038,N_1093);
or U1157 (N_1157,N_1088,N_1023);
nor U1158 (N_1158,N_1018,N_1022);
nand U1159 (N_1159,N_1021,N_1056);
or U1160 (N_1160,N_1091,N_1001);
and U1161 (N_1161,N_1039,N_1089);
xor U1162 (N_1162,N_1080,N_1036);
and U1163 (N_1163,N_1095,N_1087);
or U1164 (N_1164,N_1079,N_1097);
or U1165 (N_1165,N_1028,N_1058);
or U1166 (N_1166,N_1071,N_1088);
nor U1167 (N_1167,N_1044,N_1060);
or U1168 (N_1168,N_1093,N_1091);
nand U1169 (N_1169,N_1067,N_1083);
or U1170 (N_1170,N_1094,N_1036);
and U1171 (N_1171,N_1054,N_1066);
nor U1172 (N_1172,N_1076,N_1089);
or U1173 (N_1173,N_1045,N_1012);
nand U1174 (N_1174,N_1085,N_1038);
xnor U1175 (N_1175,N_1055,N_1097);
nor U1176 (N_1176,N_1024,N_1033);
nor U1177 (N_1177,N_1072,N_1090);
nor U1178 (N_1178,N_1065,N_1028);
or U1179 (N_1179,N_1080,N_1081);
and U1180 (N_1180,N_1014,N_1036);
and U1181 (N_1181,N_1063,N_1084);
nand U1182 (N_1182,N_1005,N_1077);
nor U1183 (N_1183,N_1030,N_1087);
and U1184 (N_1184,N_1006,N_1029);
nand U1185 (N_1185,N_1055,N_1047);
xor U1186 (N_1186,N_1032,N_1078);
or U1187 (N_1187,N_1002,N_1036);
and U1188 (N_1188,N_1090,N_1006);
nand U1189 (N_1189,N_1000,N_1012);
nand U1190 (N_1190,N_1001,N_1004);
nor U1191 (N_1191,N_1068,N_1030);
nand U1192 (N_1192,N_1078,N_1061);
and U1193 (N_1193,N_1065,N_1094);
and U1194 (N_1194,N_1063,N_1040);
and U1195 (N_1195,N_1003,N_1091);
nand U1196 (N_1196,N_1095,N_1036);
nand U1197 (N_1197,N_1069,N_1067);
or U1198 (N_1198,N_1057,N_1017);
and U1199 (N_1199,N_1001,N_1096);
xor U1200 (N_1200,N_1190,N_1177);
or U1201 (N_1201,N_1109,N_1175);
nor U1202 (N_1202,N_1164,N_1163);
and U1203 (N_1203,N_1181,N_1193);
and U1204 (N_1204,N_1130,N_1159);
or U1205 (N_1205,N_1150,N_1113);
or U1206 (N_1206,N_1155,N_1172);
nand U1207 (N_1207,N_1180,N_1171);
nand U1208 (N_1208,N_1126,N_1186);
or U1209 (N_1209,N_1120,N_1185);
nor U1210 (N_1210,N_1197,N_1161);
and U1211 (N_1211,N_1147,N_1129);
and U1212 (N_1212,N_1116,N_1145);
nor U1213 (N_1213,N_1140,N_1138);
or U1214 (N_1214,N_1187,N_1143);
or U1215 (N_1215,N_1198,N_1174);
or U1216 (N_1216,N_1112,N_1128);
nor U1217 (N_1217,N_1169,N_1142);
nor U1218 (N_1218,N_1101,N_1141);
nor U1219 (N_1219,N_1144,N_1196);
nor U1220 (N_1220,N_1139,N_1122);
xnor U1221 (N_1221,N_1157,N_1106);
nor U1222 (N_1222,N_1107,N_1132);
and U1223 (N_1223,N_1123,N_1182);
nor U1224 (N_1224,N_1184,N_1160);
nor U1225 (N_1225,N_1119,N_1158);
nand U1226 (N_1226,N_1121,N_1195);
nor U1227 (N_1227,N_1102,N_1166);
nor U1228 (N_1228,N_1194,N_1148);
nor U1229 (N_1229,N_1156,N_1191);
nand U1230 (N_1230,N_1134,N_1168);
nor U1231 (N_1231,N_1127,N_1162);
nand U1232 (N_1232,N_1173,N_1170);
nor U1233 (N_1233,N_1183,N_1110);
and U1234 (N_1234,N_1176,N_1137);
nand U1235 (N_1235,N_1146,N_1111);
and U1236 (N_1236,N_1192,N_1188);
nand U1237 (N_1237,N_1178,N_1153);
nand U1238 (N_1238,N_1189,N_1151);
nand U1239 (N_1239,N_1114,N_1199);
and U1240 (N_1240,N_1125,N_1136);
nand U1241 (N_1241,N_1100,N_1154);
or U1242 (N_1242,N_1108,N_1117);
and U1243 (N_1243,N_1124,N_1104);
nor U1244 (N_1244,N_1167,N_1149);
or U1245 (N_1245,N_1179,N_1152);
nand U1246 (N_1246,N_1131,N_1133);
xnor U1247 (N_1247,N_1115,N_1135);
and U1248 (N_1248,N_1105,N_1118);
nor U1249 (N_1249,N_1165,N_1103);
or U1250 (N_1250,N_1103,N_1161);
nor U1251 (N_1251,N_1163,N_1155);
and U1252 (N_1252,N_1186,N_1151);
nand U1253 (N_1253,N_1110,N_1137);
or U1254 (N_1254,N_1163,N_1181);
and U1255 (N_1255,N_1113,N_1186);
nor U1256 (N_1256,N_1154,N_1195);
and U1257 (N_1257,N_1178,N_1105);
xor U1258 (N_1258,N_1102,N_1138);
or U1259 (N_1259,N_1190,N_1199);
xor U1260 (N_1260,N_1189,N_1167);
and U1261 (N_1261,N_1196,N_1189);
nor U1262 (N_1262,N_1181,N_1188);
xnor U1263 (N_1263,N_1156,N_1132);
or U1264 (N_1264,N_1176,N_1157);
xor U1265 (N_1265,N_1144,N_1149);
nor U1266 (N_1266,N_1164,N_1140);
nand U1267 (N_1267,N_1184,N_1112);
nand U1268 (N_1268,N_1175,N_1121);
nand U1269 (N_1269,N_1162,N_1185);
nand U1270 (N_1270,N_1170,N_1186);
nor U1271 (N_1271,N_1128,N_1175);
nor U1272 (N_1272,N_1184,N_1161);
nor U1273 (N_1273,N_1199,N_1105);
nor U1274 (N_1274,N_1179,N_1115);
and U1275 (N_1275,N_1142,N_1128);
nor U1276 (N_1276,N_1162,N_1173);
nor U1277 (N_1277,N_1112,N_1114);
nand U1278 (N_1278,N_1133,N_1128);
or U1279 (N_1279,N_1123,N_1130);
and U1280 (N_1280,N_1169,N_1149);
xnor U1281 (N_1281,N_1123,N_1100);
or U1282 (N_1282,N_1186,N_1149);
xor U1283 (N_1283,N_1125,N_1176);
nand U1284 (N_1284,N_1178,N_1130);
or U1285 (N_1285,N_1112,N_1193);
nand U1286 (N_1286,N_1137,N_1136);
and U1287 (N_1287,N_1196,N_1139);
nor U1288 (N_1288,N_1153,N_1114);
nand U1289 (N_1289,N_1179,N_1160);
nor U1290 (N_1290,N_1130,N_1195);
and U1291 (N_1291,N_1110,N_1169);
nor U1292 (N_1292,N_1104,N_1195);
and U1293 (N_1293,N_1148,N_1175);
and U1294 (N_1294,N_1135,N_1192);
or U1295 (N_1295,N_1103,N_1143);
nand U1296 (N_1296,N_1129,N_1103);
and U1297 (N_1297,N_1144,N_1130);
or U1298 (N_1298,N_1132,N_1118);
xor U1299 (N_1299,N_1147,N_1132);
or U1300 (N_1300,N_1226,N_1299);
nor U1301 (N_1301,N_1268,N_1256);
nand U1302 (N_1302,N_1244,N_1223);
nand U1303 (N_1303,N_1251,N_1267);
or U1304 (N_1304,N_1237,N_1235);
and U1305 (N_1305,N_1273,N_1284);
and U1306 (N_1306,N_1288,N_1240);
nor U1307 (N_1307,N_1261,N_1220);
nand U1308 (N_1308,N_1266,N_1215);
and U1309 (N_1309,N_1227,N_1286);
or U1310 (N_1310,N_1278,N_1296);
xor U1311 (N_1311,N_1293,N_1243);
or U1312 (N_1312,N_1276,N_1269);
and U1313 (N_1313,N_1291,N_1208);
nand U1314 (N_1314,N_1211,N_1247);
nand U1315 (N_1315,N_1217,N_1242);
or U1316 (N_1316,N_1241,N_1230);
nor U1317 (N_1317,N_1271,N_1232);
nor U1318 (N_1318,N_1249,N_1265);
nand U1319 (N_1319,N_1287,N_1231);
or U1320 (N_1320,N_1238,N_1257);
nand U1321 (N_1321,N_1280,N_1260);
and U1322 (N_1322,N_1216,N_1283);
nand U1323 (N_1323,N_1200,N_1279);
nand U1324 (N_1324,N_1209,N_1262);
or U1325 (N_1325,N_1253,N_1203);
nor U1326 (N_1326,N_1229,N_1285);
or U1327 (N_1327,N_1206,N_1290);
nor U1328 (N_1328,N_1282,N_1221);
xor U1329 (N_1329,N_1225,N_1245);
nand U1330 (N_1330,N_1254,N_1259);
and U1331 (N_1331,N_1252,N_1246);
and U1332 (N_1332,N_1239,N_1250);
or U1333 (N_1333,N_1264,N_1201);
nor U1334 (N_1334,N_1219,N_1263);
nor U1335 (N_1335,N_1210,N_1289);
or U1336 (N_1336,N_1295,N_1272);
nand U1337 (N_1337,N_1228,N_1212);
or U1338 (N_1338,N_1204,N_1281);
nor U1339 (N_1339,N_1255,N_1202);
nand U1340 (N_1340,N_1236,N_1233);
nor U1341 (N_1341,N_1218,N_1294);
nor U1342 (N_1342,N_1224,N_1222);
nand U1343 (N_1343,N_1298,N_1274);
and U1344 (N_1344,N_1213,N_1258);
or U1345 (N_1345,N_1234,N_1270);
or U1346 (N_1346,N_1214,N_1275);
xor U1347 (N_1347,N_1248,N_1207);
xnor U1348 (N_1348,N_1297,N_1292);
and U1349 (N_1349,N_1277,N_1205);
or U1350 (N_1350,N_1243,N_1269);
and U1351 (N_1351,N_1227,N_1234);
nor U1352 (N_1352,N_1205,N_1219);
nor U1353 (N_1353,N_1203,N_1220);
and U1354 (N_1354,N_1200,N_1263);
and U1355 (N_1355,N_1258,N_1249);
nand U1356 (N_1356,N_1237,N_1231);
xor U1357 (N_1357,N_1200,N_1259);
nor U1358 (N_1358,N_1251,N_1285);
xor U1359 (N_1359,N_1208,N_1253);
and U1360 (N_1360,N_1257,N_1243);
nand U1361 (N_1361,N_1254,N_1274);
nor U1362 (N_1362,N_1271,N_1259);
nor U1363 (N_1363,N_1252,N_1214);
and U1364 (N_1364,N_1241,N_1281);
or U1365 (N_1365,N_1212,N_1205);
nor U1366 (N_1366,N_1248,N_1298);
or U1367 (N_1367,N_1233,N_1282);
nand U1368 (N_1368,N_1209,N_1223);
nor U1369 (N_1369,N_1253,N_1258);
and U1370 (N_1370,N_1216,N_1251);
nand U1371 (N_1371,N_1265,N_1241);
or U1372 (N_1372,N_1239,N_1296);
nor U1373 (N_1373,N_1203,N_1297);
nand U1374 (N_1374,N_1284,N_1282);
nand U1375 (N_1375,N_1207,N_1273);
and U1376 (N_1376,N_1270,N_1226);
nand U1377 (N_1377,N_1272,N_1260);
or U1378 (N_1378,N_1282,N_1269);
or U1379 (N_1379,N_1262,N_1283);
nor U1380 (N_1380,N_1277,N_1214);
nor U1381 (N_1381,N_1247,N_1241);
and U1382 (N_1382,N_1275,N_1233);
nand U1383 (N_1383,N_1256,N_1272);
and U1384 (N_1384,N_1268,N_1283);
nor U1385 (N_1385,N_1235,N_1266);
nor U1386 (N_1386,N_1201,N_1276);
and U1387 (N_1387,N_1250,N_1252);
nor U1388 (N_1388,N_1253,N_1256);
or U1389 (N_1389,N_1266,N_1212);
or U1390 (N_1390,N_1291,N_1235);
nand U1391 (N_1391,N_1244,N_1219);
nand U1392 (N_1392,N_1218,N_1210);
nand U1393 (N_1393,N_1248,N_1234);
nand U1394 (N_1394,N_1240,N_1276);
or U1395 (N_1395,N_1212,N_1203);
xor U1396 (N_1396,N_1276,N_1259);
or U1397 (N_1397,N_1231,N_1224);
xnor U1398 (N_1398,N_1237,N_1209);
xor U1399 (N_1399,N_1221,N_1204);
nand U1400 (N_1400,N_1334,N_1306);
and U1401 (N_1401,N_1369,N_1300);
or U1402 (N_1402,N_1387,N_1338);
nor U1403 (N_1403,N_1316,N_1314);
nand U1404 (N_1404,N_1392,N_1303);
or U1405 (N_1405,N_1361,N_1301);
or U1406 (N_1406,N_1310,N_1399);
nand U1407 (N_1407,N_1371,N_1332);
and U1408 (N_1408,N_1329,N_1370);
xor U1409 (N_1409,N_1317,N_1323);
nand U1410 (N_1410,N_1379,N_1322);
nand U1411 (N_1411,N_1360,N_1340);
nand U1412 (N_1412,N_1335,N_1354);
xnor U1413 (N_1413,N_1320,N_1385);
xor U1414 (N_1414,N_1345,N_1368);
and U1415 (N_1415,N_1365,N_1355);
nor U1416 (N_1416,N_1337,N_1367);
nand U1417 (N_1417,N_1321,N_1395);
nor U1418 (N_1418,N_1344,N_1357);
nor U1419 (N_1419,N_1394,N_1393);
and U1420 (N_1420,N_1347,N_1326);
nand U1421 (N_1421,N_1389,N_1325);
and U1422 (N_1422,N_1336,N_1311);
nand U1423 (N_1423,N_1388,N_1362);
nand U1424 (N_1424,N_1346,N_1398);
nor U1425 (N_1425,N_1312,N_1380);
or U1426 (N_1426,N_1328,N_1353);
nand U1427 (N_1427,N_1318,N_1356);
xnor U1428 (N_1428,N_1373,N_1302);
xor U1429 (N_1429,N_1330,N_1366);
nand U1430 (N_1430,N_1382,N_1339);
or U1431 (N_1431,N_1364,N_1351);
nand U1432 (N_1432,N_1341,N_1363);
nand U1433 (N_1433,N_1350,N_1324);
nor U1434 (N_1434,N_1304,N_1307);
nand U1435 (N_1435,N_1383,N_1396);
and U1436 (N_1436,N_1333,N_1359);
or U1437 (N_1437,N_1381,N_1384);
and U1438 (N_1438,N_1352,N_1331);
and U1439 (N_1439,N_1376,N_1315);
and U1440 (N_1440,N_1319,N_1313);
or U1441 (N_1441,N_1343,N_1386);
and U1442 (N_1442,N_1342,N_1358);
nor U1443 (N_1443,N_1397,N_1327);
or U1444 (N_1444,N_1375,N_1349);
xor U1445 (N_1445,N_1305,N_1390);
xnor U1446 (N_1446,N_1309,N_1372);
and U1447 (N_1447,N_1348,N_1378);
nand U1448 (N_1448,N_1374,N_1377);
or U1449 (N_1449,N_1391,N_1308);
nand U1450 (N_1450,N_1337,N_1300);
nand U1451 (N_1451,N_1385,N_1347);
nor U1452 (N_1452,N_1334,N_1394);
nor U1453 (N_1453,N_1305,N_1357);
nor U1454 (N_1454,N_1366,N_1358);
or U1455 (N_1455,N_1358,N_1354);
or U1456 (N_1456,N_1358,N_1340);
nor U1457 (N_1457,N_1310,N_1300);
and U1458 (N_1458,N_1395,N_1381);
or U1459 (N_1459,N_1334,N_1354);
and U1460 (N_1460,N_1304,N_1384);
or U1461 (N_1461,N_1361,N_1381);
nand U1462 (N_1462,N_1323,N_1395);
or U1463 (N_1463,N_1355,N_1361);
or U1464 (N_1464,N_1365,N_1316);
xor U1465 (N_1465,N_1392,N_1338);
nor U1466 (N_1466,N_1336,N_1304);
or U1467 (N_1467,N_1398,N_1331);
nand U1468 (N_1468,N_1389,N_1356);
nand U1469 (N_1469,N_1365,N_1304);
nor U1470 (N_1470,N_1333,N_1329);
nor U1471 (N_1471,N_1317,N_1392);
nor U1472 (N_1472,N_1300,N_1323);
nand U1473 (N_1473,N_1386,N_1356);
or U1474 (N_1474,N_1341,N_1322);
or U1475 (N_1475,N_1366,N_1398);
or U1476 (N_1476,N_1346,N_1370);
and U1477 (N_1477,N_1339,N_1397);
xor U1478 (N_1478,N_1349,N_1399);
nand U1479 (N_1479,N_1372,N_1398);
or U1480 (N_1480,N_1317,N_1332);
nor U1481 (N_1481,N_1344,N_1300);
nor U1482 (N_1482,N_1374,N_1310);
nand U1483 (N_1483,N_1386,N_1398);
or U1484 (N_1484,N_1302,N_1329);
xor U1485 (N_1485,N_1309,N_1365);
or U1486 (N_1486,N_1381,N_1313);
or U1487 (N_1487,N_1370,N_1369);
nand U1488 (N_1488,N_1373,N_1318);
and U1489 (N_1489,N_1378,N_1398);
or U1490 (N_1490,N_1312,N_1365);
or U1491 (N_1491,N_1399,N_1348);
nand U1492 (N_1492,N_1346,N_1317);
nor U1493 (N_1493,N_1377,N_1317);
and U1494 (N_1494,N_1379,N_1362);
nand U1495 (N_1495,N_1357,N_1312);
xnor U1496 (N_1496,N_1314,N_1353);
nor U1497 (N_1497,N_1314,N_1393);
nand U1498 (N_1498,N_1344,N_1386);
nor U1499 (N_1499,N_1359,N_1324);
and U1500 (N_1500,N_1434,N_1467);
nand U1501 (N_1501,N_1490,N_1465);
and U1502 (N_1502,N_1403,N_1404);
nand U1503 (N_1503,N_1401,N_1417);
or U1504 (N_1504,N_1469,N_1462);
nor U1505 (N_1505,N_1479,N_1489);
and U1506 (N_1506,N_1414,N_1416);
nand U1507 (N_1507,N_1487,N_1450);
nand U1508 (N_1508,N_1448,N_1423);
or U1509 (N_1509,N_1419,N_1443);
nand U1510 (N_1510,N_1494,N_1439);
nand U1511 (N_1511,N_1440,N_1485);
and U1512 (N_1512,N_1430,N_1429);
xnor U1513 (N_1513,N_1484,N_1455);
or U1514 (N_1514,N_1459,N_1413);
nand U1515 (N_1515,N_1463,N_1495);
and U1516 (N_1516,N_1402,N_1478);
nor U1517 (N_1517,N_1497,N_1405);
xor U1518 (N_1518,N_1492,N_1410);
nand U1519 (N_1519,N_1438,N_1431);
nand U1520 (N_1520,N_1436,N_1483);
xor U1521 (N_1521,N_1464,N_1482);
and U1522 (N_1522,N_1493,N_1433);
or U1523 (N_1523,N_1426,N_1421);
xor U1524 (N_1524,N_1418,N_1411);
nor U1525 (N_1525,N_1437,N_1461);
xor U1526 (N_1526,N_1488,N_1491);
xor U1527 (N_1527,N_1474,N_1468);
or U1528 (N_1528,N_1460,N_1432);
nand U1529 (N_1529,N_1452,N_1415);
nand U1530 (N_1530,N_1480,N_1466);
nor U1531 (N_1531,N_1435,N_1424);
or U1532 (N_1532,N_1451,N_1454);
xor U1533 (N_1533,N_1412,N_1473);
and U1534 (N_1534,N_1499,N_1444);
nand U1535 (N_1535,N_1445,N_1400);
or U1536 (N_1536,N_1481,N_1420);
xor U1537 (N_1537,N_1425,N_1427);
or U1538 (N_1538,N_1447,N_1476);
or U1539 (N_1539,N_1496,N_1470);
or U1540 (N_1540,N_1453,N_1408);
xnor U1541 (N_1541,N_1449,N_1486);
nand U1542 (N_1542,N_1458,N_1442);
nor U1543 (N_1543,N_1457,N_1498);
xor U1544 (N_1544,N_1477,N_1407);
nand U1545 (N_1545,N_1472,N_1441);
or U1546 (N_1546,N_1456,N_1446);
nand U1547 (N_1547,N_1422,N_1406);
or U1548 (N_1548,N_1475,N_1409);
or U1549 (N_1549,N_1428,N_1471);
or U1550 (N_1550,N_1453,N_1479);
nand U1551 (N_1551,N_1476,N_1473);
nor U1552 (N_1552,N_1442,N_1470);
or U1553 (N_1553,N_1440,N_1435);
and U1554 (N_1554,N_1413,N_1408);
and U1555 (N_1555,N_1469,N_1486);
nand U1556 (N_1556,N_1459,N_1488);
nand U1557 (N_1557,N_1430,N_1457);
nand U1558 (N_1558,N_1402,N_1492);
or U1559 (N_1559,N_1432,N_1406);
nor U1560 (N_1560,N_1449,N_1488);
and U1561 (N_1561,N_1401,N_1447);
or U1562 (N_1562,N_1462,N_1439);
xor U1563 (N_1563,N_1486,N_1413);
or U1564 (N_1564,N_1470,N_1456);
and U1565 (N_1565,N_1475,N_1415);
or U1566 (N_1566,N_1430,N_1470);
nor U1567 (N_1567,N_1475,N_1429);
nor U1568 (N_1568,N_1444,N_1492);
and U1569 (N_1569,N_1415,N_1460);
or U1570 (N_1570,N_1486,N_1466);
xnor U1571 (N_1571,N_1439,N_1466);
or U1572 (N_1572,N_1449,N_1479);
and U1573 (N_1573,N_1405,N_1483);
or U1574 (N_1574,N_1406,N_1449);
or U1575 (N_1575,N_1412,N_1417);
or U1576 (N_1576,N_1455,N_1422);
or U1577 (N_1577,N_1411,N_1468);
nor U1578 (N_1578,N_1446,N_1452);
nand U1579 (N_1579,N_1498,N_1465);
nand U1580 (N_1580,N_1474,N_1498);
nand U1581 (N_1581,N_1460,N_1442);
nand U1582 (N_1582,N_1481,N_1400);
nand U1583 (N_1583,N_1436,N_1449);
nand U1584 (N_1584,N_1489,N_1464);
and U1585 (N_1585,N_1415,N_1494);
xor U1586 (N_1586,N_1477,N_1473);
and U1587 (N_1587,N_1428,N_1409);
nand U1588 (N_1588,N_1401,N_1438);
and U1589 (N_1589,N_1437,N_1497);
xnor U1590 (N_1590,N_1400,N_1418);
nor U1591 (N_1591,N_1436,N_1462);
nor U1592 (N_1592,N_1456,N_1472);
and U1593 (N_1593,N_1467,N_1453);
nand U1594 (N_1594,N_1464,N_1406);
xnor U1595 (N_1595,N_1498,N_1488);
and U1596 (N_1596,N_1428,N_1489);
xor U1597 (N_1597,N_1491,N_1432);
nor U1598 (N_1598,N_1451,N_1446);
or U1599 (N_1599,N_1490,N_1454);
and U1600 (N_1600,N_1560,N_1556);
and U1601 (N_1601,N_1562,N_1504);
nor U1602 (N_1602,N_1518,N_1580);
or U1603 (N_1603,N_1500,N_1512);
or U1604 (N_1604,N_1584,N_1525);
and U1605 (N_1605,N_1573,N_1587);
or U1606 (N_1606,N_1506,N_1528);
or U1607 (N_1607,N_1529,N_1590);
or U1608 (N_1608,N_1521,N_1591);
nand U1609 (N_1609,N_1531,N_1585);
xnor U1610 (N_1610,N_1575,N_1565);
nor U1611 (N_1611,N_1548,N_1547);
nand U1612 (N_1612,N_1552,N_1527);
nand U1613 (N_1613,N_1576,N_1540);
xor U1614 (N_1614,N_1598,N_1596);
nand U1615 (N_1615,N_1530,N_1572);
and U1616 (N_1616,N_1559,N_1589);
nor U1617 (N_1617,N_1571,N_1520);
nor U1618 (N_1618,N_1523,N_1577);
and U1619 (N_1619,N_1526,N_1509);
or U1620 (N_1620,N_1535,N_1546);
nand U1621 (N_1621,N_1508,N_1511);
nand U1622 (N_1622,N_1564,N_1536);
and U1623 (N_1623,N_1595,N_1566);
xor U1624 (N_1624,N_1524,N_1517);
nor U1625 (N_1625,N_1594,N_1501);
and U1626 (N_1626,N_1549,N_1569);
nor U1627 (N_1627,N_1567,N_1543);
nor U1628 (N_1628,N_1545,N_1544);
or U1629 (N_1629,N_1510,N_1563);
or U1630 (N_1630,N_1561,N_1555);
nor U1631 (N_1631,N_1537,N_1574);
nor U1632 (N_1632,N_1519,N_1557);
nand U1633 (N_1633,N_1558,N_1570);
nand U1634 (N_1634,N_1515,N_1505);
nand U1635 (N_1635,N_1502,N_1532);
xor U1636 (N_1636,N_1542,N_1534);
nand U1637 (N_1637,N_1538,N_1550);
and U1638 (N_1638,N_1588,N_1581);
or U1639 (N_1639,N_1586,N_1592);
nand U1640 (N_1640,N_1507,N_1583);
and U1641 (N_1641,N_1539,N_1516);
nor U1642 (N_1642,N_1554,N_1513);
nand U1643 (N_1643,N_1503,N_1582);
nor U1644 (N_1644,N_1579,N_1514);
nand U1645 (N_1645,N_1553,N_1522);
xor U1646 (N_1646,N_1593,N_1568);
and U1647 (N_1647,N_1551,N_1599);
nor U1648 (N_1648,N_1541,N_1533);
or U1649 (N_1649,N_1578,N_1597);
nor U1650 (N_1650,N_1508,N_1565);
nor U1651 (N_1651,N_1526,N_1516);
or U1652 (N_1652,N_1592,N_1568);
or U1653 (N_1653,N_1545,N_1578);
nor U1654 (N_1654,N_1567,N_1590);
or U1655 (N_1655,N_1512,N_1513);
nand U1656 (N_1656,N_1567,N_1587);
and U1657 (N_1657,N_1524,N_1547);
xnor U1658 (N_1658,N_1583,N_1536);
or U1659 (N_1659,N_1567,N_1560);
and U1660 (N_1660,N_1588,N_1531);
nand U1661 (N_1661,N_1571,N_1599);
nand U1662 (N_1662,N_1532,N_1505);
or U1663 (N_1663,N_1591,N_1525);
nand U1664 (N_1664,N_1568,N_1543);
nand U1665 (N_1665,N_1564,N_1584);
xor U1666 (N_1666,N_1598,N_1518);
or U1667 (N_1667,N_1534,N_1564);
nand U1668 (N_1668,N_1515,N_1518);
xor U1669 (N_1669,N_1522,N_1514);
or U1670 (N_1670,N_1596,N_1521);
and U1671 (N_1671,N_1544,N_1515);
nand U1672 (N_1672,N_1571,N_1572);
and U1673 (N_1673,N_1531,N_1569);
nand U1674 (N_1674,N_1597,N_1536);
xnor U1675 (N_1675,N_1582,N_1522);
nor U1676 (N_1676,N_1549,N_1559);
nor U1677 (N_1677,N_1500,N_1502);
and U1678 (N_1678,N_1524,N_1526);
nand U1679 (N_1679,N_1578,N_1557);
nor U1680 (N_1680,N_1562,N_1515);
or U1681 (N_1681,N_1524,N_1575);
and U1682 (N_1682,N_1598,N_1513);
nand U1683 (N_1683,N_1568,N_1515);
xor U1684 (N_1684,N_1507,N_1599);
nand U1685 (N_1685,N_1549,N_1543);
or U1686 (N_1686,N_1585,N_1543);
or U1687 (N_1687,N_1525,N_1520);
nor U1688 (N_1688,N_1562,N_1581);
xnor U1689 (N_1689,N_1500,N_1515);
nor U1690 (N_1690,N_1513,N_1555);
and U1691 (N_1691,N_1587,N_1507);
nand U1692 (N_1692,N_1526,N_1557);
and U1693 (N_1693,N_1584,N_1567);
or U1694 (N_1694,N_1598,N_1555);
xnor U1695 (N_1695,N_1524,N_1504);
nor U1696 (N_1696,N_1568,N_1522);
nor U1697 (N_1697,N_1518,N_1501);
xnor U1698 (N_1698,N_1550,N_1523);
nand U1699 (N_1699,N_1589,N_1563);
or U1700 (N_1700,N_1698,N_1631);
nor U1701 (N_1701,N_1620,N_1637);
and U1702 (N_1702,N_1659,N_1670);
nor U1703 (N_1703,N_1624,N_1656);
and U1704 (N_1704,N_1613,N_1655);
xnor U1705 (N_1705,N_1671,N_1646);
or U1706 (N_1706,N_1652,N_1609);
and U1707 (N_1707,N_1642,N_1673);
and U1708 (N_1708,N_1699,N_1677);
xor U1709 (N_1709,N_1632,N_1651);
and U1710 (N_1710,N_1683,N_1663);
xor U1711 (N_1711,N_1628,N_1666);
nand U1712 (N_1712,N_1608,N_1672);
nand U1713 (N_1713,N_1629,N_1664);
or U1714 (N_1714,N_1661,N_1607);
nor U1715 (N_1715,N_1626,N_1604);
or U1716 (N_1716,N_1695,N_1687);
nor U1717 (N_1717,N_1600,N_1605);
or U1718 (N_1718,N_1616,N_1627);
and U1719 (N_1719,N_1601,N_1690);
or U1720 (N_1720,N_1693,N_1680);
nor U1721 (N_1721,N_1674,N_1612);
or U1722 (N_1722,N_1685,N_1660);
and U1723 (N_1723,N_1682,N_1619);
nor U1724 (N_1724,N_1678,N_1640);
nand U1725 (N_1725,N_1602,N_1667);
nor U1726 (N_1726,N_1668,N_1621);
nor U1727 (N_1727,N_1697,N_1603);
or U1728 (N_1728,N_1696,N_1675);
and U1729 (N_1729,N_1643,N_1662);
nor U1730 (N_1730,N_1606,N_1645);
nor U1731 (N_1731,N_1618,N_1639);
or U1732 (N_1732,N_1615,N_1694);
nor U1733 (N_1733,N_1684,N_1611);
and U1734 (N_1734,N_1622,N_1649);
or U1735 (N_1735,N_1692,N_1636);
or U1736 (N_1736,N_1686,N_1630);
and U1737 (N_1737,N_1669,N_1634);
and U1738 (N_1738,N_1648,N_1641);
nand U1739 (N_1739,N_1650,N_1681);
nor U1740 (N_1740,N_1625,N_1623);
xnor U1741 (N_1741,N_1647,N_1665);
and U1742 (N_1742,N_1676,N_1644);
xor U1743 (N_1743,N_1688,N_1654);
or U1744 (N_1744,N_1653,N_1691);
and U1745 (N_1745,N_1638,N_1658);
nor U1746 (N_1746,N_1614,N_1657);
or U1747 (N_1747,N_1633,N_1689);
and U1748 (N_1748,N_1617,N_1679);
nor U1749 (N_1749,N_1635,N_1610);
or U1750 (N_1750,N_1641,N_1653);
nand U1751 (N_1751,N_1685,N_1652);
or U1752 (N_1752,N_1670,N_1663);
xor U1753 (N_1753,N_1606,N_1626);
nand U1754 (N_1754,N_1672,N_1601);
or U1755 (N_1755,N_1666,N_1613);
or U1756 (N_1756,N_1683,N_1669);
nand U1757 (N_1757,N_1678,N_1611);
xor U1758 (N_1758,N_1696,N_1662);
nand U1759 (N_1759,N_1698,N_1646);
nand U1760 (N_1760,N_1690,N_1641);
and U1761 (N_1761,N_1660,N_1677);
nand U1762 (N_1762,N_1676,N_1692);
nand U1763 (N_1763,N_1649,N_1679);
nor U1764 (N_1764,N_1656,N_1626);
or U1765 (N_1765,N_1632,N_1650);
and U1766 (N_1766,N_1604,N_1684);
xor U1767 (N_1767,N_1623,N_1635);
or U1768 (N_1768,N_1687,N_1674);
nand U1769 (N_1769,N_1643,N_1611);
or U1770 (N_1770,N_1665,N_1602);
nand U1771 (N_1771,N_1645,N_1678);
nand U1772 (N_1772,N_1634,N_1651);
or U1773 (N_1773,N_1677,N_1661);
or U1774 (N_1774,N_1639,N_1659);
xnor U1775 (N_1775,N_1645,N_1616);
nand U1776 (N_1776,N_1619,N_1650);
nand U1777 (N_1777,N_1696,N_1697);
nor U1778 (N_1778,N_1676,N_1612);
nor U1779 (N_1779,N_1664,N_1621);
nand U1780 (N_1780,N_1626,N_1619);
nand U1781 (N_1781,N_1697,N_1691);
nor U1782 (N_1782,N_1626,N_1678);
nor U1783 (N_1783,N_1663,N_1671);
and U1784 (N_1784,N_1639,N_1636);
or U1785 (N_1785,N_1626,N_1685);
or U1786 (N_1786,N_1620,N_1600);
or U1787 (N_1787,N_1651,N_1617);
or U1788 (N_1788,N_1669,N_1662);
xor U1789 (N_1789,N_1646,N_1634);
nand U1790 (N_1790,N_1655,N_1638);
nor U1791 (N_1791,N_1670,N_1662);
nand U1792 (N_1792,N_1627,N_1688);
nor U1793 (N_1793,N_1668,N_1653);
or U1794 (N_1794,N_1602,N_1668);
and U1795 (N_1795,N_1652,N_1605);
and U1796 (N_1796,N_1641,N_1649);
nor U1797 (N_1797,N_1656,N_1651);
or U1798 (N_1798,N_1678,N_1677);
nand U1799 (N_1799,N_1687,N_1608);
and U1800 (N_1800,N_1768,N_1763);
and U1801 (N_1801,N_1753,N_1749);
xnor U1802 (N_1802,N_1783,N_1770);
nor U1803 (N_1803,N_1762,N_1713);
xor U1804 (N_1804,N_1796,N_1789);
or U1805 (N_1805,N_1797,N_1772);
and U1806 (N_1806,N_1712,N_1737);
or U1807 (N_1807,N_1727,N_1744);
and U1808 (N_1808,N_1756,N_1748);
xor U1809 (N_1809,N_1759,N_1707);
xor U1810 (N_1810,N_1765,N_1702);
or U1811 (N_1811,N_1779,N_1703);
nand U1812 (N_1812,N_1787,N_1718);
or U1813 (N_1813,N_1790,N_1751);
or U1814 (N_1814,N_1731,N_1791);
or U1815 (N_1815,N_1798,N_1777);
nand U1816 (N_1816,N_1785,N_1774);
nand U1817 (N_1817,N_1754,N_1724);
or U1818 (N_1818,N_1742,N_1704);
nor U1819 (N_1819,N_1743,N_1784);
or U1820 (N_1820,N_1795,N_1710);
nand U1821 (N_1821,N_1733,N_1781);
nor U1822 (N_1822,N_1794,N_1719);
and U1823 (N_1823,N_1700,N_1757);
nor U1824 (N_1824,N_1725,N_1705);
or U1825 (N_1825,N_1740,N_1722);
nor U1826 (N_1826,N_1788,N_1739);
or U1827 (N_1827,N_1746,N_1706);
xor U1828 (N_1828,N_1758,N_1730);
or U1829 (N_1829,N_1782,N_1764);
and U1830 (N_1830,N_1776,N_1729);
and U1831 (N_1831,N_1769,N_1752);
and U1832 (N_1832,N_1767,N_1723);
or U1833 (N_1833,N_1792,N_1735);
xor U1834 (N_1834,N_1747,N_1728);
and U1835 (N_1835,N_1738,N_1799);
and U1836 (N_1836,N_1793,N_1720);
nand U1837 (N_1837,N_1771,N_1714);
xnor U1838 (N_1838,N_1773,N_1711);
nor U1839 (N_1839,N_1780,N_1734);
xnor U1840 (N_1840,N_1755,N_1721);
nand U1841 (N_1841,N_1760,N_1775);
or U1842 (N_1842,N_1750,N_1766);
nand U1843 (N_1843,N_1709,N_1761);
and U1844 (N_1844,N_1778,N_1726);
nand U1845 (N_1845,N_1717,N_1745);
and U1846 (N_1846,N_1701,N_1741);
nand U1847 (N_1847,N_1715,N_1708);
nor U1848 (N_1848,N_1786,N_1736);
nand U1849 (N_1849,N_1716,N_1732);
or U1850 (N_1850,N_1742,N_1708);
and U1851 (N_1851,N_1745,N_1775);
and U1852 (N_1852,N_1786,N_1757);
nor U1853 (N_1853,N_1766,N_1709);
nor U1854 (N_1854,N_1709,N_1727);
or U1855 (N_1855,N_1734,N_1707);
nor U1856 (N_1856,N_1759,N_1747);
nor U1857 (N_1857,N_1717,N_1712);
or U1858 (N_1858,N_1796,N_1795);
nor U1859 (N_1859,N_1739,N_1790);
and U1860 (N_1860,N_1721,N_1740);
and U1861 (N_1861,N_1776,N_1731);
nand U1862 (N_1862,N_1788,N_1782);
or U1863 (N_1863,N_1770,N_1793);
and U1864 (N_1864,N_1736,N_1784);
xor U1865 (N_1865,N_1735,N_1788);
or U1866 (N_1866,N_1733,N_1723);
or U1867 (N_1867,N_1705,N_1769);
nor U1868 (N_1868,N_1763,N_1771);
and U1869 (N_1869,N_1725,N_1740);
xor U1870 (N_1870,N_1774,N_1780);
and U1871 (N_1871,N_1726,N_1750);
nand U1872 (N_1872,N_1740,N_1794);
nand U1873 (N_1873,N_1791,N_1729);
and U1874 (N_1874,N_1737,N_1717);
and U1875 (N_1875,N_1721,N_1756);
nor U1876 (N_1876,N_1719,N_1739);
nand U1877 (N_1877,N_1755,N_1760);
or U1878 (N_1878,N_1732,N_1795);
nor U1879 (N_1879,N_1769,N_1746);
nand U1880 (N_1880,N_1792,N_1769);
or U1881 (N_1881,N_1732,N_1709);
nand U1882 (N_1882,N_1762,N_1726);
xnor U1883 (N_1883,N_1756,N_1791);
nor U1884 (N_1884,N_1726,N_1737);
nor U1885 (N_1885,N_1745,N_1753);
nand U1886 (N_1886,N_1726,N_1771);
nor U1887 (N_1887,N_1747,N_1799);
xnor U1888 (N_1888,N_1701,N_1790);
nand U1889 (N_1889,N_1703,N_1791);
and U1890 (N_1890,N_1706,N_1736);
nor U1891 (N_1891,N_1748,N_1786);
nand U1892 (N_1892,N_1741,N_1797);
and U1893 (N_1893,N_1733,N_1774);
nor U1894 (N_1894,N_1789,N_1715);
or U1895 (N_1895,N_1729,N_1790);
or U1896 (N_1896,N_1760,N_1795);
nand U1897 (N_1897,N_1722,N_1794);
or U1898 (N_1898,N_1701,N_1735);
xnor U1899 (N_1899,N_1750,N_1707);
xor U1900 (N_1900,N_1876,N_1844);
and U1901 (N_1901,N_1837,N_1891);
nor U1902 (N_1902,N_1812,N_1817);
nor U1903 (N_1903,N_1849,N_1846);
or U1904 (N_1904,N_1867,N_1896);
and U1905 (N_1905,N_1869,N_1815);
nand U1906 (N_1906,N_1832,N_1858);
nor U1907 (N_1907,N_1879,N_1853);
nor U1908 (N_1908,N_1888,N_1873);
or U1909 (N_1909,N_1898,N_1814);
nand U1910 (N_1910,N_1866,N_1826);
nor U1911 (N_1911,N_1874,N_1882);
nor U1912 (N_1912,N_1856,N_1821);
or U1913 (N_1913,N_1813,N_1859);
xnor U1914 (N_1914,N_1822,N_1881);
or U1915 (N_1915,N_1897,N_1889);
or U1916 (N_1916,N_1841,N_1803);
and U1917 (N_1917,N_1834,N_1816);
or U1918 (N_1918,N_1852,N_1861);
nor U1919 (N_1919,N_1823,N_1833);
nand U1920 (N_1920,N_1850,N_1884);
nor U1921 (N_1921,N_1820,N_1828);
nand U1922 (N_1922,N_1827,N_1854);
or U1923 (N_1923,N_1864,N_1885);
nor U1924 (N_1924,N_1845,N_1829);
and U1925 (N_1925,N_1890,N_1801);
or U1926 (N_1926,N_1899,N_1807);
nor U1927 (N_1927,N_1848,N_1811);
and U1928 (N_1928,N_1883,N_1862);
and U1929 (N_1929,N_1808,N_1830);
nor U1930 (N_1930,N_1851,N_1831);
nand U1931 (N_1931,N_1877,N_1805);
or U1932 (N_1932,N_1868,N_1871);
nor U1933 (N_1933,N_1855,N_1886);
or U1934 (N_1934,N_1872,N_1865);
or U1935 (N_1935,N_1804,N_1847);
nand U1936 (N_1936,N_1818,N_1842);
or U1937 (N_1937,N_1894,N_1875);
nor U1938 (N_1938,N_1836,N_1819);
and U1939 (N_1939,N_1810,N_1800);
nor U1940 (N_1940,N_1802,N_1843);
nor U1941 (N_1941,N_1887,N_1860);
xnor U1942 (N_1942,N_1863,N_1870);
and U1943 (N_1943,N_1878,N_1835);
nor U1944 (N_1944,N_1806,N_1857);
or U1945 (N_1945,N_1824,N_1895);
or U1946 (N_1946,N_1892,N_1840);
nor U1947 (N_1947,N_1839,N_1893);
nand U1948 (N_1948,N_1825,N_1880);
nand U1949 (N_1949,N_1838,N_1809);
nand U1950 (N_1950,N_1821,N_1873);
nor U1951 (N_1951,N_1887,N_1853);
and U1952 (N_1952,N_1811,N_1859);
xor U1953 (N_1953,N_1820,N_1873);
nand U1954 (N_1954,N_1808,N_1850);
or U1955 (N_1955,N_1801,N_1817);
nor U1956 (N_1956,N_1853,N_1855);
and U1957 (N_1957,N_1890,N_1820);
nor U1958 (N_1958,N_1821,N_1857);
nand U1959 (N_1959,N_1825,N_1816);
and U1960 (N_1960,N_1801,N_1847);
nand U1961 (N_1961,N_1868,N_1836);
nand U1962 (N_1962,N_1856,N_1855);
and U1963 (N_1963,N_1873,N_1857);
nand U1964 (N_1964,N_1826,N_1884);
or U1965 (N_1965,N_1854,N_1820);
and U1966 (N_1966,N_1833,N_1832);
nor U1967 (N_1967,N_1835,N_1897);
nor U1968 (N_1968,N_1841,N_1887);
and U1969 (N_1969,N_1840,N_1811);
or U1970 (N_1970,N_1870,N_1808);
or U1971 (N_1971,N_1868,N_1804);
nor U1972 (N_1972,N_1835,N_1875);
xor U1973 (N_1973,N_1822,N_1841);
nor U1974 (N_1974,N_1885,N_1853);
and U1975 (N_1975,N_1834,N_1809);
nand U1976 (N_1976,N_1859,N_1856);
nor U1977 (N_1977,N_1803,N_1819);
and U1978 (N_1978,N_1880,N_1834);
xor U1979 (N_1979,N_1882,N_1830);
nor U1980 (N_1980,N_1882,N_1842);
nand U1981 (N_1981,N_1824,N_1897);
nor U1982 (N_1982,N_1823,N_1873);
xor U1983 (N_1983,N_1851,N_1829);
nand U1984 (N_1984,N_1873,N_1855);
nor U1985 (N_1985,N_1813,N_1810);
nand U1986 (N_1986,N_1861,N_1891);
nor U1987 (N_1987,N_1844,N_1808);
xnor U1988 (N_1988,N_1805,N_1867);
nand U1989 (N_1989,N_1833,N_1802);
or U1990 (N_1990,N_1824,N_1873);
or U1991 (N_1991,N_1882,N_1880);
nand U1992 (N_1992,N_1810,N_1897);
nand U1993 (N_1993,N_1834,N_1899);
or U1994 (N_1994,N_1885,N_1878);
or U1995 (N_1995,N_1853,N_1834);
nor U1996 (N_1996,N_1805,N_1853);
or U1997 (N_1997,N_1852,N_1835);
nor U1998 (N_1998,N_1807,N_1825);
nand U1999 (N_1999,N_1839,N_1821);
nor U2000 (N_2000,N_1920,N_1963);
nor U2001 (N_2001,N_1974,N_1942);
xor U2002 (N_2002,N_1934,N_1927);
and U2003 (N_2003,N_1955,N_1924);
nor U2004 (N_2004,N_1907,N_1913);
nor U2005 (N_2005,N_1958,N_1959);
or U2006 (N_2006,N_1979,N_1982);
and U2007 (N_2007,N_1964,N_1902);
nor U2008 (N_2008,N_1992,N_1944);
and U2009 (N_2009,N_1901,N_1938);
or U2010 (N_2010,N_1948,N_1922);
nor U2011 (N_2011,N_1961,N_1941);
xor U2012 (N_2012,N_1983,N_1914);
xor U2013 (N_2013,N_1939,N_1945);
nor U2014 (N_2014,N_1918,N_1912);
or U2015 (N_2015,N_1923,N_1987);
nor U2016 (N_2016,N_1910,N_1956);
or U2017 (N_2017,N_1905,N_1968);
and U2018 (N_2018,N_1976,N_1954);
xnor U2019 (N_2019,N_1921,N_1932);
nor U2020 (N_2020,N_1926,N_1925);
nor U2021 (N_2021,N_1946,N_1980);
nand U2022 (N_2022,N_1900,N_1996);
nor U2023 (N_2023,N_1940,N_1929);
nand U2024 (N_2024,N_1990,N_1951);
and U2025 (N_2025,N_1928,N_1989);
nor U2026 (N_2026,N_1933,N_1936);
nor U2027 (N_2027,N_1930,N_1911);
and U2028 (N_2028,N_1994,N_1908);
nor U2029 (N_2029,N_1967,N_1969);
nor U2030 (N_2030,N_1981,N_1986);
or U2031 (N_2031,N_1970,N_1935);
xor U2032 (N_2032,N_1943,N_1953);
and U2033 (N_2033,N_1965,N_1919);
nand U2034 (N_2034,N_1937,N_1906);
or U2035 (N_2035,N_1960,N_1998);
nor U2036 (N_2036,N_1999,N_1971);
and U2037 (N_2037,N_1972,N_1973);
nand U2038 (N_2038,N_1950,N_1957);
nor U2039 (N_2039,N_1977,N_1975);
nor U2040 (N_2040,N_1988,N_1915);
nand U2041 (N_2041,N_1949,N_1904);
or U2042 (N_2042,N_1903,N_1995);
nand U2043 (N_2043,N_1991,N_1978);
nor U2044 (N_2044,N_1962,N_1952);
nand U2045 (N_2045,N_1997,N_1984);
or U2046 (N_2046,N_1931,N_1917);
xor U2047 (N_2047,N_1947,N_1993);
or U2048 (N_2048,N_1916,N_1985);
or U2049 (N_2049,N_1909,N_1966);
or U2050 (N_2050,N_1912,N_1990);
or U2051 (N_2051,N_1986,N_1941);
nand U2052 (N_2052,N_1950,N_1942);
nor U2053 (N_2053,N_1941,N_1930);
or U2054 (N_2054,N_1980,N_1917);
or U2055 (N_2055,N_1949,N_1946);
nand U2056 (N_2056,N_1982,N_1976);
nor U2057 (N_2057,N_1976,N_1997);
nor U2058 (N_2058,N_1971,N_1927);
or U2059 (N_2059,N_1936,N_1934);
nand U2060 (N_2060,N_1950,N_1982);
nand U2061 (N_2061,N_1909,N_1942);
nand U2062 (N_2062,N_1972,N_1969);
and U2063 (N_2063,N_1953,N_1986);
and U2064 (N_2064,N_1934,N_1942);
nand U2065 (N_2065,N_1926,N_1947);
and U2066 (N_2066,N_1915,N_1967);
xor U2067 (N_2067,N_1995,N_1913);
or U2068 (N_2068,N_1983,N_1922);
and U2069 (N_2069,N_1945,N_1937);
or U2070 (N_2070,N_1923,N_1998);
nor U2071 (N_2071,N_1992,N_1977);
nor U2072 (N_2072,N_1971,N_1900);
or U2073 (N_2073,N_1983,N_1970);
xor U2074 (N_2074,N_1939,N_1996);
nor U2075 (N_2075,N_1942,N_1910);
nand U2076 (N_2076,N_1902,N_1976);
or U2077 (N_2077,N_1919,N_1930);
or U2078 (N_2078,N_1931,N_1995);
and U2079 (N_2079,N_1907,N_1968);
and U2080 (N_2080,N_1909,N_1974);
nand U2081 (N_2081,N_1974,N_1935);
and U2082 (N_2082,N_1935,N_1934);
nor U2083 (N_2083,N_1906,N_1923);
nor U2084 (N_2084,N_1952,N_1959);
or U2085 (N_2085,N_1945,N_1982);
or U2086 (N_2086,N_1987,N_1974);
and U2087 (N_2087,N_1986,N_1935);
nor U2088 (N_2088,N_1977,N_1924);
and U2089 (N_2089,N_1900,N_1974);
nand U2090 (N_2090,N_1935,N_1922);
and U2091 (N_2091,N_1969,N_1946);
or U2092 (N_2092,N_1991,N_1914);
nand U2093 (N_2093,N_1973,N_1906);
nand U2094 (N_2094,N_1965,N_1989);
xnor U2095 (N_2095,N_1911,N_1944);
or U2096 (N_2096,N_1997,N_1964);
and U2097 (N_2097,N_1936,N_1988);
nor U2098 (N_2098,N_1912,N_1913);
and U2099 (N_2099,N_1917,N_1970);
or U2100 (N_2100,N_2050,N_2041);
or U2101 (N_2101,N_2077,N_2063);
or U2102 (N_2102,N_2093,N_2091);
or U2103 (N_2103,N_2095,N_2080);
nor U2104 (N_2104,N_2021,N_2043);
or U2105 (N_2105,N_2011,N_2045);
nor U2106 (N_2106,N_2081,N_2055);
nor U2107 (N_2107,N_2074,N_2066);
nand U2108 (N_2108,N_2027,N_2002);
or U2109 (N_2109,N_2056,N_2038);
or U2110 (N_2110,N_2068,N_2008);
or U2111 (N_2111,N_2029,N_2064);
nor U2112 (N_2112,N_2046,N_2051);
or U2113 (N_2113,N_2088,N_2028);
or U2114 (N_2114,N_2015,N_2022);
nor U2115 (N_2115,N_2040,N_2042);
nand U2116 (N_2116,N_2013,N_2099);
xor U2117 (N_2117,N_2082,N_2014);
nor U2118 (N_2118,N_2019,N_2018);
or U2119 (N_2119,N_2071,N_2001);
and U2120 (N_2120,N_2098,N_2053);
nor U2121 (N_2121,N_2017,N_2078);
or U2122 (N_2122,N_2062,N_2075);
and U2123 (N_2123,N_2033,N_2058);
nand U2124 (N_2124,N_2025,N_2035);
or U2125 (N_2125,N_2039,N_2020);
and U2126 (N_2126,N_2004,N_2037);
and U2127 (N_2127,N_2034,N_2023);
nor U2128 (N_2128,N_2031,N_2084);
nand U2129 (N_2129,N_2089,N_2094);
nand U2130 (N_2130,N_2059,N_2076);
and U2131 (N_2131,N_2036,N_2079);
or U2132 (N_2132,N_2087,N_2096);
or U2133 (N_2133,N_2012,N_2005);
nand U2134 (N_2134,N_2065,N_2048);
nand U2135 (N_2135,N_2016,N_2083);
and U2136 (N_2136,N_2049,N_2054);
nor U2137 (N_2137,N_2006,N_2097);
and U2138 (N_2138,N_2057,N_2073);
nor U2139 (N_2139,N_2047,N_2067);
xor U2140 (N_2140,N_2003,N_2090);
nor U2141 (N_2141,N_2070,N_2072);
and U2142 (N_2142,N_2000,N_2060);
nand U2143 (N_2143,N_2009,N_2010);
and U2144 (N_2144,N_2030,N_2024);
and U2145 (N_2145,N_2061,N_2032);
and U2146 (N_2146,N_2086,N_2085);
nor U2147 (N_2147,N_2092,N_2069);
or U2148 (N_2148,N_2007,N_2026);
and U2149 (N_2149,N_2052,N_2044);
nand U2150 (N_2150,N_2052,N_2047);
or U2151 (N_2151,N_2089,N_2064);
and U2152 (N_2152,N_2050,N_2048);
and U2153 (N_2153,N_2081,N_2020);
nand U2154 (N_2154,N_2084,N_2065);
and U2155 (N_2155,N_2017,N_2055);
or U2156 (N_2156,N_2084,N_2080);
nor U2157 (N_2157,N_2018,N_2003);
nor U2158 (N_2158,N_2062,N_2022);
or U2159 (N_2159,N_2063,N_2099);
and U2160 (N_2160,N_2010,N_2004);
xor U2161 (N_2161,N_2057,N_2021);
nor U2162 (N_2162,N_2013,N_2030);
xor U2163 (N_2163,N_2047,N_2005);
and U2164 (N_2164,N_2005,N_2043);
nand U2165 (N_2165,N_2075,N_2005);
nor U2166 (N_2166,N_2056,N_2080);
or U2167 (N_2167,N_2019,N_2076);
nand U2168 (N_2168,N_2082,N_2091);
or U2169 (N_2169,N_2086,N_2046);
nor U2170 (N_2170,N_2026,N_2042);
xnor U2171 (N_2171,N_2076,N_2034);
and U2172 (N_2172,N_2046,N_2016);
nor U2173 (N_2173,N_2010,N_2081);
or U2174 (N_2174,N_2046,N_2022);
nand U2175 (N_2175,N_2070,N_2010);
and U2176 (N_2176,N_2075,N_2014);
nor U2177 (N_2177,N_2000,N_2088);
and U2178 (N_2178,N_2099,N_2007);
or U2179 (N_2179,N_2067,N_2039);
nor U2180 (N_2180,N_2006,N_2022);
nor U2181 (N_2181,N_2079,N_2044);
and U2182 (N_2182,N_2039,N_2000);
nand U2183 (N_2183,N_2052,N_2093);
nand U2184 (N_2184,N_2061,N_2074);
or U2185 (N_2185,N_2004,N_2066);
nor U2186 (N_2186,N_2097,N_2080);
or U2187 (N_2187,N_2047,N_2035);
nor U2188 (N_2188,N_2054,N_2023);
nor U2189 (N_2189,N_2022,N_2077);
nand U2190 (N_2190,N_2022,N_2091);
xnor U2191 (N_2191,N_2008,N_2047);
and U2192 (N_2192,N_2038,N_2034);
nor U2193 (N_2193,N_2089,N_2090);
xor U2194 (N_2194,N_2040,N_2050);
nand U2195 (N_2195,N_2038,N_2043);
nand U2196 (N_2196,N_2064,N_2085);
and U2197 (N_2197,N_2041,N_2006);
and U2198 (N_2198,N_2008,N_2002);
nand U2199 (N_2199,N_2089,N_2078);
nor U2200 (N_2200,N_2158,N_2150);
nor U2201 (N_2201,N_2132,N_2142);
or U2202 (N_2202,N_2154,N_2134);
nor U2203 (N_2203,N_2185,N_2172);
nand U2204 (N_2204,N_2110,N_2157);
or U2205 (N_2205,N_2145,N_2167);
nand U2206 (N_2206,N_2164,N_2116);
nand U2207 (N_2207,N_2143,N_2190);
nand U2208 (N_2208,N_2171,N_2114);
and U2209 (N_2209,N_2109,N_2156);
nand U2210 (N_2210,N_2181,N_2130);
and U2211 (N_2211,N_2105,N_2138);
nor U2212 (N_2212,N_2176,N_2100);
xnor U2213 (N_2213,N_2147,N_2120);
nand U2214 (N_2214,N_2146,N_2122);
and U2215 (N_2215,N_2136,N_2159);
nand U2216 (N_2216,N_2133,N_2103);
nor U2217 (N_2217,N_2177,N_2186);
nor U2218 (N_2218,N_2179,N_2151);
nor U2219 (N_2219,N_2119,N_2189);
or U2220 (N_2220,N_2187,N_2174);
or U2221 (N_2221,N_2161,N_2178);
xor U2222 (N_2222,N_2188,N_2166);
and U2223 (N_2223,N_2104,N_2125);
xor U2224 (N_2224,N_2182,N_2168);
xnor U2225 (N_2225,N_2102,N_2193);
or U2226 (N_2226,N_2123,N_2111);
and U2227 (N_2227,N_2191,N_2152);
and U2228 (N_2228,N_2131,N_2175);
and U2229 (N_2229,N_2162,N_2107);
xor U2230 (N_2230,N_2199,N_2195);
xor U2231 (N_2231,N_2196,N_2144);
nor U2232 (N_2232,N_2180,N_2140);
nand U2233 (N_2233,N_2165,N_2137);
and U2234 (N_2234,N_2197,N_2101);
nor U2235 (N_2235,N_2126,N_2192);
and U2236 (N_2236,N_2149,N_2112);
and U2237 (N_2237,N_2194,N_2198);
nand U2238 (N_2238,N_2118,N_2129);
nor U2239 (N_2239,N_2155,N_2184);
and U2240 (N_2240,N_2121,N_2106);
xnor U2241 (N_2241,N_2169,N_2139);
nand U2242 (N_2242,N_2127,N_2163);
xor U2243 (N_2243,N_2183,N_2113);
nand U2244 (N_2244,N_2148,N_2153);
nor U2245 (N_2245,N_2124,N_2160);
or U2246 (N_2246,N_2108,N_2141);
or U2247 (N_2247,N_2173,N_2170);
xnor U2248 (N_2248,N_2117,N_2115);
or U2249 (N_2249,N_2135,N_2128);
or U2250 (N_2250,N_2103,N_2182);
nor U2251 (N_2251,N_2171,N_2188);
nor U2252 (N_2252,N_2199,N_2122);
nand U2253 (N_2253,N_2139,N_2142);
and U2254 (N_2254,N_2124,N_2184);
and U2255 (N_2255,N_2127,N_2164);
nor U2256 (N_2256,N_2106,N_2189);
xnor U2257 (N_2257,N_2169,N_2126);
or U2258 (N_2258,N_2187,N_2137);
and U2259 (N_2259,N_2195,N_2151);
nand U2260 (N_2260,N_2147,N_2131);
and U2261 (N_2261,N_2130,N_2161);
and U2262 (N_2262,N_2113,N_2171);
or U2263 (N_2263,N_2143,N_2169);
nor U2264 (N_2264,N_2176,N_2106);
or U2265 (N_2265,N_2177,N_2188);
or U2266 (N_2266,N_2132,N_2124);
or U2267 (N_2267,N_2192,N_2160);
or U2268 (N_2268,N_2183,N_2114);
nand U2269 (N_2269,N_2162,N_2192);
xor U2270 (N_2270,N_2154,N_2105);
nand U2271 (N_2271,N_2186,N_2163);
and U2272 (N_2272,N_2149,N_2158);
nor U2273 (N_2273,N_2165,N_2115);
xor U2274 (N_2274,N_2128,N_2189);
nor U2275 (N_2275,N_2140,N_2125);
and U2276 (N_2276,N_2133,N_2115);
nor U2277 (N_2277,N_2193,N_2137);
nor U2278 (N_2278,N_2177,N_2190);
nand U2279 (N_2279,N_2114,N_2106);
and U2280 (N_2280,N_2161,N_2116);
nand U2281 (N_2281,N_2168,N_2132);
and U2282 (N_2282,N_2183,N_2101);
or U2283 (N_2283,N_2196,N_2145);
nor U2284 (N_2284,N_2175,N_2154);
and U2285 (N_2285,N_2104,N_2185);
nor U2286 (N_2286,N_2196,N_2151);
or U2287 (N_2287,N_2146,N_2195);
and U2288 (N_2288,N_2185,N_2181);
nor U2289 (N_2289,N_2112,N_2195);
nor U2290 (N_2290,N_2136,N_2126);
or U2291 (N_2291,N_2115,N_2191);
or U2292 (N_2292,N_2194,N_2104);
xor U2293 (N_2293,N_2134,N_2169);
and U2294 (N_2294,N_2170,N_2194);
or U2295 (N_2295,N_2172,N_2190);
xor U2296 (N_2296,N_2158,N_2122);
and U2297 (N_2297,N_2108,N_2184);
nand U2298 (N_2298,N_2177,N_2195);
nor U2299 (N_2299,N_2123,N_2115);
nor U2300 (N_2300,N_2275,N_2299);
and U2301 (N_2301,N_2253,N_2236);
or U2302 (N_2302,N_2296,N_2229);
and U2303 (N_2303,N_2242,N_2224);
and U2304 (N_2304,N_2269,N_2254);
nand U2305 (N_2305,N_2217,N_2255);
or U2306 (N_2306,N_2279,N_2225);
nor U2307 (N_2307,N_2227,N_2210);
xor U2308 (N_2308,N_2252,N_2204);
and U2309 (N_2309,N_2260,N_2277);
nor U2310 (N_2310,N_2244,N_2219);
nand U2311 (N_2311,N_2203,N_2222);
nor U2312 (N_2312,N_2286,N_2251);
nand U2313 (N_2313,N_2272,N_2215);
and U2314 (N_2314,N_2271,N_2284);
or U2315 (N_2315,N_2268,N_2274);
xnor U2316 (N_2316,N_2238,N_2276);
or U2317 (N_2317,N_2258,N_2207);
or U2318 (N_2318,N_2289,N_2265);
and U2319 (N_2319,N_2216,N_2262);
and U2320 (N_2320,N_2237,N_2200);
xnor U2321 (N_2321,N_2205,N_2283);
nor U2322 (N_2322,N_2235,N_2273);
nor U2323 (N_2323,N_2280,N_2297);
nand U2324 (N_2324,N_2292,N_2287);
nand U2325 (N_2325,N_2257,N_2298);
and U2326 (N_2326,N_2293,N_2221);
nor U2327 (N_2327,N_2202,N_2245);
nand U2328 (N_2328,N_2246,N_2208);
xnor U2329 (N_2329,N_2213,N_2256);
xor U2330 (N_2330,N_2267,N_2281);
nor U2331 (N_2331,N_2226,N_2241);
or U2332 (N_2332,N_2288,N_2201);
and U2333 (N_2333,N_2220,N_2231);
nor U2334 (N_2334,N_2206,N_2240);
or U2335 (N_2335,N_2214,N_2218);
or U2336 (N_2336,N_2212,N_2263);
nand U2337 (N_2337,N_2234,N_2295);
nand U2338 (N_2338,N_2285,N_2291);
xnor U2339 (N_2339,N_2243,N_2232);
nor U2340 (N_2340,N_2270,N_2290);
or U2341 (N_2341,N_2266,N_2250);
nor U2342 (N_2342,N_2248,N_2261);
nor U2343 (N_2343,N_2264,N_2228);
or U2344 (N_2344,N_2230,N_2278);
and U2345 (N_2345,N_2211,N_2247);
nand U2346 (N_2346,N_2239,N_2249);
nor U2347 (N_2347,N_2294,N_2223);
or U2348 (N_2348,N_2259,N_2233);
nor U2349 (N_2349,N_2282,N_2209);
or U2350 (N_2350,N_2276,N_2263);
or U2351 (N_2351,N_2284,N_2262);
or U2352 (N_2352,N_2226,N_2270);
nand U2353 (N_2353,N_2242,N_2275);
or U2354 (N_2354,N_2273,N_2279);
or U2355 (N_2355,N_2231,N_2286);
or U2356 (N_2356,N_2274,N_2276);
and U2357 (N_2357,N_2238,N_2258);
nor U2358 (N_2358,N_2239,N_2290);
or U2359 (N_2359,N_2260,N_2237);
nand U2360 (N_2360,N_2236,N_2272);
nor U2361 (N_2361,N_2255,N_2225);
and U2362 (N_2362,N_2221,N_2218);
or U2363 (N_2363,N_2274,N_2233);
and U2364 (N_2364,N_2217,N_2226);
and U2365 (N_2365,N_2203,N_2274);
nor U2366 (N_2366,N_2221,N_2271);
xnor U2367 (N_2367,N_2276,N_2212);
xnor U2368 (N_2368,N_2219,N_2278);
or U2369 (N_2369,N_2266,N_2213);
nor U2370 (N_2370,N_2278,N_2223);
nand U2371 (N_2371,N_2216,N_2201);
nor U2372 (N_2372,N_2241,N_2252);
nand U2373 (N_2373,N_2293,N_2261);
nand U2374 (N_2374,N_2249,N_2207);
nand U2375 (N_2375,N_2239,N_2208);
and U2376 (N_2376,N_2242,N_2248);
nor U2377 (N_2377,N_2204,N_2218);
nor U2378 (N_2378,N_2270,N_2232);
nand U2379 (N_2379,N_2291,N_2227);
xnor U2380 (N_2380,N_2255,N_2246);
xor U2381 (N_2381,N_2216,N_2223);
nand U2382 (N_2382,N_2234,N_2205);
or U2383 (N_2383,N_2227,N_2295);
nor U2384 (N_2384,N_2287,N_2202);
or U2385 (N_2385,N_2284,N_2248);
nor U2386 (N_2386,N_2218,N_2262);
nor U2387 (N_2387,N_2223,N_2282);
and U2388 (N_2388,N_2268,N_2217);
and U2389 (N_2389,N_2268,N_2258);
nand U2390 (N_2390,N_2241,N_2255);
xnor U2391 (N_2391,N_2259,N_2288);
and U2392 (N_2392,N_2255,N_2232);
or U2393 (N_2393,N_2239,N_2299);
or U2394 (N_2394,N_2296,N_2213);
and U2395 (N_2395,N_2248,N_2210);
nor U2396 (N_2396,N_2253,N_2279);
and U2397 (N_2397,N_2261,N_2290);
or U2398 (N_2398,N_2250,N_2247);
nor U2399 (N_2399,N_2284,N_2277);
xnor U2400 (N_2400,N_2346,N_2399);
nand U2401 (N_2401,N_2337,N_2364);
and U2402 (N_2402,N_2388,N_2344);
and U2403 (N_2403,N_2372,N_2359);
nor U2404 (N_2404,N_2378,N_2318);
xor U2405 (N_2405,N_2355,N_2377);
nor U2406 (N_2406,N_2317,N_2334);
nand U2407 (N_2407,N_2368,N_2345);
or U2408 (N_2408,N_2380,N_2312);
or U2409 (N_2409,N_2384,N_2316);
or U2410 (N_2410,N_2326,N_2349);
nand U2411 (N_2411,N_2307,N_2394);
nand U2412 (N_2412,N_2367,N_2329);
and U2413 (N_2413,N_2340,N_2308);
nand U2414 (N_2414,N_2386,N_2356);
nand U2415 (N_2415,N_2361,N_2398);
and U2416 (N_2416,N_2302,N_2374);
nor U2417 (N_2417,N_2387,N_2347);
and U2418 (N_2418,N_2351,N_2322);
nor U2419 (N_2419,N_2385,N_2338);
nand U2420 (N_2420,N_2352,N_2328);
or U2421 (N_2421,N_2323,N_2306);
nand U2422 (N_2422,N_2309,N_2301);
nor U2423 (N_2423,N_2381,N_2360);
nand U2424 (N_2424,N_2331,N_2303);
or U2425 (N_2425,N_2348,N_2300);
nor U2426 (N_2426,N_2393,N_2339);
and U2427 (N_2427,N_2350,N_2391);
or U2428 (N_2428,N_2313,N_2330);
or U2429 (N_2429,N_2343,N_2332);
nor U2430 (N_2430,N_2311,N_2319);
nor U2431 (N_2431,N_2305,N_2390);
nand U2432 (N_2432,N_2341,N_2324);
nor U2433 (N_2433,N_2358,N_2327);
or U2434 (N_2434,N_2314,N_2310);
xor U2435 (N_2435,N_2382,N_2342);
or U2436 (N_2436,N_2392,N_2396);
xor U2437 (N_2437,N_2315,N_2383);
or U2438 (N_2438,N_2365,N_2370);
nor U2439 (N_2439,N_2321,N_2366);
nand U2440 (N_2440,N_2357,N_2320);
or U2441 (N_2441,N_2373,N_2333);
nor U2442 (N_2442,N_2376,N_2395);
and U2443 (N_2443,N_2336,N_2363);
nand U2444 (N_2444,N_2389,N_2371);
nand U2445 (N_2445,N_2362,N_2375);
xor U2446 (N_2446,N_2304,N_2379);
nor U2447 (N_2447,N_2397,N_2369);
or U2448 (N_2448,N_2335,N_2325);
and U2449 (N_2449,N_2353,N_2354);
nor U2450 (N_2450,N_2361,N_2322);
nand U2451 (N_2451,N_2345,N_2309);
nand U2452 (N_2452,N_2351,N_2359);
and U2453 (N_2453,N_2347,N_2303);
nand U2454 (N_2454,N_2335,N_2377);
and U2455 (N_2455,N_2349,N_2386);
nor U2456 (N_2456,N_2377,N_2310);
and U2457 (N_2457,N_2311,N_2356);
or U2458 (N_2458,N_2386,N_2357);
nor U2459 (N_2459,N_2321,N_2330);
nand U2460 (N_2460,N_2369,N_2381);
nor U2461 (N_2461,N_2340,N_2390);
nor U2462 (N_2462,N_2343,N_2398);
xor U2463 (N_2463,N_2314,N_2379);
nand U2464 (N_2464,N_2333,N_2376);
nor U2465 (N_2465,N_2363,N_2385);
or U2466 (N_2466,N_2330,N_2379);
nand U2467 (N_2467,N_2392,N_2359);
nand U2468 (N_2468,N_2356,N_2337);
and U2469 (N_2469,N_2329,N_2309);
nand U2470 (N_2470,N_2391,N_2330);
and U2471 (N_2471,N_2369,N_2324);
and U2472 (N_2472,N_2325,N_2392);
nand U2473 (N_2473,N_2313,N_2350);
or U2474 (N_2474,N_2328,N_2318);
and U2475 (N_2475,N_2303,N_2310);
nor U2476 (N_2476,N_2370,N_2364);
nor U2477 (N_2477,N_2375,N_2310);
or U2478 (N_2478,N_2378,N_2328);
and U2479 (N_2479,N_2325,N_2316);
nand U2480 (N_2480,N_2347,N_2380);
and U2481 (N_2481,N_2379,N_2305);
nor U2482 (N_2482,N_2360,N_2304);
nand U2483 (N_2483,N_2330,N_2360);
or U2484 (N_2484,N_2346,N_2334);
nand U2485 (N_2485,N_2318,N_2373);
nor U2486 (N_2486,N_2388,N_2337);
nor U2487 (N_2487,N_2346,N_2343);
nor U2488 (N_2488,N_2388,N_2317);
nand U2489 (N_2489,N_2327,N_2308);
nand U2490 (N_2490,N_2333,N_2348);
xnor U2491 (N_2491,N_2375,N_2332);
xnor U2492 (N_2492,N_2379,N_2366);
nand U2493 (N_2493,N_2368,N_2385);
nor U2494 (N_2494,N_2308,N_2364);
and U2495 (N_2495,N_2362,N_2350);
or U2496 (N_2496,N_2306,N_2351);
and U2497 (N_2497,N_2381,N_2344);
or U2498 (N_2498,N_2350,N_2389);
nor U2499 (N_2499,N_2322,N_2353);
and U2500 (N_2500,N_2465,N_2455);
nor U2501 (N_2501,N_2490,N_2420);
xor U2502 (N_2502,N_2487,N_2468);
and U2503 (N_2503,N_2401,N_2469);
and U2504 (N_2504,N_2467,N_2452);
and U2505 (N_2505,N_2436,N_2492);
nand U2506 (N_2506,N_2471,N_2473);
nand U2507 (N_2507,N_2488,N_2418);
nor U2508 (N_2508,N_2431,N_2481);
and U2509 (N_2509,N_2447,N_2419);
nand U2510 (N_2510,N_2434,N_2493);
nor U2511 (N_2511,N_2421,N_2454);
and U2512 (N_2512,N_2402,N_2407);
nand U2513 (N_2513,N_2458,N_2445);
or U2514 (N_2514,N_2413,N_2456);
nor U2515 (N_2515,N_2426,N_2443);
nand U2516 (N_2516,N_2498,N_2477);
nor U2517 (N_2517,N_2427,N_2411);
or U2518 (N_2518,N_2404,N_2415);
xor U2519 (N_2519,N_2479,N_2430);
nor U2520 (N_2520,N_2425,N_2442);
or U2521 (N_2521,N_2408,N_2433);
nand U2522 (N_2522,N_2480,N_2414);
and U2523 (N_2523,N_2463,N_2440);
nand U2524 (N_2524,N_2476,N_2464);
nor U2525 (N_2525,N_2416,N_2475);
or U2526 (N_2526,N_2485,N_2453);
or U2527 (N_2527,N_2470,N_2429);
or U2528 (N_2528,N_2491,N_2478);
and U2529 (N_2529,N_2412,N_2400);
or U2530 (N_2530,N_2424,N_2446);
and U2531 (N_2531,N_2449,N_2457);
nand U2532 (N_2532,N_2410,N_2438);
and U2533 (N_2533,N_2496,N_2482);
xor U2534 (N_2534,N_2441,N_2461);
nor U2535 (N_2535,N_2405,N_2428);
and U2536 (N_2536,N_2448,N_2435);
or U2537 (N_2537,N_2495,N_2439);
or U2538 (N_2538,N_2432,N_2423);
nor U2539 (N_2539,N_2466,N_2489);
nor U2540 (N_2540,N_2494,N_2484);
or U2541 (N_2541,N_2472,N_2409);
and U2542 (N_2542,N_2444,N_2462);
and U2543 (N_2543,N_2406,N_2451);
and U2544 (N_2544,N_2483,N_2403);
or U2545 (N_2545,N_2422,N_2459);
nand U2546 (N_2546,N_2460,N_2499);
nand U2547 (N_2547,N_2450,N_2497);
nand U2548 (N_2548,N_2417,N_2437);
nand U2549 (N_2549,N_2474,N_2486);
and U2550 (N_2550,N_2445,N_2456);
nor U2551 (N_2551,N_2447,N_2424);
or U2552 (N_2552,N_2435,N_2463);
xor U2553 (N_2553,N_2450,N_2407);
or U2554 (N_2554,N_2458,N_2405);
nor U2555 (N_2555,N_2477,N_2404);
and U2556 (N_2556,N_2436,N_2458);
or U2557 (N_2557,N_2482,N_2429);
nor U2558 (N_2558,N_2461,N_2455);
xnor U2559 (N_2559,N_2493,N_2414);
nor U2560 (N_2560,N_2427,N_2408);
xor U2561 (N_2561,N_2491,N_2495);
nand U2562 (N_2562,N_2412,N_2442);
nor U2563 (N_2563,N_2433,N_2498);
and U2564 (N_2564,N_2493,N_2407);
nand U2565 (N_2565,N_2441,N_2460);
and U2566 (N_2566,N_2472,N_2407);
nor U2567 (N_2567,N_2427,N_2498);
nand U2568 (N_2568,N_2490,N_2457);
nand U2569 (N_2569,N_2432,N_2495);
and U2570 (N_2570,N_2428,N_2419);
or U2571 (N_2571,N_2454,N_2451);
nor U2572 (N_2572,N_2408,N_2413);
nor U2573 (N_2573,N_2402,N_2427);
or U2574 (N_2574,N_2496,N_2491);
or U2575 (N_2575,N_2424,N_2428);
nor U2576 (N_2576,N_2452,N_2426);
and U2577 (N_2577,N_2417,N_2429);
nor U2578 (N_2578,N_2457,N_2488);
nor U2579 (N_2579,N_2406,N_2412);
xnor U2580 (N_2580,N_2489,N_2433);
and U2581 (N_2581,N_2486,N_2437);
or U2582 (N_2582,N_2479,N_2411);
xnor U2583 (N_2583,N_2427,N_2461);
nand U2584 (N_2584,N_2409,N_2433);
xor U2585 (N_2585,N_2488,N_2451);
nor U2586 (N_2586,N_2460,N_2444);
nand U2587 (N_2587,N_2421,N_2488);
and U2588 (N_2588,N_2431,N_2442);
and U2589 (N_2589,N_2440,N_2438);
nor U2590 (N_2590,N_2453,N_2458);
or U2591 (N_2591,N_2417,N_2447);
or U2592 (N_2592,N_2494,N_2406);
nand U2593 (N_2593,N_2407,N_2449);
or U2594 (N_2594,N_2405,N_2498);
xnor U2595 (N_2595,N_2423,N_2485);
nand U2596 (N_2596,N_2485,N_2486);
or U2597 (N_2597,N_2466,N_2411);
and U2598 (N_2598,N_2493,N_2426);
or U2599 (N_2599,N_2436,N_2446);
or U2600 (N_2600,N_2570,N_2525);
or U2601 (N_2601,N_2582,N_2533);
nor U2602 (N_2602,N_2509,N_2562);
nand U2603 (N_2603,N_2508,N_2511);
and U2604 (N_2604,N_2578,N_2523);
nand U2605 (N_2605,N_2550,N_2530);
and U2606 (N_2606,N_2589,N_2560);
nor U2607 (N_2607,N_2527,N_2568);
and U2608 (N_2608,N_2526,N_2510);
or U2609 (N_2609,N_2536,N_2576);
nor U2610 (N_2610,N_2588,N_2518);
nor U2611 (N_2611,N_2512,N_2531);
or U2612 (N_2612,N_2524,N_2516);
nor U2613 (N_2613,N_2590,N_2599);
nand U2614 (N_2614,N_2540,N_2553);
or U2615 (N_2615,N_2547,N_2501);
xnor U2616 (N_2616,N_2554,N_2566);
and U2617 (N_2617,N_2538,N_2561);
nand U2618 (N_2618,N_2558,N_2500);
or U2619 (N_2619,N_2583,N_2544);
or U2620 (N_2620,N_2591,N_2584);
nor U2621 (N_2621,N_2571,N_2541);
and U2622 (N_2622,N_2537,N_2587);
xor U2623 (N_2623,N_2513,N_2569);
and U2624 (N_2624,N_2552,N_2595);
nand U2625 (N_2625,N_2521,N_2585);
or U2626 (N_2626,N_2594,N_2517);
and U2627 (N_2627,N_2597,N_2515);
nor U2628 (N_2628,N_2596,N_2567);
nor U2629 (N_2629,N_2563,N_2564);
nor U2630 (N_2630,N_2598,N_2586);
or U2631 (N_2631,N_2506,N_2529);
and U2632 (N_2632,N_2580,N_2575);
nand U2633 (N_2633,N_2504,N_2581);
or U2634 (N_2634,N_2551,N_2535);
nand U2635 (N_2635,N_2507,N_2545);
and U2636 (N_2636,N_2534,N_2548);
and U2637 (N_2637,N_2539,N_2573);
nand U2638 (N_2638,N_2522,N_2549);
xor U2639 (N_2639,N_2502,N_2532);
xnor U2640 (N_2640,N_2593,N_2505);
nand U2641 (N_2641,N_2514,N_2542);
and U2642 (N_2642,N_2528,N_2555);
or U2643 (N_2643,N_2519,N_2579);
xor U2644 (N_2644,N_2565,N_2556);
nand U2645 (N_2645,N_2592,N_2503);
or U2646 (N_2646,N_2559,N_2577);
nor U2647 (N_2647,N_2572,N_2574);
nor U2648 (N_2648,N_2557,N_2546);
xnor U2649 (N_2649,N_2543,N_2520);
xnor U2650 (N_2650,N_2521,N_2557);
or U2651 (N_2651,N_2562,N_2579);
nor U2652 (N_2652,N_2538,N_2576);
and U2653 (N_2653,N_2586,N_2543);
nand U2654 (N_2654,N_2547,N_2585);
or U2655 (N_2655,N_2565,N_2507);
or U2656 (N_2656,N_2545,N_2579);
nand U2657 (N_2657,N_2593,N_2550);
nand U2658 (N_2658,N_2540,N_2560);
and U2659 (N_2659,N_2587,N_2565);
nand U2660 (N_2660,N_2521,N_2536);
or U2661 (N_2661,N_2560,N_2599);
and U2662 (N_2662,N_2524,N_2542);
and U2663 (N_2663,N_2541,N_2534);
and U2664 (N_2664,N_2555,N_2545);
or U2665 (N_2665,N_2532,N_2521);
nand U2666 (N_2666,N_2516,N_2582);
nand U2667 (N_2667,N_2546,N_2525);
or U2668 (N_2668,N_2526,N_2511);
nand U2669 (N_2669,N_2574,N_2506);
or U2670 (N_2670,N_2598,N_2582);
and U2671 (N_2671,N_2541,N_2515);
nand U2672 (N_2672,N_2592,N_2575);
or U2673 (N_2673,N_2577,N_2589);
or U2674 (N_2674,N_2595,N_2555);
and U2675 (N_2675,N_2573,N_2528);
xor U2676 (N_2676,N_2566,N_2532);
or U2677 (N_2677,N_2521,N_2567);
nor U2678 (N_2678,N_2582,N_2540);
nand U2679 (N_2679,N_2552,N_2540);
xor U2680 (N_2680,N_2536,N_2511);
and U2681 (N_2681,N_2555,N_2583);
xnor U2682 (N_2682,N_2520,N_2511);
nor U2683 (N_2683,N_2558,N_2502);
or U2684 (N_2684,N_2549,N_2562);
nand U2685 (N_2685,N_2547,N_2512);
and U2686 (N_2686,N_2562,N_2536);
and U2687 (N_2687,N_2518,N_2522);
nor U2688 (N_2688,N_2555,N_2526);
nand U2689 (N_2689,N_2579,N_2593);
or U2690 (N_2690,N_2538,N_2543);
xnor U2691 (N_2691,N_2536,N_2583);
or U2692 (N_2692,N_2513,N_2519);
nand U2693 (N_2693,N_2518,N_2503);
nor U2694 (N_2694,N_2563,N_2526);
or U2695 (N_2695,N_2584,N_2571);
xor U2696 (N_2696,N_2528,N_2522);
nor U2697 (N_2697,N_2565,N_2524);
nor U2698 (N_2698,N_2564,N_2578);
or U2699 (N_2699,N_2594,N_2575);
or U2700 (N_2700,N_2610,N_2684);
nand U2701 (N_2701,N_2639,N_2627);
or U2702 (N_2702,N_2632,N_2626);
and U2703 (N_2703,N_2670,N_2604);
nor U2704 (N_2704,N_2637,N_2667);
and U2705 (N_2705,N_2659,N_2617);
or U2706 (N_2706,N_2697,N_2661);
and U2707 (N_2707,N_2668,N_2629);
and U2708 (N_2708,N_2694,N_2603);
or U2709 (N_2709,N_2631,N_2601);
and U2710 (N_2710,N_2643,N_2619);
and U2711 (N_2711,N_2647,N_2677);
or U2712 (N_2712,N_2686,N_2612);
or U2713 (N_2713,N_2696,N_2648);
nand U2714 (N_2714,N_2615,N_2663);
nor U2715 (N_2715,N_2673,N_2607);
nand U2716 (N_2716,N_2645,N_2669);
and U2717 (N_2717,N_2678,N_2693);
or U2718 (N_2718,N_2665,N_2653);
nor U2719 (N_2719,N_2606,N_2657);
or U2720 (N_2720,N_2640,N_2618);
xnor U2721 (N_2721,N_2621,N_2633);
or U2722 (N_2722,N_2680,N_2682);
and U2723 (N_2723,N_2635,N_2690);
and U2724 (N_2724,N_2600,N_2699);
xnor U2725 (N_2725,N_2660,N_2654);
or U2726 (N_2726,N_2622,N_2672);
nand U2727 (N_2727,N_2688,N_2609);
nor U2728 (N_2728,N_2681,N_2613);
and U2729 (N_2729,N_2675,N_2602);
or U2730 (N_2730,N_2646,N_2689);
nand U2731 (N_2731,N_2623,N_2664);
and U2732 (N_2732,N_2662,N_2685);
nand U2733 (N_2733,N_2634,N_2679);
or U2734 (N_2734,N_2605,N_2695);
nand U2735 (N_2735,N_2671,N_2655);
and U2736 (N_2736,N_2651,N_2649);
and U2737 (N_2737,N_2616,N_2658);
and U2738 (N_2738,N_2656,N_2638);
and U2739 (N_2739,N_2683,N_2666);
nand U2740 (N_2740,N_2636,N_2692);
nand U2741 (N_2741,N_2624,N_2644);
or U2742 (N_2742,N_2676,N_2698);
nor U2743 (N_2743,N_2642,N_2674);
nand U2744 (N_2744,N_2614,N_2641);
nor U2745 (N_2745,N_2608,N_2611);
or U2746 (N_2746,N_2650,N_2652);
and U2747 (N_2747,N_2625,N_2620);
nor U2748 (N_2748,N_2691,N_2687);
and U2749 (N_2749,N_2628,N_2630);
xnor U2750 (N_2750,N_2682,N_2630);
nand U2751 (N_2751,N_2691,N_2621);
nand U2752 (N_2752,N_2610,N_2611);
and U2753 (N_2753,N_2623,N_2650);
nor U2754 (N_2754,N_2677,N_2637);
and U2755 (N_2755,N_2623,N_2641);
or U2756 (N_2756,N_2627,N_2692);
nor U2757 (N_2757,N_2659,N_2681);
nor U2758 (N_2758,N_2679,N_2616);
xnor U2759 (N_2759,N_2670,N_2602);
and U2760 (N_2760,N_2667,N_2676);
nand U2761 (N_2761,N_2641,N_2692);
and U2762 (N_2762,N_2676,N_2605);
or U2763 (N_2763,N_2662,N_2639);
or U2764 (N_2764,N_2677,N_2680);
nor U2765 (N_2765,N_2690,N_2696);
xor U2766 (N_2766,N_2656,N_2676);
nand U2767 (N_2767,N_2608,N_2622);
nand U2768 (N_2768,N_2654,N_2689);
xor U2769 (N_2769,N_2609,N_2660);
and U2770 (N_2770,N_2633,N_2609);
nand U2771 (N_2771,N_2650,N_2644);
and U2772 (N_2772,N_2614,N_2662);
nand U2773 (N_2773,N_2659,N_2648);
nor U2774 (N_2774,N_2656,N_2607);
or U2775 (N_2775,N_2658,N_2654);
xor U2776 (N_2776,N_2638,N_2696);
nor U2777 (N_2777,N_2649,N_2672);
or U2778 (N_2778,N_2630,N_2607);
nand U2779 (N_2779,N_2635,N_2634);
or U2780 (N_2780,N_2605,N_2654);
xnor U2781 (N_2781,N_2608,N_2687);
or U2782 (N_2782,N_2648,N_2609);
nand U2783 (N_2783,N_2674,N_2677);
nand U2784 (N_2784,N_2687,N_2697);
nor U2785 (N_2785,N_2638,N_2635);
xor U2786 (N_2786,N_2662,N_2632);
nand U2787 (N_2787,N_2676,N_2621);
or U2788 (N_2788,N_2629,N_2678);
or U2789 (N_2789,N_2600,N_2668);
or U2790 (N_2790,N_2600,N_2646);
or U2791 (N_2791,N_2698,N_2658);
nor U2792 (N_2792,N_2635,N_2677);
nand U2793 (N_2793,N_2627,N_2689);
nor U2794 (N_2794,N_2600,N_2680);
or U2795 (N_2795,N_2693,N_2616);
nor U2796 (N_2796,N_2609,N_2618);
xor U2797 (N_2797,N_2679,N_2685);
nor U2798 (N_2798,N_2652,N_2667);
and U2799 (N_2799,N_2645,N_2684);
nand U2800 (N_2800,N_2757,N_2778);
nand U2801 (N_2801,N_2752,N_2797);
or U2802 (N_2802,N_2739,N_2782);
nor U2803 (N_2803,N_2776,N_2702);
nor U2804 (N_2804,N_2789,N_2783);
and U2805 (N_2805,N_2741,N_2792);
nor U2806 (N_2806,N_2750,N_2738);
nand U2807 (N_2807,N_2726,N_2799);
nor U2808 (N_2808,N_2740,N_2764);
nor U2809 (N_2809,N_2766,N_2700);
or U2810 (N_2810,N_2758,N_2705);
nand U2811 (N_2811,N_2746,N_2784);
or U2812 (N_2812,N_2703,N_2743);
and U2813 (N_2813,N_2714,N_2773);
or U2814 (N_2814,N_2785,N_2720);
nor U2815 (N_2815,N_2786,N_2775);
and U2816 (N_2816,N_2761,N_2779);
or U2817 (N_2817,N_2729,N_2755);
nor U2818 (N_2818,N_2795,N_2790);
xor U2819 (N_2819,N_2731,N_2794);
nand U2820 (N_2820,N_2718,N_2716);
nor U2821 (N_2821,N_2759,N_2765);
nand U2822 (N_2822,N_2777,N_2791);
and U2823 (N_2823,N_2732,N_2723);
or U2824 (N_2824,N_2753,N_2734);
nand U2825 (N_2825,N_2706,N_2745);
or U2826 (N_2826,N_2760,N_2737);
or U2827 (N_2827,N_2748,N_2788);
xor U2828 (N_2828,N_2715,N_2747);
nand U2829 (N_2829,N_2717,N_2735);
nor U2830 (N_2830,N_2763,N_2707);
and U2831 (N_2831,N_2711,N_2709);
xor U2832 (N_2832,N_2774,N_2751);
xnor U2833 (N_2833,N_2787,N_2724);
and U2834 (N_2834,N_2793,N_2725);
nor U2835 (N_2835,N_2772,N_2749);
or U2836 (N_2836,N_2710,N_2713);
xor U2837 (N_2837,N_2704,N_2781);
xor U2838 (N_2838,N_2798,N_2722);
xnor U2839 (N_2839,N_2762,N_2736);
or U2840 (N_2840,N_2733,N_2769);
and U2841 (N_2841,N_2768,N_2756);
and U2842 (N_2842,N_2719,N_2744);
nor U2843 (N_2843,N_2727,N_2712);
xnor U2844 (N_2844,N_2701,N_2754);
xnor U2845 (N_2845,N_2780,N_2771);
nand U2846 (N_2846,N_2721,N_2728);
and U2847 (N_2847,N_2708,N_2742);
nor U2848 (N_2848,N_2770,N_2730);
nor U2849 (N_2849,N_2767,N_2796);
or U2850 (N_2850,N_2787,N_2765);
or U2851 (N_2851,N_2788,N_2734);
nor U2852 (N_2852,N_2703,N_2791);
nand U2853 (N_2853,N_2705,N_2776);
or U2854 (N_2854,N_2790,N_2789);
nor U2855 (N_2855,N_2726,N_2768);
or U2856 (N_2856,N_2745,N_2750);
or U2857 (N_2857,N_2747,N_2728);
or U2858 (N_2858,N_2733,N_2751);
nor U2859 (N_2859,N_2718,N_2730);
nor U2860 (N_2860,N_2722,N_2793);
nor U2861 (N_2861,N_2782,N_2756);
or U2862 (N_2862,N_2765,N_2756);
nand U2863 (N_2863,N_2712,N_2707);
and U2864 (N_2864,N_2708,N_2704);
and U2865 (N_2865,N_2799,N_2771);
xnor U2866 (N_2866,N_2763,N_2713);
or U2867 (N_2867,N_2794,N_2717);
nand U2868 (N_2868,N_2786,N_2716);
nor U2869 (N_2869,N_2780,N_2785);
and U2870 (N_2870,N_2728,N_2713);
nand U2871 (N_2871,N_2753,N_2762);
nor U2872 (N_2872,N_2755,N_2701);
or U2873 (N_2873,N_2759,N_2779);
and U2874 (N_2874,N_2735,N_2773);
xor U2875 (N_2875,N_2743,N_2779);
nand U2876 (N_2876,N_2719,N_2773);
and U2877 (N_2877,N_2701,N_2757);
or U2878 (N_2878,N_2708,N_2728);
nand U2879 (N_2879,N_2746,N_2776);
nand U2880 (N_2880,N_2772,N_2709);
and U2881 (N_2881,N_2786,N_2727);
nand U2882 (N_2882,N_2744,N_2746);
or U2883 (N_2883,N_2792,N_2726);
or U2884 (N_2884,N_2761,N_2723);
nand U2885 (N_2885,N_2741,N_2799);
and U2886 (N_2886,N_2707,N_2725);
or U2887 (N_2887,N_2726,N_2718);
and U2888 (N_2888,N_2742,N_2776);
nor U2889 (N_2889,N_2738,N_2790);
nor U2890 (N_2890,N_2777,N_2782);
or U2891 (N_2891,N_2728,N_2771);
nor U2892 (N_2892,N_2769,N_2726);
xnor U2893 (N_2893,N_2721,N_2703);
or U2894 (N_2894,N_2766,N_2768);
or U2895 (N_2895,N_2722,N_2721);
or U2896 (N_2896,N_2791,N_2789);
nand U2897 (N_2897,N_2712,N_2770);
xor U2898 (N_2898,N_2734,N_2703);
nand U2899 (N_2899,N_2786,N_2789);
nor U2900 (N_2900,N_2837,N_2881);
or U2901 (N_2901,N_2858,N_2806);
and U2902 (N_2902,N_2875,N_2805);
or U2903 (N_2903,N_2895,N_2821);
and U2904 (N_2904,N_2865,N_2833);
or U2905 (N_2905,N_2886,N_2863);
and U2906 (N_2906,N_2868,N_2818);
nor U2907 (N_2907,N_2848,N_2885);
and U2908 (N_2908,N_2822,N_2864);
and U2909 (N_2909,N_2816,N_2862);
nand U2910 (N_2910,N_2870,N_2890);
nor U2911 (N_2911,N_2853,N_2819);
xor U2912 (N_2912,N_2893,N_2824);
or U2913 (N_2913,N_2874,N_2809);
and U2914 (N_2914,N_2871,N_2823);
xor U2915 (N_2915,N_2891,N_2856);
or U2916 (N_2916,N_2808,N_2873);
or U2917 (N_2917,N_2884,N_2888);
or U2918 (N_2918,N_2860,N_2845);
or U2919 (N_2919,N_2867,N_2883);
or U2920 (N_2920,N_2899,N_2817);
and U2921 (N_2921,N_2887,N_2846);
nand U2922 (N_2922,N_2829,N_2861);
nand U2923 (N_2923,N_2880,N_2843);
nand U2924 (N_2924,N_2847,N_2852);
nand U2925 (N_2925,N_2828,N_2855);
nand U2926 (N_2926,N_2892,N_2800);
nor U2927 (N_2927,N_2876,N_2878);
nand U2928 (N_2928,N_2814,N_2879);
or U2929 (N_2929,N_2834,N_2831);
nor U2930 (N_2930,N_2898,N_2811);
nor U2931 (N_2931,N_2804,N_2825);
or U2932 (N_2932,N_2872,N_2894);
and U2933 (N_2933,N_2842,N_2854);
and U2934 (N_2934,N_2840,N_2832);
nand U2935 (N_2935,N_2807,N_2810);
nor U2936 (N_2936,N_2851,N_2802);
and U2937 (N_2937,N_2813,N_2826);
nor U2938 (N_2938,N_2812,N_2803);
or U2939 (N_2939,N_2841,N_2839);
nor U2940 (N_2940,N_2896,N_2820);
nor U2941 (N_2941,N_2844,N_2801);
and U2942 (N_2942,N_2877,N_2857);
and U2943 (N_2943,N_2869,N_2835);
nor U2944 (N_2944,N_2815,N_2830);
or U2945 (N_2945,N_2850,N_2836);
nor U2946 (N_2946,N_2838,N_2827);
xor U2947 (N_2947,N_2859,N_2897);
nor U2948 (N_2948,N_2849,N_2866);
nand U2949 (N_2949,N_2882,N_2889);
and U2950 (N_2950,N_2878,N_2817);
nand U2951 (N_2951,N_2862,N_2853);
and U2952 (N_2952,N_2807,N_2803);
or U2953 (N_2953,N_2842,N_2866);
and U2954 (N_2954,N_2888,N_2827);
nor U2955 (N_2955,N_2836,N_2840);
nor U2956 (N_2956,N_2809,N_2841);
nand U2957 (N_2957,N_2823,N_2896);
nand U2958 (N_2958,N_2815,N_2878);
nor U2959 (N_2959,N_2859,N_2875);
and U2960 (N_2960,N_2846,N_2831);
nor U2961 (N_2961,N_2859,N_2820);
nor U2962 (N_2962,N_2811,N_2807);
nor U2963 (N_2963,N_2874,N_2807);
or U2964 (N_2964,N_2852,N_2862);
and U2965 (N_2965,N_2843,N_2884);
nand U2966 (N_2966,N_2854,N_2879);
and U2967 (N_2967,N_2836,N_2839);
nand U2968 (N_2968,N_2859,N_2847);
or U2969 (N_2969,N_2883,N_2838);
nand U2970 (N_2970,N_2823,N_2884);
nand U2971 (N_2971,N_2823,N_2880);
xnor U2972 (N_2972,N_2824,N_2858);
nor U2973 (N_2973,N_2881,N_2806);
xor U2974 (N_2974,N_2877,N_2851);
xor U2975 (N_2975,N_2840,N_2887);
or U2976 (N_2976,N_2813,N_2884);
or U2977 (N_2977,N_2869,N_2849);
xor U2978 (N_2978,N_2849,N_2808);
nand U2979 (N_2979,N_2881,N_2808);
and U2980 (N_2980,N_2852,N_2875);
nand U2981 (N_2981,N_2818,N_2837);
nand U2982 (N_2982,N_2829,N_2872);
or U2983 (N_2983,N_2893,N_2871);
nand U2984 (N_2984,N_2840,N_2863);
nand U2985 (N_2985,N_2876,N_2860);
nand U2986 (N_2986,N_2841,N_2824);
nand U2987 (N_2987,N_2858,N_2857);
nor U2988 (N_2988,N_2803,N_2865);
xor U2989 (N_2989,N_2833,N_2868);
nor U2990 (N_2990,N_2815,N_2885);
nand U2991 (N_2991,N_2828,N_2842);
and U2992 (N_2992,N_2845,N_2808);
or U2993 (N_2993,N_2833,N_2818);
nand U2994 (N_2994,N_2885,N_2868);
and U2995 (N_2995,N_2867,N_2833);
or U2996 (N_2996,N_2812,N_2897);
nor U2997 (N_2997,N_2852,N_2890);
nor U2998 (N_2998,N_2850,N_2823);
and U2999 (N_2999,N_2885,N_2833);
nand U3000 (N_3000,N_2954,N_2916);
xor U3001 (N_3001,N_2914,N_2977);
xnor U3002 (N_3002,N_2904,N_2943);
nor U3003 (N_3003,N_2988,N_2994);
or U3004 (N_3004,N_2956,N_2936);
or U3005 (N_3005,N_2972,N_2969);
and U3006 (N_3006,N_2929,N_2926);
nor U3007 (N_3007,N_2939,N_2983);
xnor U3008 (N_3008,N_2985,N_2951);
nor U3009 (N_3009,N_2935,N_2927);
or U3010 (N_3010,N_2975,N_2903);
or U3011 (N_3011,N_2944,N_2973);
xnor U3012 (N_3012,N_2941,N_2949);
and U3013 (N_3013,N_2992,N_2921);
or U3014 (N_3014,N_2987,N_2909);
and U3015 (N_3015,N_2947,N_2910);
and U3016 (N_3016,N_2906,N_2970);
and U3017 (N_3017,N_2980,N_2966);
or U3018 (N_3018,N_2990,N_2950);
nor U3019 (N_3019,N_2952,N_2979);
nand U3020 (N_3020,N_2942,N_2962);
and U3021 (N_3021,N_2913,N_2912);
and U3022 (N_3022,N_2997,N_2971);
xor U3023 (N_3023,N_2922,N_2945);
nor U3024 (N_3024,N_2915,N_2999);
and U3025 (N_3025,N_2981,N_2908);
or U3026 (N_3026,N_2959,N_2989);
nand U3027 (N_3027,N_2919,N_2938);
or U3028 (N_3028,N_2937,N_2976);
and U3029 (N_3029,N_2933,N_2968);
nand U3030 (N_3030,N_2900,N_2953);
and U3031 (N_3031,N_2948,N_2920);
nor U3032 (N_3032,N_2993,N_2964);
nor U3033 (N_3033,N_2925,N_2961);
or U3034 (N_3034,N_2930,N_2923);
nand U3035 (N_3035,N_2957,N_2984);
or U3036 (N_3036,N_2940,N_2911);
and U3037 (N_3037,N_2934,N_2958);
and U3038 (N_3038,N_2967,N_2932);
nor U3039 (N_3039,N_2986,N_2974);
nand U3040 (N_3040,N_2995,N_2955);
and U3041 (N_3041,N_2965,N_2946);
nand U3042 (N_3042,N_2963,N_2928);
or U3043 (N_3043,N_2982,N_2960);
nand U3044 (N_3044,N_2924,N_2917);
nor U3045 (N_3045,N_2996,N_2978);
or U3046 (N_3046,N_2907,N_2991);
or U3047 (N_3047,N_2931,N_2902);
nand U3048 (N_3048,N_2998,N_2901);
nand U3049 (N_3049,N_2905,N_2918);
nor U3050 (N_3050,N_2902,N_2945);
nand U3051 (N_3051,N_2982,N_2921);
or U3052 (N_3052,N_2950,N_2957);
and U3053 (N_3053,N_2930,N_2914);
nor U3054 (N_3054,N_2918,N_2923);
and U3055 (N_3055,N_2974,N_2948);
nand U3056 (N_3056,N_2997,N_2930);
or U3057 (N_3057,N_2972,N_2995);
or U3058 (N_3058,N_2926,N_2922);
and U3059 (N_3059,N_2958,N_2930);
nand U3060 (N_3060,N_2994,N_2981);
nand U3061 (N_3061,N_2978,N_2908);
or U3062 (N_3062,N_2957,N_2937);
nor U3063 (N_3063,N_2927,N_2988);
and U3064 (N_3064,N_2971,N_2963);
or U3065 (N_3065,N_2977,N_2921);
xnor U3066 (N_3066,N_2905,N_2993);
nor U3067 (N_3067,N_2950,N_2905);
xor U3068 (N_3068,N_2925,N_2927);
xor U3069 (N_3069,N_2934,N_2909);
and U3070 (N_3070,N_2972,N_2997);
xor U3071 (N_3071,N_2958,N_2928);
or U3072 (N_3072,N_2938,N_2936);
nand U3073 (N_3073,N_2928,N_2934);
nand U3074 (N_3074,N_2970,N_2991);
or U3075 (N_3075,N_2942,N_2958);
xnor U3076 (N_3076,N_2961,N_2938);
nand U3077 (N_3077,N_2942,N_2952);
or U3078 (N_3078,N_2948,N_2905);
or U3079 (N_3079,N_2974,N_2935);
or U3080 (N_3080,N_2901,N_2977);
or U3081 (N_3081,N_2998,N_2939);
xor U3082 (N_3082,N_2950,N_2906);
nand U3083 (N_3083,N_2953,N_2912);
and U3084 (N_3084,N_2948,N_2984);
and U3085 (N_3085,N_2901,N_2965);
xnor U3086 (N_3086,N_2984,N_2902);
xor U3087 (N_3087,N_2914,N_2964);
nor U3088 (N_3088,N_2972,N_2967);
xnor U3089 (N_3089,N_2975,N_2906);
nand U3090 (N_3090,N_2948,N_2979);
and U3091 (N_3091,N_2930,N_2920);
nor U3092 (N_3092,N_2907,N_2958);
nand U3093 (N_3093,N_2901,N_2933);
nor U3094 (N_3094,N_2934,N_2984);
or U3095 (N_3095,N_2940,N_2948);
nor U3096 (N_3096,N_2905,N_2991);
and U3097 (N_3097,N_2980,N_2906);
or U3098 (N_3098,N_2989,N_2967);
and U3099 (N_3099,N_2942,N_2933);
or U3100 (N_3100,N_3079,N_3057);
xnor U3101 (N_3101,N_3044,N_3089);
and U3102 (N_3102,N_3099,N_3038);
nor U3103 (N_3103,N_3026,N_3058);
nand U3104 (N_3104,N_3093,N_3060);
or U3105 (N_3105,N_3043,N_3080);
or U3106 (N_3106,N_3092,N_3055);
and U3107 (N_3107,N_3056,N_3039);
xnor U3108 (N_3108,N_3009,N_3000);
and U3109 (N_3109,N_3098,N_3027);
nand U3110 (N_3110,N_3001,N_3019);
nor U3111 (N_3111,N_3054,N_3049);
or U3112 (N_3112,N_3030,N_3090);
and U3113 (N_3113,N_3028,N_3025);
nand U3114 (N_3114,N_3004,N_3077);
or U3115 (N_3115,N_3081,N_3074);
or U3116 (N_3116,N_3006,N_3064);
or U3117 (N_3117,N_3033,N_3024);
and U3118 (N_3118,N_3013,N_3083);
nor U3119 (N_3119,N_3042,N_3072);
nor U3120 (N_3120,N_3011,N_3034);
nor U3121 (N_3121,N_3062,N_3040);
or U3122 (N_3122,N_3031,N_3018);
nand U3123 (N_3123,N_3005,N_3070);
nor U3124 (N_3124,N_3032,N_3085);
or U3125 (N_3125,N_3050,N_3035);
nor U3126 (N_3126,N_3088,N_3095);
or U3127 (N_3127,N_3084,N_3008);
xnor U3128 (N_3128,N_3047,N_3082);
nor U3129 (N_3129,N_3076,N_3022);
or U3130 (N_3130,N_3063,N_3037);
or U3131 (N_3131,N_3029,N_3007);
nor U3132 (N_3132,N_3065,N_3003);
nand U3133 (N_3133,N_3016,N_3052);
and U3134 (N_3134,N_3068,N_3096);
nand U3135 (N_3135,N_3071,N_3017);
nand U3136 (N_3136,N_3036,N_3002);
nand U3137 (N_3137,N_3073,N_3094);
nor U3138 (N_3138,N_3014,N_3059);
and U3139 (N_3139,N_3015,N_3010);
nor U3140 (N_3140,N_3023,N_3075);
or U3141 (N_3141,N_3087,N_3066);
nand U3142 (N_3142,N_3069,N_3053);
nor U3143 (N_3143,N_3067,N_3020);
or U3144 (N_3144,N_3091,N_3046);
nor U3145 (N_3145,N_3021,N_3045);
nand U3146 (N_3146,N_3012,N_3051);
or U3147 (N_3147,N_3078,N_3097);
nor U3148 (N_3148,N_3041,N_3086);
nor U3149 (N_3149,N_3061,N_3048);
or U3150 (N_3150,N_3003,N_3011);
nor U3151 (N_3151,N_3008,N_3098);
nand U3152 (N_3152,N_3012,N_3091);
or U3153 (N_3153,N_3030,N_3058);
nor U3154 (N_3154,N_3080,N_3062);
nor U3155 (N_3155,N_3025,N_3098);
xor U3156 (N_3156,N_3057,N_3044);
and U3157 (N_3157,N_3040,N_3087);
nor U3158 (N_3158,N_3003,N_3057);
nand U3159 (N_3159,N_3051,N_3007);
and U3160 (N_3160,N_3033,N_3087);
nor U3161 (N_3161,N_3029,N_3019);
nor U3162 (N_3162,N_3027,N_3026);
or U3163 (N_3163,N_3006,N_3072);
nand U3164 (N_3164,N_3037,N_3096);
nand U3165 (N_3165,N_3089,N_3069);
or U3166 (N_3166,N_3096,N_3029);
nor U3167 (N_3167,N_3081,N_3056);
or U3168 (N_3168,N_3099,N_3002);
nor U3169 (N_3169,N_3028,N_3089);
and U3170 (N_3170,N_3074,N_3080);
or U3171 (N_3171,N_3061,N_3028);
nand U3172 (N_3172,N_3071,N_3057);
or U3173 (N_3173,N_3082,N_3097);
nand U3174 (N_3174,N_3076,N_3030);
xnor U3175 (N_3175,N_3019,N_3097);
or U3176 (N_3176,N_3006,N_3026);
nor U3177 (N_3177,N_3040,N_3001);
nand U3178 (N_3178,N_3079,N_3056);
or U3179 (N_3179,N_3089,N_3025);
or U3180 (N_3180,N_3009,N_3037);
xor U3181 (N_3181,N_3053,N_3052);
nor U3182 (N_3182,N_3025,N_3035);
nor U3183 (N_3183,N_3070,N_3097);
and U3184 (N_3184,N_3053,N_3000);
nand U3185 (N_3185,N_3007,N_3048);
nand U3186 (N_3186,N_3077,N_3013);
nand U3187 (N_3187,N_3064,N_3001);
nor U3188 (N_3188,N_3049,N_3066);
or U3189 (N_3189,N_3079,N_3052);
nor U3190 (N_3190,N_3041,N_3087);
or U3191 (N_3191,N_3064,N_3090);
nor U3192 (N_3192,N_3042,N_3081);
and U3193 (N_3193,N_3022,N_3006);
or U3194 (N_3194,N_3037,N_3086);
nand U3195 (N_3195,N_3057,N_3048);
xnor U3196 (N_3196,N_3054,N_3087);
or U3197 (N_3197,N_3021,N_3013);
nor U3198 (N_3198,N_3034,N_3022);
nand U3199 (N_3199,N_3013,N_3022);
and U3200 (N_3200,N_3125,N_3159);
nand U3201 (N_3201,N_3114,N_3146);
or U3202 (N_3202,N_3135,N_3110);
nand U3203 (N_3203,N_3136,N_3118);
and U3204 (N_3204,N_3158,N_3105);
and U3205 (N_3205,N_3180,N_3153);
nand U3206 (N_3206,N_3113,N_3108);
or U3207 (N_3207,N_3196,N_3178);
or U3208 (N_3208,N_3124,N_3106);
nor U3209 (N_3209,N_3166,N_3170);
and U3210 (N_3210,N_3123,N_3120);
or U3211 (N_3211,N_3169,N_3149);
xor U3212 (N_3212,N_3126,N_3163);
or U3213 (N_3213,N_3117,N_3155);
or U3214 (N_3214,N_3168,N_3109);
nand U3215 (N_3215,N_3182,N_3141);
nand U3216 (N_3216,N_3176,N_3103);
nand U3217 (N_3217,N_3161,N_3165);
nand U3218 (N_3218,N_3139,N_3164);
or U3219 (N_3219,N_3107,N_3173);
nand U3220 (N_3220,N_3101,N_3185);
or U3221 (N_3221,N_3137,N_3160);
and U3222 (N_3222,N_3151,N_3157);
nand U3223 (N_3223,N_3111,N_3192);
and U3224 (N_3224,N_3188,N_3189);
nand U3225 (N_3225,N_3183,N_3131);
or U3226 (N_3226,N_3193,N_3142);
xor U3227 (N_3227,N_3134,N_3190);
xnor U3228 (N_3228,N_3184,N_3129);
nor U3229 (N_3229,N_3100,N_3148);
nand U3230 (N_3230,N_3197,N_3179);
and U3231 (N_3231,N_3115,N_3121);
xor U3232 (N_3232,N_3186,N_3104);
nand U3233 (N_3233,N_3143,N_3140);
nand U3234 (N_3234,N_3171,N_3175);
and U3235 (N_3235,N_3132,N_3128);
and U3236 (N_3236,N_3199,N_3167);
nand U3237 (N_3237,N_3102,N_3112);
nand U3238 (N_3238,N_3195,N_3122);
and U3239 (N_3239,N_3147,N_3133);
nor U3240 (N_3240,N_3174,N_3187);
nor U3241 (N_3241,N_3119,N_3150);
or U3242 (N_3242,N_3177,N_3156);
and U3243 (N_3243,N_3181,N_3144);
or U3244 (N_3244,N_3116,N_3145);
or U3245 (N_3245,N_3194,N_3154);
or U3246 (N_3246,N_3127,N_3198);
or U3247 (N_3247,N_3162,N_3138);
nor U3248 (N_3248,N_3172,N_3130);
nor U3249 (N_3249,N_3191,N_3152);
nor U3250 (N_3250,N_3121,N_3151);
nor U3251 (N_3251,N_3124,N_3143);
or U3252 (N_3252,N_3134,N_3161);
and U3253 (N_3253,N_3131,N_3185);
nand U3254 (N_3254,N_3160,N_3186);
or U3255 (N_3255,N_3189,N_3139);
nor U3256 (N_3256,N_3114,N_3116);
or U3257 (N_3257,N_3100,N_3116);
and U3258 (N_3258,N_3106,N_3186);
or U3259 (N_3259,N_3114,N_3170);
or U3260 (N_3260,N_3105,N_3128);
or U3261 (N_3261,N_3194,N_3116);
nor U3262 (N_3262,N_3145,N_3120);
xnor U3263 (N_3263,N_3198,N_3115);
nand U3264 (N_3264,N_3198,N_3101);
and U3265 (N_3265,N_3108,N_3126);
and U3266 (N_3266,N_3107,N_3124);
nand U3267 (N_3267,N_3197,N_3139);
nand U3268 (N_3268,N_3194,N_3178);
nor U3269 (N_3269,N_3122,N_3103);
or U3270 (N_3270,N_3191,N_3146);
nor U3271 (N_3271,N_3153,N_3135);
xnor U3272 (N_3272,N_3106,N_3193);
and U3273 (N_3273,N_3157,N_3108);
and U3274 (N_3274,N_3138,N_3185);
or U3275 (N_3275,N_3197,N_3173);
and U3276 (N_3276,N_3191,N_3159);
xnor U3277 (N_3277,N_3117,N_3188);
nand U3278 (N_3278,N_3109,N_3163);
or U3279 (N_3279,N_3142,N_3102);
or U3280 (N_3280,N_3118,N_3152);
or U3281 (N_3281,N_3168,N_3171);
or U3282 (N_3282,N_3161,N_3177);
or U3283 (N_3283,N_3124,N_3154);
or U3284 (N_3284,N_3173,N_3160);
nand U3285 (N_3285,N_3148,N_3184);
or U3286 (N_3286,N_3146,N_3190);
and U3287 (N_3287,N_3168,N_3146);
nor U3288 (N_3288,N_3125,N_3183);
xnor U3289 (N_3289,N_3183,N_3101);
nand U3290 (N_3290,N_3151,N_3158);
and U3291 (N_3291,N_3154,N_3113);
nand U3292 (N_3292,N_3165,N_3179);
nor U3293 (N_3293,N_3149,N_3148);
xnor U3294 (N_3294,N_3143,N_3186);
or U3295 (N_3295,N_3132,N_3149);
nand U3296 (N_3296,N_3198,N_3145);
nand U3297 (N_3297,N_3114,N_3136);
nor U3298 (N_3298,N_3191,N_3135);
xor U3299 (N_3299,N_3138,N_3140);
nand U3300 (N_3300,N_3266,N_3250);
xnor U3301 (N_3301,N_3234,N_3271);
or U3302 (N_3302,N_3257,N_3267);
and U3303 (N_3303,N_3279,N_3296);
or U3304 (N_3304,N_3225,N_3256);
xnor U3305 (N_3305,N_3275,N_3210);
xnor U3306 (N_3306,N_3219,N_3221);
or U3307 (N_3307,N_3263,N_3242);
and U3308 (N_3308,N_3274,N_3228);
and U3309 (N_3309,N_3265,N_3248);
nand U3310 (N_3310,N_3288,N_3224);
nor U3311 (N_3311,N_3273,N_3202);
nor U3312 (N_3312,N_3231,N_3277);
nand U3313 (N_3313,N_3203,N_3211);
and U3314 (N_3314,N_3284,N_3204);
xnor U3315 (N_3315,N_3258,N_3289);
nand U3316 (N_3316,N_3205,N_3217);
and U3317 (N_3317,N_3207,N_3206);
nor U3318 (N_3318,N_3264,N_3201);
or U3319 (N_3319,N_3213,N_3223);
nand U3320 (N_3320,N_3280,N_3227);
or U3321 (N_3321,N_3233,N_3230);
nand U3322 (N_3322,N_3209,N_3241);
nor U3323 (N_3323,N_3290,N_3281);
or U3324 (N_3324,N_3259,N_3208);
xnor U3325 (N_3325,N_3240,N_3283);
nor U3326 (N_3326,N_3286,N_3200);
or U3327 (N_3327,N_3272,N_3291);
and U3328 (N_3328,N_3237,N_3247);
nor U3329 (N_3329,N_3299,N_3293);
nor U3330 (N_3330,N_3239,N_3282);
xnor U3331 (N_3331,N_3246,N_3269);
and U3332 (N_3332,N_3226,N_3285);
or U3333 (N_3333,N_3297,N_3253);
and U3334 (N_3334,N_3244,N_3270);
nor U3335 (N_3335,N_3251,N_3236);
nor U3336 (N_3336,N_3243,N_3261);
xor U3337 (N_3337,N_3260,N_3294);
or U3338 (N_3338,N_3212,N_3238);
xnor U3339 (N_3339,N_3214,N_3262);
or U3340 (N_3340,N_3287,N_3215);
or U3341 (N_3341,N_3232,N_3278);
nand U3342 (N_3342,N_3254,N_3292);
and U3343 (N_3343,N_3268,N_3276);
or U3344 (N_3344,N_3218,N_3216);
or U3345 (N_3345,N_3229,N_3298);
and U3346 (N_3346,N_3252,N_3245);
or U3347 (N_3347,N_3249,N_3220);
or U3348 (N_3348,N_3222,N_3235);
nand U3349 (N_3349,N_3255,N_3295);
or U3350 (N_3350,N_3204,N_3242);
and U3351 (N_3351,N_3260,N_3241);
nand U3352 (N_3352,N_3254,N_3272);
xor U3353 (N_3353,N_3235,N_3298);
xnor U3354 (N_3354,N_3268,N_3259);
and U3355 (N_3355,N_3258,N_3281);
nor U3356 (N_3356,N_3202,N_3242);
and U3357 (N_3357,N_3228,N_3213);
and U3358 (N_3358,N_3240,N_3291);
or U3359 (N_3359,N_3205,N_3240);
nor U3360 (N_3360,N_3291,N_3298);
nor U3361 (N_3361,N_3240,N_3297);
and U3362 (N_3362,N_3288,N_3232);
or U3363 (N_3363,N_3289,N_3254);
and U3364 (N_3364,N_3295,N_3227);
and U3365 (N_3365,N_3277,N_3225);
nor U3366 (N_3366,N_3215,N_3229);
nor U3367 (N_3367,N_3285,N_3254);
nand U3368 (N_3368,N_3277,N_3219);
nand U3369 (N_3369,N_3251,N_3222);
and U3370 (N_3370,N_3219,N_3296);
nand U3371 (N_3371,N_3210,N_3242);
nor U3372 (N_3372,N_3296,N_3287);
or U3373 (N_3373,N_3250,N_3204);
nand U3374 (N_3374,N_3288,N_3215);
and U3375 (N_3375,N_3239,N_3210);
or U3376 (N_3376,N_3206,N_3232);
nand U3377 (N_3377,N_3234,N_3205);
xor U3378 (N_3378,N_3264,N_3289);
nor U3379 (N_3379,N_3287,N_3254);
xor U3380 (N_3380,N_3258,N_3229);
nor U3381 (N_3381,N_3230,N_3239);
nor U3382 (N_3382,N_3292,N_3272);
nor U3383 (N_3383,N_3222,N_3286);
nand U3384 (N_3384,N_3210,N_3278);
nor U3385 (N_3385,N_3278,N_3247);
or U3386 (N_3386,N_3217,N_3233);
or U3387 (N_3387,N_3208,N_3275);
nor U3388 (N_3388,N_3260,N_3293);
and U3389 (N_3389,N_3211,N_3213);
and U3390 (N_3390,N_3224,N_3268);
and U3391 (N_3391,N_3283,N_3246);
nand U3392 (N_3392,N_3211,N_3204);
or U3393 (N_3393,N_3200,N_3269);
xnor U3394 (N_3394,N_3289,N_3275);
nor U3395 (N_3395,N_3273,N_3248);
nor U3396 (N_3396,N_3276,N_3200);
nand U3397 (N_3397,N_3267,N_3214);
xor U3398 (N_3398,N_3299,N_3215);
and U3399 (N_3399,N_3215,N_3258);
nand U3400 (N_3400,N_3392,N_3394);
nand U3401 (N_3401,N_3308,N_3358);
or U3402 (N_3402,N_3377,N_3349);
nand U3403 (N_3403,N_3319,N_3348);
or U3404 (N_3404,N_3326,N_3332);
and U3405 (N_3405,N_3333,N_3318);
xor U3406 (N_3406,N_3301,N_3399);
and U3407 (N_3407,N_3396,N_3385);
and U3408 (N_3408,N_3309,N_3338);
xor U3409 (N_3409,N_3323,N_3398);
or U3410 (N_3410,N_3356,N_3371);
xnor U3411 (N_3411,N_3346,N_3357);
nand U3412 (N_3412,N_3312,N_3316);
nand U3413 (N_3413,N_3380,N_3317);
xnor U3414 (N_3414,N_3311,N_3328);
xnor U3415 (N_3415,N_3366,N_3372);
nor U3416 (N_3416,N_3376,N_3335);
and U3417 (N_3417,N_3369,N_3361);
xnor U3418 (N_3418,N_3324,N_3306);
and U3419 (N_3419,N_3381,N_3363);
or U3420 (N_3420,N_3345,N_3337);
nor U3421 (N_3421,N_3302,N_3327);
xor U3422 (N_3422,N_3354,N_3395);
and U3423 (N_3423,N_3362,N_3343);
xnor U3424 (N_3424,N_3303,N_3391);
xnor U3425 (N_3425,N_3360,N_3386);
and U3426 (N_3426,N_3350,N_3313);
nand U3427 (N_3427,N_3336,N_3367);
nor U3428 (N_3428,N_3382,N_3355);
xor U3429 (N_3429,N_3359,N_3390);
and U3430 (N_3430,N_3375,N_3364);
nor U3431 (N_3431,N_3300,N_3370);
and U3432 (N_3432,N_3365,N_3341);
xnor U3433 (N_3433,N_3310,N_3340);
nor U3434 (N_3434,N_3321,N_3387);
and U3435 (N_3435,N_3374,N_3388);
nor U3436 (N_3436,N_3322,N_3307);
nand U3437 (N_3437,N_3334,N_3329);
nor U3438 (N_3438,N_3368,N_3383);
nand U3439 (N_3439,N_3320,N_3378);
xnor U3440 (N_3440,N_3397,N_3314);
nor U3441 (N_3441,N_3315,N_3352);
or U3442 (N_3442,N_3330,N_3304);
or U3443 (N_3443,N_3353,N_3325);
xor U3444 (N_3444,N_3379,N_3373);
xnor U3445 (N_3445,N_3344,N_3389);
and U3446 (N_3446,N_3384,N_3339);
and U3447 (N_3447,N_3342,N_3393);
and U3448 (N_3448,N_3331,N_3351);
nand U3449 (N_3449,N_3347,N_3305);
or U3450 (N_3450,N_3376,N_3342);
xor U3451 (N_3451,N_3313,N_3393);
nand U3452 (N_3452,N_3386,N_3398);
or U3453 (N_3453,N_3387,N_3322);
and U3454 (N_3454,N_3353,N_3380);
nor U3455 (N_3455,N_3384,N_3368);
xor U3456 (N_3456,N_3348,N_3350);
nor U3457 (N_3457,N_3393,N_3325);
nand U3458 (N_3458,N_3311,N_3316);
xor U3459 (N_3459,N_3367,N_3379);
nand U3460 (N_3460,N_3306,N_3374);
or U3461 (N_3461,N_3390,N_3317);
nand U3462 (N_3462,N_3327,N_3370);
nor U3463 (N_3463,N_3302,N_3309);
nor U3464 (N_3464,N_3367,N_3311);
nor U3465 (N_3465,N_3306,N_3368);
nor U3466 (N_3466,N_3378,N_3386);
nor U3467 (N_3467,N_3384,N_3390);
nand U3468 (N_3468,N_3325,N_3373);
and U3469 (N_3469,N_3385,N_3342);
nor U3470 (N_3470,N_3346,N_3316);
nor U3471 (N_3471,N_3394,N_3303);
nor U3472 (N_3472,N_3376,N_3318);
and U3473 (N_3473,N_3314,N_3319);
nand U3474 (N_3474,N_3365,N_3359);
or U3475 (N_3475,N_3347,N_3342);
nand U3476 (N_3476,N_3307,N_3328);
nor U3477 (N_3477,N_3396,N_3352);
or U3478 (N_3478,N_3378,N_3322);
or U3479 (N_3479,N_3312,N_3369);
or U3480 (N_3480,N_3336,N_3366);
nand U3481 (N_3481,N_3378,N_3303);
or U3482 (N_3482,N_3304,N_3323);
nor U3483 (N_3483,N_3311,N_3360);
or U3484 (N_3484,N_3389,N_3319);
nand U3485 (N_3485,N_3358,N_3393);
or U3486 (N_3486,N_3380,N_3326);
or U3487 (N_3487,N_3336,N_3326);
nor U3488 (N_3488,N_3334,N_3317);
and U3489 (N_3489,N_3377,N_3392);
nand U3490 (N_3490,N_3342,N_3305);
nor U3491 (N_3491,N_3362,N_3353);
nor U3492 (N_3492,N_3357,N_3330);
nand U3493 (N_3493,N_3345,N_3323);
xnor U3494 (N_3494,N_3337,N_3374);
nor U3495 (N_3495,N_3346,N_3375);
nand U3496 (N_3496,N_3329,N_3300);
or U3497 (N_3497,N_3365,N_3372);
nor U3498 (N_3498,N_3338,N_3360);
or U3499 (N_3499,N_3350,N_3332);
nor U3500 (N_3500,N_3487,N_3482);
xor U3501 (N_3501,N_3476,N_3451);
xnor U3502 (N_3502,N_3440,N_3483);
nor U3503 (N_3503,N_3452,N_3479);
nor U3504 (N_3504,N_3418,N_3402);
xnor U3505 (N_3505,N_3414,N_3445);
or U3506 (N_3506,N_3404,N_3427);
nor U3507 (N_3507,N_3442,N_3461);
or U3508 (N_3508,N_3481,N_3462);
nor U3509 (N_3509,N_3416,N_3407);
nor U3510 (N_3510,N_3413,N_3465);
and U3511 (N_3511,N_3448,N_3454);
nand U3512 (N_3512,N_3496,N_3446);
and U3513 (N_3513,N_3463,N_3432);
and U3514 (N_3514,N_3449,N_3477);
or U3515 (N_3515,N_3457,N_3437);
nand U3516 (N_3516,N_3489,N_3439);
xor U3517 (N_3517,N_3405,N_3401);
nor U3518 (N_3518,N_3464,N_3420);
nand U3519 (N_3519,N_3472,N_3455);
nand U3520 (N_3520,N_3475,N_3434);
nand U3521 (N_3521,N_3466,N_3471);
nor U3522 (N_3522,N_3488,N_3467);
and U3523 (N_3523,N_3495,N_3491);
nor U3524 (N_3524,N_3456,N_3459);
or U3525 (N_3525,N_3441,N_3470);
nor U3526 (N_3526,N_3480,N_3403);
or U3527 (N_3527,N_3485,N_3490);
or U3528 (N_3528,N_3469,N_3433);
nor U3529 (N_3529,N_3423,N_3444);
nor U3530 (N_3530,N_3438,N_3435);
and U3531 (N_3531,N_3410,N_3417);
or U3532 (N_3532,N_3443,N_3412);
and U3533 (N_3533,N_3429,N_3478);
nor U3534 (N_3534,N_3415,N_3408);
and U3535 (N_3535,N_3424,N_3409);
or U3536 (N_3536,N_3400,N_3473);
or U3537 (N_3537,N_3468,N_3484);
and U3538 (N_3538,N_3497,N_3411);
nand U3539 (N_3539,N_3425,N_3430);
nand U3540 (N_3540,N_3499,N_3431);
and U3541 (N_3541,N_3450,N_3419);
or U3542 (N_3542,N_3406,N_3453);
nand U3543 (N_3543,N_3447,N_3422);
nor U3544 (N_3544,N_3428,N_3458);
xnor U3545 (N_3545,N_3436,N_3460);
or U3546 (N_3546,N_3492,N_3421);
nand U3547 (N_3547,N_3493,N_3498);
nor U3548 (N_3548,N_3474,N_3426);
xnor U3549 (N_3549,N_3494,N_3486);
nand U3550 (N_3550,N_3456,N_3480);
nand U3551 (N_3551,N_3499,N_3440);
or U3552 (N_3552,N_3494,N_3491);
nand U3553 (N_3553,N_3489,N_3473);
and U3554 (N_3554,N_3478,N_3426);
nor U3555 (N_3555,N_3442,N_3440);
xor U3556 (N_3556,N_3410,N_3453);
nand U3557 (N_3557,N_3495,N_3489);
xnor U3558 (N_3558,N_3448,N_3474);
and U3559 (N_3559,N_3451,N_3497);
nand U3560 (N_3560,N_3421,N_3408);
or U3561 (N_3561,N_3454,N_3492);
or U3562 (N_3562,N_3419,N_3403);
or U3563 (N_3563,N_3485,N_3412);
nand U3564 (N_3564,N_3414,N_3456);
or U3565 (N_3565,N_3462,N_3466);
nand U3566 (N_3566,N_3451,N_3453);
or U3567 (N_3567,N_3431,N_3444);
nand U3568 (N_3568,N_3485,N_3417);
nand U3569 (N_3569,N_3468,N_3434);
and U3570 (N_3570,N_3497,N_3417);
xor U3571 (N_3571,N_3419,N_3409);
or U3572 (N_3572,N_3408,N_3442);
xnor U3573 (N_3573,N_3405,N_3463);
xor U3574 (N_3574,N_3406,N_3490);
or U3575 (N_3575,N_3487,N_3401);
xnor U3576 (N_3576,N_3469,N_3430);
xnor U3577 (N_3577,N_3414,N_3422);
nor U3578 (N_3578,N_3444,N_3410);
nand U3579 (N_3579,N_3475,N_3467);
nor U3580 (N_3580,N_3457,N_3486);
or U3581 (N_3581,N_3485,N_3445);
nand U3582 (N_3582,N_3471,N_3485);
or U3583 (N_3583,N_3497,N_3434);
nand U3584 (N_3584,N_3414,N_3485);
nand U3585 (N_3585,N_3411,N_3431);
and U3586 (N_3586,N_3449,N_3401);
xor U3587 (N_3587,N_3476,N_3431);
xor U3588 (N_3588,N_3457,N_3472);
nand U3589 (N_3589,N_3438,N_3486);
and U3590 (N_3590,N_3495,N_3448);
or U3591 (N_3591,N_3490,N_3494);
or U3592 (N_3592,N_3461,N_3426);
and U3593 (N_3593,N_3468,N_3464);
nand U3594 (N_3594,N_3405,N_3432);
nand U3595 (N_3595,N_3405,N_3414);
or U3596 (N_3596,N_3486,N_3441);
and U3597 (N_3597,N_3413,N_3460);
or U3598 (N_3598,N_3434,N_3424);
nand U3599 (N_3599,N_3451,N_3450);
nand U3600 (N_3600,N_3538,N_3596);
nor U3601 (N_3601,N_3500,N_3551);
nand U3602 (N_3602,N_3549,N_3511);
nor U3603 (N_3603,N_3579,N_3541);
nand U3604 (N_3604,N_3576,N_3557);
or U3605 (N_3605,N_3542,N_3520);
xnor U3606 (N_3606,N_3507,N_3516);
nor U3607 (N_3607,N_3585,N_3593);
or U3608 (N_3608,N_3558,N_3563);
nand U3609 (N_3609,N_3577,N_3560);
or U3610 (N_3610,N_3513,N_3504);
nand U3611 (N_3611,N_3552,N_3573);
or U3612 (N_3612,N_3530,N_3581);
nand U3613 (N_3613,N_3567,N_3554);
or U3614 (N_3614,N_3578,N_3598);
nor U3615 (N_3615,N_3580,N_3570);
xnor U3616 (N_3616,N_3509,N_3582);
and U3617 (N_3617,N_3531,N_3595);
nor U3618 (N_3618,N_3571,N_3562);
nor U3619 (N_3619,N_3528,N_3532);
nor U3620 (N_3620,N_3508,N_3591);
nor U3621 (N_3621,N_3505,N_3583);
nor U3622 (N_3622,N_3574,N_3553);
and U3623 (N_3623,N_3556,N_3548);
nor U3624 (N_3624,N_3586,N_3568);
and U3625 (N_3625,N_3526,N_3565);
or U3626 (N_3626,N_3501,N_3517);
nand U3627 (N_3627,N_3540,N_3545);
nand U3628 (N_3628,N_3503,N_3555);
nor U3629 (N_3629,N_3575,N_3561);
nor U3630 (N_3630,N_3527,N_3539);
or U3631 (N_3631,N_3515,N_3535);
or U3632 (N_3632,N_3510,N_3522);
xor U3633 (N_3633,N_3521,N_3546);
xnor U3634 (N_3634,N_3572,N_3514);
nor U3635 (N_3635,N_3534,N_3523);
nand U3636 (N_3636,N_3506,N_3588);
xor U3637 (N_3637,N_3569,N_3599);
or U3638 (N_3638,N_3547,N_3519);
or U3639 (N_3639,N_3544,N_3559);
nand U3640 (N_3640,N_3594,N_3525);
and U3641 (N_3641,N_3512,N_3537);
and U3642 (N_3642,N_3589,N_3536);
nand U3643 (N_3643,N_3533,N_3566);
nor U3644 (N_3644,N_3502,N_3592);
and U3645 (N_3645,N_3584,N_3524);
nand U3646 (N_3646,N_3529,N_3550);
nor U3647 (N_3647,N_3597,N_3543);
nand U3648 (N_3648,N_3518,N_3587);
nor U3649 (N_3649,N_3564,N_3590);
nor U3650 (N_3650,N_3589,N_3548);
and U3651 (N_3651,N_3557,N_3534);
or U3652 (N_3652,N_3578,N_3551);
nand U3653 (N_3653,N_3535,N_3573);
nor U3654 (N_3654,N_3518,N_3571);
or U3655 (N_3655,N_3581,N_3584);
and U3656 (N_3656,N_3560,N_3524);
or U3657 (N_3657,N_3563,N_3590);
or U3658 (N_3658,N_3543,N_3500);
or U3659 (N_3659,N_3510,N_3580);
nand U3660 (N_3660,N_3514,N_3554);
nor U3661 (N_3661,N_3555,N_3553);
and U3662 (N_3662,N_3574,N_3507);
or U3663 (N_3663,N_3591,N_3574);
and U3664 (N_3664,N_3573,N_3570);
and U3665 (N_3665,N_3578,N_3500);
or U3666 (N_3666,N_3598,N_3585);
or U3667 (N_3667,N_3538,N_3515);
nor U3668 (N_3668,N_3502,N_3546);
nand U3669 (N_3669,N_3546,N_3540);
nand U3670 (N_3670,N_3553,N_3599);
nor U3671 (N_3671,N_3566,N_3524);
xnor U3672 (N_3672,N_3506,N_3554);
and U3673 (N_3673,N_3551,N_3525);
or U3674 (N_3674,N_3516,N_3539);
and U3675 (N_3675,N_3504,N_3536);
or U3676 (N_3676,N_3584,N_3575);
and U3677 (N_3677,N_3572,N_3524);
or U3678 (N_3678,N_3592,N_3565);
or U3679 (N_3679,N_3571,N_3583);
or U3680 (N_3680,N_3577,N_3595);
and U3681 (N_3681,N_3519,N_3574);
and U3682 (N_3682,N_3518,N_3524);
and U3683 (N_3683,N_3537,N_3538);
and U3684 (N_3684,N_3576,N_3514);
or U3685 (N_3685,N_3542,N_3540);
nand U3686 (N_3686,N_3510,N_3589);
or U3687 (N_3687,N_3507,N_3557);
or U3688 (N_3688,N_3542,N_3590);
nor U3689 (N_3689,N_3516,N_3546);
and U3690 (N_3690,N_3587,N_3569);
nor U3691 (N_3691,N_3517,N_3534);
and U3692 (N_3692,N_3564,N_3550);
and U3693 (N_3693,N_3539,N_3519);
nand U3694 (N_3694,N_3576,N_3594);
nand U3695 (N_3695,N_3539,N_3537);
nor U3696 (N_3696,N_3578,N_3573);
xnor U3697 (N_3697,N_3553,N_3548);
nand U3698 (N_3698,N_3555,N_3549);
nand U3699 (N_3699,N_3573,N_3554);
and U3700 (N_3700,N_3643,N_3692);
nor U3701 (N_3701,N_3687,N_3626);
and U3702 (N_3702,N_3657,N_3613);
nand U3703 (N_3703,N_3677,N_3612);
or U3704 (N_3704,N_3620,N_3669);
nor U3705 (N_3705,N_3607,N_3683);
and U3706 (N_3706,N_3698,N_3625);
nand U3707 (N_3707,N_3618,N_3637);
xor U3708 (N_3708,N_3651,N_3655);
and U3709 (N_3709,N_3686,N_3697);
nand U3710 (N_3710,N_3617,N_3601);
nand U3711 (N_3711,N_3689,N_3634);
nor U3712 (N_3712,N_3659,N_3631);
nand U3713 (N_3713,N_3662,N_3636);
and U3714 (N_3714,N_3647,N_3656);
or U3715 (N_3715,N_3638,N_3609);
xor U3716 (N_3716,N_3600,N_3693);
xor U3717 (N_3717,N_3621,N_3660);
nand U3718 (N_3718,N_3652,N_3681);
or U3719 (N_3719,N_3673,N_3679);
and U3720 (N_3720,N_3688,N_3629);
nor U3721 (N_3721,N_3653,N_3696);
nand U3722 (N_3722,N_3684,N_3602);
nand U3723 (N_3723,N_3658,N_3603);
nand U3724 (N_3724,N_3667,N_3666);
nand U3725 (N_3725,N_3690,N_3604);
nor U3726 (N_3726,N_3699,N_3668);
and U3727 (N_3727,N_3644,N_3615);
or U3728 (N_3728,N_3624,N_3676);
xnor U3729 (N_3729,N_3691,N_3645);
nor U3730 (N_3730,N_3642,N_3680);
nand U3731 (N_3731,N_3606,N_3635);
and U3732 (N_3732,N_3640,N_3611);
nor U3733 (N_3733,N_3619,N_3616);
and U3734 (N_3734,N_3622,N_3685);
or U3735 (N_3735,N_3646,N_3661);
and U3736 (N_3736,N_3608,N_3641);
and U3737 (N_3737,N_3665,N_3605);
nand U3738 (N_3738,N_3663,N_3610);
nor U3739 (N_3739,N_3633,N_3627);
xnor U3740 (N_3740,N_3654,N_3649);
nor U3741 (N_3741,N_3623,N_3664);
and U3742 (N_3742,N_3672,N_3678);
nand U3743 (N_3743,N_3671,N_3614);
xor U3744 (N_3744,N_3639,N_3650);
or U3745 (N_3745,N_3648,N_3694);
and U3746 (N_3746,N_3632,N_3670);
and U3747 (N_3747,N_3675,N_3695);
nand U3748 (N_3748,N_3630,N_3674);
nor U3749 (N_3749,N_3682,N_3628);
and U3750 (N_3750,N_3697,N_3677);
nor U3751 (N_3751,N_3603,N_3639);
or U3752 (N_3752,N_3686,N_3635);
nand U3753 (N_3753,N_3627,N_3650);
or U3754 (N_3754,N_3604,N_3616);
or U3755 (N_3755,N_3680,N_3695);
or U3756 (N_3756,N_3658,N_3694);
nand U3757 (N_3757,N_3601,N_3629);
and U3758 (N_3758,N_3683,N_3641);
and U3759 (N_3759,N_3632,N_3630);
or U3760 (N_3760,N_3601,N_3683);
nand U3761 (N_3761,N_3638,N_3651);
nor U3762 (N_3762,N_3627,N_3651);
or U3763 (N_3763,N_3637,N_3681);
and U3764 (N_3764,N_3640,N_3620);
nand U3765 (N_3765,N_3655,N_3668);
nand U3766 (N_3766,N_3698,N_3687);
nor U3767 (N_3767,N_3684,N_3650);
nand U3768 (N_3768,N_3620,N_3683);
or U3769 (N_3769,N_3691,N_3636);
and U3770 (N_3770,N_3643,N_3608);
and U3771 (N_3771,N_3689,N_3674);
or U3772 (N_3772,N_3676,N_3622);
nor U3773 (N_3773,N_3650,N_3624);
or U3774 (N_3774,N_3674,N_3650);
xor U3775 (N_3775,N_3687,N_3657);
xor U3776 (N_3776,N_3657,N_3661);
nand U3777 (N_3777,N_3643,N_3682);
nor U3778 (N_3778,N_3638,N_3669);
xnor U3779 (N_3779,N_3692,N_3649);
nor U3780 (N_3780,N_3633,N_3640);
nand U3781 (N_3781,N_3647,N_3640);
and U3782 (N_3782,N_3603,N_3685);
or U3783 (N_3783,N_3626,N_3611);
and U3784 (N_3784,N_3604,N_3655);
nand U3785 (N_3785,N_3653,N_3672);
nand U3786 (N_3786,N_3618,N_3671);
and U3787 (N_3787,N_3643,N_3647);
nand U3788 (N_3788,N_3677,N_3606);
or U3789 (N_3789,N_3614,N_3672);
nand U3790 (N_3790,N_3671,N_3617);
and U3791 (N_3791,N_3647,N_3637);
nor U3792 (N_3792,N_3613,N_3601);
nor U3793 (N_3793,N_3628,N_3616);
nor U3794 (N_3794,N_3644,N_3635);
and U3795 (N_3795,N_3621,N_3611);
and U3796 (N_3796,N_3694,N_3652);
xnor U3797 (N_3797,N_3657,N_3697);
xnor U3798 (N_3798,N_3622,N_3696);
or U3799 (N_3799,N_3696,N_3646);
nor U3800 (N_3800,N_3761,N_3702);
or U3801 (N_3801,N_3707,N_3797);
nor U3802 (N_3802,N_3794,N_3737);
nor U3803 (N_3803,N_3791,N_3785);
nor U3804 (N_3804,N_3728,N_3734);
nor U3805 (N_3805,N_3710,N_3742);
nand U3806 (N_3806,N_3744,N_3721);
or U3807 (N_3807,N_3780,N_3774);
nand U3808 (N_3808,N_3775,N_3783);
nor U3809 (N_3809,N_3747,N_3724);
nand U3810 (N_3810,N_3701,N_3757);
and U3811 (N_3811,N_3723,N_3764);
and U3812 (N_3812,N_3756,N_3735);
nor U3813 (N_3813,N_3795,N_3799);
nand U3814 (N_3814,N_3787,N_3739);
nand U3815 (N_3815,N_3700,N_3726);
nor U3816 (N_3816,N_3712,N_3762);
and U3817 (N_3817,N_3748,N_3778);
and U3818 (N_3818,N_3760,N_3770);
nand U3819 (N_3819,N_3705,N_3773);
or U3820 (N_3820,N_3715,N_3740);
or U3821 (N_3821,N_3751,N_3713);
nand U3822 (N_3822,N_3792,N_3754);
xnor U3823 (N_3823,N_3703,N_3714);
nand U3824 (N_3824,N_3769,N_3746);
or U3825 (N_3825,N_3759,N_3772);
or U3826 (N_3826,N_3750,N_3709);
nor U3827 (N_3827,N_3716,N_3763);
xnor U3828 (N_3828,N_3736,N_3755);
or U3829 (N_3829,N_3720,N_3765);
nor U3830 (N_3830,N_3786,N_3768);
nor U3831 (N_3831,N_3781,N_3771);
nand U3832 (N_3832,N_3790,N_3719);
or U3833 (N_3833,N_3796,N_3708);
nand U3834 (N_3834,N_3745,N_3706);
and U3835 (N_3835,N_3766,N_3733);
nor U3836 (N_3836,N_3704,N_3718);
nand U3837 (N_3837,N_3731,N_3788);
nor U3838 (N_3838,N_3749,N_3782);
nand U3839 (N_3839,N_3730,N_3741);
nor U3840 (N_3840,N_3779,N_3743);
nand U3841 (N_3841,N_3725,N_3722);
and U3842 (N_3842,N_3798,N_3711);
nand U3843 (N_3843,N_3789,N_3727);
or U3844 (N_3844,N_3793,N_3753);
and U3845 (N_3845,N_3776,N_3752);
nor U3846 (N_3846,N_3738,N_3784);
nand U3847 (N_3847,N_3717,N_3758);
or U3848 (N_3848,N_3732,N_3777);
and U3849 (N_3849,N_3729,N_3767);
and U3850 (N_3850,N_3716,N_3725);
xor U3851 (N_3851,N_3793,N_3786);
or U3852 (N_3852,N_3721,N_3789);
nor U3853 (N_3853,N_3701,N_3764);
and U3854 (N_3854,N_3772,N_3732);
and U3855 (N_3855,N_3776,N_3795);
nand U3856 (N_3856,N_3775,N_3719);
nand U3857 (N_3857,N_3777,N_3760);
nand U3858 (N_3858,N_3782,N_3716);
or U3859 (N_3859,N_3784,N_3754);
or U3860 (N_3860,N_3734,N_3767);
nor U3861 (N_3861,N_3782,N_3700);
or U3862 (N_3862,N_3748,N_3745);
or U3863 (N_3863,N_3731,N_3764);
nand U3864 (N_3864,N_3776,N_3784);
or U3865 (N_3865,N_3709,N_3749);
nand U3866 (N_3866,N_3726,N_3777);
nor U3867 (N_3867,N_3757,N_3730);
nand U3868 (N_3868,N_3721,N_3703);
nand U3869 (N_3869,N_3788,N_3701);
nand U3870 (N_3870,N_3780,N_3711);
nor U3871 (N_3871,N_3787,N_3711);
and U3872 (N_3872,N_3744,N_3795);
or U3873 (N_3873,N_3776,N_3728);
nand U3874 (N_3874,N_3738,N_3787);
nand U3875 (N_3875,N_3738,N_3749);
nor U3876 (N_3876,N_3728,N_3789);
nor U3877 (N_3877,N_3785,N_3781);
nand U3878 (N_3878,N_3737,N_3716);
nor U3879 (N_3879,N_3750,N_3777);
or U3880 (N_3880,N_3795,N_3715);
nor U3881 (N_3881,N_3789,N_3739);
or U3882 (N_3882,N_3706,N_3771);
and U3883 (N_3883,N_3768,N_3799);
nor U3884 (N_3884,N_3713,N_3766);
or U3885 (N_3885,N_3716,N_3722);
nor U3886 (N_3886,N_3797,N_3736);
nor U3887 (N_3887,N_3719,N_3789);
nor U3888 (N_3888,N_3771,N_3798);
and U3889 (N_3889,N_3748,N_3707);
and U3890 (N_3890,N_3756,N_3709);
and U3891 (N_3891,N_3778,N_3737);
or U3892 (N_3892,N_3712,N_3769);
and U3893 (N_3893,N_3732,N_3754);
nor U3894 (N_3894,N_3714,N_3787);
nand U3895 (N_3895,N_3788,N_3726);
xor U3896 (N_3896,N_3738,N_3706);
and U3897 (N_3897,N_3796,N_3760);
nor U3898 (N_3898,N_3729,N_3779);
nand U3899 (N_3899,N_3707,N_3737);
nor U3900 (N_3900,N_3862,N_3802);
nor U3901 (N_3901,N_3889,N_3849);
nand U3902 (N_3902,N_3846,N_3803);
xor U3903 (N_3903,N_3817,N_3820);
nand U3904 (N_3904,N_3872,N_3855);
and U3905 (N_3905,N_3808,N_3809);
and U3906 (N_3906,N_3813,N_3891);
nor U3907 (N_3907,N_3870,N_3888);
nor U3908 (N_3908,N_3871,N_3859);
nand U3909 (N_3909,N_3860,N_3829);
or U3910 (N_3910,N_3822,N_3895);
or U3911 (N_3911,N_3818,N_3836);
and U3912 (N_3912,N_3801,N_3816);
or U3913 (N_3913,N_3831,N_3805);
or U3914 (N_3914,N_3876,N_3841);
nand U3915 (N_3915,N_3812,N_3847);
xnor U3916 (N_3916,N_3873,N_3894);
or U3917 (N_3917,N_3807,N_3844);
nand U3918 (N_3918,N_3858,N_3877);
and U3919 (N_3919,N_3857,N_3887);
or U3920 (N_3920,N_3897,N_3842);
or U3921 (N_3921,N_3845,N_3843);
or U3922 (N_3922,N_3806,N_3875);
nor U3923 (N_3923,N_3800,N_3821);
nand U3924 (N_3924,N_3838,N_3856);
or U3925 (N_3925,N_3825,N_3810);
or U3926 (N_3926,N_3832,N_3835);
nand U3927 (N_3927,N_3882,N_3861);
and U3928 (N_3928,N_3823,N_3826);
and U3929 (N_3929,N_3828,N_3804);
and U3930 (N_3930,N_3839,N_3898);
nor U3931 (N_3931,N_3881,N_3886);
nor U3932 (N_3932,N_3853,N_3884);
nor U3933 (N_3933,N_3830,N_3892);
nor U3934 (N_3934,N_3878,N_3852);
nor U3935 (N_3935,N_3867,N_3850);
nand U3936 (N_3936,N_3851,N_3854);
xor U3937 (N_3937,N_3814,N_3834);
or U3938 (N_3938,N_3883,N_3879);
nor U3939 (N_3939,N_3819,N_3874);
nand U3940 (N_3940,N_3893,N_3840);
nand U3941 (N_3941,N_3815,N_3869);
or U3942 (N_3942,N_3880,N_3827);
or U3943 (N_3943,N_3824,N_3899);
nand U3944 (N_3944,N_3885,N_3896);
and U3945 (N_3945,N_3833,N_3866);
or U3946 (N_3946,N_3890,N_3868);
xor U3947 (N_3947,N_3837,N_3864);
and U3948 (N_3948,N_3863,N_3865);
and U3949 (N_3949,N_3811,N_3848);
nor U3950 (N_3950,N_3866,N_3874);
and U3951 (N_3951,N_3813,N_3810);
and U3952 (N_3952,N_3869,N_3800);
xor U3953 (N_3953,N_3821,N_3824);
nor U3954 (N_3954,N_3883,N_3840);
or U3955 (N_3955,N_3860,N_3898);
or U3956 (N_3956,N_3864,N_3876);
nand U3957 (N_3957,N_3891,N_3821);
or U3958 (N_3958,N_3895,N_3880);
nand U3959 (N_3959,N_3860,N_3899);
nor U3960 (N_3960,N_3887,N_3897);
nand U3961 (N_3961,N_3823,N_3883);
and U3962 (N_3962,N_3828,N_3809);
nor U3963 (N_3963,N_3850,N_3848);
nor U3964 (N_3964,N_3818,N_3891);
and U3965 (N_3965,N_3891,N_3834);
and U3966 (N_3966,N_3877,N_3884);
or U3967 (N_3967,N_3862,N_3861);
nor U3968 (N_3968,N_3836,N_3876);
xnor U3969 (N_3969,N_3810,N_3853);
or U3970 (N_3970,N_3830,N_3836);
nand U3971 (N_3971,N_3870,N_3869);
or U3972 (N_3972,N_3842,N_3817);
nor U3973 (N_3973,N_3839,N_3881);
or U3974 (N_3974,N_3811,N_3851);
and U3975 (N_3975,N_3871,N_3848);
or U3976 (N_3976,N_3827,N_3845);
nor U3977 (N_3977,N_3854,N_3866);
nand U3978 (N_3978,N_3826,N_3889);
and U3979 (N_3979,N_3844,N_3870);
nand U3980 (N_3980,N_3840,N_3881);
and U3981 (N_3981,N_3894,N_3863);
xor U3982 (N_3982,N_3871,N_3893);
nand U3983 (N_3983,N_3810,N_3803);
and U3984 (N_3984,N_3813,N_3847);
or U3985 (N_3985,N_3821,N_3817);
xnor U3986 (N_3986,N_3813,N_3896);
nor U3987 (N_3987,N_3826,N_3834);
nor U3988 (N_3988,N_3871,N_3820);
nor U3989 (N_3989,N_3841,N_3816);
and U3990 (N_3990,N_3885,N_3898);
nor U3991 (N_3991,N_3899,N_3893);
or U3992 (N_3992,N_3821,N_3881);
nor U3993 (N_3993,N_3868,N_3843);
or U3994 (N_3994,N_3861,N_3899);
nor U3995 (N_3995,N_3834,N_3858);
nor U3996 (N_3996,N_3821,N_3804);
and U3997 (N_3997,N_3831,N_3890);
or U3998 (N_3998,N_3859,N_3806);
and U3999 (N_3999,N_3818,N_3831);
nand U4000 (N_4000,N_3905,N_3978);
nor U4001 (N_4001,N_3907,N_3968);
nand U4002 (N_4002,N_3982,N_3931);
nand U4003 (N_4003,N_3949,N_3997);
nand U4004 (N_4004,N_3952,N_3993);
xnor U4005 (N_4005,N_3918,N_3954);
nor U4006 (N_4006,N_3950,N_3937);
or U4007 (N_4007,N_3960,N_3924);
or U4008 (N_4008,N_3955,N_3929);
or U4009 (N_4009,N_3930,N_3974);
and U4010 (N_4010,N_3919,N_3958);
or U4011 (N_4011,N_3951,N_3987);
nor U4012 (N_4012,N_3983,N_3944);
or U4013 (N_4013,N_3957,N_3956);
nor U4014 (N_4014,N_3946,N_3995);
nand U4015 (N_4015,N_3922,N_3981);
xnor U4016 (N_4016,N_3940,N_3991);
and U4017 (N_4017,N_3994,N_3965);
xor U4018 (N_4018,N_3900,N_3909);
or U4019 (N_4019,N_3923,N_3904);
nor U4020 (N_4020,N_3917,N_3935);
nor U4021 (N_4021,N_3962,N_3986);
and U4022 (N_4022,N_3976,N_3925);
or U4023 (N_4023,N_3933,N_3927);
nand U4024 (N_4024,N_3911,N_3953);
nand U4025 (N_4025,N_3912,N_3926);
nor U4026 (N_4026,N_3967,N_3932);
or U4027 (N_4027,N_3998,N_3945);
nand U4028 (N_4028,N_3969,N_3902);
and U4029 (N_4029,N_3910,N_3939);
and U4030 (N_4030,N_3990,N_3914);
and U4031 (N_4031,N_3943,N_3988);
nor U4032 (N_4032,N_3915,N_3948);
nand U4033 (N_4033,N_3947,N_3928);
nand U4034 (N_4034,N_3996,N_3984);
nand U4035 (N_4035,N_3979,N_3985);
xnor U4036 (N_4036,N_3973,N_3999);
and U4037 (N_4037,N_3916,N_3920);
nand U4038 (N_4038,N_3959,N_3961);
xnor U4039 (N_4039,N_3975,N_3906);
xnor U4040 (N_4040,N_3992,N_3964);
and U4041 (N_4041,N_3980,N_3941);
nand U4042 (N_4042,N_3942,N_3989);
or U4043 (N_4043,N_3903,N_3913);
or U4044 (N_4044,N_3977,N_3901);
nand U4045 (N_4045,N_3963,N_3966);
nor U4046 (N_4046,N_3934,N_3921);
nand U4047 (N_4047,N_3908,N_3938);
or U4048 (N_4048,N_3970,N_3972);
or U4049 (N_4049,N_3936,N_3971);
nor U4050 (N_4050,N_3932,N_3920);
nand U4051 (N_4051,N_3944,N_3900);
nor U4052 (N_4052,N_3921,N_3995);
and U4053 (N_4053,N_3909,N_3925);
nor U4054 (N_4054,N_3987,N_3972);
and U4055 (N_4055,N_3938,N_3983);
nand U4056 (N_4056,N_3990,N_3909);
nor U4057 (N_4057,N_3976,N_3932);
nor U4058 (N_4058,N_3976,N_3945);
nand U4059 (N_4059,N_3956,N_3959);
nor U4060 (N_4060,N_3933,N_3975);
and U4061 (N_4061,N_3959,N_3995);
nand U4062 (N_4062,N_3974,N_3941);
nor U4063 (N_4063,N_3953,N_3903);
nand U4064 (N_4064,N_3954,N_3930);
and U4065 (N_4065,N_3948,N_3958);
nand U4066 (N_4066,N_3937,N_3934);
xor U4067 (N_4067,N_3981,N_3982);
xnor U4068 (N_4068,N_3937,N_3956);
or U4069 (N_4069,N_3911,N_3944);
nand U4070 (N_4070,N_3943,N_3976);
and U4071 (N_4071,N_3998,N_3905);
nand U4072 (N_4072,N_3926,N_3955);
nand U4073 (N_4073,N_3993,N_3907);
nor U4074 (N_4074,N_3985,N_3933);
nor U4075 (N_4075,N_3911,N_3957);
or U4076 (N_4076,N_3953,N_3995);
or U4077 (N_4077,N_3910,N_3997);
nor U4078 (N_4078,N_3969,N_3938);
and U4079 (N_4079,N_3983,N_3955);
and U4080 (N_4080,N_3910,N_3917);
and U4081 (N_4081,N_3945,N_3982);
and U4082 (N_4082,N_3994,N_3980);
or U4083 (N_4083,N_3998,N_3974);
nand U4084 (N_4084,N_3990,N_3910);
or U4085 (N_4085,N_3907,N_3965);
nand U4086 (N_4086,N_3915,N_3952);
nand U4087 (N_4087,N_3908,N_3946);
nor U4088 (N_4088,N_3946,N_3909);
or U4089 (N_4089,N_3922,N_3908);
or U4090 (N_4090,N_3965,N_3998);
nor U4091 (N_4091,N_3981,N_3907);
xor U4092 (N_4092,N_3924,N_3995);
nor U4093 (N_4093,N_3914,N_3931);
or U4094 (N_4094,N_3908,N_3984);
xor U4095 (N_4095,N_3980,N_3954);
nand U4096 (N_4096,N_3958,N_3988);
xnor U4097 (N_4097,N_3904,N_3984);
and U4098 (N_4098,N_3996,N_3907);
nor U4099 (N_4099,N_3902,N_3952);
nand U4100 (N_4100,N_4028,N_4020);
and U4101 (N_4101,N_4009,N_4039);
or U4102 (N_4102,N_4018,N_4015);
nor U4103 (N_4103,N_4070,N_4002);
xnor U4104 (N_4104,N_4060,N_4030);
or U4105 (N_4105,N_4025,N_4029);
nand U4106 (N_4106,N_4097,N_4095);
and U4107 (N_4107,N_4023,N_4014);
nand U4108 (N_4108,N_4036,N_4048);
or U4109 (N_4109,N_4057,N_4092);
and U4110 (N_4110,N_4037,N_4049);
nand U4111 (N_4111,N_4019,N_4050);
nor U4112 (N_4112,N_4079,N_4027);
and U4113 (N_4113,N_4081,N_4006);
and U4114 (N_4114,N_4098,N_4089);
or U4115 (N_4115,N_4091,N_4063);
or U4116 (N_4116,N_4088,N_4004);
nand U4117 (N_4117,N_4040,N_4044);
nand U4118 (N_4118,N_4072,N_4033);
or U4119 (N_4119,N_4055,N_4064);
or U4120 (N_4120,N_4077,N_4061);
nor U4121 (N_4121,N_4065,N_4071);
nor U4122 (N_4122,N_4052,N_4085);
nand U4123 (N_4123,N_4068,N_4035);
nor U4124 (N_4124,N_4042,N_4096);
and U4125 (N_4125,N_4007,N_4086);
nand U4126 (N_4126,N_4026,N_4008);
nor U4127 (N_4127,N_4032,N_4003);
nor U4128 (N_4128,N_4001,N_4093);
and U4129 (N_4129,N_4075,N_4038);
nand U4130 (N_4130,N_4056,N_4021);
nor U4131 (N_4131,N_4012,N_4046);
or U4132 (N_4132,N_4067,N_4066);
and U4133 (N_4133,N_4087,N_4054);
or U4134 (N_4134,N_4078,N_4094);
nor U4135 (N_4135,N_4047,N_4041);
or U4136 (N_4136,N_4045,N_4069);
nand U4137 (N_4137,N_4031,N_4090);
nor U4138 (N_4138,N_4043,N_4010);
or U4139 (N_4139,N_4011,N_4082);
nor U4140 (N_4140,N_4034,N_4051);
xor U4141 (N_4141,N_4080,N_4053);
and U4142 (N_4142,N_4059,N_4013);
and U4143 (N_4143,N_4062,N_4076);
xor U4144 (N_4144,N_4000,N_4024);
or U4145 (N_4145,N_4073,N_4058);
nor U4146 (N_4146,N_4084,N_4099);
xnor U4147 (N_4147,N_4083,N_4016);
nor U4148 (N_4148,N_4017,N_4022);
and U4149 (N_4149,N_4005,N_4074);
nor U4150 (N_4150,N_4044,N_4052);
and U4151 (N_4151,N_4046,N_4083);
and U4152 (N_4152,N_4040,N_4006);
and U4153 (N_4153,N_4045,N_4034);
and U4154 (N_4154,N_4043,N_4068);
or U4155 (N_4155,N_4052,N_4088);
nor U4156 (N_4156,N_4045,N_4003);
and U4157 (N_4157,N_4090,N_4049);
and U4158 (N_4158,N_4066,N_4056);
or U4159 (N_4159,N_4087,N_4022);
nand U4160 (N_4160,N_4005,N_4011);
nand U4161 (N_4161,N_4060,N_4049);
nand U4162 (N_4162,N_4011,N_4074);
and U4163 (N_4163,N_4006,N_4059);
and U4164 (N_4164,N_4058,N_4022);
xor U4165 (N_4165,N_4034,N_4032);
nor U4166 (N_4166,N_4074,N_4036);
nand U4167 (N_4167,N_4067,N_4008);
or U4168 (N_4168,N_4013,N_4073);
nand U4169 (N_4169,N_4055,N_4003);
or U4170 (N_4170,N_4091,N_4078);
nor U4171 (N_4171,N_4004,N_4086);
nor U4172 (N_4172,N_4040,N_4063);
nor U4173 (N_4173,N_4019,N_4033);
and U4174 (N_4174,N_4081,N_4016);
nand U4175 (N_4175,N_4036,N_4056);
nor U4176 (N_4176,N_4040,N_4056);
xor U4177 (N_4177,N_4029,N_4018);
and U4178 (N_4178,N_4056,N_4016);
nor U4179 (N_4179,N_4084,N_4002);
nor U4180 (N_4180,N_4053,N_4074);
nand U4181 (N_4181,N_4050,N_4013);
nand U4182 (N_4182,N_4075,N_4080);
nand U4183 (N_4183,N_4037,N_4097);
or U4184 (N_4184,N_4007,N_4000);
or U4185 (N_4185,N_4009,N_4049);
or U4186 (N_4186,N_4073,N_4050);
nor U4187 (N_4187,N_4030,N_4012);
or U4188 (N_4188,N_4042,N_4008);
nor U4189 (N_4189,N_4029,N_4076);
or U4190 (N_4190,N_4052,N_4043);
xor U4191 (N_4191,N_4039,N_4043);
nand U4192 (N_4192,N_4067,N_4016);
xnor U4193 (N_4193,N_4091,N_4050);
nor U4194 (N_4194,N_4055,N_4043);
nor U4195 (N_4195,N_4037,N_4058);
nor U4196 (N_4196,N_4075,N_4032);
or U4197 (N_4197,N_4096,N_4012);
and U4198 (N_4198,N_4014,N_4040);
xor U4199 (N_4199,N_4044,N_4084);
nand U4200 (N_4200,N_4165,N_4179);
xnor U4201 (N_4201,N_4146,N_4128);
xor U4202 (N_4202,N_4185,N_4175);
nand U4203 (N_4203,N_4178,N_4142);
or U4204 (N_4204,N_4139,N_4169);
or U4205 (N_4205,N_4123,N_4158);
and U4206 (N_4206,N_4120,N_4137);
nand U4207 (N_4207,N_4188,N_4162);
and U4208 (N_4208,N_4184,N_4148);
or U4209 (N_4209,N_4134,N_4144);
nor U4210 (N_4210,N_4180,N_4107);
nor U4211 (N_4211,N_4164,N_4135);
or U4212 (N_4212,N_4122,N_4194);
and U4213 (N_4213,N_4112,N_4125);
or U4214 (N_4214,N_4102,N_4159);
or U4215 (N_4215,N_4132,N_4190);
nor U4216 (N_4216,N_4171,N_4111);
nand U4217 (N_4217,N_4105,N_4174);
nand U4218 (N_4218,N_4108,N_4183);
and U4219 (N_4219,N_4193,N_4197);
or U4220 (N_4220,N_4116,N_4104);
nor U4221 (N_4221,N_4155,N_4191);
nor U4222 (N_4222,N_4189,N_4126);
nor U4223 (N_4223,N_4152,N_4121);
xor U4224 (N_4224,N_4196,N_4109);
nand U4225 (N_4225,N_4172,N_4115);
nor U4226 (N_4226,N_4161,N_4127);
nor U4227 (N_4227,N_4100,N_4129);
nor U4228 (N_4228,N_4182,N_4198);
or U4229 (N_4229,N_4150,N_4143);
nand U4230 (N_4230,N_4199,N_4176);
nand U4231 (N_4231,N_4140,N_4149);
and U4232 (N_4232,N_4101,N_4173);
nand U4233 (N_4233,N_4130,N_4136);
or U4234 (N_4234,N_4181,N_4145);
nand U4235 (N_4235,N_4157,N_4113);
and U4236 (N_4236,N_4156,N_4151);
or U4237 (N_4237,N_4118,N_4153);
nor U4238 (N_4238,N_4163,N_4187);
nand U4239 (N_4239,N_4154,N_4160);
or U4240 (N_4240,N_4114,N_4166);
or U4241 (N_4241,N_4141,N_4119);
nor U4242 (N_4242,N_4131,N_4147);
or U4243 (N_4243,N_4170,N_4195);
nor U4244 (N_4244,N_4106,N_4124);
and U4245 (N_4245,N_4138,N_4177);
nor U4246 (N_4246,N_4117,N_4186);
nor U4247 (N_4247,N_4103,N_4168);
or U4248 (N_4248,N_4167,N_4110);
and U4249 (N_4249,N_4192,N_4133);
nand U4250 (N_4250,N_4165,N_4158);
and U4251 (N_4251,N_4145,N_4126);
and U4252 (N_4252,N_4152,N_4101);
nor U4253 (N_4253,N_4114,N_4103);
nand U4254 (N_4254,N_4139,N_4146);
or U4255 (N_4255,N_4113,N_4148);
and U4256 (N_4256,N_4156,N_4127);
or U4257 (N_4257,N_4124,N_4100);
or U4258 (N_4258,N_4104,N_4192);
nand U4259 (N_4259,N_4111,N_4113);
nor U4260 (N_4260,N_4168,N_4136);
and U4261 (N_4261,N_4132,N_4163);
nor U4262 (N_4262,N_4104,N_4141);
and U4263 (N_4263,N_4139,N_4116);
or U4264 (N_4264,N_4178,N_4189);
or U4265 (N_4265,N_4117,N_4127);
and U4266 (N_4266,N_4150,N_4128);
nor U4267 (N_4267,N_4129,N_4111);
nand U4268 (N_4268,N_4162,N_4132);
nor U4269 (N_4269,N_4161,N_4104);
xor U4270 (N_4270,N_4112,N_4163);
xor U4271 (N_4271,N_4111,N_4182);
or U4272 (N_4272,N_4162,N_4147);
or U4273 (N_4273,N_4197,N_4186);
nand U4274 (N_4274,N_4137,N_4149);
xor U4275 (N_4275,N_4186,N_4165);
xor U4276 (N_4276,N_4178,N_4190);
and U4277 (N_4277,N_4113,N_4105);
nor U4278 (N_4278,N_4156,N_4174);
nand U4279 (N_4279,N_4191,N_4154);
nor U4280 (N_4280,N_4110,N_4116);
and U4281 (N_4281,N_4164,N_4114);
nor U4282 (N_4282,N_4140,N_4196);
and U4283 (N_4283,N_4112,N_4175);
nand U4284 (N_4284,N_4108,N_4135);
nor U4285 (N_4285,N_4104,N_4131);
nor U4286 (N_4286,N_4104,N_4196);
nor U4287 (N_4287,N_4190,N_4109);
and U4288 (N_4288,N_4103,N_4178);
nand U4289 (N_4289,N_4106,N_4164);
nor U4290 (N_4290,N_4187,N_4101);
nor U4291 (N_4291,N_4145,N_4103);
or U4292 (N_4292,N_4136,N_4141);
nor U4293 (N_4293,N_4186,N_4169);
nor U4294 (N_4294,N_4171,N_4107);
nor U4295 (N_4295,N_4193,N_4181);
nor U4296 (N_4296,N_4133,N_4128);
and U4297 (N_4297,N_4197,N_4168);
and U4298 (N_4298,N_4112,N_4122);
or U4299 (N_4299,N_4106,N_4121);
nand U4300 (N_4300,N_4293,N_4299);
nor U4301 (N_4301,N_4296,N_4294);
and U4302 (N_4302,N_4262,N_4210);
nor U4303 (N_4303,N_4255,N_4241);
or U4304 (N_4304,N_4284,N_4274);
or U4305 (N_4305,N_4251,N_4295);
or U4306 (N_4306,N_4283,N_4235);
nor U4307 (N_4307,N_4245,N_4277);
and U4308 (N_4308,N_4271,N_4227);
and U4309 (N_4309,N_4263,N_4261);
and U4310 (N_4310,N_4268,N_4289);
and U4311 (N_4311,N_4240,N_4265);
nor U4312 (N_4312,N_4228,N_4202);
or U4313 (N_4313,N_4288,N_4249);
nor U4314 (N_4314,N_4282,N_4244);
nor U4315 (N_4315,N_4243,N_4290);
nand U4316 (N_4316,N_4220,N_4231);
and U4317 (N_4317,N_4211,N_4232);
and U4318 (N_4318,N_4256,N_4205);
or U4319 (N_4319,N_4246,N_4201);
nor U4320 (N_4320,N_4209,N_4203);
or U4321 (N_4321,N_4258,N_4229);
or U4322 (N_4322,N_4272,N_4225);
nand U4323 (N_4323,N_4221,N_4242);
and U4324 (N_4324,N_4279,N_4212);
or U4325 (N_4325,N_4219,N_4257);
nor U4326 (N_4326,N_4286,N_4238);
or U4327 (N_4327,N_4234,N_4208);
or U4328 (N_4328,N_4278,N_4247);
xnor U4329 (N_4329,N_4207,N_4236);
nor U4330 (N_4330,N_4269,N_4204);
nor U4331 (N_4331,N_4291,N_4224);
and U4332 (N_4332,N_4270,N_4285);
nand U4333 (N_4333,N_4200,N_4223);
nand U4334 (N_4334,N_4267,N_4217);
or U4335 (N_4335,N_4297,N_4287);
nor U4336 (N_4336,N_4233,N_4275);
xor U4337 (N_4337,N_4266,N_4213);
nand U4338 (N_4338,N_4248,N_4298);
or U4339 (N_4339,N_4254,N_4215);
nor U4340 (N_4340,N_4218,N_4264);
nand U4341 (N_4341,N_4281,N_4206);
or U4342 (N_4342,N_4259,N_4280);
and U4343 (N_4343,N_4226,N_4292);
or U4344 (N_4344,N_4216,N_4260);
nand U4345 (N_4345,N_4239,N_4273);
and U4346 (N_4346,N_4252,N_4250);
nor U4347 (N_4347,N_4253,N_4222);
or U4348 (N_4348,N_4237,N_4276);
nor U4349 (N_4349,N_4214,N_4230);
and U4350 (N_4350,N_4262,N_4252);
nand U4351 (N_4351,N_4271,N_4294);
nor U4352 (N_4352,N_4210,N_4277);
and U4353 (N_4353,N_4243,N_4236);
or U4354 (N_4354,N_4235,N_4297);
and U4355 (N_4355,N_4278,N_4255);
nor U4356 (N_4356,N_4237,N_4233);
nor U4357 (N_4357,N_4293,N_4289);
xnor U4358 (N_4358,N_4203,N_4284);
or U4359 (N_4359,N_4231,N_4257);
nor U4360 (N_4360,N_4210,N_4285);
nand U4361 (N_4361,N_4256,N_4206);
or U4362 (N_4362,N_4240,N_4274);
nor U4363 (N_4363,N_4288,N_4279);
nand U4364 (N_4364,N_4290,N_4220);
nand U4365 (N_4365,N_4233,N_4299);
or U4366 (N_4366,N_4246,N_4248);
nand U4367 (N_4367,N_4285,N_4278);
and U4368 (N_4368,N_4284,N_4264);
or U4369 (N_4369,N_4237,N_4260);
and U4370 (N_4370,N_4227,N_4222);
xnor U4371 (N_4371,N_4265,N_4299);
xnor U4372 (N_4372,N_4229,N_4250);
nor U4373 (N_4373,N_4257,N_4286);
nor U4374 (N_4374,N_4249,N_4214);
xor U4375 (N_4375,N_4237,N_4274);
nand U4376 (N_4376,N_4224,N_4289);
nor U4377 (N_4377,N_4299,N_4228);
and U4378 (N_4378,N_4256,N_4274);
or U4379 (N_4379,N_4283,N_4231);
xnor U4380 (N_4380,N_4201,N_4234);
nand U4381 (N_4381,N_4210,N_4201);
and U4382 (N_4382,N_4210,N_4293);
and U4383 (N_4383,N_4295,N_4247);
nand U4384 (N_4384,N_4205,N_4295);
and U4385 (N_4385,N_4297,N_4242);
xor U4386 (N_4386,N_4260,N_4217);
nand U4387 (N_4387,N_4250,N_4271);
or U4388 (N_4388,N_4206,N_4291);
and U4389 (N_4389,N_4263,N_4223);
and U4390 (N_4390,N_4280,N_4249);
nand U4391 (N_4391,N_4265,N_4221);
nand U4392 (N_4392,N_4201,N_4203);
or U4393 (N_4393,N_4223,N_4213);
and U4394 (N_4394,N_4287,N_4286);
and U4395 (N_4395,N_4230,N_4272);
nand U4396 (N_4396,N_4253,N_4245);
nor U4397 (N_4397,N_4238,N_4259);
nand U4398 (N_4398,N_4211,N_4240);
and U4399 (N_4399,N_4216,N_4206);
or U4400 (N_4400,N_4349,N_4384);
xor U4401 (N_4401,N_4320,N_4371);
nor U4402 (N_4402,N_4387,N_4385);
nor U4403 (N_4403,N_4375,N_4309);
nor U4404 (N_4404,N_4302,N_4393);
xor U4405 (N_4405,N_4350,N_4382);
nand U4406 (N_4406,N_4333,N_4397);
and U4407 (N_4407,N_4368,N_4334);
nand U4408 (N_4408,N_4359,N_4342);
and U4409 (N_4409,N_4327,N_4366);
and U4410 (N_4410,N_4300,N_4325);
nand U4411 (N_4411,N_4391,N_4328);
nor U4412 (N_4412,N_4311,N_4389);
and U4413 (N_4413,N_4338,N_4316);
nor U4414 (N_4414,N_4326,N_4318);
nand U4415 (N_4415,N_4360,N_4364);
or U4416 (N_4416,N_4345,N_4352);
and U4417 (N_4417,N_4370,N_4329);
or U4418 (N_4418,N_4388,N_4337);
or U4419 (N_4419,N_4357,N_4324);
or U4420 (N_4420,N_4367,N_4376);
and U4421 (N_4421,N_4390,N_4344);
nand U4422 (N_4422,N_4336,N_4301);
nor U4423 (N_4423,N_4373,N_4378);
or U4424 (N_4424,N_4340,N_4358);
and U4425 (N_4425,N_4335,N_4396);
nand U4426 (N_4426,N_4313,N_4395);
nor U4427 (N_4427,N_4322,N_4317);
and U4428 (N_4428,N_4372,N_4305);
nand U4429 (N_4429,N_4381,N_4347);
and U4430 (N_4430,N_4374,N_4356);
or U4431 (N_4431,N_4380,N_4392);
nor U4432 (N_4432,N_4399,N_4304);
nand U4433 (N_4433,N_4343,N_4383);
or U4434 (N_4434,N_4323,N_4361);
or U4435 (N_4435,N_4353,N_4354);
or U4436 (N_4436,N_4306,N_4348);
nor U4437 (N_4437,N_4310,N_4346);
and U4438 (N_4438,N_4362,N_4312);
nor U4439 (N_4439,N_4369,N_4330);
and U4440 (N_4440,N_4365,N_4351);
or U4441 (N_4441,N_4339,N_4331);
nor U4442 (N_4442,N_4314,N_4363);
nor U4443 (N_4443,N_4307,N_4394);
and U4444 (N_4444,N_4379,N_4321);
and U4445 (N_4445,N_4315,N_4355);
and U4446 (N_4446,N_4386,N_4303);
or U4447 (N_4447,N_4319,N_4341);
nand U4448 (N_4448,N_4308,N_4377);
nor U4449 (N_4449,N_4332,N_4398);
xnor U4450 (N_4450,N_4303,N_4367);
xor U4451 (N_4451,N_4396,N_4325);
or U4452 (N_4452,N_4357,N_4399);
nor U4453 (N_4453,N_4315,N_4344);
or U4454 (N_4454,N_4329,N_4312);
nand U4455 (N_4455,N_4380,N_4315);
or U4456 (N_4456,N_4374,N_4365);
nand U4457 (N_4457,N_4389,N_4387);
nor U4458 (N_4458,N_4305,N_4366);
nor U4459 (N_4459,N_4356,N_4332);
nand U4460 (N_4460,N_4351,N_4310);
xor U4461 (N_4461,N_4316,N_4311);
xnor U4462 (N_4462,N_4346,N_4380);
nor U4463 (N_4463,N_4314,N_4386);
nor U4464 (N_4464,N_4360,N_4314);
or U4465 (N_4465,N_4314,N_4326);
or U4466 (N_4466,N_4366,N_4344);
nor U4467 (N_4467,N_4319,N_4356);
nor U4468 (N_4468,N_4316,N_4367);
or U4469 (N_4469,N_4362,N_4395);
nor U4470 (N_4470,N_4385,N_4355);
nand U4471 (N_4471,N_4321,N_4332);
nand U4472 (N_4472,N_4316,N_4344);
and U4473 (N_4473,N_4301,N_4395);
xor U4474 (N_4474,N_4300,N_4370);
nor U4475 (N_4475,N_4304,N_4387);
nor U4476 (N_4476,N_4342,N_4307);
or U4477 (N_4477,N_4399,N_4385);
and U4478 (N_4478,N_4383,N_4395);
nand U4479 (N_4479,N_4366,N_4390);
or U4480 (N_4480,N_4350,N_4371);
and U4481 (N_4481,N_4339,N_4388);
xnor U4482 (N_4482,N_4346,N_4303);
nor U4483 (N_4483,N_4300,N_4354);
nand U4484 (N_4484,N_4397,N_4347);
nor U4485 (N_4485,N_4349,N_4393);
nor U4486 (N_4486,N_4309,N_4329);
nor U4487 (N_4487,N_4382,N_4321);
or U4488 (N_4488,N_4342,N_4312);
or U4489 (N_4489,N_4339,N_4314);
nor U4490 (N_4490,N_4317,N_4348);
nor U4491 (N_4491,N_4302,N_4335);
or U4492 (N_4492,N_4304,N_4346);
nand U4493 (N_4493,N_4353,N_4385);
xnor U4494 (N_4494,N_4342,N_4341);
or U4495 (N_4495,N_4326,N_4306);
or U4496 (N_4496,N_4304,N_4362);
nor U4497 (N_4497,N_4332,N_4394);
nand U4498 (N_4498,N_4330,N_4353);
and U4499 (N_4499,N_4341,N_4311);
nand U4500 (N_4500,N_4429,N_4406);
or U4501 (N_4501,N_4421,N_4495);
and U4502 (N_4502,N_4449,N_4424);
xor U4503 (N_4503,N_4401,N_4482);
and U4504 (N_4504,N_4445,N_4480);
and U4505 (N_4505,N_4461,N_4439);
and U4506 (N_4506,N_4434,N_4441);
nand U4507 (N_4507,N_4436,N_4426);
or U4508 (N_4508,N_4454,N_4417);
nand U4509 (N_4509,N_4452,N_4438);
and U4510 (N_4510,N_4492,N_4405);
and U4511 (N_4511,N_4412,N_4404);
and U4512 (N_4512,N_4494,N_4464);
nand U4513 (N_4513,N_4456,N_4423);
nand U4514 (N_4514,N_4428,N_4422);
and U4515 (N_4515,N_4444,N_4443);
nand U4516 (N_4516,N_4447,N_4458);
nand U4517 (N_4517,N_4498,N_4446);
nand U4518 (N_4518,N_4431,N_4471);
or U4519 (N_4519,N_4460,N_4453);
and U4520 (N_4520,N_4437,N_4465);
and U4521 (N_4521,N_4468,N_4408);
or U4522 (N_4522,N_4493,N_4470);
and U4523 (N_4523,N_4466,N_4425);
nand U4524 (N_4524,N_4488,N_4403);
or U4525 (N_4525,N_4472,N_4467);
nand U4526 (N_4526,N_4400,N_4486);
nor U4527 (N_4527,N_4418,N_4407);
nand U4528 (N_4528,N_4442,N_4419);
nor U4529 (N_4529,N_4415,N_4410);
nand U4530 (N_4530,N_4451,N_4499);
or U4531 (N_4531,N_4420,N_4490);
or U4532 (N_4532,N_4477,N_4496);
xor U4533 (N_4533,N_4432,N_4416);
nand U4534 (N_4534,N_4459,N_4440);
nor U4535 (N_4535,N_4487,N_4489);
and U4536 (N_4536,N_4473,N_4484);
and U4537 (N_4537,N_4435,N_4474);
nor U4538 (N_4538,N_4491,N_4483);
or U4539 (N_4539,N_4450,N_4476);
nand U4540 (N_4540,N_4462,N_4463);
and U4541 (N_4541,N_4485,N_4448);
nor U4542 (N_4542,N_4455,N_4402);
or U4543 (N_4543,N_4457,N_4413);
or U4544 (N_4544,N_4430,N_4497);
and U4545 (N_4545,N_4481,N_4411);
and U4546 (N_4546,N_4478,N_4427);
or U4547 (N_4547,N_4414,N_4409);
xor U4548 (N_4548,N_4433,N_4469);
or U4549 (N_4549,N_4475,N_4479);
nor U4550 (N_4550,N_4445,N_4493);
nor U4551 (N_4551,N_4457,N_4469);
nand U4552 (N_4552,N_4403,N_4424);
nor U4553 (N_4553,N_4421,N_4485);
or U4554 (N_4554,N_4450,N_4489);
nand U4555 (N_4555,N_4498,N_4481);
or U4556 (N_4556,N_4475,N_4400);
nand U4557 (N_4557,N_4483,N_4470);
nand U4558 (N_4558,N_4478,N_4443);
or U4559 (N_4559,N_4420,N_4436);
xnor U4560 (N_4560,N_4457,N_4448);
or U4561 (N_4561,N_4452,N_4491);
nor U4562 (N_4562,N_4475,N_4469);
xnor U4563 (N_4563,N_4445,N_4453);
and U4564 (N_4564,N_4474,N_4494);
and U4565 (N_4565,N_4427,N_4464);
nand U4566 (N_4566,N_4451,N_4427);
nor U4567 (N_4567,N_4423,N_4466);
or U4568 (N_4568,N_4498,N_4486);
nor U4569 (N_4569,N_4464,N_4415);
nand U4570 (N_4570,N_4427,N_4457);
or U4571 (N_4571,N_4438,N_4444);
nand U4572 (N_4572,N_4475,N_4444);
xnor U4573 (N_4573,N_4464,N_4418);
nand U4574 (N_4574,N_4418,N_4406);
and U4575 (N_4575,N_4481,N_4432);
nand U4576 (N_4576,N_4487,N_4442);
nor U4577 (N_4577,N_4447,N_4488);
nor U4578 (N_4578,N_4440,N_4404);
nand U4579 (N_4579,N_4420,N_4469);
xnor U4580 (N_4580,N_4446,N_4416);
nand U4581 (N_4581,N_4478,N_4459);
and U4582 (N_4582,N_4487,N_4420);
nor U4583 (N_4583,N_4441,N_4459);
nor U4584 (N_4584,N_4427,N_4473);
or U4585 (N_4585,N_4493,N_4451);
or U4586 (N_4586,N_4492,N_4444);
or U4587 (N_4587,N_4439,N_4401);
and U4588 (N_4588,N_4427,N_4498);
nor U4589 (N_4589,N_4472,N_4446);
and U4590 (N_4590,N_4458,N_4411);
or U4591 (N_4591,N_4490,N_4404);
nor U4592 (N_4592,N_4445,N_4483);
nand U4593 (N_4593,N_4466,N_4405);
and U4594 (N_4594,N_4448,N_4429);
xnor U4595 (N_4595,N_4455,N_4459);
or U4596 (N_4596,N_4461,N_4450);
and U4597 (N_4597,N_4430,N_4492);
or U4598 (N_4598,N_4493,N_4408);
nor U4599 (N_4599,N_4447,N_4414);
nor U4600 (N_4600,N_4509,N_4520);
and U4601 (N_4601,N_4586,N_4566);
xnor U4602 (N_4602,N_4594,N_4523);
nand U4603 (N_4603,N_4541,N_4505);
and U4604 (N_4604,N_4512,N_4536);
nor U4605 (N_4605,N_4560,N_4576);
nand U4606 (N_4606,N_4574,N_4588);
nor U4607 (N_4607,N_4501,N_4545);
nand U4608 (N_4608,N_4521,N_4587);
nand U4609 (N_4609,N_4514,N_4510);
xor U4610 (N_4610,N_4506,N_4518);
nor U4611 (N_4611,N_4579,N_4556);
or U4612 (N_4612,N_4583,N_4548);
nand U4613 (N_4613,N_4559,N_4546);
nor U4614 (N_4614,N_4567,N_4551);
or U4615 (N_4615,N_4504,N_4511);
and U4616 (N_4616,N_4530,N_4585);
and U4617 (N_4617,N_4584,N_4565);
nor U4618 (N_4618,N_4571,N_4543);
and U4619 (N_4619,N_4528,N_4570);
or U4620 (N_4620,N_4581,N_4508);
or U4621 (N_4621,N_4589,N_4533);
nand U4622 (N_4622,N_4593,N_4526);
nand U4623 (N_4623,N_4500,N_4544);
and U4624 (N_4624,N_4519,N_4539);
and U4625 (N_4625,N_4564,N_4580);
or U4626 (N_4626,N_4557,N_4569);
nand U4627 (N_4627,N_4590,N_4524);
xnor U4628 (N_4628,N_4563,N_4540);
nand U4629 (N_4629,N_4535,N_4527);
and U4630 (N_4630,N_4575,N_4542);
or U4631 (N_4631,N_4578,N_4529);
nand U4632 (N_4632,N_4522,N_4547);
and U4633 (N_4633,N_4553,N_4532);
or U4634 (N_4634,N_4513,N_4549);
nor U4635 (N_4635,N_4507,N_4537);
nor U4636 (N_4636,N_4561,N_4515);
and U4637 (N_4637,N_4525,N_4502);
nor U4638 (N_4638,N_4597,N_4531);
or U4639 (N_4639,N_4555,N_4573);
nand U4640 (N_4640,N_4552,N_4503);
nor U4641 (N_4641,N_4572,N_4596);
or U4642 (N_4642,N_4562,N_4534);
and U4643 (N_4643,N_4598,N_4558);
xnor U4644 (N_4644,N_4550,N_4599);
xor U4645 (N_4645,N_4538,N_4568);
nor U4646 (N_4646,N_4516,N_4554);
or U4647 (N_4647,N_4591,N_4577);
or U4648 (N_4648,N_4595,N_4592);
or U4649 (N_4649,N_4517,N_4582);
nor U4650 (N_4650,N_4530,N_4587);
and U4651 (N_4651,N_4589,N_4596);
and U4652 (N_4652,N_4523,N_4589);
nand U4653 (N_4653,N_4528,N_4537);
nand U4654 (N_4654,N_4519,N_4573);
nand U4655 (N_4655,N_4570,N_4541);
or U4656 (N_4656,N_4545,N_4508);
or U4657 (N_4657,N_4572,N_4553);
nor U4658 (N_4658,N_4531,N_4599);
or U4659 (N_4659,N_4540,N_4596);
nand U4660 (N_4660,N_4524,N_4553);
and U4661 (N_4661,N_4518,N_4519);
nand U4662 (N_4662,N_4501,N_4502);
and U4663 (N_4663,N_4561,N_4518);
or U4664 (N_4664,N_4552,N_4594);
or U4665 (N_4665,N_4521,N_4598);
nand U4666 (N_4666,N_4558,N_4591);
nand U4667 (N_4667,N_4571,N_4539);
nand U4668 (N_4668,N_4550,N_4585);
nor U4669 (N_4669,N_4581,N_4587);
and U4670 (N_4670,N_4513,N_4528);
or U4671 (N_4671,N_4568,N_4588);
nand U4672 (N_4672,N_4510,N_4554);
nor U4673 (N_4673,N_4567,N_4555);
or U4674 (N_4674,N_4580,N_4533);
or U4675 (N_4675,N_4553,N_4501);
xor U4676 (N_4676,N_4561,N_4519);
or U4677 (N_4677,N_4536,N_4565);
and U4678 (N_4678,N_4526,N_4517);
nor U4679 (N_4679,N_4516,N_4555);
nor U4680 (N_4680,N_4507,N_4577);
or U4681 (N_4681,N_4562,N_4567);
nand U4682 (N_4682,N_4501,N_4527);
nor U4683 (N_4683,N_4502,N_4507);
nor U4684 (N_4684,N_4580,N_4510);
and U4685 (N_4685,N_4512,N_4505);
and U4686 (N_4686,N_4598,N_4520);
and U4687 (N_4687,N_4583,N_4557);
xor U4688 (N_4688,N_4571,N_4589);
nor U4689 (N_4689,N_4526,N_4534);
or U4690 (N_4690,N_4539,N_4597);
nand U4691 (N_4691,N_4573,N_4533);
nand U4692 (N_4692,N_4539,N_4547);
nor U4693 (N_4693,N_4563,N_4556);
nor U4694 (N_4694,N_4524,N_4567);
and U4695 (N_4695,N_4510,N_4539);
xor U4696 (N_4696,N_4588,N_4561);
and U4697 (N_4697,N_4587,N_4538);
nor U4698 (N_4698,N_4598,N_4551);
or U4699 (N_4699,N_4508,N_4589);
xor U4700 (N_4700,N_4672,N_4641);
nor U4701 (N_4701,N_4658,N_4686);
nor U4702 (N_4702,N_4628,N_4639);
nand U4703 (N_4703,N_4695,N_4643);
or U4704 (N_4704,N_4619,N_4629);
nand U4705 (N_4705,N_4683,N_4656);
nor U4706 (N_4706,N_4687,N_4652);
nand U4707 (N_4707,N_4657,N_4671);
xor U4708 (N_4708,N_4689,N_4668);
and U4709 (N_4709,N_4644,N_4670);
and U4710 (N_4710,N_4616,N_4623);
nand U4711 (N_4711,N_4609,N_4667);
nor U4712 (N_4712,N_4621,N_4648);
nand U4713 (N_4713,N_4693,N_4655);
and U4714 (N_4714,N_4692,N_4622);
nor U4715 (N_4715,N_4696,N_4605);
or U4716 (N_4716,N_4649,N_4633);
and U4717 (N_4717,N_4646,N_4624);
or U4718 (N_4718,N_4614,N_4676);
nand U4719 (N_4719,N_4678,N_4602);
or U4720 (N_4720,N_4613,N_4675);
nor U4721 (N_4721,N_4680,N_4679);
or U4722 (N_4722,N_4632,N_4610);
xor U4723 (N_4723,N_4640,N_4663);
nor U4724 (N_4724,N_4688,N_4631);
nor U4725 (N_4725,N_4625,N_4669);
or U4726 (N_4726,N_4664,N_4603);
xnor U4727 (N_4727,N_4608,N_4682);
and U4728 (N_4728,N_4665,N_4626);
or U4729 (N_4729,N_4691,N_4637);
nor U4730 (N_4730,N_4650,N_4677);
and U4731 (N_4731,N_4674,N_4666);
nor U4732 (N_4732,N_4636,N_4660);
xor U4733 (N_4733,N_4698,N_4654);
nor U4734 (N_4734,N_4617,N_4630);
xnor U4735 (N_4735,N_4647,N_4627);
and U4736 (N_4736,N_4635,N_4673);
xor U4737 (N_4737,N_4653,N_4634);
nand U4738 (N_4738,N_4651,N_4685);
and U4739 (N_4739,N_4618,N_4638);
nor U4740 (N_4740,N_4681,N_4694);
or U4741 (N_4741,N_4684,N_4607);
xnor U4742 (N_4742,N_4600,N_4642);
nor U4743 (N_4743,N_4659,N_4604);
and U4744 (N_4744,N_4601,N_4699);
nor U4745 (N_4745,N_4615,N_4662);
and U4746 (N_4746,N_4620,N_4661);
and U4747 (N_4747,N_4697,N_4611);
and U4748 (N_4748,N_4612,N_4645);
and U4749 (N_4749,N_4606,N_4690);
nor U4750 (N_4750,N_4651,N_4637);
nor U4751 (N_4751,N_4608,N_4612);
nand U4752 (N_4752,N_4691,N_4622);
nor U4753 (N_4753,N_4678,N_4622);
nor U4754 (N_4754,N_4698,N_4643);
xor U4755 (N_4755,N_4681,N_4672);
and U4756 (N_4756,N_4643,N_4682);
or U4757 (N_4757,N_4685,N_4691);
nor U4758 (N_4758,N_4677,N_4694);
nand U4759 (N_4759,N_4609,N_4605);
nor U4760 (N_4760,N_4667,N_4658);
or U4761 (N_4761,N_4630,N_4607);
and U4762 (N_4762,N_4651,N_4667);
or U4763 (N_4763,N_4697,N_4604);
nand U4764 (N_4764,N_4685,N_4695);
and U4765 (N_4765,N_4680,N_4637);
nor U4766 (N_4766,N_4654,N_4625);
and U4767 (N_4767,N_4691,N_4635);
and U4768 (N_4768,N_4687,N_4670);
and U4769 (N_4769,N_4665,N_4605);
nand U4770 (N_4770,N_4653,N_4668);
and U4771 (N_4771,N_4669,N_4696);
nand U4772 (N_4772,N_4615,N_4696);
nand U4773 (N_4773,N_4657,N_4689);
xor U4774 (N_4774,N_4672,N_4625);
nor U4775 (N_4775,N_4639,N_4689);
nand U4776 (N_4776,N_4621,N_4600);
nor U4777 (N_4777,N_4650,N_4619);
nand U4778 (N_4778,N_4657,N_4603);
xnor U4779 (N_4779,N_4625,N_4651);
nor U4780 (N_4780,N_4660,N_4613);
or U4781 (N_4781,N_4674,N_4697);
and U4782 (N_4782,N_4664,N_4648);
or U4783 (N_4783,N_4681,N_4628);
or U4784 (N_4784,N_4675,N_4684);
xor U4785 (N_4785,N_4621,N_4603);
nor U4786 (N_4786,N_4640,N_4627);
and U4787 (N_4787,N_4605,N_4682);
and U4788 (N_4788,N_4685,N_4648);
nand U4789 (N_4789,N_4666,N_4637);
nand U4790 (N_4790,N_4687,N_4641);
or U4791 (N_4791,N_4636,N_4624);
nor U4792 (N_4792,N_4629,N_4660);
or U4793 (N_4793,N_4687,N_4609);
nand U4794 (N_4794,N_4640,N_4646);
and U4795 (N_4795,N_4640,N_4691);
and U4796 (N_4796,N_4689,N_4665);
xor U4797 (N_4797,N_4692,N_4694);
nand U4798 (N_4798,N_4689,N_4675);
and U4799 (N_4799,N_4679,N_4647);
and U4800 (N_4800,N_4724,N_4740);
or U4801 (N_4801,N_4760,N_4731);
nand U4802 (N_4802,N_4704,N_4776);
nand U4803 (N_4803,N_4784,N_4748);
or U4804 (N_4804,N_4737,N_4793);
nand U4805 (N_4805,N_4723,N_4735);
or U4806 (N_4806,N_4712,N_4791);
nor U4807 (N_4807,N_4769,N_4759);
xnor U4808 (N_4808,N_4774,N_4715);
and U4809 (N_4809,N_4753,N_4746);
and U4810 (N_4810,N_4777,N_4703);
nand U4811 (N_4811,N_4750,N_4734);
xnor U4812 (N_4812,N_4782,N_4743);
xor U4813 (N_4813,N_4721,N_4718);
and U4814 (N_4814,N_4755,N_4739);
or U4815 (N_4815,N_4716,N_4762);
nand U4816 (N_4816,N_4745,N_4781);
and U4817 (N_4817,N_4742,N_4770);
xor U4818 (N_4818,N_4756,N_4713);
or U4819 (N_4819,N_4780,N_4727);
xor U4820 (N_4820,N_4797,N_4720);
or U4821 (N_4821,N_4796,N_4729);
nor U4822 (N_4822,N_4763,N_4767);
nand U4823 (N_4823,N_4794,N_4786);
nor U4824 (N_4824,N_4709,N_4736);
or U4825 (N_4825,N_4701,N_4717);
nor U4826 (N_4826,N_4772,N_4741);
and U4827 (N_4827,N_4757,N_4700);
nor U4828 (N_4828,N_4738,N_4788);
nor U4829 (N_4829,N_4771,N_4726);
and U4830 (N_4830,N_4725,N_4768);
or U4831 (N_4831,N_4744,N_4752);
or U4832 (N_4832,N_4706,N_4778);
or U4833 (N_4833,N_4758,N_4775);
nand U4834 (N_4834,N_4730,N_4708);
nand U4835 (N_4835,N_4714,N_4785);
and U4836 (N_4836,N_4719,N_4789);
and U4837 (N_4837,N_4799,N_4798);
nand U4838 (N_4838,N_4732,N_4761);
nand U4839 (N_4839,N_4783,N_4705);
nand U4840 (N_4840,N_4765,N_4792);
nor U4841 (N_4841,N_4766,N_4728);
and U4842 (N_4842,N_4779,N_4795);
or U4843 (N_4843,N_4722,N_4749);
xnor U4844 (N_4844,N_4733,N_4773);
nor U4845 (N_4845,N_4702,N_4747);
nand U4846 (N_4846,N_4711,N_4764);
nand U4847 (N_4847,N_4787,N_4707);
nor U4848 (N_4848,N_4710,N_4751);
and U4849 (N_4849,N_4754,N_4790);
nand U4850 (N_4850,N_4755,N_4793);
and U4851 (N_4851,N_4707,N_4724);
and U4852 (N_4852,N_4728,N_4794);
or U4853 (N_4853,N_4738,N_4772);
and U4854 (N_4854,N_4715,N_4767);
nor U4855 (N_4855,N_4784,N_4722);
xor U4856 (N_4856,N_4787,N_4772);
and U4857 (N_4857,N_4734,N_4784);
nor U4858 (N_4858,N_4717,N_4762);
or U4859 (N_4859,N_4774,N_4796);
and U4860 (N_4860,N_4766,N_4747);
xnor U4861 (N_4861,N_4788,N_4789);
or U4862 (N_4862,N_4725,N_4750);
xor U4863 (N_4863,N_4723,N_4761);
or U4864 (N_4864,N_4702,N_4785);
nor U4865 (N_4865,N_4799,N_4775);
or U4866 (N_4866,N_4793,N_4760);
nor U4867 (N_4867,N_4731,N_4745);
and U4868 (N_4868,N_4759,N_4755);
nand U4869 (N_4869,N_4703,N_4707);
nand U4870 (N_4870,N_4727,N_4711);
nand U4871 (N_4871,N_4738,N_4700);
nor U4872 (N_4872,N_4742,N_4700);
nor U4873 (N_4873,N_4703,N_4766);
and U4874 (N_4874,N_4766,N_4780);
or U4875 (N_4875,N_4713,N_4754);
and U4876 (N_4876,N_4724,N_4705);
or U4877 (N_4877,N_4772,N_4759);
nor U4878 (N_4878,N_4727,N_4794);
or U4879 (N_4879,N_4736,N_4752);
and U4880 (N_4880,N_4769,N_4721);
nand U4881 (N_4881,N_4729,N_4721);
nor U4882 (N_4882,N_4700,N_4747);
and U4883 (N_4883,N_4741,N_4703);
and U4884 (N_4884,N_4713,N_4744);
nand U4885 (N_4885,N_4712,N_4714);
or U4886 (N_4886,N_4752,N_4742);
nor U4887 (N_4887,N_4753,N_4750);
nand U4888 (N_4888,N_4785,N_4777);
or U4889 (N_4889,N_4786,N_4779);
nand U4890 (N_4890,N_4770,N_4713);
nor U4891 (N_4891,N_4736,N_4747);
and U4892 (N_4892,N_4724,N_4782);
xnor U4893 (N_4893,N_4722,N_4743);
nor U4894 (N_4894,N_4707,N_4734);
nor U4895 (N_4895,N_4742,N_4749);
and U4896 (N_4896,N_4700,N_4714);
or U4897 (N_4897,N_4753,N_4795);
nor U4898 (N_4898,N_4729,N_4791);
nand U4899 (N_4899,N_4750,N_4798);
nor U4900 (N_4900,N_4863,N_4888);
nand U4901 (N_4901,N_4803,N_4894);
nor U4902 (N_4902,N_4866,N_4800);
xor U4903 (N_4903,N_4857,N_4886);
or U4904 (N_4904,N_4835,N_4841);
nor U4905 (N_4905,N_4865,N_4873);
nand U4906 (N_4906,N_4860,N_4870);
and U4907 (N_4907,N_4819,N_4817);
nor U4908 (N_4908,N_4878,N_4869);
or U4909 (N_4909,N_4896,N_4809);
or U4910 (N_4910,N_4864,N_4899);
nor U4911 (N_4911,N_4858,N_4887);
or U4912 (N_4912,N_4832,N_4859);
and U4913 (N_4913,N_4845,N_4823);
nor U4914 (N_4914,N_4893,N_4812);
and U4915 (N_4915,N_4884,N_4880);
or U4916 (N_4916,N_4808,N_4848);
and U4917 (N_4917,N_4871,N_4862);
nor U4918 (N_4918,N_4889,N_4810);
nand U4919 (N_4919,N_4892,N_4822);
or U4920 (N_4920,N_4801,N_4851);
nor U4921 (N_4921,N_4806,N_4849);
nand U4922 (N_4922,N_4831,N_4853);
and U4923 (N_4923,N_4842,N_4883);
nor U4924 (N_4924,N_4839,N_4890);
and U4925 (N_4925,N_4818,N_4898);
xnor U4926 (N_4926,N_4885,N_4837);
and U4927 (N_4927,N_4847,N_4824);
and U4928 (N_4928,N_4850,N_4821);
and U4929 (N_4929,N_4879,N_4895);
xnor U4930 (N_4930,N_4833,N_4867);
nand U4931 (N_4931,N_4874,N_4852);
xnor U4932 (N_4932,N_4811,N_4876);
nand U4933 (N_4933,N_4827,N_4813);
nand U4934 (N_4934,N_4814,N_4844);
or U4935 (N_4935,N_4897,N_4882);
or U4936 (N_4936,N_4825,N_4820);
or U4937 (N_4937,N_4802,N_4861);
nand U4938 (N_4938,N_4881,N_4816);
and U4939 (N_4939,N_4834,N_4891);
nor U4940 (N_4940,N_4828,N_4826);
and U4941 (N_4941,N_4846,N_4843);
nand U4942 (N_4942,N_4836,N_4804);
xor U4943 (N_4943,N_4854,N_4875);
nand U4944 (N_4944,N_4877,N_4807);
or U4945 (N_4945,N_4838,N_4868);
xor U4946 (N_4946,N_4829,N_4830);
nor U4947 (N_4947,N_4856,N_4840);
and U4948 (N_4948,N_4872,N_4855);
nor U4949 (N_4949,N_4805,N_4815);
and U4950 (N_4950,N_4801,N_4809);
nor U4951 (N_4951,N_4859,N_4834);
and U4952 (N_4952,N_4898,N_4840);
nand U4953 (N_4953,N_4826,N_4831);
nor U4954 (N_4954,N_4899,N_4866);
nor U4955 (N_4955,N_4858,N_4831);
xnor U4956 (N_4956,N_4823,N_4873);
or U4957 (N_4957,N_4857,N_4829);
or U4958 (N_4958,N_4811,N_4856);
or U4959 (N_4959,N_4893,N_4825);
nand U4960 (N_4960,N_4840,N_4804);
nand U4961 (N_4961,N_4870,N_4886);
nand U4962 (N_4962,N_4843,N_4856);
and U4963 (N_4963,N_4812,N_4849);
or U4964 (N_4964,N_4808,N_4822);
xor U4965 (N_4965,N_4817,N_4839);
nand U4966 (N_4966,N_4891,N_4865);
nand U4967 (N_4967,N_4867,N_4815);
or U4968 (N_4968,N_4840,N_4870);
nor U4969 (N_4969,N_4836,N_4851);
and U4970 (N_4970,N_4842,N_4833);
and U4971 (N_4971,N_4851,N_4879);
or U4972 (N_4972,N_4821,N_4882);
and U4973 (N_4973,N_4853,N_4805);
or U4974 (N_4974,N_4875,N_4876);
and U4975 (N_4975,N_4897,N_4865);
nand U4976 (N_4976,N_4812,N_4867);
and U4977 (N_4977,N_4824,N_4859);
and U4978 (N_4978,N_4854,N_4831);
nor U4979 (N_4979,N_4839,N_4885);
and U4980 (N_4980,N_4811,N_4847);
nand U4981 (N_4981,N_4899,N_4813);
nor U4982 (N_4982,N_4871,N_4802);
nand U4983 (N_4983,N_4871,N_4846);
and U4984 (N_4984,N_4871,N_4870);
nand U4985 (N_4985,N_4812,N_4857);
nor U4986 (N_4986,N_4848,N_4844);
nand U4987 (N_4987,N_4817,N_4838);
nand U4988 (N_4988,N_4808,N_4897);
and U4989 (N_4989,N_4868,N_4819);
nand U4990 (N_4990,N_4866,N_4810);
or U4991 (N_4991,N_4898,N_4826);
and U4992 (N_4992,N_4817,N_4872);
xor U4993 (N_4993,N_4812,N_4807);
and U4994 (N_4994,N_4891,N_4828);
nand U4995 (N_4995,N_4855,N_4894);
nand U4996 (N_4996,N_4854,N_4841);
or U4997 (N_4997,N_4849,N_4814);
or U4998 (N_4998,N_4836,N_4865);
or U4999 (N_4999,N_4882,N_4841);
xor U5000 (N_5000,N_4970,N_4919);
and U5001 (N_5001,N_4986,N_4905);
xor U5002 (N_5002,N_4983,N_4985);
nor U5003 (N_5003,N_4994,N_4922);
nor U5004 (N_5004,N_4920,N_4929);
or U5005 (N_5005,N_4987,N_4947);
and U5006 (N_5006,N_4921,N_4961);
or U5007 (N_5007,N_4950,N_4954);
nor U5008 (N_5008,N_4923,N_4917);
or U5009 (N_5009,N_4981,N_4984);
or U5010 (N_5010,N_4907,N_4980);
xor U5011 (N_5011,N_4932,N_4924);
and U5012 (N_5012,N_4957,N_4912);
and U5013 (N_5013,N_4992,N_4995);
and U5014 (N_5014,N_4925,N_4900);
nor U5015 (N_5015,N_4903,N_4938);
or U5016 (N_5016,N_4951,N_4944);
nand U5017 (N_5017,N_4963,N_4931);
and U5018 (N_5018,N_4936,N_4955);
nand U5019 (N_5019,N_4967,N_4909);
nand U5020 (N_5020,N_4948,N_4916);
and U5021 (N_5021,N_4974,N_4962);
nor U5022 (N_5022,N_4959,N_4915);
or U5023 (N_5023,N_4953,N_4945);
xor U5024 (N_5024,N_4940,N_4952);
nor U5025 (N_5025,N_4902,N_4941);
nor U5026 (N_5026,N_4949,N_4906);
and U5027 (N_5027,N_4937,N_4979);
and U5028 (N_5028,N_4911,N_4930);
xor U5029 (N_5029,N_4966,N_4965);
nor U5030 (N_5030,N_4989,N_4998);
nor U5031 (N_5031,N_4914,N_4960);
nand U5032 (N_5032,N_4972,N_4934);
nand U5033 (N_5033,N_4964,N_4997);
nand U5034 (N_5034,N_4975,N_4993);
nand U5035 (N_5035,N_4928,N_4976);
nand U5036 (N_5036,N_4926,N_4996);
nand U5037 (N_5037,N_4956,N_4904);
and U5038 (N_5038,N_4910,N_4978);
xor U5039 (N_5039,N_4933,N_4935);
xor U5040 (N_5040,N_4918,N_4943);
and U5041 (N_5041,N_4968,N_4969);
and U5042 (N_5042,N_4913,N_4999);
or U5043 (N_5043,N_4908,N_4927);
nand U5044 (N_5044,N_4982,N_4971);
nand U5045 (N_5045,N_4977,N_4990);
xnor U5046 (N_5046,N_4988,N_4946);
nand U5047 (N_5047,N_4991,N_4973);
xor U5048 (N_5048,N_4958,N_4942);
or U5049 (N_5049,N_4901,N_4939);
nand U5050 (N_5050,N_4961,N_4993);
nand U5051 (N_5051,N_4964,N_4904);
and U5052 (N_5052,N_4938,N_4934);
nand U5053 (N_5053,N_4967,N_4948);
or U5054 (N_5054,N_4978,N_4934);
nor U5055 (N_5055,N_4984,N_4941);
or U5056 (N_5056,N_4952,N_4916);
nor U5057 (N_5057,N_4904,N_4937);
and U5058 (N_5058,N_4912,N_4981);
or U5059 (N_5059,N_4915,N_4963);
or U5060 (N_5060,N_4926,N_4974);
or U5061 (N_5061,N_4934,N_4908);
nor U5062 (N_5062,N_4952,N_4958);
or U5063 (N_5063,N_4981,N_4920);
and U5064 (N_5064,N_4998,N_4913);
nand U5065 (N_5065,N_4969,N_4941);
nor U5066 (N_5066,N_4981,N_4902);
nand U5067 (N_5067,N_4975,N_4905);
nand U5068 (N_5068,N_4975,N_4979);
and U5069 (N_5069,N_4982,N_4958);
nor U5070 (N_5070,N_4929,N_4938);
nand U5071 (N_5071,N_4919,N_4989);
and U5072 (N_5072,N_4988,N_4926);
nor U5073 (N_5073,N_4927,N_4968);
or U5074 (N_5074,N_4951,N_4933);
and U5075 (N_5075,N_4926,N_4946);
and U5076 (N_5076,N_4920,N_4931);
and U5077 (N_5077,N_4953,N_4955);
nor U5078 (N_5078,N_4925,N_4905);
xor U5079 (N_5079,N_4942,N_4931);
and U5080 (N_5080,N_4989,N_4937);
nor U5081 (N_5081,N_4925,N_4914);
or U5082 (N_5082,N_4922,N_4911);
or U5083 (N_5083,N_4920,N_4968);
or U5084 (N_5084,N_4934,N_4918);
or U5085 (N_5085,N_4967,N_4990);
nand U5086 (N_5086,N_4970,N_4976);
nor U5087 (N_5087,N_4915,N_4923);
xnor U5088 (N_5088,N_4961,N_4900);
nor U5089 (N_5089,N_4922,N_4996);
or U5090 (N_5090,N_4994,N_4906);
nand U5091 (N_5091,N_4990,N_4931);
nand U5092 (N_5092,N_4991,N_4988);
and U5093 (N_5093,N_4903,N_4936);
and U5094 (N_5094,N_4921,N_4944);
or U5095 (N_5095,N_4927,N_4958);
or U5096 (N_5096,N_4942,N_4914);
or U5097 (N_5097,N_4907,N_4979);
nand U5098 (N_5098,N_4958,N_4916);
nor U5099 (N_5099,N_4947,N_4979);
nor U5100 (N_5100,N_5053,N_5018);
nand U5101 (N_5101,N_5007,N_5095);
or U5102 (N_5102,N_5063,N_5036);
or U5103 (N_5103,N_5049,N_5017);
and U5104 (N_5104,N_5052,N_5088);
nor U5105 (N_5105,N_5026,N_5070);
and U5106 (N_5106,N_5084,N_5065);
nand U5107 (N_5107,N_5034,N_5091);
xor U5108 (N_5108,N_5081,N_5093);
nor U5109 (N_5109,N_5069,N_5031);
xnor U5110 (N_5110,N_5032,N_5048);
nand U5111 (N_5111,N_5020,N_5011);
and U5112 (N_5112,N_5012,N_5074);
and U5113 (N_5113,N_5078,N_5073);
xnor U5114 (N_5114,N_5046,N_5077);
nor U5115 (N_5115,N_5066,N_5056);
or U5116 (N_5116,N_5006,N_5042);
nand U5117 (N_5117,N_5089,N_5039);
or U5118 (N_5118,N_5086,N_5041);
and U5119 (N_5119,N_5071,N_5055);
nor U5120 (N_5120,N_5067,N_5044);
or U5121 (N_5121,N_5021,N_5057);
nor U5122 (N_5122,N_5075,N_5000);
and U5123 (N_5123,N_5085,N_5094);
nand U5124 (N_5124,N_5099,N_5019);
nor U5125 (N_5125,N_5028,N_5054);
or U5126 (N_5126,N_5016,N_5090);
and U5127 (N_5127,N_5029,N_5058);
nand U5128 (N_5128,N_5047,N_5037);
and U5129 (N_5129,N_5083,N_5022);
xor U5130 (N_5130,N_5009,N_5072);
nand U5131 (N_5131,N_5061,N_5015);
nand U5132 (N_5132,N_5033,N_5064);
or U5133 (N_5133,N_5024,N_5035);
nor U5134 (N_5134,N_5003,N_5027);
nor U5135 (N_5135,N_5025,N_5051);
and U5136 (N_5136,N_5087,N_5068);
and U5137 (N_5137,N_5043,N_5045);
nor U5138 (N_5138,N_5040,N_5038);
xor U5139 (N_5139,N_5098,N_5013);
xnor U5140 (N_5140,N_5097,N_5010);
and U5141 (N_5141,N_5002,N_5023);
or U5142 (N_5142,N_5080,N_5030);
xor U5143 (N_5143,N_5008,N_5092);
nand U5144 (N_5144,N_5004,N_5062);
nand U5145 (N_5145,N_5059,N_5082);
nand U5146 (N_5146,N_5060,N_5014);
and U5147 (N_5147,N_5050,N_5001);
or U5148 (N_5148,N_5096,N_5005);
or U5149 (N_5149,N_5076,N_5079);
nor U5150 (N_5150,N_5048,N_5051);
and U5151 (N_5151,N_5056,N_5071);
nor U5152 (N_5152,N_5092,N_5065);
and U5153 (N_5153,N_5039,N_5045);
nand U5154 (N_5154,N_5003,N_5079);
nor U5155 (N_5155,N_5026,N_5099);
and U5156 (N_5156,N_5099,N_5028);
nand U5157 (N_5157,N_5042,N_5057);
nand U5158 (N_5158,N_5095,N_5010);
xor U5159 (N_5159,N_5090,N_5052);
and U5160 (N_5160,N_5018,N_5008);
or U5161 (N_5161,N_5083,N_5072);
xor U5162 (N_5162,N_5038,N_5003);
xor U5163 (N_5163,N_5033,N_5044);
xor U5164 (N_5164,N_5042,N_5000);
nand U5165 (N_5165,N_5040,N_5056);
or U5166 (N_5166,N_5089,N_5054);
and U5167 (N_5167,N_5095,N_5009);
and U5168 (N_5168,N_5028,N_5014);
nand U5169 (N_5169,N_5047,N_5086);
nor U5170 (N_5170,N_5082,N_5024);
nor U5171 (N_5171,N_5056,N_5004);
nand U5172 (N_5172,N_5022,N_5028);
nand U5173 (N_5173,N_5003,N_5076);
or U5174 (N_5174,N_5071,N_5025);
or U5175 (N_5175,N_5080,N_5042);
and U5176 (N_5176,N_5044,N_5097);
xor U5177 (N_5177,N_5036,N_5017);
or U5178 (N_5178,N_5015,N_5007);
or U5179 (N_5179,N_5096,N_5091);
nor U5180 (N_5180,N_5028,N_5078);
and U5181 (N_5181,N_5084,N_5073);
nor U5182 (N_5182,N_5004,N_5064);
or U5183 (N_5183,N_5058,N_5086);
nor U5184 (N_5184,N_5085,N_5064);
xor U5185 (N_5185,N_5047,N_5026);
nor U5186 (N_5186,N_5011,N_5079);
xnor U5187 (N_5187,N_5036,N_5064);
and U5188 (N_5188,N_5046,N_5076);
and U5189 (N_5189,N_5047,N_5076);
xnor U5190 (N_5190,N_5024,N_5089);
and U5191 (N_5191,N_5077,N_5072);
or U5192 (N_5192,N_5036,N_5079);
nand U5193 (N_5193,N_5021,N_5051);
or U5194 (N_5194,N_5080,N_5096);
or U5195 (N_5195,N_5046,N_5078);
nand U5196 (N_5196,N_5017,N_5032);
xnor U5197 (N_5197,N_5009,N_5064);
and U5198 (N_5198,N_5011,N_5004);
or U5199 (N_5199,N_5044,N_5086);
nor U5200 (N_5200,N_5130,N_5152);
nor U5201 (N_5201,N_5172,N_5164);
xnor U5202 (N_5202,N_5188,N_5122);
nand U5203 (N_5203,N_5192,N_5197);
and U5204 (N_5204,N_5183,N_5180);
nor U5205 (N_5205,N_5105,N_5115);
xor U5206 (N_5206,N_5133,N_5198);
and U5207 (N_5207,N_5142,N_5110);
xnor U5208 (N_5208,N_5193,N_5141);
nor U5209 (N_5209,N_5127,N_5145);
nand U5210 (N_5210,N_5167,N_5182);
or U5211 (N_5211,N_5171,N_5153);
and U5212 (N_5212,N_5104,N_5162);
and U5213 (N_5213,N_5157,N_5111);
and U5214 (N_5214,N_5113,N_5136);
nand U5215 (N_5215,N_5199,N_5149);
or U5216 (N_5216,N_5100,N_5120);
xor U5217 (N_5217,N_5139,N_5150);
and U5218 (N_5218,N_5119,N_5109);
and U5219 (N_5219,N_5160,N_5117);
or U5220 (N_5220,N_5102,N_5179);
or U5221 (N_5221,N_5163,N_5135);
or U5222 (N_5222,N_5118,N_5176);
nor U5223 (N_5223,N_5155,N_5191);
nor U5224 (N_5224,N_5126,N_5121);
nand U5225 (N_5225,N_5187,N_5156);
nor U5226 (N_5226,N_5181,N_5114);
nand U5227 (N_5227,N_5124,N_5147);
nand U5228 (N_5228,N_5194,N_5103);
and U5229 (N_5229,N_5144,N_5196);
and U5230 (N_5230,N_5148,N_5169);
xnor U5231 (N_5231,N_5108,N_5184);
and U5232 (N_5232,N_5189,N_5175);
and U5233 (N_5233,N_5174,N_5161);
and U5234 (N_5234,N_5132,N_5101);
nor U5235 (N_5235,N_5154,N_5166);
and U5236 (N_5236,N_5178,N_5106);
nor U5237 (N_5237,N_5146,N_5190);
nand U5238 (N_5238,N_5151,N_5125);
xnor U5239 (N_5239,N_5129,N_5134);
or U5240 (N_5240,N_5143,N_5112);
nand U5241 (N_5241,N_5173,N_5128);
nor U5242 (N_5242,N_5165,N_5158);
and U5243 (N_5243,N_5116,N_5168);
or U5244 (N_5244,N_5140,N_5137);
or U5245 (N_5245,N_5131,N_5107);
nand U5246 (N_5246,N_5123,N_5177);
nor U5247 (N_5247,N_5159,N_5195);
nand U5248 (N_5248,N_5185,N_5186);
or U5249 (N_5249,N_5170,N_5138);
nor U5250 (N_5250,N_5101,N_5131);
nor U5251 (N_5251,N_5107,N_5150);
xnor U5252 (N_5252,N_5142,N_5161);
or U5253 (N_5253,N_5123,N_5193);
nand U5254 (N_5254,N_5146,N_5120);
and U5255 (N_5255,N_5131,N_5185);
and U5256 (N_5256,N_5170,N_5123);
or U5257 (N_5257,N_5145,N_5199);
or U5258 (N_5258,N_5144,N_5164);
and U5259 (N_5259,N_5154,N_5144);
or U5260 (N_5260,N_5190,N_5103);
nor U5261 (N_5261,N_5151,N_5199);
nor U5262 (N_5262,N_5127,N_5121);
and U5263 (N_5263,N_5196,N_5124);
or U5264 (N_5264,N_5144,N_5178);
or U5265 (N_5265,N_5121,N_5130);
nor U5266 (N_5266,N_5191,N_5174);
nor U5267 (N_5267,N_5158,N_5186);
nor U5268 (N_5268,N_5119,N_5177);
or U5269 (N_5269,N_5161,N_5114);
xor U5270 (N_5270,N_5104,N_5173);
nor U5271 (N_5271,N_5140,N_5123);
xor U5272 (N_5272,N_5187,N_5199);
nor U5273 (N_5273,N_5165,N_5193);
and U5274 (N_5274,N_5107,N_5161);
nand U5275 (N_5275,N_5135,N_5187);
and U5276 (N_5276,N_5138,N_5129);
and U5277 (N_5277,N_5151,N_5123);
xnor U5278 (N_5278,N_5113,N_5165);
xnor U5279 (N_5279,N_5157,N_5110);
or U5280 (N_5280,N_5137,N_5109);
or U5281 (N_5281,N_5137,N_5199);
nand U5282 (N_5282,N_5110,N_5160);
nor U5283 (N_5283,N_5145,N_5118);
or U5284 (N_5284,N_5120,N_5114);
or U5285 (N_5285,N_5139,N_5172);
or U5286 (N_5286,N_5106,N_5193);
and U5287 (N_5287,N_5151,N_5113);
nor U5288 (N_5288,N_5134,N_5115);
nand U5289 (N_5289,N_5142,N_5114);
and U5290 (N_5290,N_5112,N_5156);
and U5291 (N_5291,N_5125,N_5102);
nand U5292 (N_5292,N_5158,N_5195);
nor U5293 (N_5293,N_5147,N_5141);
nor U5294 (N_5294,N_5167,N_5136);
nand U5295 (N_5295,N_5107,N_5134);
xor U5296 (N_5296,N_5107,N_5132);
and U5297 (N_5297,N_5151,N_5171);
xor U5298 (N_5298,N_5187,N_5144);
and U5299 (N_5299,N_5140,N_5198);
nand U5300 (N_5300,N_5201,N_5233);
or U5301 (N_5301,N_5208,N_5299);
nor U5302 (N_5302,N_5273,N_5282);
and U5303 (N_5303,N_5207,N_5231);
xor U5304 (N_5304,N_5206,N_5245);
nor U5305 (N_5305,N_5287,N_5286);
or U5306 (N_5306,N_5218,N_5203);
and U5307 (N_5307,N_5292,N_5276);
nor U5308 (N_5308,N_5227,N_5283);
nand U5309 (N_5309,N_5280,N_5272);
or U5310 (N_5310,N_5220,N_5252);
or U5311 (N_5311,N_5253,N_5250);
and U5312 (N_5312,N_5248,N_5297);
nor U5313 (N_5313,N_5260,N_5288);
nand U5314 (N_5314,N_5275,N_5232);
nor U5315 (N_5315,N_5298,N_5284);
nand U5316 (N_5316,N_5238,N_5263);
or U5317 (N_5317,N_5211,N_5237);
nor U5318 (N_5318,N_5224,N_5285);
and U5319 (N_5319,N_5223,N_5225);
or U5320 (N_5320,N_5230,N_5217);
nor U5321 (N_5321,N_5226,N_5246);
nand U5322 (N_5322,N_5251,N_5258);
or U5323 (N_5323,N_5210,N_5289);
and U5324 (N_5324,N_5254,N_5242);
and U5325 (N_5325,N_5271,N_5236);
nor U5326 (N_5326,N_5267,N_5257);
nor U5327 (N_5327,N_5239,N_5255);
nor U5328 (N_5328,N_5249,N_5274);
and U5329 (N_5329,N_5200,N_5202);
nand U5330 (N_5330,N_5214,N_5216);
nor U5331 (N_5331,N_5243,N_5295);
or U5332 (N_5332,N_5229,N_5265);
nand U5333 (N_5333,N_5247,N_5240);
and U5334 (N_5334,N_5256,N_5215);
nand U5335 (N_5335,N_5278,N_5266);
or U5336 (N_5336,N_5279,N_5294);
and U5337 (N_5337,N_5221,N_5228);
nand U5338 (N_5338,N_5261,N_5291);
nand U5339 (N_5339,N_5204,N_5269);
xnor U5340 (N_5340,N_5219,N_5293);
or U5341 (N_5341,N_5213,N_5205);
or U5342 (N_5342,N_5235,N_5212);
nor U5343 (N_5343,N_5244,N_5222);
nand U5344 (N_5344,N_5277,N_5264);
and U5345 (N_5345,N_5268,N_5290);
or U5346 (N_5346,N_5241,N_5296);
and U5347 (N_5347,N_5281,N_5209);
nand U5348 (N_5348,N_5259,N_5262);
nor U5349 (N_5349,N_5234,N_5270);
and U5350 (N_5350,N_5247,N_5252);
xnor U5351 (N_5351,N_5252,N_5202);
nor U5352 (N_5352,N_5293,N_5215);
nor U5353 (N_5353,N_5262,N_5235);
nor U5354 (N_5354,N_5225,N_5203);
and U5355 (N_5355,N_5232,N_5285);
nor U5356 (N_5356,N_5276,N_5267);
xor U5357 (N_5357,N_5241,N_5216);
or U5358 (N_5358,N_5253,N_5262);
nor U5359 (N_5359,N_5291,N_5278);
xor U5360 (N_5360,N_5211,N_5274);
and U5361 (N_5361,N_5293,N_5226);
and U5362 (N_5362,N_5271,N_5231);
or U5363 (N_5363,N_5202,N_5201);
xor U5364 (N_5364,N_5233,N_5242);
nor U5365 (N_5365,N_5206,N_5228);
and U5366 (N_5366,N_5210,N_5281);
nand U5367 (N_5367,N_5265,N_5236);
or U5368 (N_5368,N_5294,N_5280);
and U5369 (N_5369,N_5227,N_5292);
nor U5370 (N_5370,N_5257,N_5225);
and U5371 (N_5371,N_5237,N_5217);
nor U5372 (N_5372,N_5288,N_5290);
or U5373 (N_5373,N_5222,N_5257);
nand U5374 (N_5374,N_5290,N_5235);
nand U5375 (N_5375,N_5216,N_5279);
nor U5376 (N_5376,N_5209,N_5255);
nor U5377 (N_5377,N_5229,N_5297);
nand U5378 (N_5378,N_5200,N_5223);
and U5379 (N_5379,N_5229,N_5278);
nor U5380 (N_5380,N_5221,N_5270);
or U5381 (N_5381,N_5279,N_5204);
or U5382 (N_5382,N_5283,N_5212);
or U5383 (N_5383,N_5295,N_5290);
or U5384 (N_5384,N_5201,N_5225);
or U5385 (N_5385,N_5204,N_5222);
nand U5386 (N_5386,N_5288,N_5263);
or U5387 (N_5387,N_5200,N_5264);
xnor U5388 (N_5388,N_5248,N_5296);
nor U5389 (N_5389,N_5295,N_5251);
or U5390 (N_5390,N_5268,N_5278);
nor U5391 (N_5391,N_5203,N_5271);
and U5392 (N_5392,N_5296,N_5275);
or U5393 (N_5393,N_5223,N_5282);
and U5394 (N_5394,N_5298,N_5274);
or U5395 (N_5395,N_5273,N_5202);
xor U5396 (N_5396,N_5250,N_5275);
nand U5397 (N_5397,N_5214,N_5258);
and U5398 (N_5398,N_5230,N_5218);
nor U5399 (N_5399,N_5216,N_5260);
nor U5400 (N_5400,N_5327,N_5308);
nand U5401 (N_5401,N_5348,N_5349);
and U5402 (N_5402,N_5391,N_5351);
and U5403 (N_5403,N_5360,N_5377);
and U5404 (N_5404,N_5330,N_5352);
nor U5405 (N_5405,N_5369,N_5301);
nand U5406 (N_5406,N_5346,N_5316);
and U5407 (N_5407,N_5373,N_5309);
or U5408 (N_5408,N_5324,N_5367);
and U5409 (N_5409,N_5300,N_5393);
and U5410 (N_5410,N_5399,N_5315);
nor U5411 (N_5411,N_5338,N_5374);
or U5412 (N_5412,N_5313,N_5341);
nor U5413 (N_5413,N_5368,N_5325);
and U5414 (N_5414,N_5333,N_5382);
or U5415 (N_5415,N_5331,N_5385);
xor U5416 (N_5416,N_5305,N_5302);
and U5417 (N_5417,N_5372,N_5356);
and U5418 (N_5418,N_5342,N_5317);
nor U5419 (N_5419,N_5355,N_5370);
nor U5420 (N_5420,N_5397,N_5335);
or U5421 (N_5421,N_5311,N_5303);
nor U5422 (N_5422,N_5319,N_5321);
or U5423 (N_5423,N_5304,N_5354);
or U5424 (N_5424,N_5396,N_5379);
nor U5425 (N_5425,N_5318,N_5326);
and U5426 (N_5426,N_5376,N_5340);
nor U5427 (N_5427,N_5386,N_5362);
or U5428 (N_5428,N_5345,N_5357);
or U5429 (N_5429,N_5371,N_5389);
and U5430 (N_5430,N_5388,N_5334);
nand U5431 (N_5431,N_5358,N_5332);
nand U5432 (N_5432,N_5322,N_5329);
or U5433 (N_5433,N_5390,N_5384);
or U5434 (N_5434,N_5353,N_5380);
nand U5435 (N_5435,N_5310,N_5387);
nor U5436 (N_5436,N_5361,N_5395);
or U5437 (N_5437,N_5398,N_5314);
or U5438 (N_5438,N_5366,N_5392);
or U5439 (N_5439,N_5339,N_5320);
and U5440 (N_5440,N_5378,N_5365);
xnor U5441 (N_5441,N_5375,N_5381);
or U5442 (N_5442,N_5344,N_5336);
nand U5443 (N_5443,N_5383,N_5328);
nor U5444 (N_5444,N_5343,N_5364);
and U5445 (N_5445,N_5363,N_5337);
or U5446 (N_5446,N_5307,N_5323);
nor U5447 (N_5447,N_5347,N_5312);
or U5448 (N_5448,N_5394,N_5306);
and U5449 (N_5449,N_5359,N_5350);
nor U5450 (N_5450,N_5387,N_5344);
and U5451 (N_5451,N_5342,N_5352);
nor U5452 (N_5452,N_5323,N_5380);
nand U5453 (N_5453,N_5392,N_5390);
nor U5454 (N_5454,N_5358,N_5368);
nor U5455 (N_5455,N_5398,N_5321);
or U5456 (N_5456,N_5354,N_5344);
nor U5457 (N_5457,N_5372,N_5333);
nand U5458 (N_5458,N_5391,N_5397);
xnor U5459 (N_5459,N_5373,N_5352);
or U5460 (N_5460,N_5390,N_5369);
or U5461 (N_5461,N_5311,N_5342);
or U5462 (N_5462,N_5392,N_5300);
and U5463 (N_5463,N_5331,N_5366);
xor U5464 (N_5464,N_5355,N_5315);
nor U5465 (N_5465,N_5372,N_5353);
nand U5466 (N_5466,N_5312,N_5384);
or U5467 (N_5467,N_5334,N_5372);
and U5468 (N_5468,N_5319,N_5375);
or U5469 (N_5469,N_5391,N_5377);
nor U5470 (N_5470,N_5318,N_5310);
nor U5471 (N_5471,N_5327,N_5303);
or U5472 (N_5472,N_5362,N_5385);
and U5473 (N_5473,N_5360,N_5365);
and U5474 (N_5474,N_5316,N_5309);
or U5475 (N_5475,N_5358,N_5379);
nor U5476 (N_5476,N_5360,N_5374);
and U5477 (N_5477,N_5362,N_5356);
and U5478 (N_5478,N_5362,N_5336);
nor U5479 (N_5479,N_5322,N_5312);
nand U5480 (N_5480,N_5359,N_5387);
or U5481 (N_5481,N_5380,N_5384);
nand U5482 (N_5482,N_5385,N_5306);
nor U5483 (N_5483,N_5345,N_5379);
and U5484 (N_5484,N_5346,N_5371);
or U5485 (N_5485,N_5394,N_5305);
nand U5486 (N_5486,N_5380,N_5316);
nand U5487 (N_5487,N_5360,N_5359);
and U5488 (N_5488,N_5393,N_5380);
and U5489 (N_5489,N_5322,N_5343);
or U5490 (N_5490,N_5304,N_5331);
or U5491 (N_5491,N_5392,N_5334);
and U5492 (N_5492,N_5321,N_5301);
or U5493 (N_5493,N_5315,N_5391);
nand U5494 (N_5494,N_5379,N_5394);
nand U5495 (N_5495,N_5325,N_5362);
nor U5496 (N_5496,N_5329,N_5327);
xor U5497 (N_5497,N_5381,N_5367);
xor U5498 (N_5498,N_5370,N_5354);
and U5499 (N_5499,N_5361,N_5389);
nand U5500 (N_5500,N_5456,N_5431);
nor U5501 (N_5501,N_5423,N_5477);
or U5502 (N_5502,N_5458,N_5471);
nor U5503 (N_5503,N_5454,N_5427);
or U5504 (N_5504,N_5416,N_5468);
and U5505 (N_5505,N_5404,N_5415);
and U5506 (N_5506,N_5465,N_5474);
and U5507 (N_5507,N_5446,N_5450);
and U5508 (N_5508,N_5401,N_5435);
and U5509 (N_5509,N_5410,N_5473);
nand U5510 (N_5510,N_5455,N_5438);
or U5511 (N_5511,N_5461,N_5491);
or U5512 (N_5512,N_5443,N_5400);
nor U5513 (N_5513,N_5439,N_5428);
or U5514 (N_5514,N_5492,N_5434);
nand U5515 (N_5515,N_5463,N_5424);
and U5516 (N_5516,N_5483,N_5405);
nor U5517 (N_5517,N_5498,N_5490);
xnor U5518 (N_5518,N_5476,N_5420);
nor U5519 (N_5519,N_5496,N_5499);
nor U5520 (N_5520,N_5494,N_5480);
xnor U5521 (N_5521,N_5408,N_5460);
nor U5522 (N_5522,N_5429,N_5479);
and U5523 (N_5523,N_5421,N_5444);
nand U5524 (N_5524,N_5464,N_5478);
nor U5525 (N_5525,N_5412,N_5436);
nor U5526 (N_5526,N_5486,N_5487);
nand U5527 (N_5527,N_5488,N_5469);
or U5528 (N_5528,N_5467,N_5406);
nand U5529 (N_5529,N_5472,N_5448);
nand U5530 (N_5530,N_5413,N_5445);
nand U5531 (N_5531,N_5419,N_5481);
nand U5532 (N_5532,N_5457,N_5430);
nand U5533 (N_5533,N_5470,N_5422);
nand U5534 (N_5534,N_5449,N_5437);
and U5535 (N_5535,N_5462,N_5453);
and U5536 (N_5536,N_5484,N_5426);
or U5537 (N_5537,N_5459,N_5452);
nor U5538 (N_5538,N_5418,N_5414);
or U5539 (N_5539,N_5407,N_5495);
and U5540 (N_5540,N_5442,N_5440);
and U5541 (N_5541,N_5482,N_5417);
xor U5542 (N_5542,N_5489,N_5432);
nand U5543 (N_5543,N_5447,N_5451);
and U5544 (N_5544,N_5441,N_5466);
or U5545 (N_5545,N_5403,N_5475);
nand U5546 (N_5546,N_5485,N_5497);
and U5547 (N_5547,N_5425,N_5409);
xor U5548 (N_5548,N_5493,N_5433);
nand U5549 (N_5549,N_5411,N_5402);
and U5550 (N_5550,N_5470,N_5464);
and U5551 (N_5551,N_5438,N_5463);
nand U5552 (N_5552,N_5415,N_5446);
xnor U5553 (N_5553,N_5446,N_5400);
nor U5554 (N_5554,N_5450,N_5425);
nor U5555 (N_5555,N_5471,N_5450);
nand U5556 (N_5556,N_5456,N_5461);
and U5557 (N_5557,N_5467,N_5409);
or U5558 (N_5558,N_5429,N_5409);
xnor U5559 (N_5559,N_5491,N_5444);
nor U5560 (N_5560,N_5413,N_5477);
or U5561 (N_5561,N_5416,N_5497);
or U5562 (N_5562,N_5409,N_5438);
nor U5563 (N_5563,N_5463,N_5437);
nor U5564 (N_5564,N_5492,N_5456);
nor U5565 (N_5565,N_5452,N_5406);
and U5566 (N_5566,N_5449,N_5412);
xor U5567 (N_5567,N_5419,N_5443);
nor U5568 (N_5568,N_5487,N_5466);
and U5569 (N_5569,N_5475,N_5420);
nor U5570 (N_5570,N_5441,N_5493);
nand U5571 (N_5571,N_5448,N_5429);
or U5572 (N_5572,N_5472,N_5430);
and U5573 (N_5573,N_5487,N_5498);
nor U5574 (N_5574,N_5423,N_5435);
nand U5575 (N_5575,N_5456,N_5409);
or U5576 (N_5576,N_5487,N_5439);
and U5577 (N_5577,N_5412,N_5418);
nand U5578 (N_5578,N_5418,N_5475);
or U5579 (N_5579,N_5412,N_5429);
or U5580 (N_5580,N_5473,N_5408);
or U5581 (N_5581,N_5442,N_5449);
nor U5582 (N_5582,N_5420,N_5471);
nor U5583 (N_5583,N_5478,N_5400);
nand U5584 (N_5584,N_5429,N_5437);
and U5585 (N_5585,N_5470,N_5499);
or U5586 (N_5586,N_5466,N_5446);
or U5587 (N_5587,N_5480,N_5405);
xnor U5588 (N_5588,N_5406,N_5411);
and U5589 (N_5589,N_5400,N_5405);
xnor U5590 (N_5590,N_5422,N_5406);
nand U5591 (N_5591,N_5449,N_5455);
or U5592 (N_5592,N_5411,N_5486);
or U5593 (N_5593,N_5443,N_5454);
and U5594 (N_5594,N_5453,N_5455);
nand U5595 (N_5595,N_5497,N_5434);
nor U5596 (N_5596,N_5431,N_5443);
nor U5597 (N_5597,N_5490,N_5464);
nor U5598 (N_5598,N_5461,N_5478);
and U5599 (N_5599,N_5499,N_5498);
nor U5600 (N_5600,N_5595,N_5581);
or U5601 (N_5601,N_5530,N_5582);
nor U5602 (N_5602,N_5571,N_5562);
and U5603 (N_5603,N_5587,N_5500);
xnor U5604 (N_5604,N_5533,N_5560);
nor U5605 (N_5605,N_5550,N_5516);
and U5606 (N_5606,N_5537,N_5545);
nor U5607 (N_5607,N_5589,N_5548);
and U5608 (N_5608,N_5578,N_5523);
and U5609 (N_5609,N_5549,N_5544);
or U5610 (N_5610,N_5592,N_5577);
or U5611 (N_5611,N_5555,N_5520);
and U5612 (N_5612,N_5506,N_5569);
nor U5613 (N_5613,N_5513,N_5501);
or U5614 (N_5614,N_5558,N_5510);
and U5615 (N_5615,N_5524,N_5594);
nor U5616 (N_5616,N_5504,N_5542);
nand U5617 (N_5617,N_5538,N_5591);
or U5618 (N_5618,N_5547,N_5575);
nor U5619 (N_5619,N_5597,N_5528);
nor U5620 (N_5620,N_5599,N_5598);
xnor U5621 (N_5621,N_5509,N_5573);
and U5622 (N_5622,N_5563,N_5565);
nand U5623 (N_5623,N_5588,N_5572);
xor U5624 (N_5624,N_5559,N_5593);
or U5625 (N_5625,N_5505,N_5564);
or U5626 (N_5626,N_5580,N_5526);
nor U5627 (N_5627,N_5532,N_5566);
or U5628 (N_5628,N_5574,N_5517);
and U5629 (N_5629,N_5596,N_5521);
nor U5630 (N_5630,N_5515,N_5568);
nand U5631 (N_5631,N_5585,N_5514);
or U5632 (N_5632,N_5512,N_5586);
or U5633 (N_5633,N_5519,N_5546);
nor U5634 (N_5634,N_5552,N_5556);
nor U5635 (N_5635,N_5557,N_5525);
nand U5636 (N_5636,N_5534,N_5527);
nand U5637 (N_5637,N_5579,N_5554);
or U5638 (N_5638,N_5503,N_5561);
and U5639 (N_5639,N_5584,N_5570);
nor U5640 (N_5640,N_5536,N_5541);
nor U5641 (N_5641,N_5576,N_5590);
nor U5642 (N_5642,N_5518,N_5553);
and U5643 (N_5643,N_5567,N_5522);
and U5644 (N_5644,N_5529,N_5535);
nand U5645 (N_5645,N_5583,N_5508);
and U5646 (N_5646,N_5507,N_5539);
xor U5647 (N_5647,N_5531,N_5551);
nand U5648 (N_5648,N_5502,N_5540);
and U5649 (N_5649,N_5543,N_5511);
xnor U5650 (N_5650,N_5503,N_5559);
nand U5651 (N_5651,N_5566,N_5520);
and U5652 (N_5652,N_5564,N_5587);
and U5653 (N_5653,N_5546,N_5595);
nand U5654 (N_5654,N_5500,N_5595);
nand U5655 (N_5655,N_5554,N_5514);
nand U5656 (N_5656,N_5588,N_5599);
nand U5657 (N_5657,N_5567,N_5525);
xor U5658 (N_5658,N_5500,N_5519);
and U5659 (N_5659,N_5562,N_5540);
or U5660 (N_5660,N_5546,N_5540);
or U5661 (N_5661,N_5501,N_5579);
nand U5662 (N_5662,N_5574,N_5594);
or U5663 (N_5663,N_5502,N_5533);
and U5664 (N_5664,N_5505,N_5563);
and U5665 (N_5665,N_5571,N_5578);
nor U5666 (N_5666,N_5588,N_5529);
xnor U5667 (N_5667,N_5529,N_5539);
and U5668 (N_5668,N_5544,N_5533);
nand U5669 (N_5669,N_5589,N_5557);
nand U5670 (N_5670,N_5571,N_5508);
or U5671 (N_5671,N_5527,N_5506);
nor U5672 (N_5672,N_5536,N_5565);
and U5673 (N_5673,N_5589,N_5556);
and U5674 (N_5674,N_5562,N_5579);
nand U5675 (N_5675,N_5516,N_5509);
or U5676 (N_5676,N_5575,N_5536);
and U5677 (N_5677,N_5581,N_5549);
nor U5678 (N_5678,N_5547,N_5574);
xor U5679 (N_5679,N_5512,N_5528);
or U5680 (N_5680,N_5583,N_5567);
xor U5681 (N_5681,N_5530,N_5567);
nor U5682 (N_5682,N_5573,N_5523);
nor U5683 (N_5683,N_5566,N_5585);
nand U5684 (N_5684,N_5514,N_5568);
and U5685 (N_5685,N_5594,N_5529);
nand U5686 (N_5686,N_5588,N_5521);
and U5687 (N_5687,N_5589,N_5506);
and U5688 (N_5688,N_5572,N_5536);
and U5689 (N_5689,N_5526,N_5555);
or U5690 (N_5690,N_5524,N_5523);
nor U5691 (N_5691,N_5562,N_5519);
nand U5692 (N_5692,N_5560,N_5519);
nand U5693 (N_5693,N_5512,N_5592);
nand U5694 (N_5694,N_5567,N_5518);
and U5695 (N_5695,N_5568,N_5545);
nand U5696 (N_5696,N_5598,N_5585);
and U5697 (N_5697,N_5502,N_5585);
or U5698 (N_5698,N_5508,N_5599);
xor U5699 (N_5699,N_5535,N_5549);
or U5700 (N_5700,N_5610,N_5644);
or U5701 (N_5701,N_5645,N_5665);
or U5702 (N_5702,N_5615,N_5603);
nor U5703 (N_5703,N_5678,N_5676);
nor U5704 (N_5704,N_5607,N_5663);
or U5705 (N_5705,N_5680,N_5621);
nor U5706 (N_5706,N_5655,N_5652);
nor U5707 (N_5707,N_5662,N_5668);
and U5708 (N_5708,N_5618,N_5630);
xor U5709 (N_5709,N_5691,N_5654);
nor U5710 (N_5710,N_5642,N_5604);
nand U5711 (N_5711,N_5685,N_5656);
nor U5712 (N_5712,N_5650,N_5627);
nand U5713 (N_5713,N_5692,N_5602);
nand U5714 (N_5714,N_5631,N_5647);
or U5715 (N_5715,N_5622,N_5646);
nand U5716 (N_5716,N_5689,N_5682);
or U5717 (N_5717,N_5675,N_5632);
and U5718 (N_5718,N_5601,N_5612);
nand U5719 (N_5719,N_5697,N_5693);
or U5720 (N_5720,N_5683,N_5684);
nand U5721 (N_5721,N_5611,N_5677);
and U5722 (N_5722,N_5616,N_5628);
and U5723 (N_5723,N_5688,N_5671);
and U5724 (N_5724,N_5657,N_5613);
nand U5725 (N_5725,N_5661,N_5670);
and U5726 (N_5726,N_5651,N_5643);
nor U5727 (N_5727,N_5629,N_5617);
nand U5728 (N_5728,N_5687,N_5669);
xor U5729 (N_5729,N_5625,N_5698);
nor U5730 (N_5730,N_5659,N_5624);
nor U5731 (N_5731,N_5620,N_5696);
xor U5732 (N_5732,N_5639,N_5653);
or U5733 (N_5733,N_5633,N_5672);
and U5734 (N_5734,N_5667,N_5623);
or U5735 (N_5735,N_5626,N_5679);
nand U5736 (N_5736,N_5673,N_5666);
or U5737 (N_5737,N_5686,N_5606);
nor U5738 (N_5738,N_5600,N_5649);
nand U5739 (N_5739,N_5614,N_5681);
or U5740 (N_5740,N_5635,N_5648);
nor U5741 (N_5741,N_5658,N_5608);
nand U5742 (N_5742,N_5699,N_5674);
and U5743 (N_5743,N_5637,N_5641);
or U5744 (N_5744,N_5695,N_5664);
nor U5745 (N_5745,N_5636,N_5638);
nand U5746 (N_5746,N_5634,N_5640);
nand U5747 (N_5747,N_5694,N_5605);
xnor U5748 (N_5748,N_5660,N_5690);
xnor U5749 (N_5749,N_5619,N_5609);
nand U5750 (N_5750,N_5627,N_5616);
nor U5751 (N_5751,N_5606,N_5691);
nand U5752 (N_5752,N_5683,N_5648);
nand U5753 (N_5753,N_5699,N_5601);
and U5754 (N_5754,N_5614,N_5628);
nand U5755 (N_5755,N_5688,N_5689);
nand U5756 (N_5756,N_5682,N_5639);
nand U5757 (N_5757,N_5637,N_5666);
nor U5758 (N_5758,N_5699,N_5684);
nand U5759 (N_5759,N_5603,N_5698);
nor U5760 (N_5760,N_5619,N_5664);
or U5761 (N_5761,N_5648,N_5629);
or U5762 (N_5762,N_5601,N_5678);
or U5763 (N_5763,N_5609,N_5688);
nand U5764 (N_5764,N_5675,N_5611);
or U5765 (N_5765,N_5679,N_5663);
or U5766 (N_5766,N_5695,N_5613);
nor U5767 (N_5767,N_5690,N_5649);
or U5768 (N_5768,N_5661,N_5608);
nor U5769 (N_5769,N_5637,N_5603);
nor U5770 (N_5770,N_5675,N_5654);
or U5771 (N_5771,N_5694,N_5678);
or U5772 (N_5772,N_5699,N_5663);
nor U5773 (N_5773,N_5605,N_5602);
or U5774 (N_5774,N_5601,N_5640);
or U5775 (N_5775,N_5618,N_5693);
nor U5776 (N_5776,N_5663,N_5698);
xnor U5777 (N_5777,N_5644,N_5614);
and U5778 (N_5778,N_5645,N_5671);
and U5779 (N_5779,N_5686,N_5619);
xor U5780 (N_5780,N_5613,N_5615);
or U5781 (N_5781,N_5657,N_5681);
xnor U5782 (N_5782,N_5698,N_5635);
nor U5783 (N_5783,N_5612,N_5640);
or U5784 (N_5784,N_5629,N_5667);
xnor U5785 (N_5785,N_5671,N_5628);
nand U5786 (N_5786,N_5688,N_5683);
nand U5787 (N_5787,N_5639,N_5618);
nand U5788 (N_5788,N_5666,N_5694);
and U5789 (N_5789,N_5659,N_5655);
or U5790 (N_5790,N_5642,N_5677);
nor U5791 (N_5791,N_5687,N_5600);
and U5792 (N_5792,N_5609,N_5672);
nand U5793 (N_5793,N_5618,N_5628);
and U5794 (N_5794,N_5615,N_5605);
nand U5795 (N_5795,N_5601,N_5639);
and U5796 (N_5796,N_5628,N_5610);
and U5797 (N_5797,N_5635,N_5657);
nand U5798 (N_5798,N_5673,N_5662);
and U5799 (N_5799,N_5616,N_5600);
nand U5800 (N_5800,N_5770,N_5704);
nor U5801 (N_5801,N_5783,N_5715);
and U5802 (N_5802,N_5757,N_5764);
nor U5803 (N_5803,N_5740,N_5797);
xor U5804 (N_5804,N_5779,N_5734);
nor U5805 (N_5805,N_5778,N_5781);
nor U5806 (N_5806,N_5726,N_5753);
nand U5807 (N_5807,N_5744,N_5701);
or U5808 (N_5808,N_5713,N_5794);
nand U5809 (N_5809,N_5774,N_5745);
xor U5810 (N_5810,N_5709,N_5760);
nand U5811 (N_5811,N_5790,N_5748);
or U5812 (N_5812,N_5749,N_5799);
nor U5813 (N_5813,N_5763,N_5756);
nand U5814 (N_5814,N_5736,N_5703);
or U5815 (N_5815,N_5705,N_5751);
nor U5816 (N_5816,N_5771,N_5729);
nand U5817 (N_5817,N_5784,N_5766);
nor U5818 (N_5818,N_5732,N_5711);
or U5819 (N_5819,N_5792,N_5742);
nand U5820 (N_5820,N_5777,N_5727);
and U5821 (N_5821,N_5718,N_5793);
and U5822 (N_5822,N_5752,N_5707);
xnor U5823 (N_5823,N_5785,N_5786);
and U5824 (N_5824,N_5787,N_5731);
nand U5825 (N_5825,N_5758,N_5720);
and U5826 (N_5826,N_5712,N_5741);
nand U5827 (N_5827,N_5733,N_5722);
nand U5828 (N_5828,N_5743,N_5719);
nor U5829 (N_5829,N_5798,N_5788);
nand U5830 (N_5830,N_5772,N_5702);
nand U5831 (N_5831,N_5761,N_5700);
and U5832 (N_5832,N_5780,N_5795);
and U5833 (N_5833,N_5754,N_5796);
nand U5834 (N_5834,N_5730,N_5747);
nand U5835 (N_5835,N_5735,N_5737);
nor U5836 (N_5836,N_5773,N_5725);
nand U5837 (N_5837,N_5723,N_5762);
or U5838 (N_5838,N_5759,N_5724);
or U5839 (N_5839,N_5768,N_5755);
nor U5840 (N_5840,N_5765,N_5750);
xnor U5841 (N_5841,N_5716,N_5738);
nor U5842 (N_5842,N_5769,N_5767);
and U5843 (N_5843,N_5728,N_5782);
and U5844 (N_5844,N_5708,N_5714);
or U5845 (N_5845,N_5721,N_5710);
and U5846 (N_5846,N_5775,N_5746);
nor U5847 (N_5847,N_5776,N_5789);
nand U5848 (N_5848,N_5706,N_5791);
nor U5849 (N_5849,N_5717,N_5739);
xor U5850 (N_5850,N_5748,N_5734);
nand U5851 (N_5851,N_5756,N_5728);
and U5852 (N_5852,N_5787,N_5767);
nor U5853 (N_5853,N_5796,N_5726);
or U5854 (N_5854,N_5749,N_5766);
nand U5855 (N_5855,N_5756,N_5708);
or U5856 (N_5856,N_5745,N_5735);
or U5857 (N_5857,N_5729,N_5798);
nor U5858 (N_5858,N_5799,N_5797);
and U5859 (N_5859,N_5707,N_5700);
or U5860 (N_5860,N_5703,N_5758);
or U5861 (N_5861,N_5735,N_5780);
nand U5862 (N_5862,N_5770,N_5796);
nor U5863 (N_5863,N_5727,N_5730);
nand U5864 (N_5864,N_5751,N_5734);
nand U5865 (N_5865,N_5725,N_5753);
or U5866 (N_5866,N_5769,N_5706);
nand U5867 (N_5867,N_5783,N_5781);
nand U5868 (N_5868,N_5775,N_5774);
nand U5869 (N_5869,N_5720,N_5724);
and U5870 (N_5870,N_5779,N_5789);
and U5871 (N_5871,N_5765,N_5705);
or U5872 (N_5872,N_5709,N_5718);
nor U5873 (N_5873,N_5797,N_5775);
nand U5874 (N_5874,N_5700,N_5734);
and U5875 (N_5875,N_5703,N_5754);
xnor U5876 (N_5876,N_5779,N_5764);
nand U5877 (N_5877,N_5716,N_5714);
or U5878 (N_5878,N_5743,N_5704);
nor U5879 (N_5879,N_5757,N_5742);
nor U5880 (N_5880,N_5712,N_5747);
and U5881 (N_5881,N_5766,N_5731);
or U5882 (N_5882,N_5736,N_5797);
or U5883 (N_5883,N_5776,N_5796);
nand U5884 (N_5884,N_5718,N_5720);
nand U5885 (N_5885,N_5715,N_5784);
and U5886 (N_5886,N_5712,N_5795);
nand U5887 (N_5887,N_5776,N_5729);
nor U5888 (N_5888,N_5791,N_5782);
nand U5889 (N_5889,N_5758,N_5786);
or U5890 (N_5890,N_5750,N_5746);
nor U5891 (N_5891,N_5728,N_5730);
or U5892 (N_5892,N_5763,N_5751);
and U5893 (N_5893,N_5759,N_5739);
nor U5894 (N_5894,N_5776,N_5739);
nand U5895 (N_5895,N_5736,N_5743);
nand U5896 (N_5896,N_5790,N_5755);
and U5897 (N_5897,N_5703,N_5767);
nor U5898 (N_5898,N_5792,N_5746);
or U5899 (N_5899,N_5751,N_5744);
and U5900 (N_5900,N_5853,N_5897);
nor U5901 (N_5901,N_5862,N_5895);
nor U5902 (N_5902,N_5811,N_5830);
and U5903 (N_5903,N_5803,N_5832);
nand U5904 (N_5904,N_5839,N_5849);
or U5905 (N_5905,N_5842,N_5857);
and U5906 (N_5906,N_5879,N_5899);
nand U5907 (N_5907,N_5872,N_5861);
nor U5908 (N_5908,N_5801,N_5874);
or U5909 (N_5909,N_5813,N_5898);
and U5910 (N_5910,N_5847,N_5825);
nor U5911 (N_5911,N_5894,N_5806);
and U5912 (N_5912,N_5829,N_5884);
or U5913 (N_5913,N_5869,N_5812);
nor U5914 (N_5914,N_5864,N_5877);
nand U5915 (N_5915,N_5802,N_5840);
nand U5916 (N_5916,N_5836,N_5881);
or U5917 (N_5917,N_5875,N_5833);
nor U5918 (N_5918,N_5854,N_5863);
or U5919 (N_5919,N_5824,N_5819);
nand U5920 (N_5920,N_5868,N_5883);
nor U5921 (N_5921,N_5826,N_5835);
nand U5922 (N_5922,N_5844,N_5858);
nand U5923 (N_5923,N_5821,N_5887);
or U5924 (N_5924,N_5804,N_5817);
and U5925 (N_5925,N_5888,N_5891);
and U5926 (N_5926,N_5831,N_5866);
or U5927 (N_5927,N_5892,N_5838);
nand U5928 (N_5928,N_5889,N_5896);
nor U5929 (N_5929,N_5827,N_5846);
xnor U5930 (N_5930,N_5870,N_5890);
nor U5931 (N_5931,N_5823,N_5865);
and U5932 (N_5932,N_5818,N_5851);
or U5933 (N_5933,N_5809,N_5814);
xnor U5934 (N_5934,N_5860,N_5880);
and U5935 (N_5935,N_5878,N_5855);
and U5936 (N_5936,N_5820,N_5882);
or U5937 (N_5937,N_5815,N_5841);
xor U5938 (N_5938,N_5859,N_5850);
nor U5939 (N_5939,N_5871,N_5834);
or U5940 (N_5940,N_5805,N_5816);
nor U5941 (N_5941,N_5873,N_5886);
nor U5942 (N_5942,N_5828,N_5843);
nor U5943 (N_5943,N_5810,N_5893);
and U5944 (N_5944,N_5800,N_5837);
nor U5945 (N_5945,N_5807,N_5845);
nand U5946 (N_5946,N_5822,N_5808);
nand U5947 (N_5947,N_5856,N_5867);
nor U5948 (N_5948,N_5848,N_5885);
nand U5949 (N_5949,N_5876,N_5852);
nor U5950 (N_5950,N_5843,N_5845);
nor U5951 (N_5951,N_5801,N_5876);
nand U5952 (N_5952,N_5835,N_5804);
nor U5953 (N_5953,N_5862,N_5868);
nand U5954 (N_5954,N_5806,N_5883);
nand U5955 (N_5955,N_5885,N_5894);
nand U5956 (N_5956,N_5876,N_5808);
or U5957 (N_5957,N_5836,N_5824);
nor U5958 (N_5958,N_5848,N_5825);
nand U5959 (N_5959,N_5843,N_5818);
nand U5960 (N_5960,N_5873,N_5861);
xnor U5961 (N_5961,N_5805,N_5869);
xnor U5962 (N_5962,N_5851,N_5855);
xnor U5963 (N_5963,N_5832,N_5885);
nand U5964 (N_5964,N_5802,N_5847);
or U5965 (N_5965,N_5868,N_5872);
nor U5966 (N_5966,N_5834,N_5853);
nor U5967 (N_5967,N_5890,N_5894);
nand U5968 (N_5968,N_5844,N_5872);
or U5969 (N_5969,N_5812,N_5809);
nor U5970 (N_5970,N_5832,N_5880);
or U5971 (N_5971,N_5840,N_5819);
or U5972 (N_5972,N_5857,N_5873);
nor U5973 (N_5973,N_5821,N_5837);
nor U5974 (N_5974,N_5872,N_5883);
nor U5975 (N_5975,N_5838,N_5879);
xor U5976 (N_5976,N_5846,N_5854);
nand U5977 (N_5977,N_5818,N_5844);
nor U5978 (N_5978,N_5876,N_5819);
and U5979 (N_5979,N_5890,N_5848);
or U5980 (N_5980,N_5818,N_5817);
nor U5981 (N_5981,N_5830,N_5886);
nor U5982 (N_5982,N_5822,N_5804);
or U5983 (N_5983,N_5864,N_5815);
nor U5984 (N_5984,N_5823,N_5864);
nor U5985 (N_5985,N_5820,N_5894);
nand U5986 (N_5986,N_5868,N_5825);
or U5987 (N_5987,N_5840,N_5871);
or U5988 (N_5988,N_5851,N_5826);
or U5989 (N_5989,N_5848,N_5827);
or U5990 (N_5990,N_5820,N_5886);
and U5991 (N_5991,N_5851,N_5811);
nor U5992 (N_5992,N_5837,N_5827);
xnor U5993 (N_5993,N_5845,N_5839);
xor U5994 (N_5994,N_5847,N_5868);
nand U5995 (N_5995,N_5806,N_5820);
nand U5996 (N_5996,N_5875,N_5869);
nor U5997 (N_5997,N_5867,N_5815);
xor U5998 (N_5998,N_5886,N_5834);
nand U5999 (N_5999,N_5846,N_5835);
nand U6000 (N_6000,N_5993,N_5983);
and U6001 (N_6001,N_5978,N_5962);
nand U6002 (N_6002,N_5988,N_5965);
or U6003 (N_6003,N_5959,N_5975);
or U6004 (N_6004,N_5932,N_5987);
and U6005 (N_6005,N_5955,N_5985);
nor U6006 (N_6006,N_5951,N_5940);
nor U6007 (N_6007,N_5925,N_5904);
nor U6008 (N_6008,N_5977,N_5930);
nand U6009 (N_6009,N_5922,N_5907);
and U6010 (N_6010,N_5918,N_5969);
nand U6011 (N_6011,N_5994,N_5928);
nor U6012 (N_6012,N_5924,N_5926);
nand U6013 (N_6013,N_5917,N_5900);
or U6014 (N_6014,N_5982,N_5938);
and U6015 (N_6015,N_5948,N_5903);
and U6016 (N_6016,N_5967,N_5943);
nor U6017 (N_6017,N_5915,N_5960);
nor U6018 (N_6018,N_5992,N_5990);
or U6019 (N_6019,N_5952,N_5968);
and U6020 (N_6020,N_5939,N_5923);
nand U6021 (N_6021,N_5979,N_5991);
nor U6022 (N_6022,N_5950,N_5913);
and U6023 (N_6023,N_5998,N_5901);
nor U6024 (N_6024,N_5947,N_5970);
or U6025 (N_6025,N_5956,N_5966);
or U6026 (N_6026,N_5984,N_5909);
or U6027 (N_6027,N_5937,N_5963);
or U6028 (N_6028,N_5905,N_5972);
nor U6029 (N_6029,N_5954,N_5980);
nand U6030 (N_6030,N_5931,N_5961);
and U6031 (N_6031,N_5958,N_5941);
nor U6032 (N_6032,N_5914,N_5976);
nand U6033 (N_6033,N_5912,N_5908);
or U6034 (N_6034,N_5910,N_5919);
nor U6035 (N_6035,N_5953,N_5945);
or U6036 (N_6036,N_5921,N_5986);
nor U6037 (N_6037,N_5906,N_5973);
or U6038 (N_6038,N_5942,N_5949);
and U6039 (N_6039,N_5927,N_5902);
nor U6040 (N_6040,N_5989,N_5934);
and U6041 (N_6041,N_5974,N_5929);
or U6042 (N_6042,N_5933,N_5936);
nand U6043 (N_6043,N_5957,N_5935);
nor U6044 (N_6044,N_5964,N_5995);
or U6045 (N_6045,N_5911,N_5997);
xnor U6046 (N_6046,N_5944,N_5916);
nand U6047 (N_6047,N_5920,N_5999);
nand U6048 (N_6048,N_5981,N_5971);
xnor U6049 (N_6049,N_5996,N_5946);
nand U6050 (N_6050,N_5997,N_5982);
and U6051 (N_6051,N_5908,N_5952);
or U6052 (N_6052,N_5956,N_5900);
and U6053 (N_6053,N_5901,N_5905);
nor U6054 (N_6054,N_5975,N_5936);
and U6055 (N_6055,N_5999,N_5963);
and U6056 (N_6056,N_5933,N_5970);
and U6057 (N_6057,N_5973,N_5949);
and U6058 (N_6058,N_5985,N_5979);
nand U6059 (N_6059,N_5977,N_5968);
nand U6060 (N_6060,N_5965,N_5967);
and U6061 (N_6061,N_5913,N_5977);
nor U6062 (N_6062,N_5964,N_5935);
xnor U6063 (N_6063,N_5955,N_5904);
xnor U6064 (N_6064,N_5936,N_5946);
nand U6065 (N_6065,N_5938,N_5960);
and U6066 (N_6066,N_5934,N_5930);
nor U6067 (N_6067,N_5952,N_5935);
and U6068 (N_6068,N_5935,N_5977);
nand U6069 (N_6069,N_5919,N_5994);
nand U6070 (N_6070,N_5919,N_5908);
nor U6071 (N_6071,N_5921,N_5973);
or U6072 (N_6072,N_5971,N_5937);
nor U6073 (N_6073,N_5986,N_5976);
and U6074 (N_6074,N_5900,N_5978);
or U6075 (N_6075,N_5994,N_5988);
nand U6076 (N_6076,N_5940,N_5907);
or U6077 (N_6077,N_5901,N_5939);
nor U6078 (N_6078,N_5924,N_5953);
and U6079 (N_6079,N_5982,N_5907);
and U6080 (N_6080,N_5910,N_5941);
and U6081 (N_6081,N_5917,N_5919);
nand U6082 (N_6082,N_5956,N_5995);
or U6083 (N_6083,N_5962,N_5970);
and U6084 (N_6084,N_5931,N_5938);
or U6085 (N_6085,N_5989,N_5992);
nor U6086 (N_6086,N_5938,N_5972);
nor U6087 (N_6087,N_5936,N_5965);
nand U6088 (N_6088,N_5913,N_5995);
or U6089 (N_6089,N_5923,N_5904);
and U6090 (N_6090,N_5904,N_5940);
or U6091 (N_6091,N_5976,N_5921);
nor U6092 (N_6092,N_5969,N_5900);
nand U6093 (N_6093,N_5920,N_5942);
xnor U6094 (N_6094,N_5963,N_5943);
and U6095 (N_6095,N_5945,N_5986);
nor U6096 (N_6096,N_5944,N_5990);
nand U6097 (N_6097,N_5975,N_5958);
or U6098 (N_6098,N_5927,N_5960);
and U6099 (N_6099,N_5989,N_5940);
and U6100 (N_6100,N_6065,N_6049);
xor U6101 (N_6101,N_6005,N_6082);
nand U6102 (N_6102,N_6004,N_6087);
nand U6103 (N_6103,N_6092,N_6026);
or U6104 (N_6104,N_6001,N_6089);
nand U6105 (N_6105,N_6090,N_6095);
xnor U6106 (N_6106,N_6024,N_6050);
and U6107 (N_6107,N_6073,N_6056);
nor U6108 (N_6108,N_6091,N_6014);
or U6109 (N_6109,N_6036,N_6039);
and U6110 (N_6110,N_6054,N_6068);
nand U6111 (N_6111,N_6029,N_6031);
and U6112 (N_6112,N_6063,N_6017);
or U6113 (N_6113,N_6083,N_6012);
and U6114 (N_6114,N_6081,N_6066);
nor U6115 (N_6115,N_6030,N_6098);
xor U6116 (N_6116,N_6022,N_6040);
nor U6117 (N_6117,N_6008,N_6042);
and U6118 (N_6118,N_6055,N_6086);
or U6119 (N_6119,N_6067,N_6070);
and U6120 (N_6120,N_6009,N_6011);
nor U6121 (N_6121,N_6080,N_6006);
nand U6122 (N_6122,N_6019,N_6069);
nand U6123 (N_6123,N_6043,N_6044);
nand U6124 (N_6124,N_6046,N_6077);
and U6125 (N_6125,N_6059,N_6058);
or U6126 (N_6126,N_6051,N_6076);
nor U6127 (N_6127,N_6045,N_6041);
and U6128 (N_6128,N_6015,N_6037);
nand U6129 (N_6129,N_6003,N_6057);
and U6130 (N_6130,N_6062,N_6075);
nor U6131 (N_6131,N_6016,N_6020);
nor U6132 (N_6132,N_6033,N_6074);
or U6133 (N_6133,N_6052,N_6034);
and U6134 (N_6134,N_6002,N_6023);
or U6135 (N_6135,N_6053,N_6084);
and U6136 (N_6136,N_6097,N_6013);
nor U6137 (N_6137,N_6071,N_6010);
and U6138 (N_6138,N_6099,N_6027);
and U6139 (N_6139,N_6032,N_6093);
or U6140 (N_6140,N_6038,N_6021);
nand U6141 (N_6141,N_6018,N_6025);
xor U6142 (N_6142,N_6048,N_6079);
and U6143 (N_6143,N_6072,N_6028);
or U6144 (N_6144,N_6061,N_6064);
and U6145 (N_6145,N_6094,N_6007);
nand U6146 (N_6146,N_6096,N_6078);
xnor U6147 (N_6147,N_6088,N_6060);
nand U6148 (N_6148,N_6047,N_6035);
nor U6149 (N_6149,N_6000,N_6085);
and U6150 (N_6150,N_6031,N_6094);
and U6151 (N_6151,N_6063,N_6051);
and U6152 (N_6152,N_6057,N_6015);
nor U6153 (N_6153,N_6050,N_6051);
nor U6154 (N_6154,N_6057,N_6096);
nand U6155 (N_6155,N_6098,N_6062);
xnor U6156 (N_6156,N_6089,N_6009);
nor U6157 (N_6157,N_6020,N_6072);
nor U6158 (N_6158,N_6054,N_6029);
or U6159 (N_6159,N_6024,N_6089);
nor U6160 (N_6160,N_6086,N_6031);
nor U6161 (N_6161,N_6014,N_6066);
or U6162 (N_6162,N_6062,N_6021);
xor U6163 (N_6163,N_6099,N_6046);
or U6164 (N_6164,N_6025,N_6023);
nor U6165 (N_6165,N_6092,N_6066);
nand U6166 (N_6166,N_6045,N_6024);
nor U6167 (N_6167,N_6063,N_6078);
or U6168 (N_6168,N_6016,N_6035);
nand U6169 (N_6169,N_6029,N_6021);
nand U6170 (N_6170,N_6085,N_6028);
xnor U6171 (N_6171,N_6099,N_6030);
or U6172 (N_6172,N_6079,N_6053);
and U6173 (N_6173,N_6011,N_6029);
xor U6174 (N_6174,N_6040,N_6019);
and U6175 (N_6175,N_6046,N_6078);
or U6176 (N_6176,N_6079,N_6003);
nor U6177 (N_6177,N_6041,N_6030);
or U6178 (N_6178,N_6001,N_6004);
and U6179 (N_6179,N_6035,N_6009);
xnor U6180 (N_6180,N_6017,N_6005);
xnor U6181 (N_6181,N_6003,N_6032);
xnor U6182 (N_6182,N_6082,N_6086);
nand U6183 (N_6183,N_6082,N_6017);
and U6184 (N_6184,N_6087,N_6091);
nand U6185 (N_6185,N_6045,N_6092);
or U6186 (N_6186,N_6071,N_6034);
or U6187 (N_6187,N_6000,N_6065);
or U6188 (N_6188,N_6002,N_6070);
and U6189 (N_6189,N_6048,N_6056);
nand U6190 (N_6190,N_6025,N_6075);
nand U6191 (N_6191,N_6018,N_6000);
nor U6192 (N_6192,N_6091,N_6017);
or U6193 (N_6193,N_6004,N_6035);
or U6194 (N_6194,N_6078,N_6009);
or U6195 (N_6195,N_6017,N_6068);
and U6196 (N_6196,N_6012,N_6088);
nor U6197 (N_6197,N_6012,N_6090);
and U6198 (N_6198,N_6054,N_6022);
nand U6199 (N_6199,N_6006,N_6037);
and U6200 (N_6200,N_6120,N_6169);
xor U6201 (N_6201,N_6103,N_6195);
xor U6202 (N_6202,N_6166,N_6144);
and U6203 (N_6203,N_6127,N_6184);
or U6204 (N_6204,N_6198,N_6113);
nor U6205 (N_6205,N_6128,N_6160);
nor U6206 (N_6206,N_6119,N_6190);
and U6207 (N_6207,N_6162,N_6147);
nor U6208 (N_6208,N_6180,N_6176);
nor U6209 (N_6209,N_6197,N_6131);
and U6210 (N_6210,N_6199,N_6112);
and U6211 (N_6211,N_6177,N_6109);
nand U6212 (N_6212,N_6181,N_6172);
and U6213 (N_6213,N_6114,N_6105);
and U6214 (N_6214,N_6121,N_6111);
nand U6215 (N_6215,N_6106,N_6187);
nor U6216 (N_6216,N_6107,N_6149);
or U6217 (N_6217,N_6173,N_6179);
xor U6218 (N_6218,N_6185,N_6145);
xor U6219 (N_6219,N_6125,N_6135);
and U6220 (N_6220,N_6182,N_6159);
nand U6221 (N_6221,N_6102,N_6118);
xnor U6222 (N_6222,N_6164,N_6194);
or U6223 (N_6223,N_6139,N_6117);
and U6224 (N_6224,N_6189,N_6115);
and U6225 (N_6225,N_6192,N_6154);
nand U6226 (N_6226,N_6170,N_6146);
nand U6227 (N_6227,N_6126,N_6168);
and U6228 (N_6228,N_6140,N_6150);
nor U6229 (N_6229,N_6110,N_6123);
nand U6230 (N_6230,N_6153,N_6174);
nor U6231 (N_6231,N_6171,N_6100);
and U6232 (N_6232,N_6186,N_6148);
and U6233 (N_6233,N_6183,N_6116);
nor U6234 (N_6234,N_6167,N_6191);
or U6235 (N_6235,N_6155,N_6132);
xor U6236 (N_6236,N_6196,N_6161);
and U6237 (N_6237,N_6143,N_6129);
xnor U6238 (N_6238,N_6141,N_6157);
or U6239 (N_6239,N_6158,N_6175);
nor U6240 (N_6240,N_6101,N_6137);
nand U6241 (N_6241,N_6178,N_6124);
or U6242 (N_6242,N_6165,N_6142);
and U6243 (N_6243,N_6134,N_6188);
and U6244 (N_6244,N_6163,N_6152);
or U6245 (N_6245,N_6108,N_6151);
nor U6246 (N_6246,N_6104,N_6136);
and U6247 (N_6247,N_6133,N_6193);
nor U6248 (N_6248,N_6122,N_6156);
nor U6249 (N_6249,N_6130,N_6138);
xor U6250 (N_6250,N_6178,N_6164);
nand U6251 (N_6251,N_6172,N_6155);
nor U6252 (N_6252,N_6197,N_6185);
xor U6253 (N_6253,N_6189,N_6102);
xnor U6254 (N_6254,N_6162,N_6131);
and U6255 (N_6255,N_6117,N_6111);
or U6256 (N_6256,N_6169,N_6131);
nand U6257 (N_6257,N_6151,N_6171);
and U6258 (N_6258,N_6143,N_6118);
xnor U6259 (N_6259,N_6146,N_6113);
or U6260 (N_6260,N_6186,N_6138);
or U6261 (N_6261,N_6106,N_6126);
nand U6262 (N_6262,N_6171,N_6142);
or U6263 (N_6263,N_6118,N_6137);
and U6264 (N_6264,N_6166,N_6132);
xnor U6265 (N_6265,N_6146,N_6111);
and U6266 (N_6266,N_6155,N_6123);
nor U6267 (N_6267,N_6107,N_6190);
nand U6268 (N_6268,N_6114,N_6140);
and U6269 (N_6269,N_6170,N_6134);
nor U6270 (N_6270,N_6173,N_6177);
nand U6271 (N_6271,N_6197,N_6139);
and U6272 (N_6272,N_6199,N_6162);
and U6273 (N_6273,N_6100,N_6132);
and U6274 (N_6274,N_6140,N_6189);
nand U6275 (N_6275,N_6139,N_6110);
nor U6276 (N_6276,N_6196,N_6172);
nor U6277 (N_6277,N_6111,N_6104);
and U6278 (N_6278,N_6194,N_6197);
nor U6279 (N_6279,N_6135,N_6142);
nor U6280 (N_6280,N_6159,N_6199);
nor U6281 (N_6281,N_6106,N_6154);
or U6282 (N_6282,N_6198,N_6189);
and U6283 (N_6283,N_6153,N_6167);
nand U6284 (N_6284,N_6159,N_6165);
nand U6285 (N_6285,N_6173,N_6180);
nor U6286 (N_6286,N_6136,N_6197);
or U6287 (N_6287,N_6163,N_6120);
nand U6288 (N_6288,N_6194,N_6125);
or U6289 (N_6289,N_6148,N_6184);
and U6290 (N_6290,N_6132,N_6152);
or U6291 (N_6291,N_6164,N_6131);
xor U6292 (N_6292,N_6147,N_6177);
and U6293 (N_6293,N_6101,N_6150);
nor U6294 (N_6294,N_6128,N_6170);
or U6295 (N_6295,N_6140,N_6192);
xnor U6296 (N_6296,N_6174,N_6150);
nand U6297 (N_6297,N_6128,N_6186);
and U6298 (N_6298,N_6196,N_6189);
or U6299 (N_6299,N_6190,N_6121);
and U6300 (N_6300,N_6254,N_6286);
or U6301 (N_6301,N_6202,N_6241);
nor U6302 (N_6302,N_6265,N_6267);
or U6303 (N_6303,N_6278,N_6288);
nor U6304 (N_6304,N_6205,N_6252);
or U6305 (N_6305,N_6204,N_6226);
nor U6306 (N_6306,N_6280,N_6219);
and U6307 (N_6307,N_6208,N_6245);
nor U6308 (N_6308,N_6238,N_6274);
nand U6309 (N_6309,N_6213,N_6218);
and U6310 (N_6310,N_6221,N_6269);
nand U6311 (N_6311,N_6246,N_6292);
and U6312 (N_6312,N_6264,N_6227);
nor U6313 (N_6313,N_6201,N_6212);
nor U6314 (N_6314,N_6249,N_6247);
or U6315 (N_6315,N_6279,N_6299);
and U6316 (N_6316,N_6203,N_6257);
and U6317 (N_6317,N_6253,N_6216);
xnor U6318 (N_6318,N_6282,N_6200);
nor U6319 (N_6319,N_6211,N_6281);
nand U6320 (N_6320,N_6232,N_6234);
or U6321 (N_6321,N_6296,N_6258);
or U6322 (N_6322,N_6271,N_6285);
nand U6323 (N_6323,N_6291,N_6295);
or U6324 (N_6324,N_6225,N_6284);
or U6325 (N_6325,N_6289,N_6236);
nor U6326 (N_6326,N_6250,N_6260);
or U6327 (N_6327,N_6266,N_6229);
or U6328 (N_6328,N_6293,N_6268);
or U6329 (N_6329,N_6228,N_6215);
xnor U6330 (N_6330,N_6210,N_6263);
and U6331 (N_6331,N_6237,N_6275);
and U6332 (N_6332,N_6242,N_6244);
and U6333 (N_6333,N_6270,N_6220);
nand U6334 (N_6334,N_6223,N_6243);
nand U6335 (N_6335,N_6273,N_6240);
nor U6336 (N_6336,N_6248,N_6230);
or U6337 (N_6337,N_6297,N_6233);
nor U6338 (N_6338,N_6207,N_6209);
and U6339 (N_6339,N_6222,N_6235);
nand U6340 (N_6340,N_6239,N_6287);
nor U6341 (N_6341,N_6255,N_6259);
xor U6342 (N_6342,N_6294,N_6217);
and U6343 (N_6343,N_6276,N_6256);
nor U6344 (N_6344,N_6277,N_6231);
nand U6345 (N_6345,N_6224,N_6261);
and U6346 (N_6346,N_6272,N_6290);
nand U6347 (N_6347,N_6214,N_6298);
and U6348 (N_6348,N_6262,N_6251);
xnor U6349 (N_6349,N_6283,N_6206);
or U6350 (N_6350,N_6248,N_6219);
nand U6351 (N_6351,N_6208,N_6220);
nand U6352 (N_6352,N_6203,N_6278);
nand U6353 (N_6353,N_6247,N_6285);
xnor U6354 (N_6354,N_6205,N_6280);
nor U6355 (N_6355,N_6279,N_6273);
nand U6356 (N_6356,N_6245,N_6240);
nand U6357 (N_6357,N_6291,N_6293);
or U6358 (N_6358,N_6278,N_6264);
or U6359 (N_6359,N_6260,N_6271);
xnor U6360 (N_6360,N_6282,N_6295);
or U6361 (N_6361,N_6206,N_6241);
nor U6362 (N_6362,N_6221,N_6289);
nor U6363 (N_6363,N_6280,N_6282);
nand U6364 (N_6364,N_6285,N_6259);
nor U6365 (N_6365,N_6294,N_6210);
nand U6366 (N_6366,N_6241,N_6291);
nor U6367 (N_6367,N_6269,N_6207);
nand U6368 (N_6368,N_6259,N_6296);
xnor U6369 (N_6369,N_6231,N_6240);
or U6370 (N_6370,N_6240,N_6275);
nand U6371 (N_6371,N_6290,N_6246);
and U6372 (N_6372,N_6299,N_6252);
and U6373 (N_6373,N_6244,N_6289);
nor U6374 (N_6374,N_6225,N_6292);
and U6375 (N_6375,N_6274,N_6277);
xor U6376 (N_6376,N_6293,N_6263);
nor U6377 (N_6377,N_6228,N_6298);
and U6378 (N_6378,N_6283,N_6200);
xor U6379 (N_6379,N_6204,N_6283);
and U6380 (N_6380,N_6221,N_6265);
nand U6381 (N_6381,N_6287,N_6298);
nand U6382 (N_6382,N_6298,N_6212);
nand U6383 (N_6383,N_6237,N_6271);
xnor U6384 (N_6384,N_6296,N_6208);
and U6385 (N_6385,N_6220,N_6247);
nand U6386 (N_6386,N_6220,N_6224);
or U6387 (N_6387,N_6265,N_6219);
nor U6388 (N_6388,N_6224,N_6210);
nor U6389 (N_6389,N_6253,N_6250);
or U6390 (N_6390,N_6205,N_6219);
nor U6391 (N_6391,N_6289,N_6217);
xor U6392 (N_6392,N_6293,N_6238);
nand U6393 (N_6393,N_6225,N_6246);
xnor U6394 (N_6394,N_6235,N_6262);
xnor U6395 (N_6395,N_6278,N_6214);
nor U6396 (N_6396,N_6282,N_6288);
nand U6397 (N_6397,N_6244,N_6219);
and U6398 (N_6398,N_6249,N_6286);
nor U6399 (N_6399,N_6243,N_6215);
and U6400 (N_6400,N_6363,N_6396);
nand U6401 (N_6401,N_6354,N_6324);
and U6402 (N_6402,N_6344,N_6378);
nor U6403 (N_6403,N_6362,N_6311);
and U6404 (N_6404,N_6361,N_6377);
nand U6405 (N_6405,N_6350,N_6372);
xor U6406 (N_6406,N_6321,N_6318);
and U6407 (N_6407,N_6374,N_6368);
and U6408 (N_6408,N_6371,N_6348);
xor U6409 (N_6409,N_6383,N_6369);
and U6410 (N_6410,N_6323,N_6390);
or U6411 (N_6411,N_6341,N_6335);
nor U6412 (N_6412,N_6375,N_6313);
nor U6413 (N_6413,N_6360,N_6366);
or U6414 (N_6414,N_6316,N_6302);
nor U6415 (N_6415,N_6336,N_6340);
or U6416 (N_6416,N_6346,N_6339);
and U6417 (N_6417,N_6388,N_6385);
and U6418 (N_6418,N_6317,N_6320);
nand U6419 (N_6419,N_6325,N_6329);
and U6420 (N_6420,N_6355,N_6391);
nor U6421 (N_6421,N_6330,N_6386);
or U6422 (N_6422,N_6334,N_6310);
or U6423 (N_6423,N_6387,N_6301);
nand U6424 (N_6424,N_6352,N_6376);
nor U6425 (N_6425,N_6309,N_6398);
nand U6426 (N_6426,N_6359,N_6364);
nand U6427 (N_6427,N_6342,N_6379);
nor U6428 (N_6428,N_6300,N_6326);
nor U6429 (N_6429,N_6338,N_6382);
xor U6430 (N_6430,N_6380,N_6343);
and U6431 (N_6431,N_6347,N_6351);
or U6432 (N_6432,N_6337,N_6367);
and U6433 (N_6433,N_6392,N_6381);
nand U6434 (N_6434,N_6365,N_6393);
and U6435 (N_6435,N_6395,N_6332);
xnor U6436 (N_6436,N_6327,N_6315);
nand U6437 (N_6437,N_6357,N_6345);
and U6438 (N_6438,N_6389,N_6307);
nand U6439 (N_6439,N_6370,N_6331);
nand U6440 (N_6440,N_6306,N_6394);
nand U6441 (N_6441,N_6304,N_6328);
or U6442 (N_6442,N_6384,N_6399);
and U6443 (N_6443,N_6303,N_6322);
or U6444 (N_6444,N_6356,N_6353);
and U6445 (N_6445,N_6314,N_6349);
and U6446 (N_6446,N_6308,N_6312);
or U6447 (N_6447,N_6319,N_6397);
nor U6448 (N_6448,N_6358,N_6373);
and U6449 (N_6449,N_6305,N_6333);
xnor U6450 (N_6450,N_6369,N_6346);
or U6451 (N_6451,N_6323,N_6306);
and U6452 (N_6452,N_6314,N_6331);
xnor U6453 (N_6453,N_6396,N_6312);
or U6454 (N_6454,N_6371,N_6355);
and U6455 (N_6455,N_6308,N_6396);
or U6456 (N_6456,N_6310,N_6317);
and U6457 (N_6457,N_6319,N_6318);
or U6458 (N_6458,N_6394,N_6391);
or U6459 (N_6459,N_6346,N_6311);
or U6460 (N_6460,N_6370,N_6328);
or U6461 (N_6461,N_6350,N_6371);
or U6462 (N_6462,N_6393,N_6301);
nand U6463 (N_6463,N_6341,N_6391);
nand U6464 (N_6464,N_6314,N_6315);
and U6465 (N_6465,N_6308,N_6368);
xnor U6466 (N_6466,N_6325,N_6344);
and U6467 (N_6467,N_6379,N_6314);
and U6468 (N_6468,N_6389,N_6393);
nor U6469 (N_6469,N_6337,N_6348);
nor U6470 (N_6470,N_6311,N_6328);
nand U6471 (N_6471,N_6374,N_6385);
and U6472 (N_6472,N_6376,N_6325);
nand U6473 (N_6473,N_6336,N_6369);
or U6474 (N_6474,N_6342,N_6331);
nand U6475 (N_6475,N_6348,N_6321);
xor U6476 (N_6476,N_6392,N_6368);
and U6477 (N_6477,N_6322,N_6348);
nor U6478 (N_6478,N_6381,N_6346);
nand U6479 (N_6479,N_6389,N_6334);
nor U6480 (N_6480,N_6315,N_6376);
nor U6481 (N_6481,N_6354,N_6369);
or U6482 (N_6482,N_6366,N_6396);
nand U6483 (N_6483,N_6353,N_6324);
nor U6484 (N_6484,N_6317,N_6328);
nand U6485 (N_6485,N_6308,N_6348);
nand U6486 (N_6486,N_6310,N_6307);
or U6487 (N_6487,N_6328,N_6389);
or U6488 (N_6488,N_6324,N_6386);
or U6489 (N_6489,N_6348,N_6398);
and U6490 (N_6490,N_6338,N_6360);
or U6491 (N_6491,N_6316,N_6359);
or U6492 (N_6492,N_6399,N_6346);
nor U6493 (N_6493,N_6383,N_6358);
xnor U6494 (N_6494,N_6379,N_6306);
nor U6495 (N_6495,N_6350,N_6383);
nand U6496 (N_6496,N_6399,N_6381);
nor U6497 (N_6497,N_6336,N_6387);
or U6498 (N_6498,N_6311,N_6352);
nand U6499 (N_6499,N_6395,N_6303);
nor U6500 (N_6500,N_6440,N_6401);
xnor U6501 (N_6501,N_6420,N_6461);
nor U6502 (N_6502,N_6428,N_6435);
nand U6503 (N_6503,N_6452,N_6439);
nor U6504 (N_6504,N_6432,N_6414);
nor U6505 (N_6505,N_6489,N_6474);
and U6506 (N_6506,N_6426,N_6406);
and U6507 (N_6507,N_6448,N_6485);
nor U6508 (N_6508,N_6445,N_6421);
or U6509 (N_6509,N_6433,N_6457);
or U6510 (N_6510,N_6478,N_6492);
nor U6511 (N_6511,N_6484,N_6480);
nand U6512 (N_6512,N_6447,N_6427);
nor U6513 (N_6513,N_6412,N_6493);
or U6514 (N_6514,N_6466,N_6405);
and U6515 (N_6515,N_6419,N_6418);
nor U6516 (N_6516,N_6410,N_6455);
nand U6517 (N_6517,N_6472,N_6402);
and U6518 (N_6518,N_6425,N_6486);
nand U6519 (N_6519,N_6459,N_6430);
nor U6520 (N_6520,N_6483,N_6449);
nor U6521 (N_6521,N_6404,N_6496);
or U6522 (N_6522,N_6434,N_6479);
nand U6523 (N_6523,N_6495,N_6437);
nand U6524 (N_6524,N_6403,N_6456);
nor U6525 (N_6525,N_6475,N_6499);
xnor U6526 (N_6526,N_6429,N_6488);
and U6527 (N_6527,N_6481,N_6491);
nand U6528 (N_6528,N_6465,N_6422);
nand U6529 (N_6529,N_6464,N_6409);
or U6530 (N_6530,N_6498,N_6408);
nand U6531 (N_6531,N_6468,N_6454);
and U6532 (N_6532,N_6460,N_6443);
and U6533 (N_6533,N_6423,N_6494);
and U6534 (N_6534,N_6431,N_6467);
nor U6535 (N_6535,N_6446,N_6470);
xnor U6536 (N_6536,N_6413,N_6450);
xnor U6537 (N_6537,N_6444,N_6497);
nand U6538 (N_6538,N_6469,N_6417);
or U6539 (N_6539,N_6451,N_6462);
or U6540 (N_6540,N_6442,N_6416);
and U6541 (N_6541,N_6438,N_6473);
nor U6542 (N_6542,N_6400,N_6487);
nand U6543 (N_6543,N_6490,N_6471);
xor U6544 (N_6544,N_6458,N_6411);
and U6545 (N_6545,N_6482,N_6477);
nor U6546 (N_6546,N_6436,N_6441);
and U6547 (N_6547,N_6415,N_6476);
nor U6548 (N_6548,N_6407,N_6453);
nor U6549 (N_6549,N_6463,N_6424);
nand U6550 (N_6550,N_6409,N_6418);
nor U6551 (N_6551,N_6464,N_6449);
xnor U6552 (N_6552,N_6480,N_6465);
or U6553 (N_6553,N_6402,N_6497);
or U6554 (N_6554,N_6461,N_6403);
xor U6555 (N_6555,N_6481,N_6402);
or U6556 (N_6556,N_6406,N_6493);
nor U6557 (N_6557,N_6454,N_6464);
nand U6558 (N_6558,N_6484,N_6489);
xnor U6559 (N_6559,N_6499,N_6408);
xnor U6560 (N_6560,N_6429,N_6448);
or U6561 (N_6561,N_6413,N_6436);
nand U6562 (N_6562,N_6479,N_6486);
and U6563 (N_6563,N_6435,N_6421);
nor U6564 (N_6564,N_6456,N_6477);
xnor U6565 (N_6565,N_6468,N_6439);
or U6566 (N_6566,N_6429,N_6446);
and U6567 (N_6567,N_6406,N_6407);
and U6568 (N_6568,N_6490,N_6485);
or U6569 (N_6569,N_6445,N_6410);
nand U6570 (N_6570,N_6498,N_6458);
or U6571 (N_6571,N_6488,N_6417);
nand U6572 (N_6572,N_6446,N_6423);
and U6573 (N_6573,N_6444,N_6447);
or U6574 (N_6574,N_6445,N_6449);
nor U6575 (N_6575,N_6425,N_6419);
nand U6576 (N_6576,N_6490,N_6452);
nor U6577 (N_6577,N_6469,N_6413);
nand U6578 (N_6578,N_6452,N_6457);
and U6579 (N_6579,N_6429,N_6434);
and U6580 (N_6580,N_6486,N_6407);
or U6581 (N_6581,N_6471,N_6476);
nand U6582 (N_6582,N_6445,N_6455);
and U6583 (N_6583,N_6474,N_6422);
nand U6584 (N_6584,N_6440,N_6448);
nand U6585 (N_6585,N_6458,N_6408);
nor U6586 (N_6586,N_6424,N_6419);
or U6587 (N_6587,N_6411,N_6493);
nand U6588 (N_6588,N_6460,N_6435);
nor U6589 (N_6589,N_6467,N_6409);
nand U6590 (N_6590,N_6438,N_6443);
or U6591 (N_6591,N_6468,N_6415);
nor U6592 (N_6592,N_6466,N_6423);
or U6593 (N_6593,N_6409,N_6469);
and U6594 (N_6594,N_6427,N_6414);
nand U6595 (N_6595,N_6428,N_6452);
nor U6596 (N_6596,N_6467,N_6470);
nand U6597 (N_6597,N_6470,N_6402);
xor U6598 (N_6598,N_6449,N_6417);
and U6599 (N_6599,N_6454,N_6416);
and U6600 (N_6600,N_6597,N_6542);
and U6601 (N_6601,N_6522,N_6512);
or U6602 (N_6602,N_6536,N_6503);
and U6603 (N_6603,N_6587,N_6531);
and U6604 (N_6604,N_6546,N_6589);
and U6605 (N_6605,N_6583,N_6550);
nor U6606 (N_6606,N_6501,N_6596);
nor U6607 (N_6607,N_6560,N_6518);
xor U6608 (N_6608,N_6580,N_6572);
and U6609 (N_6609,N_6566,N_6573);
nand U6610 (N_6610,N_6571,N_6544);
and U6611 (N_6611,N_6561,N_6593);
nor U6612 (N_6612,N_6506,N_6591);
or U6613 (N_6613,N_6562,N_6568);
and U6614 (N_6614,N_6590,N_6570);
nor U6615 (N_6615,N_6535,N_6509);
nand U6616 (N_6616,N_6564,N_6552);
or U6617 (N_6617,N_6599,N_6526);
nand U6618 (N_6618,N_6505,N_6557);
and U6619 (N_6619,N_6534,N_6543);
xnor U6620 (N_6620,N_6515,N_6537);
nand U6621 (N_6621,N_6521,N_6559);
and U6622 (N_6622,N_6548,N_6581);
nor U6623 (N_6623,N_6510,N_6516);
nand U6624 (N_6624,N_6528,N_6539);
and U6625 (N_6625,N_6530,N_6595);
xor U6626 (N_6626,N_6598,N_6567);
or U6627 (N_6627,N_6577,N_6579);
nand U6628 (N_6628,N_6549,N_6563);
nor U6629 (N_6629,N_6565,N_6533);
or U6630 (N_6630,N_6517,N_6584);
nor U6631 (N_6631,N_6578,N_6500);
nor U6632 (N_6632,N_6532,N_6553);
nor U6633 (N_6633,N_6558,N_6523);
and U6634 (N_6634,N_6527,N_6520);
or U6635 (N_6635,N_6519,N_6576);
or U6636 (N_6636,N_6547,N_6555);
and U6637 (N_6637,N_6524,N_6538);
or U6638 (N_6638,N_6575,N_6556);
and U6639 (N_6639,N_6545,N_6551);
and U6640 (N_6640,N_6504,N_6513);
or U6641 (N_6641,N_6529,N_6507);
and U6642 (N_6642,N_6541,N_6514);
or U6643 (N_6643,N_6554,N_6511);
and U6644 (N_6644,N_6586,N_6508);
or U6645 (N_6645,N_6588,N_6574);
nor U6646 (N_6646,N_6585,N_6525);
nor U6647 (N_6647,N_6582,N_6594);
and U6648 (N_6648,N_6540,N_6592);
or U6649 (N_6649,N_6569,N_6502);
or U6650 (N_6650,N_6544,N_6586);
or U6651 (N_6651,N_6531,N_6577);
or U6652 (N_6652,N_6533,N_6521);
nand U6653 (N_6653,N_6556,N_6576);
and U6654 (N_6654,N_6576,N_6591);
nor U6655 (N_6655,N_6588,N_6518);
nor U6656 (N_6656,N_6568,N_6540);
xor U6657 (N_6657,N_6524,N_6514);
or U6658 (N_6658,N_6544,N_6501);
nand U6659 (N_6659,N_6536,N_6507);
nand U6660 (N_6660,N_6526,N_6562);
or U6661 (N_6661,N_6563,N_6530);
and U6662 (N_6662,N_6554,N_6579);
and U6663 (N_6663,N_6598,N_6547);
and U6664 (N_6664,N_6563,N_6508);
nand U6665 (N_6665,N_6581,N_6529);
and U6666 (N_6666,N_6525,N_6587);
nand U6667 (N_6667,N_6589,N_6501);
and U6668 (N_6668,N_6583,N_6588);
and U6669 (N_6669,N_6573,N_6589);
nor U6670 (N_6670,N_6584,N_6567);
and U6671 (N_6671,N_6592,N_6520);
or U6672 (N_6672,N_6528,N_6508);
xor U6673 (N_6673,N_6507,N_6546);
or U6674 (N_6674,N_6506,N_6522);
nand U6675 (N_6675,N_6523,N_6530);
nor U6676 (N_6676,N_6587,N_6574);
or U6677 (N_6677,N_6508,N_6594);
nor U6678 (N_6678,N_6563,N_6579);
or U6679 (N_6679,N_6540,N_6563);
and U6680 (N_6680,N_6585,N_6528);
nor U6681 (N_6681,N_6535,N_6554);
or U6682 (N_6682,N_6531,N_6528);
nor U6683 (N_6683,N_6520,N_6573);
xor U6684 (N_6684,N_6547,N_6561);
or U6685 (N_6685,N_6520,N_6536);
or U6686 (N_6686,N_6559,N_6525);
nand U6687 (N_6687,N_6521,N_6503);
or U6688 (N_6688,N_6551,N_6567);
or U6689 (N_6689,N_6532,N_6542);
nand U6690 (N_6690,N_6540,N_6534);
and U6691 (N_6691,N_6589,N_6540);
and U6692 (N_6692,N_6515,N_6539);
or U6693 (N_6693,N_6570,N_6542);
or U6694 (N_6694,N_6511,N_6570);
nor U6695 (N_6695,N_6500,N_6562);
nor U6696 (N_6696,N_6597,N_6598);
and U6697 (N_6697,N_6541,N_6524);
or U6698 (N_6698,N_6574,N_6547);
or U6699 (N_6699,N_6538,N_6549);
or U6700 (N_6700,N_6662,N_6641);
or U6701 (N_6701,N_6649,N_6628);
or U6702 (N_6702,N_6679,N_6698);
nand U6703 (N_6703,N_6626,N_6687);
nor U6704 (N_6704,N_6684,N_6686);
or U6705 (N_6705,N_6619,N_6602);
xor U6706 (N_6706,N_6689,N_6657);
nor U6707 (N_6707,N_6648,N_6697);
xor U6708 (N_6708,N_6677,N_6609);
and U6709 (N_6709,N_6694,N_6681);
or U6710 (N_6710,N_6636,N_6646);
and U6711 (N_6711,N_6661,N_6673);
xnor U6712 (N_6712,N_6650,N_6604);
and U6713 (N_6713,N_6645,N_6635);
or U6714 (N_6714,N_6692,N_6659);
and U6715 (N_6715,N_6699,N_6654);
nor U6716 (N_6716,N_6680,N_6618);
nand U6717 (N_6717,N_6642,N_6613);
or U6718 (N_6718,N_6653,N_6615);
and U6719 (N_6719,N_6605,N_6608);
or U6720 (N_6720,N_6601,N_6647);
or U6721 (N_6721,N_6607,N_6663);
nand U6722 (N_6722,N_6665,N_6678);
and U6723 (N_6723,N_6629,N_6693);
nor U6724 (N_6724,N_6644,N_6671);
nor U6725 (N_6725,N_6603,N_6633);
nor U6726 (N_6726,N_6625,N_6612);
nor U6727 (N_6727,N_6621,N_6658);
nor U6728 (N_6728,N_6664,N_6672);
or U6729 (N_6729,N_6616,N_6634);
nor U6730 (N_6730,N_6674,N_6652);
nand U6731 (N_6731,N_6614,N_6667);
nand U6732 (N_6732,N_6651,N_6688);
or U6733 (N_6733,N_6696,N_6655);
or U6734 (N_6734,N_6695,N_6669);
xor U6735 (N_6735,N_6623,N_6637);
and U6736 (N_6736,N_6617,N_6622);
nand U6737 (N_6737,N_6640,N_6656);
and U6738 (N_6738,N_6660,N_6620);
and U6739 (N_6739,N_6606,N_6643);
and U6740 (N_6740,N_6638,N_6627);
nor U6741 (N_6741,N_6668,N_6632);
nand U6742 (N_6742,N_6624,N_6639);
or U6743 (N_6743,N_6600,N_6683);
nand U6744 (N_6744,N_6611,N_6670);
nor U6745 (N_6745,N_6691,N_6630);
and U6746 (N_6746,N_6690,N_6666);
or U6747 (N_6747,N_6685,N_6610);
nand U6748 (N_6748,N_6631,N_6675);
nor U6749 (N_6749,N_6682,N_6676);
nand U6750 (N_6750,N_6655,N_6601);
nand U6751 (N_6751,N_6683,N_6693);
nor U6752 (N_6752,N_6640,N_6632);
or U6753 (N_6753,N_6684,N_6680);
nor U6754 (N_6754,N_6600,N_6676);
nand U6755 (N_6755,N_6611,N_6613);
nand U6756 (N_6756,N_6663,N_6683);
nand U6757 (N_6757,N_6612,N_6656);
or U6758 (N_6758,N_6632,N_6663);
nand U6759 (N_6759,N_6691,N_6649);
nor U6760 (N_6760,N_6682,N_6638);
nor U6761 (N_6761,N_6619,N_6607);
xor U6762 (N_6762,N_6692,N_6607);
nor U6763 (N_6763,N_6669,N_6683);
or U6764 (N_6764,N_6618,N_6628);
nand U6765 (N_6765,N_6689,N_6692);
or U6766 (N_6766,N_6605,N_6626);
and U6767 (N_6767,N_6601,N_6654);
xor U6768 (N_6768,N_6653,N_6648);
nor U6769 (N_6769,N_6602,N_6635);
or U6770 (N_6770,N_6606,N_6603);
xnor U6771 (N_6771,N_6629,N_6644);
and U6772 (N_6772,N_6670,N_6620);
nor U6773 (N_6773,N_6644,N_6657);
nor U6774 (N_6774,N_6622,N_6609);
and U6775 (N_6775,N_6659,N_6628);
and U6776 (N_6776,N_6609,N_6657);
nand U6777 (N_6777,N_6658,N_6602);
and U6778 (N_6778,N_6644,N_6610);
nor U6779 (N_6779,N_6688,N_6685);
and U6780 (N_6780,N_6600,N_6644);
or U6781 (N_6781,N_6668,N_6678);
and U6782 (N_6782,N_6629,N_6681);
nand U6783 (N_6783,N_6643,N_6623);
nor U6784 (N_6784,N_6690,N_6633);
nand U6785 (N_6785,N_6678,N_6659);
or U6786 (N_6786,N_6664,N_6669);
and U6787 (N_6787,N_6613,N_6680);
nand U6788 (N_6788,N_6648,N_6683);
xnor U6789 (N_6789,N_6650,N_6622);
nor U6790 (N_6790,N_6674,N_6693);
xor U6791 (N_6791,N_6653,N_6612);
or U6792 (N_6792,N_6675,N_6663);
and U6793 (N_6793,N_6664,N_6654);
nor U6794 (N_6794,N_6656,N_6663);
nor U6795 (N_6795,N_6683,N_6673);
or U6796 (N_6796,N_6626,N_6682);
nand U6797 (N_6797,N_6683,N_6626);
and U6798 (N_6798,N_6657,N_6683);
nand U6799 (N_6799,N_6688,N_6617);
nand U6800 (N_6800,N_6785,N_6723);
nand U6801 (N_6801,N_6729,N_6731);
nand U6802 (N_6802,N_6747,N_6760);
nor U6803 (N_6803,N_6701,N_6776);
and U6804 (N_6804,N_6728,N_6740);
and U6805 (N_6805,N_6725,N_6761);
and U6806 (N_6806,N_6704,N_6734);
nand U6807 (N_6807,N_6771,N_6773);
nand U6808 (N_6808,N_6781,N_6719);
nand U6809 (N_6809,N_6778,N_6744);
nand U6810 (N_6810,N_6741,N_6767);
nand U6811 (N_6811,N_6790,N_6799);
or U6812 (N_6812,N_6739,N_6764);
nor U6813 (N_6813,N_6768,N_6758);
nand U6814 (N_6814,N_6779,N_6718);
or U6815 (N_6815,N_6753,N_6711);
and U6816 (N_6816,N_6757,N_6705);
nand U6817 (N_6817,N_6749,N_6796);
nand U6818 (N_6818,N_6724,N_6722);
nor U6819 (N_6819,N_6737,N_6792);
nor U6820 (N_6820,N_6702,N_6791);
nor U6821 (N_6821,N_6795,N_6775);
nand U6822 (N_6822,N_6794,N_6726);
nor U6823 (N_6823,N_6709,N_6780);
nor U6824 (N_6824,N_6735,N_6754);
and U6825 (N_6825,N_6772,N_6721);
and U6826 (N_6826,N_6708,N_6742);
nor U6827 (N_6827,N_6706,N_6703);
or U6828 (N_6828,N_6762,N_6748);
or U6829 (N_6829,N_6769,N_6786);
and U6830 (N_6830,N_6710,N_6715);
nand U6831 (N_6831,N_6745,N_6738);
xor U6832 (N_6832,N_6713,N_6777);
or U6833 (N_6833,N_6755,N_6720);
nor U6834 (N_6834,N_6770,N_6712);
and U6835 (N_6835,N_6732,N_6787);
or U6836 (N_6836,N_6736,N_6717);
nor U6837 (N_6837,N_6783,N_6759);
nand U6838 (N_6838,N_6746,N_6730);
and U6839 (N_6839,N_6727,N_6750);
or U6840 (N_6840,N_6716,N_6707);
xor U6841 (N_6841,N_6766,N_6793);
or U6842 (N_6842,N_6743,N_6797);
nor U6843 (N_6843,N_6751,N_6756);
nand U6844 (N_6844,N_6765,N_6752);
or U6845 (N_6845,N_6788,N_6733);
and U6846 (N_6846,N_6789,N_6700);
or U6847 (N_6847,N_6782,N_6714);
or U6848 (N_6848,N_6763,N_6784);
and U6849 (N_6849,N_6798,N_6774);
and U6850 (N_6850,N_6785,N_6709);
nand U6851 (N_6851,N_6798,N_6764);
nor U6852 (N_6852,N_6743,N_6760);
nand U6853 (N_6853,N_6705,N_6748);
and U6854 (N_6854,N_6735,N_6730);
nand U6855 (N_6855,N_6712,N_6732);
nor U6856 (N_6856,N_6750,N_6716);
or U6857 (N_6857,N_6783,N_6702);
nand U6858 (N_6858,N_6724,N_6787);
and U6859 (N_6859,N_6760,N_6777);
or U6860 (N_6860,N_6772,N_6717);
nor U6861 (N_6861,N_6700,N_6717);
nor U6862 (N_6862,N_6771,N_6754);
nor U6863 (N_6863,N_6754,N_6797);
and U6864 (N_6864,N_6700,N_6795);
nand U6865 (N_6865,N_6763,N_6748);
nor U6866 (N_6866,N_6756,N_6724);
and U6867 (N_6867,N_6734,N_6718);
nor U6868 (N_6868,N_6778,N_6796);
xnor U6869 (N_6869,N_6741,N_6751);
nand U6870 (N_6870,N_6750,N_6717);
nand U6871 (N_6871,N_6797,N_6716);
nor U6872 (N_6872,N_6742,N_6741);
and U6873 (N_6873,N_6781,N_6701);
nand U6874 (N_6874,N_6746,N_6741);
nor U6875 (N_6875,N_6775,N_6790);
nor U6876 (N_6876,N_6768,N_6752);
nand U6877 (N_6877,N_6725,N_6748);
xor U6878 (N_6878,N_6789,N_6704);
xnor U6879 (N_6879,N_6719,N_6770);
or U6880 (N_6880,N_6722,N_6706);
nor U6881 (N_6881,N_6723,N_6753);
xor U6882 (N_6882,N_6750,N_6772);
nor U6883 (N_6883,N_6737,N_6719);
or U6884 (N_6884,N_6773,N_6768);
xor U6885 (N_6885,N_6746,N_6727);
and U6886 (N_6886,N_6731,N_6724);
and U6887 (N_6887,N_6703,N_6715);
nand U6888 (N_6888,N_6718,N_6702);
and U6889 (N_6889,N_6727,N_6705);
nor U6890 (N_6890,N_6760,N_6789);
and U6891 (N_6891,N_6787,N_6740);
and U6892 (N_6892,N_6731,N_6783);
nor U6893 (N_6893,N_6738,N_6741);
and U6894 (N_6894,N_6788,N_6750);
and U6895 (N_6895,N_6709,N_6798);
xor U6896 (N_6896,N_6795,N_6707);
or U6897 (N_6897,N_6773,N_6739);
and U6898 (N_6898,N_6720,N_6718);
nor U6899 (N_6899,N_6716,N_6760);
and U6900 (N_6900,N_6830,N_6840);
xnor U6901 (N_6901,N_6816,N_6884);
nor U6902 (N_6902,N_6838,N_6834);
or U6903 (N_6903,N_6837,N_6890);
or U6904 (N_6904,N_6820,N_6801);
nand U6905 (N_6905,N_6876,N_6808);
and U6906 (N_6906,N_6802,N_6885);
nand U6907 (N_6907,N_6863,N_6864);
nand U6908 (N_6908,N_6815,N_6877);
and U6909 (N_6909,N_6882,N_6818);
nand U6910 (N_6910,N_6855,N_6868);
and U6911 (N_6911,N_6805,N_6897);
nor U6912 (N_6912,N_6860,N_6874);
or U6913 (N_6913,N_6851,N_6873);
nor U6914 (N_6914,N_6888,N_6862);
nor U6915 (N_6915,N_6829,N_6866);
xnor U6916 (N_6916,N_6879,N_6894);
or U6917 (N_6917,N_6883,N_6887);
xnor U6918 (N_6918,N_6853,N_6861);
or U6919 (N_6919,N_6803,N_6847);
or U6920 (N_6920,N_6806,N_6835);
nand U6921 (N_6921,N_6854,N_6831);
and U6922 (N_6922,N_6881,N_6895);
or U6923 (N_6923,N_6899,N_6844);
nand U6924 (N_6924,N_6822,N_6824);
and U6925 (N_6925,N_6892,N_6836);
nor U6926 (N_6926,N_6880,N_6823);
or U6927 (N_6927,N_6843,N_6800);
nor U6928 (N_6928,N_6869,N_6845);
nand U6929 (N_6929,N_6870,N_6848);
nand U6930 (N_6930,N_6807,N_6842);
xor U6931 (N_6931,N_6893,N_6841);
nor U6932 (N_6932,N_6809,N_6878);
nor U6933 (N_6933,N_6865,N_6886);
nand U6934 (N_6934,N_6898,N_6846);
nand U6935 (N_6935,N_6858,N_6833);
or U6936 (N_6936,N_6819,N_6826);
nor U6937 (N_6937,N_6889,N_6859);
and U6938 (N_6938,N_6821,N_6839);
and U6939 (N_6939,N_6891,N_6813);
or U6940 (N_6940,N_6849,N_6871);
and U6941 (N_6941,N_6856,N_6810);
or U6942 (N_6942,N_6825,N_6817);
and U6943 (N_6943,N_6804,N_6850);
or U6944 (N_6944,N_6867,N_6828);
nor U6945 (N_6945,N_6832,N_6857);
nand U6946 (N_6946,N_6852,N_6811);
nand U6947 (N_6947,N_6812,N_6872);
and U6948 (N_6948,N_6896,N_6875);
nand U6949 (N_6949,N_6827,N_6814);
or U6950 (N_6950,N_6833,N_6887);
nor U6951 (N_6951,N_6871,N_6844);
and U6952 (N_6952,N_6840,N_6814);
or U6953 (N_6953,N_6815,N_6818);
or U6954 (N_6954,N_6808,N_6882);
nor U6955 (N_6955,N_6868,N_6833);
and U6956 (N_6956,N_6849,N_6815);
nor U6957 (N_6957,N_6885,N_6868);
nor U6958 (N_6958,N_6849,N_6888);
xor U6959 (N_6959,N_6822,N_6868);
or U6960 (N_6960,N_6805,N_6819);
and U6961 (N_6961,N_6823,N_6834);
nand U6962 (N_6962,N_6858,N_6863);
or U6963 (N_6963,N_6811,N_6833);
nand U6964 (N_6964,N_6880,N_6810);
and U6965 (N_6965,N_6862,N_6832);
or U6966 (N_6966,N_6889,N_6846);
nor U6967 (N_6967,N_6837,N_6817);
xnor U6968 (N_6968,N_6845,N_6877);
or U6969 (N_6969,N_6846,N_6840);
nand U6970 (N_6970,N_6892,N_6816);
nand U6971 (N_6971,N_6852,N_6884);
nor U6972 (N_6972,N_6802,N_6849);
nor U6973 (N_6973,N_6818,N_6895);
or U6974 (N_6974,N_6804,N_6854);
nor U6975 (N_6975,N_6814,N_6874);
or U6976 (N_6976,N_6879,N_6814);
nand U6977 (N_6977,N_6857,N_6813);
nand U6978 (N_6978,N_6852,N_6830);
or U6979 (N_6979,N_6810,N_6822);
or U6980 (N_6980,N_6822,N_6830);
nor U6981 (N_6981,N_6820,N_6872);
and U6982 (N_6982,N_6813,N_6806);
or U6983 (N_6983,N_6867,N_6878);
or U6984 (N_6984,N_6849,N_6844);
nand U6985 (N_6985,N_6878,N_6831);
or U6986 (N_6986,N_6872,N_6857);
and U6987 (N_6987,N_6887,N_6815);
nor U6988 (N_6988,N_6888,N_6833);
nand U6989 (N_6989,N_6808,N_6831);
and U6990 (N_6990,N_6878,N_6816);
and U6991 (N_6991,N_6844,N_6819);
nand U6992 (N_6992,N_6803,N_6831);
or U6993 (N_6993,N_6882,N_6871);
nor U6994 (N_6994,N_6830,N_6841);
or U6995 (N_6995,N_6848,N_6836);
nand U6996 (N_6996,N_6806,N_6872);
or U6997 (N_6997,N_6852,N_6802);
nor U6998 (N_6998,N_6816,N_6864);
or U6999 (N_6999,N_6830,N_6823);
nand U7000 (N_7000,N_6984,N_6951);
nor U7001 (N_7001,N_6983,N_6913);
nand U7002 (N_7002,N_6971,N_6967);
nor U7003 (N_7003,N_6991,N_6904);
or U7004 (N_7004,N_6969,N_6938);
nand U7005 (N_7005,N_6908,N_6995);
nand U7006 (N_7006,N_6903,N_6920);
or U7007 (N_7007,N_6902,N_6941);
or U7008 (N_7008,N_6990,N_6932);
and U7009 (N_7009,N_6911,N_6923);
nand U7010 (N_7010,N_6975,N_6963);
nor U7011 (N_7011,N_6968,N_6929);
or U7012 (N_7012,N_6985,N_6940);
and U7013 (N_7013,N_6974,N_6996);
nand U7014 (N_7014,N_6988,N_6964);
or U7015 (N_7015,N_6958,N_6981);
or U7016 (N_7016,N_6935,N_6979);
and U7017 (N_7017,N_6942,N_6922);
or U7018 (N_7018,N_6926,N_6909);
nor U7019 (N_7019,N_6978,N_6918);
nor U7020 (N_7020,N_6930,N_6960);
and U7021 (N_7021,N_6924,N_6966);
nor U7022 (N_7022,N_6961,N_6928);
and U7023 (N_7023,N_6970,N_6916);
nand U7024 (N_7024,N_6956,N_6933);
or U7025 (N_7025,N_6947,N_6954);
nor U7026 (N_7026,N_6999,N_6936);
xnor U7027 (N_7027,N_6914,N_6915);
and U7028 (N_7028,N_6986,N_6997);
and U7029 (N_7029,N_6994,N_6927);
and U7030 (N_7030,N_6931,N_6989);
nor U7031 (N_7031,N_6907,N_6982);
or U7032 (N_7032,N_6917,N_6937);
nand U7033 (N_7033,N_6921,N_6976);
nand U7034 (N_7034,N_6950,N_6925);
nand U7035 (N_7035,N_6912,N_6919);
nand U7036 (N_7036,N_6993,N_6901);
or U7037 (N_7037,N_6949,N_6906);
or U7038 (N_7038,N_6944,N_6953);
and U7039 (N_7039,N_6905,N_6910);
and U7040 (N_7040,N_6957,N_6945);
or U7041 (N_7041,N_6992,N_6977);
or U7042 (N_7042,N_6980,N_6948);
and U7043 (N_7043,N_6998,N_6955);
nand U7044 (N_7044,N_6946,N_6952);
or U7045 (N_7045,N_6987,N_6959);
nor U7046 (N_7046,N_6900,N_6939);
nor U7047 (N_7047,N_6972,N_6965);
nand U7048 (N_7048,N_6934,N_6973);
nand U7049 (N_7049,N_6943,N_6962);
nor U7050 (N_7050,N_6933,N_6912);
nor U7051 (N_7051,N_6920,N_6969);
or U7052 (N_7052,N_6909,N_6923);
or U7053 (N_7053,N_6956,N_6973);
xor U7054 (N_7054,N_6907,N_6992);
and U7055 (N_7055,N_6928,N_6958);
nand U7056 (N_7056,N_6996,N_6913);
or U7057 (N_7057,N_6998,N_6935);
nand U7058 (N_7058,N_6952,N_6906);
or U7059 (N_7059,N_6949,N_6955);
or U7060 (N_7060,N_6961,N_6983);
or U7061 (N_7061,N_6940,N_6993);
nand U7062 (N_7062,N_6939,N_6921);
xnor U7063 (N_7063,N_6970,N_6991);
nand U7064 (N_7064,N_6908,N_6928);
nor U7065 (N_7065,N_6907,N_6963);
or U7066 (N_7066,N_6910,N_6936);
nor U7067 (N_7067,N_6993,N_6902);
or U7068 (N_7068,N_6966,N_6973);
nor U7069 (N_7069,N_6930,N_6957);
or U7070 (N_7070,N_6970,N_6932);
nand U7071 (N_7071,N_6997,N_6940);
nand U7072 (N_7072,N_6957,N_6978);
nand U7073 (N_7073,N_6912,N_6961);
and U7074 (N_7074,N_6945,N_6952);
nor U7075 (N_7075,N_6902,N_6995);
xnor U7076 (N_7076,N_6952,N_6938);
nand U7077 (N_7077,N_6988,N_6998);
nand U7078 (N_7078,N_6981,N_6952);
and U7079 (N_7079,N_6985,N_6918);
or U7080 (N_7080,N_6956,N_6925);
and U7081 (N_7081,N_6940,N_6903);
nand U7082 (N_7082,N_6994,N_6940);
or U7083 (N_7083,N_6958,N_6944);
and U7084 (N_7084,N_6990,N_6968);
and U7085 (N_7085,N_6981,N_6997);
nor U7086 (N_7086,N_6904,N_6940);
or U7087 (N_7087,N_6911,N_6984);
nand U7088 (N_7088,N_6960,N_6962);
nor U7089 (N_7089,N_6962,N_6949);
xnor U7090 (N_7090,N_6905,N_6985);
nand U7091 (N_7091,N_6977,N_6912);
nor U7092 (N_7092,N_6977,N_6914);
nand U7093 (N_7093,N_6908,N_6951);
xnor U7094 (N_7094,N_6918,N_6996);
and U7095 (N_7095,N_6981,N_6975);
nand U7096 (N_7096,N_6904,N_6983);
xor U7097 (N_7097,N_6991,N_6962);
xnor U7098 (N_7098,N_6902,N_6903);
or U7099 (N_7099,N_6976,N_6978);
nor U7100 (N_7100,N_7008,N_7028);
and U7101 (N_7101,N_7025,N_7075);
or U7102 (N_7102,N_7094,N_7045);
nand U7103 (N_7103,N_7030,N_7013);
xnor U7104 (N_7104,N_7050,N_7082);
and U7105 (N_7105,N_7073,N_7044);
nor U7106 (N_7106,N_7080,N_7038);
nand U7107 (N_7107,N_7079,N_7029);
nor U7108 (N_7108,N_7003,N_7012);
and U7109 (N_7109,N_7043,N_7061);
nor U7110 (N_7110,N_7014,N_7084);
or U7111 (N_7111,N_7034,N_7037);
and U7112 (N_7112,N_7086,N_7048);
nor U7113 (N_7113,N_7058,N_7076);
or U7114 (N_7114,N_7059,N_7054);
and U7115 (N_7115,N_7021,N_7002);
nand U7116 (N_7116,N_7060,N_7085);
nand U7117 (N_7117,N_7062,N_7067);
nor U7118 (N_7118,N_7066,N_7052);
nor U7119 (N_7119,N_7032,N_7091);
and U7120 (N_7120,N_7063,N_7007);
nor U7121 (N_7121,N_7026,N_7078);
nand U7122 (N_7122,N_7024,N_7023);
xnor U7123 (N_7123,N_7020,N_7031);
nand U7124 (N_7124,N_7036,N_7047);
or U7125 (N_7125,N_7088,N_7069);
xor U7126 (N_7126,N_7055,N_7015);
nor U7127 (N_7127,N_7046,N_7017);
nor U7128 (N_7128,N_7099,N_7033);
nor U7129 (N_7129,N_7097,N_7090);
and U7130 (N_7130,N_7089,N_7081);
nand U7131 (N_7131,N_7018,N_7065);
nor U7132 (N_7132,N_7000,N_7006);
nand U7133 (N_7133,N_7016,N_7077);
nor U7134 (N_7134,N_7001,N_7022);
nor U7135 (N_7135,N_7041,N_7083);
and U7136 (N_7136,N_7049,N_7098);
xnor U7137 (N_7137,N_7072,N_7064);
xnor U7138 (N_7138,N_7068,N_7053);
nor U7139 (N_7139,N_7035,N_7096);
nand U7140 (N_7140,N_7074,N_7071);
xnor U7141 (N_7141,N_7005,N_7010);
nor U7142 (N_7142,N_7095,N_7087);
and U7143 (N_7143,N_7093,N_7057);
nand U7144 (N_7144,N_7042,N_7039);
xor U7145 (N_7145,N_7092,N_7011);
nor U7146 (N_7146,N_7019,N_7004);
and U7147 (N_7147,N_7027,N_7056);
and U7148 (N_7148,N_7040,N_7009);
nand U7149 (N_7149,N_7070,N_7051);
or U7150 (N_7150,N_7031,N_7091);
nand U7151 (N_7151,N_7002,N_7095);
or U7152 (N_7152,N_7063,N_7075);
nor U7153 (N_7153,N_7075,N_7086);
nand U7154 (N_7154,N_7084,N_7026);
nor U7155 (N_7155,N_7078,N_7096);
or U7156 (N_7156,N_7074,N_7082);
nand U7157 (N_7157,N_7031,N_7008);
nor U7158 (N_7158,N_7073,N_7091);
nor U7159 (N_7159,N_7047,N_7067);
nor U7160 (N_7160,N_7000,N_7095);
or U7161 (N_7161,N_7046,N_7090);
nand U7162 (N_7162,N_7025,N_7079);
nand U7163 (N_7163,N_7085,N_7023);
nor U7164 (N_7164,N_7004,N_7094);
xor U7165 (N_7165,N_7082,N_7087);
nand U7166 (N_7166,N_7021,N_7027);
nor U7167 (N_7167,N_7035,N_7078);
nand U7168 (N_7168,N_7082,N_7046);
xnor U7169 (N_7169,N_7091,N_7025);
nor U7170 (N_7170,N_7055,N_7083);
or U7171 (N_7171,N_7080,N_7056);
or U7172 (N_7172,N_7013,N_7053);
or U7173 (N_7173,N_7075,N_7049);
nor U7174 (N_7174,N_7058,N_7019);
or U7175 (N_7175,N_7091,N_7043);
or U7176 (N_7176,N_7025,N_7063);
and U7177 (N_7177,N_7061,N_7044);
nand U7178 (N_7178,N_7087,N_7046);
and U7179 (N_7179,N_7040,N_7043);
and U7180 (N_7180,N_7010,N_7038);
nor U7181 (N_7181,N_7071,N_7066);
nand U7182 (N_7182,N_7059,N_7001);
and U7183 (N_7183,N_7053,N_7094);
nor U7184 (N_7184,N_7028,N_7038);
nand U7185 (N_7185,N_7070,N_7025);
or U7186 (N_7186,N_7095,N_7052);
nand U7187 (N_7187,N_7097,N_7046);
or U7188 (N_7188,N_7058,N_7090);
nand U7189 (N_7189,N_7077,N_7021);
or U7190 (N_7190,N_7032,N_7048);
nor U7191 (N_7191,N_7058,N_7078);
nand U7192 (N_7192,N_7027,N_7096);
nand U7193 (N_7193,N_7046,N_7066);
and U7194 (N_7194,N_7028,N_7014);
nor U7195 (N_7195,N_7084,N_7064);
nor U7196 (N_7196,N_7069,N_7037);
nor U7197 (N_7197,N_7032,N_7061);
and U7198 (N_7198,N_7057,N_7013);
and U7199 (N_7199,N_7065,N_7006);
nor U7200 (N_7200,N_7181,N_7171);
and U7201 (N_7201,N_7138,N_7102);
nor U7202 (N_7202,N_7199,N_7169);
nor U7203 (N_7203,N_7185,N_7120);
or U7204 (N_7204,N_7127,N_7198);
xnor U7205 (N_7205,N_7117,N_7148);
nand U7206 (N_7206,N_7136,N_7108);
nand U7207 (N_7207,N_7168,N_7130);
nand U7208 (N_7208,N_7112,N_7144);
or U7209 (N_7209,N_7167,N_7143);
and U7210 (N_7210,N_7128,N_7179);
nand U7211 (N_7211,N_7101,N_7182);
and U7212 (N_7212,N_7170,N_7116);
or U7213 (N_7213,N_7105,N_7135);
nor U7214 (N_7214,N_7115,N_7165);
or U7215 (N_7215,N_7114,N_7146);
or U7216 (N_7216,N_7190,N_7154);
and U7217 (N_7217,N_7149,N_7188);
xnor U7218 (N_7218,N_7109,N_7133);
or U7219 (N_7219,N_7160,N_7129);
nand U7220 (N_7220,N_7172,N_7163);
and U7221 (N_7221,N_7192,N_7174);
and U7222 (N_7222,N_7140,N_7161);
or U7223 (N_7223,N_7113,N_7123);
xnor U7224 (N_7224,N_7141,N_7156);
nor U7225 (N_7225,N_7111,N_7139);
nor U7226 (N_7226,N_7193,N_7106);
or U7227 (N_7227,N_7152,N_7189);
or U7228 (N_7228,N_7159,N_7166);
and U7229 (N_7229,N_7187,N_7178);
nand U7230 (N_7230,N_7175,N_7126);
or U7231 (N_7231,N_7103,N_7158);
nor U7232 (N_7232,N_7176,N_7191);
nor U7233 (N_7233,N_7132,N_7197);
or U7234 (N_7234,N_7150,N_7153);
nor U7235 (N_7235,N_7110,N_7155);
and U7236 (N_7236,N_7184,N_7162);
or U7237 (N_7237,N_7134,N_7121);
nand U7238 (N_7238,N_7151,N_7137);
nand U7239 (N_7239,N_7180,N_7124);
nor U7240 (N_7240,N_7195,N_7122);
xnor U7241 (N_7241,N_7173,N_7104);
and U7242 (N_7242,N_7157,N_7194);
or U7243 (N_7243,N_7196,N_7142);
or U7244 (N_7244,N_7100,N_7118);
and U7245 (N_7245,N_7177,N_7186);
xnor U7246 (N_7246,N_7107,N_7183);
or U7247 (N_7247,N_7145,N_7131);
xor U7248 (N_7248,N_7147,N_7164);
and U7249 (N_7249,N_7119,N_7125);
nand U7250 (N_7250,N_7147,N_7188);
and U7251 (N_7251,N_7194,N_7107);
and U7252 (N_7252,N_7155,N_7112);
nor U7253 (N_7253,N_7184,N_7120);
nor U7254 (N_7254,N_7135,N_7147);
nand U7255 (N_7255,N_7186,N_7112);
and U7256 (N_7256,N_7148,N_7182);
and U7257 (N_7257,N_7116,N_7136);
nand U7258 (N_7258,N_7126,N_7137);
and U7259 (N_7259,N_7120,N_7104);
nand U7260 (N_7260,N_7114,N_7144);
nand U7261 (N_7261,N_7148,N_7186);
nand U7262 (N_7262,N_7103,N_7117);
or U7263 (N_7263,N_7149,N_7178);
and U7264 (N_7264,N_7177,N_7100);
nor U7265 (N_7265,N_7166,N_7106);
nor U7266 (N_7266,N_7148,N_7175);
nor U7267 (N_7267,N_7168,N_7194);
nor U7268 (N_7268,N_7108,N_7127);
nor U7269 (N_7269,N_7182,N_7143);
nor U7270 (N_7270,N_7107,N_7118);
and U7271 (N_7271,N_7109,N_7160);
or U7272 (N_7272,N_7187,N_7119);
nand U7273 (N_7273,N_7133,N_7163);
nor U7274 (N_7274,N_7176,N_7175);
and U7275 (N_7275,N_7159,N_7100);
and U7276 (N_7276,N_7137,N_7161);
nand U7277 (N_7277,N_7189,N_7188);
or U7278 (N_7278,N_7173,N_7123);
nor U7279 (N_7279,N_7192,N_7177);
nor U7280 (N_7280,N_7153,N_7143);
xnor U7281 (N_7281,N_7160,N_7193);
nand U7282 (N_7282,N_7171,N_7128);
xor U7283 (N_7283,N_7139,N_7142);
and U7284 (N_7284,N_7155,N_7118);
nand U7285 (N_7285,N_7132,N_7112);
or U7286 (N_7286,N_7181,N_7183);
and U7287 (N_7287,N_7113,N_7195);
nor U7288 (N_7288,N_7155,N_7124);
and U7289 (N_7289,N_7164,N_7130);
nand U7290 (N_7290,N_7181,N_7144);
and U7291 (N_7291,N_7186,N_7154);
xor U7292 (N_7292,N_7143,N_7109);
nand U7293 (N_7293,N_7178,N_7174);
and U7294 (N_7294,N_7151,N_7153);
or U7295 (N_7295,N_7127,N_7101);
and U7296 (N_7296,N_7187,N_7197);
xnor U7297 (N_7297,N_7185,N_7130);
nand U7298 (N_7298,N_7110,N_7193);
nor U7299 (N_7299,N_7163,N_7181);
and U7300 (N_7300,N_7234,N_7295);
nor U7301 (N_7301,N_7238,N_7253);
xnor U7302 (N_7302,N_7200,N_7248);
nor U7303 (N_7303,N_7288,N_7212);
and U7304 (N_7304,N_7239,N_7289);
nor U7305 (N_7305,N_7259,N_7230);
nor U7306 (N_7306,N_7222,N_7271);
or U7307 (N_7307,N_7270,N_7293);
nand U7308 (N_7308,N_7286,N_7284);
nand U7309 (N_7309,N_7294,N_7243);
or U7310 (N_7310,N_7206,N_7258);
or U7311 (N_7311,N_7240,N_7266);
nand U7312 (N_7312,N_7292,N_7250);
nand U7313 (N_7313,N_7268,N_7201);
nand U7314 (N_7314,N_7287,N_7281);
and U7315 (N_7315,N_7247,N_7299);
or U7316 (N_7316,N_7257,N_7296);
or U7317 (N_7317,N_7209,N_7254);
nand U7318 (N_7318,N_7226,N_7211);
nor U7319 (N_7319,N_7261,N_7231);
and U7320 (N_7320,N_7237,N_7213);
nor U7321 (N_7321,N_7275,N_7262);
or U7322 (N_7322,N_7256,N_7273);
and U7323 (N_7323,N_7251,N_7279);
xnor U7324 (N_7324,N_7214,N_7208);
and U7325 (N_7325,N_7227,N_7219);
and U7326 (N_7326,N_7265,N_7267);
xnor U7327 (N_7327,N_7210,N_7260);
and U7328 (N_7328,N_7205,N_7229);
or U7329 (N_7329,N_7244,N_7221);
nor U7330 (N_7330,N_7235,N_7297);
and U7331 (N_7331,N_7218,N_7216);
or U7332 (N_7332,N_7272,N_7291);
and U7333 (N_7333,N_7277,N_7278);
xor U7334 (N_7334,N_7241,N_7249);
nor U7335 (N_7335,N_7246,N_7220);
nand U7336 (N_7336,N_7263,N_7252);
and U7337 (N_7337,N_7282,N_7285);
and U7338 (N_7338,N_7245,N_7276);
nor U7339 (N_7339,N_7274,N_7280);
and U7340 (N_7340,N_7290,N_7236);
nand U7341 (N_7341,N_7255,N_7264);
and U7342 (N_7342,N_7228,N_7223);
and U7343 (N_7343,N_7224,N_7283);
and U7344 (N_7344,N_7204,N_7269);
nand U7345 (N_7345,N_7232,N_7207);
and U7346 (N_7346,N_7203,N_7225);
and U7347 (N_7347,N_7202,N_7242);
or U7348 (N_7348,N_7298,N_7217);
or U7349 (N_7349,N_7233,N_7215);
nand U7350 (N_7350,N_7279,N_7255);
and U7351 (N_7351,N_7219,N_7279);
and U7352 (N_7352,N_7212,N_7202);
or U7353 (N_7353,N_7215,N_7259);
and U7354 (N_7354,N_7250,N_7296);
xor U7355 (N_7355,N_7231,N_7271);
or U7356 (N_7356,N_7241,N_7233);
or U7357 (N_7357,N_7216,N_7204);
and U7358 (N_7358,N_7298,N_7210);
nor U7359 (N_7359,N_7229,N_7264);
nor U7360 (N_7360,N_7270,N_7209);
xnor U7361 (N_7361,N_7241,N_7217);
and U7362 (N_7362,N_7246,N_7264);
or U7363 (N_7363,N_7247,N_7251);
xnor U7364 (N_7364,N_7256,N_7249);
or U7365 (N_7365,N_7279,N_7224);
nand U7366 (N_7366,N_7265,N_7271);
nand U7367 (N_7367,N_7220,N_7274);
nand U7368 (N_7368,N_7267,N_7258);
xnor U7369 (N_7369,N_7251,N_7263);
nand U7370 (N_7370,N_7274,N_7287);
or U7371 (N_7371,N_7252,N_7288);
nor U7372 (N_7372,N_7223,N_7264);
or U7373 (N_7373,N_7253,N_7284);
or U7374 (N_7374,N_7235,N_7225);
xor U7375 (N_7375,N_7241,N_7268);
xor U7376 (N_7376,N_7257,N_7238);
nand U7377 (N_7377,N_7205,N_7283);
or U7378 (N_7378,N_7262,N_7283);
and U7379 (N_7379,N_7281,N_7232);
nor U7380 (N_7380,N_7273,N_7206);
or U7381 (N_7381,N_7202,N_7265);
and U7382 (N_7382,N_7210,N_7255);
nor U7383 (N_7383,N_7206,N_7209);
nor U7384 (N_7384,N_7268,N_7243);
or U7385 (N_7385,N_7243,N_7229);
nand U7386 (N_7386,N_7202,N_7201);
xor U7387 (N_7387,N_7274,N_7288);
and U7388 (N_7388,N_7200,N_7206);
and U7389 (N_7389,N_7292,N_7235);
nor U7390 (N_7390,N_7225,N_7243);
nor U7391 (N_7391,N_7229,N_7265);
or U7392 (N_7392,N_7217,N_7201);
nor U7393 (N_7393,N_7223,N_7217);
xor U7394 (N_7394,N_7248,N_7254);
or U7395 (N_7395,N_7239,N_7236);
or U7396 (N_7396,N_7283,N_7218);
and U7397 (N_7397,N_7280,N_7293);
and U7398 (N_7398,N_7228,N_7273);
and U7399 (N_7399,N_7259,N_7251);
nand U7400 (N_7400,N_7346,N_7349);
and U7401 (N_7401,N_7393,N_7300);
and U7402 (N_7402,N_7344,N_7358);
nor U7403 (N_7403,N_7312,N_7397);
nor U7404 (N_7404,N_7305,N_7382);
xnor U7405 (N_7405,N_7374,N_7377);
or U7406 (N_7406,N_7335,N_7354);
or U7407 (N_7407,N_7310,N_7304);
or U7408 (N_7408,N_7330,N_7329);
xnor U7409 (N_7409,N_7359,N_7372);
nor U7410 (N_7410,N_7315,N_7367);
xnor U7411 (N_7411,N_7398,N_7353);
xor U7412 (N_7412,N_7301,N_7325);
nor U7413 (N_7413,N_7386,N_7326);
nor U7414 (N_7414,N_7342,N_7340);
nor U7415 (N_7415,N_7396,N_7362);
and U7416 (N_7416,N_7323,N_7373);
xor U7417 (N_7417,N_7316,N_7306);
nand U7418 (N_7418,N_7389,N_7348);
nand U7419 (N_7419,N_7357,N_7395);
and U7420 (N_7420,N_7366,N_7332);
or U7421 (N_7421,N_7363,N_7341);
nor U7422 (N_7422,N_7334,N_7385);
nand U7423 (N_7423,N_7369,N_7364);
nor U7424 (N_7424,N_7392,N_7338);
or U7425 (N_7425,N_7380,N_7322);
nand U7426 (N_7426,N_7317,N_7303);
or U7427 (N_7427,N_7390,N_7352);
xnor U7428 (N_7428,N_7351,N_7319);
xnor U7429 (N_7429,N_7333,N_7324);
and U7430 (N_7430,N_7331,N_7307);
nand U7431 (N_7431,N_7314,N_7378);
and U7432 (N_7432,N_7391,N_7355);
nor U7433 (N_7433,N_7360,N_7350);
or U7434 (N_7434,N_7376,N_7343);
and U7435 (N_7435,N_7361,N_7368);
and U7436 (N_7436,N_7387,N_7347);
and U7437 (N_7437,N_7381,N_7383);
and U7438 (N_7438,N_7356,N_7309);
nor U7439 (N_7439,N_7375,N_7365);
xor U7440 (N_7440,N_7302,N_7379);
nor U7441 (N_7441,N_7336,N_7388);
nor U7442 (N_7442,N_7318,N_7327);
nand U7443 (N_7443,N_7313,N_7320);
nand U7444 (N_7444,N_7337,N_7321);
or U7445 (N_7445,N_7311,N_7339);
nor U7446 (N_7446,N_7399,N_7371);
nand U7447 (N_7447,N_7328,N_7345);
xnor U7448 (N_7448,N_7370,N_7308);
and U7449 (N_7449,N_7394,N_7384);
or U7450 (N_7450,N_7340,N_7382);
nor U7451 (N_7451,N_7387,N_7318);
nand U7452 (N_7452,N_7301,N_7338);
or U7453 (N_7453,N_7332,N_7310);
xnor U7454 (N_7454,N_7372,N_7336);
nor U7455 (N_7455,N_7380,N_7311);
nand U7456 (N_7456,N_7341,N_7376);
and U7457 (N_7457,N_7310,N_7394);
nor U7458 (N_7458,N_7366,N_7328);
and U7459 (N_7459,N_7368,N_7351);
and U7460 (N_7460,N_7382,N_7323);
nand U7461 (N_7461,N_7339,N_7337);
nand U7462 (N_7462,N_7305,N_7398);
nand U7463 (N_7463,N_7368,N_7376);
or U7464 (N_7464,N_7337,N_7335);
xor U7465 (N_7465,N_7348,N_7330);
nor U7466 (N_7466,N_7363,N_7325);
and U7467 (N_7467,N_7309,N_7353);
nor U7468 (N_7468,N_7324,N_7317);
xnor U7469 (N_7469,N_7368,N_7355);
xnor U7470 (N_7470,N_7377,N_7335);
nor U7471 (N_7471,N_7316,N_7305);
xnor U7472 (N_7472,N_7312,N_7365);
and U7473 (N_7473,N_7370,N_7328);
nor U7474 (N_7474,N_7375,N_7305);
nor U7475 (N_7475,N_7304,N_7351);
nand U7476 (N_7476,N_7369,N_7359);
or U7477 (N_7477,N_7303,N_7327);
or U7478 (N_7478,N_7330,N_7336);
or U7479 (N_7479,N_7305,N_7387);
or U7480 (N_7480,N_7384,N_7375);
or U7481 (N_7481,N_7315,N_7347);
or U7482 (N_7482,N_7372,N_7328);
or U7483 (N_7483,N_7339,N_7322);
nor U7484 (N_7484,N_7383,N_7370);
nand U7485 (N_7485,N_7371,N_7353);
and U7486 (N_7486,N_7389,N_7376);
and U7487 (N_7487,N_7364,N_7308);
and U7488 (N_7488,N_7305,N_7385);
nand U7489 (N_7489,N_7361,N_7335);
xnor U7490 (N_7490,N_7326,N_7398);
or U7491 (N_7491,N_7387,N_7370);
xnor U7492 (N_7492,N_7366,N_7320);
nor U7493 (N_7493,N_7304,N_7331);
nor U7494 (N_7494,N_7321,N_7370);
or U7495 (N_7495,N_7302,N_7318);
or U7496 (N_7496,N_7318,N_7346);
nand U7497 (N_7497,N_7361,N_7309);
or U7498 (N_7498,N_7366,N_7364);
or U7499 (N_7499,N_7323,N_7349);
and U7500 (N_7500,N_7471,N_7486);
or U7501 (N_7501,N_7414,N_7485);
or U7502 (N_7502,N_7404,N_7449);
nand U7503 (N_7503,N_7417,N_7427);
or U7504 (N_7504,N_7400,N_7407);
xnor U7505 (N_7505,N_7453,N_7478);
nor U7506 (N_7506,N_7461,N_7422);
and U7507 (N_7507,N_7423,N_7480);
and U7508 (N_7508,N_7476,N_7432);
and U7509 (N_7509,N_7412,N_7466);
or U7510 (N_7510,N_7488,N_7439);
nand U7511 (N_7511,N_7489,N_7415);
nand U7512 (N_7512,N_7413,N_7483);
nand U7513 (N_7513,N_7473,N_7429);
nand U7514 (N_7514,N_7443,N_7438);
and U7515 (N_7515,N_7440,N_7497);
or U7516 (N_7516,N_7482,N_7479);
xnor U7517 (N_7517,N_7465,N_7454);
nand U7518 (N_7518,N_7475,N_7484);
nor U7519 (N_7519,N_7469,N_7499);
nand U7520 (N_7520,N_7464,N_7460);
xor U7521 (N_7521,N_7421,N_7472);
or U7522 (N_7522,N_7444,N_7491);
xor U7523 (N_7523,N_7448,N_7446);
nand U7524 (N_7524,N_7487,N_7434);
or U7525 (N_7525,N_7433,N_7474);
or U7526 (N_7526,N_7492,N_7458);
and U7527 (N_7527,N_7467,N_7463);
xor U7528 (N_7528,N_7428,N_7435);
nand U7529 (N_7529,N_7455,N_7442);
nor U7530 (N_7530,N_7436,N_7403);
and U7531 (N_7531,N_7405,N_7452);
xor U7532 (N_7532,N_7426,N_7418);
nor U7533 (N_7533,N_7470,N_7445);
nand U7534 (N_7534,N_7437,N_7425);
nand U7535 (N_7535,N_7498,N_7457);
nand U7536 (N_7536,N_7459,N_7450);
xnor U7537 (N_7537,N_7409,N_7424);
nand U7538 (N_7538,N_7441,N_7451);
nand U7539 (N_7539,N_7462,N_7419);
or U7540 (N_7540,N_7493,N_7490);
or U7541 (N_7541,N_7406,N_7408);
nand U7542 (N_7542,N_7477,N_7401);
and U7543 (N_7543,N_7495,N_7468);
nor U7544 (N_7544,N_7402,N_7410);
or U7545 (N_7545,N_7420,N_7481);
nor U7546 (N_7546,N_7411,N_7456);
nor U7547 (N_7547,N_7431,N_7447);
and U7548 (N_7548,N_7494,N_7416);
xnor U7549 (N_7549,N_7430,N_7496);
nor U7550 (N_7550,N_7448,N_7417);
nand U7551 (N_7551,N_7491,N_7420);
nor U7552 (N_7552,N_7457,N_7418);
and U7553 (N_7553,N_7424,N_7480);
or U7554 (N_7554,N_7484,N_7441);
nor U7555 (N_7555,N_7477,N_7426);
nand U7556 (N_7556,N_7449,N_7452);
or U7557 (N_7557,N_7466,N_7445);
xnor U7558 (N_7558,N_7429,N_7463);
nand U7559 (N_7559,N_7468,N_7445);
or U7560 (N_7560,N_7470,N_7471);
nor U7561 (N_7561,N_7449,N_7411);
nor U7562 (N_7562,N_7478,N_7483);
or U7563 (N_7563,N_7423,N_7475);
nand U7564 (N_7564,N_7424,N_7489);
and U7565 (N_7565,N_7479,N_7427);
xnor U7566 (N_7566,N_7462,N_7430);
nor U7567 (N_7567,N_7429,N_7443);
nor U7568 (N_7568,N_7418,N_7456);
nor U7569 (N_7569,N_7408,N_7458);
nor U7570 (N_7570,N_7455,N_7410);
nand U7571 (N_7571,N_7410,N_7473);
or U7572 (N_7572,N_7468,N_7400);
or U7573 (N_7573,N_7445,N_7462);
or U7574 (N_7574,N_7417,N_7435);
nand U7575 (N_7575,N_7406,N_7482);
xor U7576 (N_7576,N_7458,N_7424);
xnor U7577 (N_7577,N_7431,N_7422);
or U7578 (N_7578,N_7411,N_7407);
nor U7579 (N_7579,N_7438,N_7419);
or U7580 (N_7580,N_7440,N_7412);
nor U7581 (N_7581,N_7455,N_7430);
nand U7582 (N_7582,N_7468,N_7486);
and U7583 (N_7583,N_7442,N_7440);
nor U7584 (N_7584,N_7441,N_7448);
nor U7585 (N_7585,N_7414,N_7457);
nor U7586 (N_7586,N_7438,N_7420);
and U7587 (N_7587,N_7492,N_7443);
or U7588 (N_7588,N_7425,N_7431);
or U7589 (N_7589,N_7429,N_7413);
nand U7590 (N_7590,N_7466,N_7420);
nor U7591 (N_7591,N_7446,N_7499);
and U7592 (N_7592,N_7486,N_7457);
and U7593 (N_7593,N_7441,N_7463);
or U7594 (N_7594,N_7474,N_7481);
nor U7595 (N_7595,N_7401,N_7468);
or U7596 (N_7596,N_7430,N_7439);
nand U7597 (N_7597,N_7432,N_7477);
and U7598 (N_7598,N_7430,N_7410);
and U7599 (N_7599,N_7446,N_7407);
nor U7600 (N_7600,N_7539,N_7560);
nand U7601 (N_7601,N_7584,N_7525);
nor U7602 (N_7602,N_7587,N_7599);
nor U7603 (N_7603,N_7578,N_7597);
and U7604 (N_7604,N_7582,N_7534);
and U7605 (N_7605,N_7522,N_7570);
nor U7606 (N_7606,N_7524,N_7555);
or U7607 (N_7607,N_7576,N_7501);
nand U7608 (N_7608,N_7523,N_7574);
xnor U7609 (N_7609,N_7579,N_7551);
or U7610 (N_7610,N_7583,N_7530);
xnor U7611 (N_7611,N_7543,N_7589);
nor U7612 (N_7612,N_7598,N_7558);
and U7613 (N_7613,N_7561,N_7503);
xor U7614 (N_7614,N_7519,N_7575);
and U7615 (N_7615,N_7509,N_7580);
or U7616 (N_7616,N_7564,N_7529);
nor U7617 (N_7617,N_7514,N_7557);
nand U7618 (N_7618,N_7553,N_7517);
xnor U7619 (N_7619,N_7565,N_7506);
and U7620 (N_7620,N_7544,N_7556);
nand U7621 (N_7621,N_7549,N_7567);
and U7622 (N_7622,N_7596,N_7581);
or U7623 (N_7623,N_7520,N_7526);
or U7624 (N_7624,N_7577,N_7593);
and U7625 (N_7625,N_7592,N_7508);
nor U7626 (N_7626,N_7535,N_7568);
or U7627 (N_7627,N_7518,N_7541);
xnor U7628 (N_7628,N_7510,N_7516);
and U7629 (N_7629,N_7562,N_7511);
nor U7630 (N_7630,N_7548,N_7528);
nor U7631 (N_7631,N_7566,N_7573);
and U7632 (N_7632,N_7594,N_7500);
nor U7633 (N_7633,N_7527,N_7546);
nor U7634 (N_7634,N_7547,N_7513);
nor U7635 (N_7635,N_7538,N_7502);
nand U7636 (N_7636,N_7505,N_7591);
nand U7637 (N_7637,N_7590,N_7532);
nand U7638 (N_7638,N_7540,N_7533);
or U7639 (N_7639,N_7586,N_7536);
nand U7640 (N_7640,N_7559,N_7595);
nand U7641 (N_7641,N_7572,N_7585);
nor U7642 (N_7642,N_7569,N_7550);
nor U7643 (N_7643,N_7531,N_7563);
and U7644 (N_7644,N_7512,N_7571);
nand U7645 (N_7645,N_7545,N_7554);
nand U7646 (N_7646,N_7552,N_7537);
nor U7647 (N_7647,N_7542,N_7521);
nor U7648 (N_7648,N_7507,N_7515);
nand U7649 (N_7649,N_7588,N_7504);
xor U7650 (N_7650,N_7524,N_7560);
nor U7651 (N_7651,N_7523,N_7559);
nand U7652 (N_7652,N_7517,N_7566);
and U7653 (N_7653,N_7594,N_7556);
or U7654 (N_7654,N_7568,N_7578);
nor U7655 (N_7655,N_7557,N_7569);
nor U7656 (N_7656,N_7551,N_7543);
nand U7657 (N_7657,N_7524,N_7515);
nand U7658 (N_7658,N_7536,N_7549);
nor U7659 (N_7659,N_7519,N_7550);
or U7660 (N_7660,N_7506,N_7588);
or U7661 (N_7661,N_7531,N_7597);
nor U7662 (N_7662,N_7571,N_7536);
nor U7663 (N_7663,N_7573,N_7542);
or U7664 (N_7664,N_7577,N_7514);
xnor U7665 (N_7665,N_7511,N_7565);
nor U7666 (N_7666,N_7553,N_7584);
xor U7667 (N_7667,N_7598,N_7542);
nand U7668 (N_7668,N_7599,N_7561);
nor U7669 (N_7669,N_7519,N_7592);
nand U7670 (N_7670,N_7581,N_7598);
and U7671 (N_7671,N_7588,N_7583);
xor U7672 (N_7672,N_7519,N_7556);
or U7673 (N_7673,N_7534,N_7506);
xor U7674 (N_7674,N_7522,N_7536);
or U7675 (N_7675,N_7518,N_7507);
xor U7676 (N_7676,N_7510,N_7599);
or U7677 (N_7677,N_7500,N_7552);
and U7678 (N_7678,N_7543,N_7549);
nor U7679 (N_7679,N_7536,N_7563);
nand U7680 (N_7680,N_7501,N_7529);
and U7681 (N_7681,N_7501,N_7548);
or U7682 (N_7682,N_7503,N_7507);
nand U7683 (N_7683,N_7552,N_7584);
xor U7684 (N_7684,N_7585,N_7522);
and U7685 (N_7685,N_7566,N_7542);
nor U7686 (N_7686,N_7517,N_7595);
and U7687 (N_7687,N_7501,N_7583);
nor U7688 (N_7688,N_7579,N_7539);
and U7689 (N_7689,N_7518,N_7504);
nor U7690 (N_7690,N_7526,N_7500);
nor U7691 (N_7691,N_7536,N_7533);
nor U7692 (N_7692,N_7552,N_7597);
nor U7693 (N_7693,N_7502,N_7517);
and U7694 (N_7694,N_7582,N_7555);
and U7695 (N_7695,N_7557,N_7583);
or U7696 (N_7696,N_7566,N_7553);
and U7697 (N_7697,N_7587,N_7591);
xnor U7698 (N_7698,N_7502,N_7520);
nand U7699 (N_7699,N_7512,N_7532);
and U7700 (N_7700,N_7646,N_7629);
nand U7701 (N_7701,N_7666,N_7689);
or U7702 (N_7702,N_7640,N_7643);
nand U7703 (N_7703,N_7676,N_7606);
nor U7704 (N_7704,N_7677,N_7697);
or U7705 (N_7705,N_7639,N_7653);
and U7706 (N_7706,N_7616,N_7652);
nand U7707 (N_7707,N_7601,N_7612);
and U7708 (N_7708,N_7656,N_7634);
nand U7709 (N_7709,N_7602,N_7624);
nand U7710 (N_7710,N_7607,N_7663);
nand U7711 (N_7711,N_7665,N_7649);
nor U7712 (N_7712,N_7675,N_7654);
and U7713 (N_7713,N_7690,N_7614);
or U7714 (N_7714,N_7625,N_7678);
xnor U7715 (N_7715,N_7635,N_7645);
nand U7716 (N_7716,N_7620,N_7695);
nor U7717 (N_7717,N_7600,N_7605);
nand U7718 (N_7718,N_7683,N_7685);
nand U7719 (N_7719,N_7642,N_7694);
xor U7720 (N_7720,N_7662,N_7641);
xnor U7721 (N_7721,N_7650,N_7619);
or U7722 (N_7722,N_7687,N_7603);
nor U7723 (N_7723,N_7632,N_7648);
and U7724 (N_7724,N_7658,N_7672);
nand U7725 (N_7725,N_7604,N_7674);
and U7726 (N_7726,N_7644,N_7659);
nor U7727 (N_7727,N_7628,N_7637);
or U7728 (N_7728,N_7626,N_7684);
and U7729 (N_7729,N_7623,N_7613);
and U7730 (N_7730,N_7610,N_7647);
and U7731 (N_7731,N_7673,N_7671);
and U7732 (N_7732,N_7696,N_7655);
nand U7733 (N_7733,N_7638,N_7692);
or U7734 (N_7734,N_7636,N_7617);
xnor U7735 (N_7735,N_7698,N_7679);
or U7736 (N_7736,N_7668,N_7631);
nand U7737 (N_7737,N_7669,N_7630);
xor U7738 (N_7738,N_7699,N_7621);
nor U7739 (N_7739,N_7670,N_7633);
or U7740 (N_7740,N_7615,N_7622);
nand U7741 (N_7741,N_7609,N_7680);
nor U7742 (N_7742,N_7651,N_7660);
nor U7743 (N_7743,N_7691,N_7686);
nand U7744 (N_7744,N_7618,N_7682);
nand U7745 (N_7745,N_7667,N_7661);
and U7746 (N_7746,N_7693,N_7657);
nor U7747 (N_7747,N_7611,N_7608);
or U7748 (N_7748,N_7688,N_7681);
and U7749 (N_7749,N_7627,N_7664);
nor U7750 (N_7750,N_7699,N_7689);
and U7751 (N_7751,N_7607,N_7633);
and U7752 (N_7752,N_7687,N_7667);
or U7753 (N_7753,N_7608,N_7695);
or U7754 (N_7754,N_7665,N_7617);
xnor U7755 (N_7755,N_7681,N_7693);
xor U7756 (N_7756,N_7673,N_7658);
or U7757 (N_7757,N_7690,N_7600);
or U7758 (N_7758,N_7688,N_7628);
nand U7759 (N_7759,N_7651,N_7696);
and U7760 (N_7760,N_7632,N_7644);
nor U7761 (N_7761,N_7648,N_7614);
nand U7762 (N_7762,N_7695,N_7627);
or U7763 (N_7763,N_7627,N_7694);
or U7764 (N_7764,N_7623,N_7621);
nand U7765 (N_7765,N_7659,N_7667);
and U7766 (N_7766,N_7663,N_7678);
nor U7767 (N_7767,N_7603,N_7623);
nor U7768 (N_7768,N_7682,N_7637);
or U7769 (N_7769,N_7634,N_7609);
and U7770 (N_7770,N_7680,N_7614);
xnor U7771 (N_7771,N_7681,N_7611);
and U7772 (N_7772,N_7646,N_7650);
nand U7773 (N_7773,N_7601,N_7655);
and U7774 (N_7774,N_7684,N_7625);
nor U7775 (N_7775,N_7660,N_7678);
and U7776 (N_7776,N_7622,N_7620);
nor U7777 (N_7777,N_7644,N_7609);
xnor U7778 (N_7778,N_7613,N_7667);
and U7779 (N_7779,N_7692,N_7610);
and U7780 (N_7780,N_7666,N_7690);
or U7781 (N_7781,N_7674,N_7627);
nand U7782 (N_7782,N_7693,N_7614);
nand U7783 (N_7783,N_7654,N_7607);
or U7784 (N_7784,N_7657,N_7690);
nand U7785 (N_7785,N_7626,N_7656);
and U7786 (N_7786,N_7606,N_7684);
or U7787 (N_7787,N_7652,N_7630);
xor U7788 (N_7788,N_7637,N_7636);
xnor U7789 (N_7789,N_7639,N_7631);
nor U7790 (N_7790,N_7659,N_7679);
nand U7791 (N_7791,N_7679,N_7661);
and U7792 (N_7792,N_7640,N_7660);
nand U7793 (N_7793,N_7673,N_7649);
or U7794 (N_7794,N_7697,N_7600);
nor U7795 (N_7795,N_7683,N_7612);
or U7796 (N_7796,N_7652,N_7655);
nor U7797 (N_7797,N_7687,N_7617);
nor U7798 (N_7798,N_7636,N_7644);
and U7799 (N_7799,N_7670,N_7650);
nor U7800 (N_7800,N_7726,N_7755);
or U7801 (N_7801,N_7714,N_7701);
xor U7802 (N_7802,N_7749,N_7772);
or U7803 (N_7803,N_7773,N_7710);
or U7804 (N_7804,N_7715,N_7712);
nor U7805 (N_7805,N_7737,N_7708);
or U7806 (N_7806,N_7730,N_7783);
nor U7807 (N_7807,N_7721,N_7763);
nand U7808 (N_7808,N_7787,N_7790);
or U7809 (N_7809,N_7724,N_7762);
nor U7810 (N_7810,N_7704,N_7741);
and U7811 (N_7811,N_7743,N_7778);
xnor U7812 (N_7812,N_7754,N_7742);
or U7813 (N_7813,N_7700,N_7770);
nand U7814 (N_7814,N_7767,N_7748);
xnor U7815 (N_7815,N_7798,N_7738);
or U7816 (N_7816,N_7791,N_7744);
xor U7817 (N_7817,N_7745,N_7761);
nand U7818 (N_7818,N_7792,N_7718);
or U7819 (N_7819,N_7766,N_7747);
nor U7820 (N_7820,N_7784,N_7746);
nand U7821 (N_7821,N_7727,N_7775);
xnor U7822 (N_7822,N_7733,N_7785);
nor U7823 (N_7823,N_7723,N_7765);
or U7824 (N_7824,N_7757,N_7789);
nor U7825 (N_7825,N_7768,N_7706);
and U7826 (N_7826,N_7777,N_7758);
nand U7827 (N_7827,N_7703,N_7702);
nand U7828 (N_7828,N_7799,N_7705);
xnor U7829 (N_7829,N_7797,N_7756);
nor U7830 (N_7830,N_7795,N_7760);
or U7831 (N_7831,N_7728,N_7776);
nor U7832 (N_7832,N_7740,N_7736);
nor U7833 (N_7833,N_7732,N_7774);
xor U7834 (N_7834,N_7750,N_7781);
or U7835 (N_7835,N_7722,N_7725);
and U7836 (N_7836,N_7707,N_7759);
nor U7837 (N_7837,N_7779,N_7717);
nor U7838 (N_7838,N_7751,N_7729);
or U7839 (N_7839,N_7731,N_7716);
nand U7840 (N_7840,N_7753,N_7764);
nand U7841 (N_7841,N_7735,N_7739);
nor U7842 (N_7842,N_7752,N_7713);
nor U7843 (N_7843,N_7771,N_7734);
xor U7844 (N_7844,N_7786,N_7788);
nand U7845 (N_7845,N_7720,N_7709);
nand U7846 (N_7846,N_7780,N_7719);
nor U7847 (N_7847,N_7793,N_7794);
xor U7848 (N_7848,N_7782,N_7711);
nand U7849 (N_7849,N_7796,N_7769);
or U7850 (N_7850,N_7767,N_7740);
nor U7851 (N_7851,N_7761,N_7733);
nand U7852 (N_7852,N_7705,N_7725);
and U7853 (N_7853,N_7740,N_7788);
xnor U7854 (N_7854,N_7740,N_7742);
xor U7855 (N_7855,N_7706,N_7727);
nor U7856 (N_7856,N_7724,N_7760);
and U7857 (N_7857,N_7740,N_7786);
and U7858 (N_7858,N_7797,N_7794);
nand U7859 (N_7859,N_7712,N_7739);
or U7860 (N_7860,N_7792,N_7756);
nand U7861 (N_7861,N_7730,N_7727);
and U7862 (N_7862,N_7737,N_7724);
nor U7863 (N_7863,N_7728,N_7785);
or U7864 (N_7864,N_7792,N_7787);
and U7865 (N_7865,N_7733,N_7788);
nand U7866 (N_7866,N_7743,N_7700);
nor U7867 (N_7867,N_7755,N_7720);
and U7868 (N_7868,N_7719,N_7766);
xnor U7869 (N_7869,N_7763,N_7732);
nor U7870 (N_7870,N_7774,N_7747);
nand U7871 (N_7871,N_7785,N_7771);
or U7872 (N_7872,N_7749,N_7757);
and U7873 (N_7873,N_7795,N_7710);
or U7874 (N_7874,N_7727,N_7783);
and U7875 (N_7875,N_7798,N_7769);
or U7876 (N_7876,N_7751,N_7730);
and U7877 (N_7877,N_7789,N_7793);
nor U7878 (N_7878,N_7749,N_7794);
nand U7879 (N_7879,N_7714,N_7731);
xor U7880 (N_7880,N_7744,N_7714);
nand U7881 (N_7881,N_7747,N_7783);
nand U7882 (N_7882,N_7784,N_7770);
nand U7883 (N_7883,N_7702,N_7743);
or U7884 (N_7884,N_7743,N_7764);
or U7885 (N_7885,N_7739,N_7794);
or U7886 (N_7886,N_7714,N_7792);
and U7887 (N_7887,N_7740,N_7713);
xnor U7888 (N_7888,N_7792,N_7771);
or U7889 (N_7889,N_7794,N_7707);
xnor U7890 (N_7890,N_7791,N_7723);
nor U7891 (N_7891,N_7707,N_7709);
and U7892 (N_7892,N_7705,N_7756);
and U7893 (N_7893,N_7738,N_7716);
xnor U7894 (N_7894,N_7787,N_7732);
xnor U7895 (N_7895,N_7761,N_7771);
nand U7896 (N_7896,N_7743,N_7748);
and U7897 (N_7897,N_7728,N_7726);
nor U7898 (N_7898,N_7780,N_7703);
nor U7899 (N_7899,N_7797,N_7780);
or U7900 (N_7900,N_7861,N_7834);
nand U7901 (N_7901,N_7802,N_7816);
or U7902 (N_7902,N_7850,N_7820);
nor U7903 (N_7903,N_7869,N_7822);
nor U7904 (N_7904,N_7847,N_7866);
or U7905 (N_7905,N_7848,N_7836);
or U7906 (N_7906,N_7823,N_7831);
nand U7907 (N_7907,N_7846,N_7898);
or U7908 (N_7908,N_7843,N_7880);
nand U7909 (N_7909,N_7805,N_7809);
xnor U7910 (N_7910,N_7810,N_7878);
nor U7911 (N_7911,N_7854,N_7873);
or U7912 (N_7912,N_7872,N_7899);
or U7913 (N_7913,N_7807,N_7895);
nand U7914 (N_7914,N_7864,N_7833);
xnor U7915 (N_7915,N_7835,N_7825);
or U7916 (N_7916,N_7859,N_7885);
nand U7917 (N_7917,N_7891,N_7841);
nand U7918 (N_7918,N_7887,N_7881);
xor U7919 (N_7919,N_7804,N_7883);
or U7920 (N_7920,N_7828,N_7829);
nand U7921 (N_7921,N_7840,N_7855);
and U7922 (N_7922,N_7868,N_7875);
or U7923 (N_7923,N_7877,N_7824);
and U7924 (N_7924,N_7842,N_7874);
nand U7925 (N_7925,N_7801,N_7879);
nand U7926 (N_7926,N_7860,N_7892);
xor U7927 (N_7927,N_7871,N_7811);
and U7928 (N_7928,N_7853,N_7890);
or U7929 (N_7929,N_7800,N_7812);
and U7930 (N_7930,N_7827,N_7826);
nand U7931 (N_7931,N_7882,N_7803);
and U7932 (N_7932,N_7806,N_7857);
and U7933 (N_7933,N_7889,N_7870);
xor U7934 (N_7934,N_7830,N_7894);
nor U7935 (N_7935,N_7896,N_7865);
nor U7936 (N_7936,N_7808,N_7851);
or U7937 (N_7937,N_7814,N_7856);
nand U7938 (N_7938,N_7821,N_7838);
and U7939 (N_7939,N_7867,N_7845);
nand U7940 (N_7940,N_7837,N_7817);
or U7941 (N_7941,N_7839,N_7876);
and U7942 (N_7942,N_7863,N_7862);
nand U7943 (N_7943,N_7858,N_7844);
or U7944 (N_7944,N_7819,N_7852);
nand U7945 (N_7945,N_7813,N_7886);
or U7946 (N_7946,N_7897,N_7815);
nand U7947 (N_7947,N_7884,N_7832);
and U7948 (N_7948,N_7818,N_7888);
xor U7949 (N_7949,N_7849,N_7893);
nor U7950 (N_7950,N_7802,N_7833);
or U7951 (N_7951,N_7811,N_7819);
nand U7952 (N_7952,N_7807,N_7828);
or U7953 (N_7953,N_7828,N_7887);
and U7954 (N_7954,N_7879,N_7854);
and U7955 (N_7955,N_7847,N_7886);
nand U7956 (N_7956,N_7850,N_7807);
or U7957 (N_7957,N_7847,N_7818);
and U7958 (N_7958,N_7855,N_7882);
or U7959 (N_7959,N_7817,N_7851);
and U7960 (N_7960,N_7833,N_7899);
and U7961 (N_7961,N_7895,N_7806);
nor U7962 (N_7962,N_7826,N_7836);
nor U7963 (N_7963,N_7827,N_7846);
nand U7964 (N_7964,N_7835,N_7862);
nor U7965 (N_7965,N_7855,N_7831);
or U7966 (N_7966,N_7862,N_7854);
nor U7967 (N_7967,N_7831,N_7842);
or U7968 (N_7968,N_7897,N_7869);
nand U7969 (N_7969,N_7816,N_7889);
nand U7970 (N_7970,N_7899,N_7889);
or U7971 (N_7971,N_7869,N_7817);
nor U7972 (N_7972,N_7880,N_7833);
or U7973 (N_7973,N_7891,N_7837);
nor U7974 (N_7974,N_7822,N_7852);
or U7975 (N_7975,N_7816,N_7852);
nand U7976 (N_7976,N_7812,N_7836);
nand U7977 (N_7977,N_7862,N_7857);
and U7978 (N_7978,N_7857,N_7843);
or U7979 (N_7979,N_7842,N_7807);
nand U7980 (N_7980,N_7813,N_7892);
xor U7981 (N_7981,N_7875,N_7845);
or U7982 (N_7982,N_7863,N_7864);
nand U7983 (N_7983,N_7821,N_7818);
and U7984 (N_7984,N_7826,N_7894);
nand U7985 (N_7985,N_7881,N_7872);
or U7986 (N_7986,N_7851,N_7878);
nand U7987 (N_7987,N_7887,N_7806);
xnor U7988 (N_7988,N_7857,N_7863);
xor U7989 (N_7989,N_7832,N_7878);
nor U7990 (N_7990,N_7852,N_7809);
nand U7991 (N_7991,N_7877,N_7871);
or U7992 (N_7992,N_7826,N_7864);
nand U7993 (N_7993,N_7814,N_7891);
nand U7994 (N_7994,N_7808,N_7828);
or U7995 (N_7995,N_7868,N_7819);
or U7996 (N_7996,N_7805,N_7861);
or U7997 (N_7997,N_7858,N_7800);
nor U7998 (N_7998,N_7889,N_7880);
nor U7999 (N_7999,N_7829,N_7885);
nor U8000 (N_8000,N_7952,N_7984);
nor U8001 (N_8001,N_7937,N_7920);
nand U8002 (N_8002,N_7902,N_7942);
and U8003 (N_8003,N_7948,N_7989);
and U8004 (N_8004,N_7901,N_7986);
xnor U8005 (N_8005,N_7940,N_7968);
and U8006 (N_8006,N_7999,N_7945);
nor U8007 (N_8007,N_7998,N_7979);
xnor U8008 (N_8008,N_7935,N_7947);
and U8009 (N_8009,N_7980,N_7971);
nand U8010 (N_8010,N_7991,N_7927);
nor U8011 (N_8011,N_7904,N_7957);
nor U8012 (N_8012,N_7933,N_7916);
and U8013 (N_8013,N_7954,N_7964);
and U8014 (N_8014,N_7946,N_7930);
or U8015 (N_8015,N_7963,N_7965);
nor U8016 (N_8016,N_7977,N_7978);
and U8017 (N_8017,N_7912,N_7974);
xnor U8018 (N_8018,N_7938,N_7985);
xnor U8019 (N_8019,N_7939,N_7924);
nor U8020 (N_8020,N_7911,N_7909);
and U8021 (N_8021,N_7915,N_7981);
and U8022 (N_8022,N_7982,N_7919);
and U8023 (N_8023,N_7997,N_7914);
nor U8024 (N_8024,N_7926,N_7959);
nor U8025 (N_8025,N_7961,N_7944);
and U8026 (N_8026,N_7956,N_7921);
and U8027 (N_8027,N_7905,N_7962);
nor U8028 (N_8028,N_7922,N_7988);
nand U8029 (N_8029,N_7993,N_7975);
or U8030 (N_8030,N_7929,N_7970);
and U8031 (N_8031,N_7906,N_7925);
nor U8032 (N_8032,N_7917,N_7943);
or U8033 (N_8033,N_7931,N_7967);
xor U8034 (N_8034,N_7941,N_7966);
or U8035 (N_8035,N_7918,N_7950);
and U8036 (N_8036,N_7983,N_7910);
nand U8037 (N_8037,N_7932,N_7953);
nor U8038 (N_8038,N_7913,N_7990);
or U8039 (N_8039,N_7987,N_7955);
xnor U8040 (N_8040,N_7972,N_7996);
nor U8041 (N_8041,N_7936,N_7958);
and U8042 (N_8042,N_7934,N_7995);
and U8043 (N_8043,N_7969,N_7903);
nand U8044 (N_8044,N_7973,N_7960);
and U8045 (N_8045,N_7923,N_7928);
xnor U8046 (N_8046,N_7949,N_7992);
nor U8047 (N_8047,N_7976,N_7907);
xor U8048 (N_8048,N_7994,N_7908);
or U8049 (N_8049,N_7900,N_7951);
nand U8050 (N_8050,N_7926,N_7919);
nor U8051 (N_8051,N_7993,N_7987);
and U8052 (N_8052,N_7979,N_7910);
and U8053 (N_8053,N_7984,N_7911);
and U8054 (N_8054,N_7962,N_7969);
nand U8055 (N_8055,N_7950,N_7910);
and U8056 (N_8056,N_7960,N_7988);
nor U8057 (N_8057,N_7909,N_7966);
and U8058 (N_8058,N_7997,N_7918);
nor U8059 (N_8059,N_7933,N_7967);
or U8060 (N_8060,N_7964,N_7928);
nor U8061 (N_8061,N_7937,N_7955);
nor U8062 (N_8062,N_7976,N_7991);
nand U8063 (N_8063,N_7929,N_7983);
nand U8064 (N_8064,N_7909,N_7953);
or U8065 (N_8065,N_7969,N_7945);
and U8066 (N_8066,N_7928,N_7927);
xor U8067 (N_8067,N_7934,N_7940);
nor U8068 (N_8068,N_7991,N_7912);
nand U8069 (N_8069,N_7990,N_7984);
nor U8070 (N_8070,N_7988,N_7915);
nor U8071 (N_8071,N_7979,N_7964);
or U8072 (N_8072,N_7947,N_7919);
nor U8073 (N_8073,N_7966,N_7944);
nor U8074 (N_8074,N_7974,N_7972);
or U8075 (N_8075,N_7973,N_7961);
nor U8076 (N_8076,N_7959,N_7943);
and U8077 (N_8077,N_7996,N_7933);
nand U8078 (N_8078,N_7974,N_7940);
and U8079 (N_8079,N_7961,N_7918);
nor U8080 (N_8080,N_7950,N_7934);
and U8081 (N_8081,N_7981,N_7959);
and U8082 (N_8082,N_7901,N_7931);
or U8083 (N_8083,N_7900,N_7929);
nor U8084 (N_8084,N_7981,N_7975);
and U8085 (N_8085,N_7963,N_7975);
and U8086 (N_8086,N_7988,N_7977);
nor U8087 (N_8087,N_7974,N_7955);
and U8088 (N_8088,N_7914,N_7928);
nand U8089 (N_8089,N_7925,N_7926);
nor U8090 (N_8090,N_7935,N_7928);
and U8091 (N_8091,N_7937,N_7976);
or U8092 (N_8092,N_7974,N_7950);
nor U8093 (N_8093,N_7956,N_7933);
xor U8094 (N_8094,N_7982,N_7937);
nor U8095 (N_8095,N_7964,N_7907);
nor U8096 (N_8096,N_7938,N_7940);
or U8097 (N_8097,N_7950,N_7984);
nand U8098 (N_8098,N_7930,N_7919);
nand U8099 (N_8099,N_7921,N_7965);
nand U8100 (N_8100,N_8007,N_8046);
nor U8101 (N_8101,N_8079,N_8084);
and U8102 (N_8102,N_8043,N_8042);
or U8103 (N_8103,N_8088,N_8013);
nor U8104 (N_8104,N_8037,N_8064);
and U8105 (N_8105,N_8022,N_8092);
nand U8106 (N_8106,N_8024,N_8067);
nand U8107 (N_8107,N_8026,N_8047);
or U8108 (N_8108,N_8000,N_8020);
or U8109 (N_8109,N_8053,N_8070);
or U8110 (N_8110,N_8089,N_8005);
xor U8111 (N_8111,N_8017,N_8019);
nor U8112 (N_8112,N_8008,N_8069);
and U8113 (N_8113,N_8057,N_8091);
or U8114 (N_8114,N_8058,N_8015);
and U8115 (N_8115,N_8096,N_8031);
nor U8116 (N_8116,N_8074,N_8083);
nand U8117 (N_8117,N_8029,N_8059);
nand U8118 (N_8118,N_8068,N_8023);
and U8119 (N_8119,N_8062,N_8048);
nor U8120 (N_8120,N_8010,N_8061);
nor U8121 (N_8121,N_8054,N_8098);
nand U8122 (N_8122,N_8006,N_8049);
nand U8123 (N_8123,N_8027,N_8063);
nand U8124 (N_8124,N_8094,N_8078);
and U8125 (N_8125,N_8076,N_8009);
and U8126 (N_8126,N_8001,N_8052);
nand U8127 (N_8127,N_8090,N_8075);
or U8128 (N_8128,N_8066,N_8033);
nand U8129 (N_8129,N_8087,N_8097);
xnor U8130 (N_8130,N_8003,N_8093);
xnor U8131 (N_8131,N_8014,N_8086);
or U8132 (N_8132,N_8032,N_8012);
and U8133 (N_8133,N_8081,N_8050);
nor U8134 (N_8134,N_8021,N_8018);
nand U8135 (N_8135,N_8065,N_8071);
or U8136 (N_8136,N_8034,N_8060);
nor U8137 (N_8137,N_8011,N_8002);
or U8138 (N_8138,N_8040,N_8004);
xnor U8139 (N_8139,N_8077,N_8030);
nand U8140 (N_8140,N_8039,N_8055);
xnor U8141 (N_8141,N_8036,N_8025);
and U8142 (N_8142,N_8035,N_8044);
and U8143 (N_8143,N_8028,N_8080);
and U8144 (N_8144,N_8056,N_8072);
nand U8145 (N_8145,N_8095,N_8051);
and U8146 (N_8146,N_8016,N_8082);
xnor U8147 (N_8147,N_8045,N_8073);
or U8148 (N_8148,N_8041,N_8038);
or U8149 (N_8149,N_8099,N_8085);
xnor U8150 (N_8150,N_8077,N_8062);
nor U8151 (N_8151,N_8027,N_8071);
xor U8152 (N_8152,N_8069,N_8059);
nand U8153 (N_8153,N_8043,N_8027);
nand U8154 (N_8154,N_8083,N_8006);
nor U8155 (N_8155,N_8041,N_8021);
nand U8156 (N_8156,N_8078,N_8099);
and U8157 (N_8157,N_8009,N_8082);
nor U8158 (N_8158,N_8021,N_8035);
nor U8159 (N_8159,N_8003,N_8052);
and U8160 (N_8160,N_8024,N_8008);
or U8161 (N_8161,N_8066,N_8030);
nand U8162 (N_8162,N_8094,N_8052);
and U8163 (N_8163,N_8073,N_8026);
nand U8164 (N_8164,N_8005,N_8037);
nor U8165 (N_8165,N_8025,N_8009);
and U8166 (N_8166,N_8036,N_8066);
and U8167 (N_8167,N_8041,N_8091);
xor U8168 (N_8168,N_8078,N_8028);
nor U8169 (N_8169,N_8077,N_8080);
nor U8170 (N_8170,N_8062,N_8019);
and U8171 (N_8171,N_8034,N_8076);
or U8172 (N_8172,N_8044,N_8055);
and U8173 (N_8173,N_8036,N_8060);
or U8174 (N_8174,N_8076,N_8096);
or U8175 (N_8175,N_8057,N_8009);
nor U8176 (N_8176,N_8020,N_8066);
nor U8177 (N_8177,N_8057,N_8089);
nor U8178 (N_8178,N_8079,N_8087);
nand U8179 (N_8179,N_8053,N_8008);
or U8180 (N_8180,N_8020,N_8018);
xor U8181 (N_8181,N_8067,N_8050);
and U8182 (N_8182,N_8036,N_8081);
xnor U8183 (N_8183,N_8033,N_8065);
nor U8184 (N_8184,N_8048,N_8035);
or U8185 (N_8185,N_8090,N_8098);
nor U8186 (N_8186,N_8051,N_8062);
or U8187 (N_8187,N_8039,N_8075);
nor U8188 (N_8188,N_8044,N_8008);
nor U8189 (N_8189,N_8091,N_8088);
nor U8190 (N_8190,N_8095,N_8026);
nor U8191 (N_8191,N_8003,N_8032);
or U8192 (N_8192,N_8061,N_8069);
and U8193 (N_8193,N_8057,N_8014);
nand U8194 (N_8194,N_8070,N_8024);
nor U8195 (N_8195,N_8027,N_8038);
nor U8196 (N_8196,N_8056,N_8045);
nand U8197 (N_8197,N_8026,N_8069);
xor U8198 (N_8198,N_8098,N_8007);
and U8199 (N_8199,N_8006,N_8058);
nor U8200 (N_8200,N_8192,N_8126);
or U8201 (N_8201,N_8152,N_8108);
nand U8202 (N_8202,N_8101,N_8153);
and U8203 (N_8203,N_8155,N_8184);
nor U8204 (N_8204,N_8168,N_8198);
nor U8205 (N_8205,N_8118,N_8119);
nand U8206 (N_8206,N_8161,N_8127);
and U8207 (N_8207,N_8115,N_8160);
nand U8208 (N_8208,N_8129,N_8142);
nor U8209 (N_8209,N_8171,N_8162);
and U8210 (N_8210,N_8185,N_8141);
and U8211 (N_8211,N_8172,N_8116);
xnor U8212 (N_8212,N_8132,N_8159);
and U8213 (N_8213,N_8174,N_8169);
or U8214 (N_8214,N_8110,N_8177);
and U8215 (N_8215,N_8156,N_8187);
and U8216 (N_8216,N_8196,N_8128);
or U8217 (N_8217,N_8191,N_8122);
xor U8218 (N_8218,N_8102,N_8123);
and U8219 (N_8219,N_8113,N_8131);
or U8220 (N_8220,N_8100,N_8107);
nand U8221 (N_8221,N_8181,N_8151);
and U8222 (N_8222,N_8158,N_8165);
nand U8223 (N_8223,N_8133,N_8167);
nor U8224 (N_8224,N_8144,N_8112);
nand U8225 (N_8225,N_8199,N_8189);
and U8226 (N_8226,N_8175,N_8178);
nand U8227 (N_8227,N_8180,N_8170);
and U8228 (N_8228,N_8106,N_8105);
or U8229 (N_8229,N_8173,N_8121);
and U8230 (N_8230,N_8188,N_8164);
xor U8231 (N_8231,N_8117,N_8145);
nor U8232 (N_8232,N_8114,N_8124);
and U8233 (N_8233,N_8140,N_8195);
nand U8234 (N_8234,N_8186,N_8139);
nand U8235 (N_8235,N_8104,N_8193);
and U8236 (N_8236,N_8134,N_8154);
nand U8237 (N_8237,N_8149,N_8138);
or U8238 (N_8238,N_8179,N_8137);
xor U8239 (N_8239,N_8183,N_8148);
and U8240 (N_8240,N_8109,N_8194);
and U8241 (N_8241,N_8147,N_8146);
nand U8242 (N_8242,N_8130,N_8150);
or U8243 (N_8243,N_8176,N_8111);
nor U8244 (N_8244,N_8197,N_8166);
nand U8245 (N_8245,N_8157,N_8163);
nor U8246 (N_8246,N_8136,N_8182);
or U8247 (N_8247,N_8143,N_8125);
nor U8248 (N_8248,N_8120,N_8190);
nand U8249 (N_8249,N_8103,N_8135);
nand U8250 (N_8250,N_8134,N_8117);
and U8251 (N_8251,N_8143,N_8180);
xor U8252 (N_8252,N_8175,N_8189);
xnor U8253 (N_8253,N_8177,N_8199);
nand U8254 (N_8254,N_8134,N_8161);
nor U8255 (N_8255,N_8194,N_8158);
and U8256 (N_8256,N_8193,N_8179);
nand U8257 (N_8257,N_8192,N_8133);
or U8258 (N_8258,N_8145,N_8176);
nor U8259 (N_8259,N_8187,N_8126);
or U8260 (N_8260,N_8136,N_8126);
nor U8261 (N_8261,N_8134,N_8121);
nand U8262 (N_8262,N_8165,N_8178);
and U8263 (N_8263,N_8174,N_8121);
and U8264 (N_8264,N_8113,N_8182);
and U8265 (N_8265,N_8113,N_8186);
nor U8266 (N_8266,N_8178,N_8102);
nand U8267 (N_8267,N_8157,N_8147);
and U8268 (N_8268,N_8161,N_8114);
and U8269 (N_8269,N_8183,N_8115);
or U8270 (N_8270,N_8104,N_8111);
and U8271 (N_8271,N_8158,N_8109);
nand U8272 (N_8272,N_8111,N_8177);
or U8273 (N_8273,N_8133,N_8145);
and U8274 (N_8274,N_8155,N_8105);
nor U8275 (N_8275,N_8118,N_8140);
nand U8276 (N_8276,N_8120,N_8114);
and U8277 (N_8277,N_8191,N_8142);
nor U8278 (N_8278,N_8114,N_8185);
nand U8279 (N_8279,N_8112,N_8129);
or U8280 (N_8280,N_8121,N_8101);
nand U8281 (N_8281,N_8163,N_8126);
or U8282 (N_8282,N_8113,N_8141);
xnor U8283 (N_8283,N_8140,N_8110);
or U8284 (N_8284,N_8145,N_8164);
xnor U8285 (N_8285,N_8173,N_8191);
or U8286 (N_8286,N_8153,N_8103);
and U8287 (N_8287,N_8117,N_8110);
nand U8288 (N_8288,N_8145,N_8124);
nor U8289 (N_8289,N_8115,N_8192);
nand U8290 (N_8290,N_8173,N_8169);
nand U8291 (N_8291,N_8177,N_8139);
nor U8292 (N_8292,N_8163,N_8189);
nor U8293 (N_8293,N_8155,N_8149);
nand U8294 (N_8294,N_8191,N_8134);
and U8295 (N_8295,N_8100,N_8157);
and U8296 (N_8296,N_8151,N_8130);
and U8297 (N_8297,N_8160,N_8179);
and U8298 (N_8298,N_8183,N_8118);
nand U8299 (N_8299,N_8169,N_8155);
nand U8300 (N_8300,N_8225,N_8224);
xnor U8301 (N_8301,N_8222,N_8292);
nor U8302 (N_8302,N_8206,N_8205);
and U8303 (N_8303,N_8231,N_8277);
or U8304 (N_8304,N_8212,N_8243);
xor U8305 (N_8305,N_8207,N_8271);
nand U8306 (N_8306,N_8215,N_8202);
nor U8307 (N_8307,N_8294,N_8252);
and U8308 (N_8308,N_8286,N_8265);
nor U8309 (N_8309,N_8299,N_8240);
and U8310 (N_8310,N_8213,N_8236);
nand U8311 (N_8311,N_8208,N_8250);
or U8312 (N_8312,N_8278,N_8264);
and U8313 (N_8313,N_8296,N_8219);
nand U8314 (N_8314,N_8221,N_8217);
nor U8315 (N_8315,N_8248,N_8262);
nand U8316 (N_8316,N_8238,N_8256);
nand U8317 (N_8317,N_8283,N_8298);
or U8318 (N_8318,N_8239,N_8209);
nand U8319 (N_8319,N_8263,N_8241);
nand U8320 (N_8320,N_8266,N_8251);
or U8321 (N_8321,N_8290,N_8285);
or U8322 (N_8322,N_8279,N_8280);
or U8323 (N_8323,N_8200,N_8274);
and U8324 (N_8324,N_8249,N_8273);
nor U8325 (N_8325,N_8247,N_8242);
nand U8326 (N_8326,N_8218,N_8201);
nand U8327 (N_8327,N_8293,N_8275);
nor U8328 (N_8328,N_8258,N_8244);
and U8329 (N_8329,N_8287,N_8226);
and U8330 (N_8330,N_8269,N_8253);
or U8331 (N_8331,N_8204,N_8237);
or U8332 (N_8332,N_8284,N_8255);
nand U8333 (N_8333,N_8295,N_8214);
nor U8334 (N_8334,N_8230,N_8228);
or U8335 (N_8335,N_8289,N_8234);
nor U8336 (N_8336,N_8267,N_8297);
and U8337 (N_8337,N_8227,N_8254);
and U8338 (N_8338,N_8216,N_8261);
and U8339 (N_8339,N_8246,N_8272);
xor U8340 (N_8340,N_8259,N_8233);
xor U8341 (N_8341,N_8291,N_8211);
xnor U8342 (N_8342,N_8229,N_8268);
xnor U8343 (N_8343,N_8232,N_8210);
nand U8344 (N_8344,N_8257,N_8282);
nand U8345 (N_8345,N_8281,N_8270);
or U8346 (N_8346,N_8288,N_8223);
or U8347 (N_8347,N_8276,N_8245);
or U8348 (N_8348,N_8260,N_8203);
nor U8349 (N_8349,N_8220,N_8235);
nor U8350 (N_8350,N_8279,N_8256);
nand U8351 (N_8351,N_8277,N_8220);
and U8352 (N_8352,N_8233,N_8242);
nor U8353 (N_8353,N_8266,N_8205);
nor U8354 (N_8354,N_8284,N_8245);
and U8355 (N_8355,N_8243,N_8214);
nor U8356 (N_8356,N_8253,N_8250);
or U8357 (N_8357,N_8243,N_8251);
and U8358 (N_8358,N_8267,N_8251);
nand U8359 (N_8359,N_8265,N_8282);
nor U8360 (N_8360,N_8266,N_8238);
nor U8361 (N_8361,N_8237,N_8292);
xor U8362 (N_8362,N_8204,N_8216);
and U8363 (N_8363,N_8219,N_8243);
and U8364 (N_8364,N_8210,N_8297);
and U8365 (N_8365,N_8213,N_8261);
nor U8366 (N_8366,N_8254,N_8247);
nand U8367 (N_8367,N_8297,N_8237);
and U8368 (N_8368,N_8242,N_8252);
or U8369 (N_8369,N_8232,N_8271);
or U8370 (N_8370,N_8282,N_8280);
or U8371 (N_8371,N_8226,N_8273);
nand U8372 (N_8372,N_8235,N_8268);
and U8373 (N_8373,N_8225,N_8252);
and U8374 (N_8374,N_8267,N_8260);
nand U8375 (N_8375,N_8274,N_8265);
nand U8376 (N_8376,N_8222,N_8286);
nand U8377 (N_8377,N_8264,N_8231);
nand U8378 (N_8378,N_8200,N_8273);
nand U8379 (N_8379,N_8291,N_8267);
and U8380 (N_8380,N_8246,N_8222);
nand U8381 (N_8381,N_8295,N_8252);
and U8382 (N_8382,N_8219,N_8201);
xnor U8383 (N_8383,N_8289,N_8207);
and U8384 (N_8384,N_8213,N_8249);
nor U8385 (N_8385,N_8279,N_8261);
and U8386 (N_8386,N_8206,N_8275);
or U8387 (N_8387,N_8200,N_8275);
or U8388 (N_8388,N_8228,N_8219);
or U8389 (N_8389,N_8200,N_8292);
xnor U8390 (N_8390,N_8255,N_8259);
or U8391 (N_8391,N_8219,N_8209);
or U8392 (N_8392,N_8232,N_8256);
nor U8393 (N_8393,N_8268,N_8289);
or U8394 (N_8394,N_8228,N_8286);
nor U8395 (N_8395,N_8262,N_8258);
and U8396 (N_8396,N_8272,N_8230);
nor U8397 (N_8397,N_8291,N_8284);
and U8398 (N_8398,N_8217,N_8226);
nand U8399 (N_8399,N_8255,N_8245);
and U8400 (N_8400,N_8328,N_8301);
and U8401 (N_8401,N_8309,N_8321);
nand U8402 (N_8402,N_8354,N_8361);
or U8403 (N_8403,N_8329,N_8338);
nand U8404 (N_8404,N_8377,N_8394);
nor U8405 (N_8405,N_8306,N_8355);
and U8406 (N_8406,N_8332,N_8366);
and U8407 (N_8407,N_8388,N_8305);
nand U8408 (N_8408,N_8390,N_8304);
and U8409 (N_8409,N_8356,N_8324);
nand U8410 (N_8410,N_8308,N_8364);
and U8411 (N_8411,N_8399,N_8345);
or U8412 (N_8412,N_8363,N_8373);
nor U8413 (N_8413,N_8351,N_8331);
or U8414 (N_8414,N_8311,N_8319);
and U8415 (N_8415,N_8317,N_8362);
nor U8416 (N_8416,N_8387,N_8349);
or U8417 (N_8417,N_8303,N_8320);
or U8418 (N_8418,N_8312,N_8313);
nand U8419 (N_8419,N_8371,N_8344);
or U8420 (N_8420,N_8360,N_8310);
nor U8421 (N_8421,N_8392,N_8381);
nor U8422 (N_8422,N_8322,N_8323);
or U8423 (N_8423,N_8342,N_8396);
nand U8424 (N_8424,N_8382,N_8359);
and U8425 (N_8425,N_8340,N_8358);
and U8426 (N_8426,N_8343,N_8302);
xnor U8427 (N_8427,N_8380,N_8389);
nand U8428 (N_8428,N_8352,N_8325);
nand U8429 (N_8429,N_8333,N_8353);
or U8430 (N_8430,N_8346,N_8386);
or U8431 (N_8431,N_8385,N_8327);
or U8432 (N_8432,N_8347,N_8336);
nand U8433 (N_8433,N_8307,N_8395);
or U8434 (N_8434,N_8367,N_8339);
or U8435 (N_8435,N_8383,N_8393);
or U8436 (N_8436,N_8376,N_8397);
and U8437 (N_8437,N_8314,N_8372);
nor U8438 (N_8438,N_8398,N_8300);
and U8439 (N_8439,N_8334,N_8370);
or U8440 (N_8440,N_8326,N_8316);
xnor U8441 (N_8441,N_8318,N_8315);
or U8442 (N_8442,N_8391,N_8335);
nor U8443 (N_8443,N_8374,N_8330);
nor U8444 (N_8444,N_8369,N_8379);
nor U8445 (N_8445,N_8378,N_8365);
or U8446 (N_8446,N_8341,N_8384);
and U8447 (N_8447,N_8357,N_8337);
nor U8448 (N_8448,N_8350,N_8348);
or U8449 (N_8449,N_8368,N_8375);
and U8450 (N_8450,N_8387,N_8344);
nor U8451 (N_8451,N_8399,N_8358);
nand U8452 (N_8452,N_8321,N_8351);
nor U8453 (N_8453,N_8311,N_8307);
or U8454 (N_8454,N_8369,N_8376);
or U8455 (N_8455,N_8338,N_8326);
or U8456 (N_8456,N_8333,N_8301);
or U8457 (N_8457,N_8359,N_8367);
nor U8458 (N_8458,N_8310,N_8352);
or U8459 (N_8459,N_8330,N_8354);
and U8460 (N_8460,N_8365,N_8396);
or U8461 (N_8461,N_8379,N_8389);
nor U8462 (N_8462,N_8363,N_8359);
or U8463 (N_8463,N_8395,N_8308);
nand U8464 (N_8464,N_8348,N_8369);
or U8465 (N_8465,N_8319,N_8365);
or U8466 (N_8466,N_8374,N_8311);
and U8467 (N_8467,N_8329,N_8303);
and U8468 (N_8468,N_8362,N_8351);
nand U8469 (N_8469,N_8336,N_8304);
or U8470 (N_8470,N_8345,N_8325);
and U8471 (N_8471,N_8346,N_8348);
nor U8472 (N_8472,N_8356,N_8336);
nor U8473 (N_8473,N_8322,N_8381);
xor U8474 (N_8474,N_8324,N_8361);
nor U8475 (N_8475,N_8384,N_8379);
and U8476 (N_8476,N_8392,N_8312);
xnor U8477 (N_8477,N_8397,N_8317);
and U8478 (N_8478,N_8304,N_8381);
xnor U8479 (N_8479,N_8336,N_8300);
nor U8480 (N_8480,N_8370,N_8328);
and U8481 (N_8481,N_8355,N_8327);
and U8482 (N_8482,N_8316,N_8370);
nor U8483 (N_8483,N_8317,N_8381);
nand U8484 (N_8484,N_8354,N_8367);
and U8485 (N_8485,N_8336,N_8331);
nand U8486 (N_8486,N_8306,N_8376);
and U8487 (N_8487,N_8320,N_8375);
nand U8488 (N_8488,N_8389,N_8304);
and U8489 (N_8489,N_8357,N_8377);
nand U8490 (N_8490,N_8347,N_8388);
or U8491 (N_8491,N_8309,N_8376);
nor U8492 (N_8492,N_8388,N_8385);
nand U8493 (N_8493,N_8350,N_8362);
nor U8494 (N_8494,N_8350,N_8369);
nor U8495 (N_8495,N_8381,N_8393);
nor U8496 (N_8496,N_8316,N_8365);
xnor U8497 (N_8497,N_8335,N_8352);
and U8498 (N_8498,N_8352,N_8368);
or U8499 (N_8499,N_8309,N_8384);
nand U8500 (N_8500,N_8497,N_8478);
nand U8501 (N_8501,N_8433,N_8437);
xor U8502 (N_8502,N_8457,N_8406);
xor U8503 (N_8503,N_8498,N_8450);
nand U8504 (N_8504,N_8487,N_8464);
nor U8505 (N_8505,N_8456,N_8455);
or U8506 (N_8506,N_8407,N_8440);
or U8507 (N_8507,N_8405,N_8494);
and U8508 (N_8508,N_8454,N_8479);
and U8509 (N_8509,N_8473,N_8428);
nor U8510 (N_8510,N_8417,N_8400);
nor U8511 (N_8511,N_8490,N_8442);
nand U8512 (N_8512,N_8410,N_8480);
and U8513 (N_8513,N_8481,N_8409);
or U8514 (N_8514,N_8418,N_8416);
and U8515 (N_8515,N_8436,N_8491);
or U8516 (N_8516,N_8439,N_8484);
nand U8517 (N_8517,N_8447,N_8415);
nand U8518 (N_8518,N_8486,N_8458);
nand U8519 (N_8519,N_8476,N_8424);
nand U8520 (N_8520,N_8493,N_8492);
or U8521 (N_8521,N_8448,N_8445);
nand U8522 (N_8522,N_8488,N_8438);
nand U8523 (N_8523,N_8462,N_8443);
xnor U8524 (N_8524,N_8441,N_8470);
xnor U8525 (N_8525,N_8496,N_8475);
and U8526 (N_8526,N_8423,N_8446);
nand U8527 (N_8527,N_8422,N_8465);
nor U8528 (N_8528,N_8474,N_8477);
and U8529 (N_8529,N_8435,N_8430);
or U8530 (N_8530,N_8420,N_8467);
xor U8531 (N_8531,N_8472,N_8463);
and U8532 (N_8532,N_8434,N_8469);
nor U8533 (N_8533,N_8461,N_8468);
nor U8534 (N_8534,N_8431,N_8444);
and U8535 (N_8535,N_8412,N_8408);
or U8536 (N_8536,N_8452,N_8427);
and U8537 (N_8537,N_8432,N_8471);
or U8538 (N_8538,N_8401,N_8426);
nand U8539 (N_8539,N_8499,N_8425);
nand U8540 (N_8540,N_8404,N_8459);
nand U8541 (N_8541,N_8460,N_8466);
xor U8542 (N_8542,N_8453,N_8414);
and U8543 (N_8543,N_8485,N_8483);
nand U8544 (N_8544,N_8421,N_8489);
nand U8545 (N_8545,N_8402,N_8403);
nor U8546 (N_8546,N_8411,N_8482);
nand U8547 (N_8547,N_8449,N_8451);
and U8548 (N_8548,N_8419,N_8429);
or U8549 (N_8549,N_8495,N_8413);
or U8550 (N_8550,N_8425,N_8417);
or U8551 (N_8551,N_8450,N_8442);
or U8552 (N_8552,N_8422,N_8424);
nor U8553 (N_8553,N_8435,N_8473);
and U8554 (N_8554,N_8482,N_8450);
or U8555 (N_8555,N_8497,N_8435);
nand U8556 (N_8556,N_8427,N_8451);
or U8557 (N_8557,N_8452,N_8494);
and U8558 (N_8558,N_8465,N_8495);
and U8559 (N_8559,N_8415,N_8475);
nand U8560 (N_8560,N_8453,N_8435);
and U8561 (N_8561,N_8434,N_8441);
nor U8562 (N_8562,N_8497,N_8483);
nor U8563 (N_8563,N_8434,N_8444);
and U8564 (N_8564,N_8456,N_8458);
or U8565 (N_8565,N_8418,N_8472);
or U8566 (N_8566,N_8494,N_8498);
or U8567 (N_8567,N_8445,N_8464);
nor U8568 (N_8568,N_8451,N_8461);
or U8569 (N_8569,N_8408,N_8462);
nand U8570 (N_8570,N_8491,N_8425);
nor U8571 (N_8571,N_8463,N_8404);
nor U8572 (N_8572,N_8486,N_8449);
or U8573 (N_8573,N_8428,N_8421);
xnor U8574 (N_8574,N_8470,N_8452);
and U8575 (N_8575,N_8485,N_8400);
nand U8576 (N_8576,N_8413,N_8494);
nand U8577 (N_8577,N_8443,N_8453);
and U8578 (N_8578,N_8463,N_8473);
nor U8579 (N_8579,N_8412,N_8446);
nand U8580 (N_8580,N_8469,N_8497);
and U8581 (N_8581,N_8478,N_8484);
xnor U8582 (N_8582,N_8498,N_8445);
nor U8583 (N_8583,N_8436,N_8470);
nor U8584 (N_8584,N_8409,N_8422);
xnor U8585 (N_8585,N_8408,N_8447);
or U8586 (N_8586,N_8414,N_8424);
nand U8587 (N_8587,N_8496,N_8419);
xor U8588 (N_8588,N_8495,N_8416);
nand U8589 (N_8589,N_8491,N_8499);
nor U8590 (N_8590,N_8400,N_8420);
and U8591 (N_8591,N_8445,N_8463);
nand U8592 (N_8592,N_8463,N_8405);
and U8593 (N_8593,N_8472,N_8454);
nand U8594 (N_8594,N_8488,N_8415);
nand U8595 (N_8595,N_8420,N_8405);
nor U8596 (N_8596,N_8438,N_8411);
nand U8597 (N_8597,N_8449,N_8492);
nor U8598 (N_8598,N_8430,N_8409);
or U8599 (N_8599,N_8473,N_8446);
nand U8600 (N_8600,N_8505,N_8592);
nand U8601 (N_8601,N_8532,N_8515);
or U8602 (N_8602,N_8590,N_8583);
xnor U8603 (N_8603,N_8543,N_8513);
xor U8604 (N_8604,N_8584,N_8569);
and U8605 (N_8605,N_8525,N_8550);
or U8606 (N_8606,N_8599,N_8574);
xor U8607 (N_8607,N_8597,N_8549);
nand U8608 (N_8608,N_8510,N_8572);
or U8609 (N_8609,N_8500,N_8552);
or U8610 (N_8610,N_8524,N_8537);
xnor U8611 (N_8611,N_8531,N_8553);
and U8612 (N_8612,N_8521,N_8534);
and U8613 (N_8613,N_8581,N_8563);
nor U8614 (N_8614,N_8507,N_8544);
and U8615 (N_8615,N_8579,N_8506);
nand U8616 (N_8616,N_8539,N_8588);
nand U8617 (N_8617,N_8547,N_8522);
and U8618 (N_8618,N_8591,N_8512);
nor U8619 (N_8619,N_8554,N_8538);
xnor U8620 (N_8620,N_8567,N_8586);
and U8621 (N_8621,N_8551,N_8565);
nand U8622 (N_8622,N_8557,N_8523);
or U8623 (N_8623,N_8566,N_8529);
and U8624 (N_8624,N_8502,N_8578);
nand U8625 (N_8625,N_8540,N_8535);
nand U8626 (N_8626,N_8514,N_8585);
nor U8627 (N_8627,N_8501,N_8541);
or U8628 (N_8628,N_8589,N_8561);
or U8629 (N_8629,N_8517,N_8577);
nor U8630 (N_8630,N_8536,N_8573);
xnor U8631 (N_8631,N_8555,N_8568);
nand U8632 (N_8632,N_8526,N_8508);
xor U8633 (N_8633,N_8575,N_8559);
or U8634 (N_8634,N_8504,N_8598);
or U8635 (N_8635,N_8560,N_8520);
nand U8636 (N_8636,N_8582,N_8503);
or U8637 (N_8637,N_8570,N_8527);
nand U8638 (N_8638,N_8518,N_8546);
nand U8639 (N_8639,N_8571,N_8548);
and U8640 (N_8640,N_8596,N_8528);
nand U8641 (N_8641,N_8530,N_8509);
and U8642 (N_8642,N_8587,N_8564);
nand U8643 (N_8643,N_8542,N_8516);
and U8644 (N_8644,N_8558,N_8545);
nand U8645 (N_8645,N_8594,N_8576);
nor U8646 (N_8646,N_8519,N_8595);
or U8647 (N_8647,N_8511,N_8580);
and U8648 (N_8648,N_8533,N_8556);
nor U8649 (N_8649,N_8562,N_8593);
or U8650 (N_8650,N_8528,N_8506);
or U8651 (N_8651,N_8508,N_8524);
or U8652 (N_8652,N_8508,N_8570);
and U8653 (N_8653,N_8587,N_8598);
nor U8654 (N_8654,N_8556,N_8590);
or U8655 (N_8655,N_8530,N_8515);
nor U8656 (N_8656,N_8556,N_8592);
nor U8657 (N_8657,N_8586,N_8561);
and U8658 (N_8658,N_8593,N_8597);
or U8659 (N_8659,N_8506,N_8543);
and U8660 (N_8660,N_8560,N_8524);
xor U8661 (N_8661,N_8503,N_8518);
or U8662 (N_8662,N_8585,N_8509);
nand U8663 (N_8663,N_8561,N_8563);
xor U8664 (N_8664,N_8501,N_8581);
nor U8665 (N_8665,N_8541,N_8532);
and U8666 (N_8666,N_8544,N_8567);
and U8667 (N_8667,N_8584,N_8574);
nand U8668 (N_8668,N_8558,N_8562);
or U8669 (N_8669,N_8533,N_8574);
or U8670 (N_8670,N_8593,N_8511);
nand U8671 (N_8671,N_8562,N_8525);
or U8672 (N_8672,N_8532,N_8517);
nand U8673 (N_8673,N_8557,N_8594);
nand U8674 (N_8674,N_8531,N_8510);
and U8675 (N_8675,N_8522,N_8501);
and U8676 (N_8676,N_8591,N_8527);
nor U8677 (N_8677,N_8587,N_8560);
or U8678 (N_8678,N_8581,N_8580);
xor U8679 (N_8679,N_8538,N_8586);
and U8680 (N_8680,N_8506,N_8522);
and U8681 (N_8681,N_8551,N_8518);
or U8682 (N_8682,N_8563,N_8584);
and U8683 (N_8683,N_8575,N_8592);
or U8684 (N_8684,N_8504,N_8546);
or U8685 (N_8685,N_8585,N_8552);
nand U8686 (N_8686,N_8554,N_8536);
or U8687 (N_8687,N_8555,N_8564);
and U8688 (N_8688,N_8592,N_8535);
or U8689 (N_8689,N_8571,N_8514);
and U8690 (N_8690,N_8510,N_8594);
nand U8691 (N_8691,N_8523,N_8521);
or U8692 (N_8692,N_8540,N_8503);
nand U8693 (N_8693,N_8549,N_8577);
nand U8694 (N_8694,N_8555,N_8507);
nand U8695 (N_8695,N_8599,N_8542);
nor U8696 (N_8696,N_8540,N_8580);
nor U8697 (N_8697,N_8508,N_8597);
or U8698 (N_8698,N_8541,N_8518);
nor U8699 (N_8699,N_8564,N_8530);
or U8700 (N_8700,N_8610,N_8654);
and U8701 (N_8701,N_8622,N_8618);
nand U8702 (N_8702,N_8609,N_8650);
and U8703 (N_8703,N_8644,N_8660);
and U8704 (N_8704,N_8630,N_8670);
nand U8705 (N_8705,N_8646,N_8689);
nor U8706 (N_8706,N_8664,N_8603);
nand U8707 (N_8707,N_8645,N_8693);
or U8708 (N_8708,N_8671,N_8686);
nand U8709 (N_8709,N_8631,N_8651);
and U8710 (N_8710,N_8649,N_8697);
nor U8711 (N_8711,N_8612,N_8659);
nor U8712 (N_8712,N_8602,N_8632);
and U8713 (N_8713,N_8696,N_8617);
and U8714 (N_8714,N_8685,N_8698);
and U8715 (N_8715,N_8613,N_8667);
nand U8716 (N_8716,N_8604,N_8624);
and U8717 (N_8717,N_8680,N_8611);
nor U8718 (N_8718,N_8626,N_8691);
nor U8719 (N_8719,N_8669,N_8681);
or U8720 (N_8720,N_8627,N_8661);
or U8721 (N_8721,N_8658,N_8665);
nor U8722 (N_8722,N_8687,N_8699);
nand U8723 (N_8723,N_8642,N_8621);
xor U8724 (N_8724,N_8655,N_8676);
or U8725 (N_8725,N_8688,N_8607);
nor U8726 (N_8726,N_8690,N_8633);
nor U8727 (N_8727,N_8694,N_8648);
or U8728 (N_8728,N_8637,N_8636);
nor U8729 (N_8729,N_8619,N_8616);
and U8730 (N_8730,N_8666,N_8640);
and U8731 (N_8731,N_8601,N_8653);
and U8732 (N_8732,N_8656,N_8641);
nand U8733 (N_8733,N_8639,N_8673);
nand U8734 (N_8734,N_8692,N_8635);
or U8735 (N_8735,N_8620,N_8623);
nand U8736 (N_8736,N_8679,N_8675);
nor U8737 (N_8737,N_8643,N_8672);
nor U8738 (N_8738,N_8605,N_8668);
and U8739 (N_8739,N_8614,N_8683);
and U8740 (N_8740,N_8606,N_8600);
or U8741 (N_8741,N_8657,N_8629);
nor U8742 (N_8742,N_8628,N_8608);
and U8743 (N_8743,N_8615,N_8682);
or U8744 (N_8744,N_8674,N_8638);
and U8745 (N_8745,N_8678,N_8684);
nand U8746 (N_8746,N_8695,N_8625);
nand U8747 (N_8747,N_8662,N_8677);
and U8748 (N_8748,N_8634,N_8663);
nor U8749 (N_8749,N_8647,N_8652);
or U8750 (N_8750,N_8627,N_8640);
and U8751 (N_8751,N_8614,N_8681);
nand U8752 (N_8752,N_8684,N_8633);
nor U8753 (N_8753,N_8628,N_8638);
xor U8754 (N_8754,N_8644,N_8618);
and U8755 (N_8755,N_8688,N_8670);
and U8756 (N_8756,N_8652,N_8615);
and U8757 (N_8757,N_8621,N_8695);
nor U8758 (N_8758,N_8684,N_8676);
and U8759 (N_8759,N_8653,N_8628);
nand U8760 (N_8760,N_8673,N_8649);
and U8761 (N_8761,N_8668,N_8689);
or U8762 (N_8762,N_8608,N_8670);
nor U8763 (N_8763,N_8629,N_8614);
and U8764 (N_8764,N_8618,N_8603);
and U8765 (N_8765,N_8676,N_8629);
nor U8766 (N_8766,N_8604,N_8692);
xor U8767 (N_8767,N_8622,N_8617);
nor U8768 (N_8768,N_8659,N_8663);
and U8769 (N_8769,N_8618,N_8692);
and U8770 (N_8770,N_8603,N_8627);
and U8771 (N_8771,N_8689,N_8678);
nand U8772 (N_8772,N_8640,N_8619);
nor U8773 (N_8773,N_8622,N_8696);
and U8774 (N_8774,N_8648,N_8675);
xor U8775 (N_8775,N_8674,N_8671);
nand U8776 (N_8776,N_8695,N_8663);
and U8777 (N_8777,N_8666,N_8665);
and U8778 (N_8778,N_8634,N_8662);
or U8779 (N_8779,N_8665,N_8661);
nand U8780 (N_8780,N_8685,N_8659);
and U8781 (N_8781,N_8676,N_8607);
or U8782 (N_8782,N_8665,N_8627);
or U8783 (N_8783,N_8610,N_8644);
nand U8784 (N_8784,N_8600,N_8641);
nor U8785 (N_8785,N_8666,N_8610);
nor U8786 (N_8786,N_8631,N_8621);
nand U8787 (N_8787,N_8614,N_8620);
nand U8788 (N_8788,N_8662,N_8617);
or U8789 (N_8789,N_8683,N_8681);
and U8790 (N_8790,N_8650,N_8622);
xnor U8791 (N_8791,N_8665,N_8689);
xnor U8792 (N_8792,N_8663,N_8609);
nand U8793 (N_8793,N_8682,N_8698);
nor U8794 (N_8794,N_8607,N_8604);
nand U8795 (N_8795,N_8615,N_8667);
nor U8796 (N_8796,N_8662,N_8638);
or U8797 (N_8797,N_8685,N_8662);
or U8798 (N_8798,N_8653,N_8640);
nor U8799 (N_8799,N_8642,N_8666);
and U8800 (N_8800,N_8732,N_8725);
or U8801 (N_8801,N_8722,N_8777);
nor U8802 (N_8802,N_8705,N_8782);
and U8803 (N_8803,N_8723,N_8798);
nor U8804 (N_8804,N_8772,N_8774);
nor U8805 (N_8805,N_8726,N_8717);
xnor U8806 (N_8806,N_8754,N_8767);
or U8807 (N_8807,N_8775,N_8734);
or U8808 (N_8808,N_8728,N_8793);
and U8809 (N_8809,N_8721,N_8785);
or U8810 (N_8810,N_8704,N_8736);
nor U8811 (N_8811,N_8759,N_8766);
nor U8812 (N_8812,N_8724,N_8770);
nor U8813 (N_8813,N_8792,N_8791);
nor U8814 (N_8814,N_8750,N_8742);
nand U8815 (N_8815,N_8790,N_8749);
xor U8816 (N_8816,N_8753,N_8762);
or U8817 (N_8817,N_8748,N_8768);
nor U8818 (N_8818,N_8714,N_8729);
nor U8819 (N_8819,N_8715,N_8780);
nand U8820 (N_8820,N_8781,N_8743);
nor U8821 (N_8821,N_8769,N_8703);
nor U8822 (N_8822,N_8708,N_8707);
and U8823 (N_8823,N_8794,N_8706);
nand U8824 (N_8824,N_8756,N_8713);
nor U8825 (N_8825,N_8702,N_8740);
nand U8826 (N_8826,N_8716,N_8752);
nor U8827 (N_8827,N_8757,N_8739);
nand U8828 (N_8828,N_8758,N_8738);
and U8829 (N_8829,N_8733,N_8778);
nor U8830 (N_8830,N_8773,N_8788);
nand U8831 (N_8831,N_8797,N_8711);
and U8832 (N_8832,N_8718,N_8735);
nor U8833 (N_8833,N_8737,N_8764);
nor U8834 (N_8834,N_8731,N_8763);
or U8835 (N_8835,N_8701,N_8787);
nor U8836 (N_8836,N_8761,N_8765);
or U8837 (N_8837,N_8727,N_8784);
and U8838 (N_8838,N_8744,N_8796);
or U8839 (N_8839,N_8799,N_8789);
xnor U8840 (N_8840,N_8747,N_8710);
or U8841 (N_8841,N_8760,N_8720);
nand U8842 (N_8842,N_8741,N_8745);
nand U8843 (N_8843,N_8719,N_8746);
nor U8844 (N_8844,N_8755,N_8700);
nand U8845 (N_8845,N_8776,N_8795);
and U8846 (N_8846,N_8779,N_8786);
or U8847 (N_8847,N_8709,N_8712);
and U8848 (N_8848,N_8751,N_8730);
or U8849 (N_8849,N_8783,N_8771);
xor U8850 (N_8850,N_8728,N_8754);
nor U8851 (N_8851,N_8782,N_8799);
nand U8852 (N_8852,N_8794,N_8716);
nand U8853 (N_8853,N_8703,N_8777);
and U8854 (N_8854,N_8798,N_8726);
and U8855 (N_8855,N_8734,N_8745);
and U8856 (N_8856,N_8725,N_8744);
and U8857 (N_8857,N_8720,N_8741);
and U8858 (N_8858,N_8775,N_8796);
or U8859 (N_8859,N_8729,N_8751);
or U8860 (N_8860,N_8715,N_8757);
nand U8861 (N_8861,N_8735,N_8741);
nor U8862 (N_8862,N_8795,N_8799);
and U8863 (N_8863,N_8782,N_8762);
nand U8864 (N_8864,N_8746,N_8765);
or U8865 (N_8865,N_8711,N_8721);
nand U8866 (N_8866,N_8759,N_8775);
nand U8867 (N_8867,N_8772,N_8732);
nand U8868 (N_8868,N_8726,N_8741);
and U8869 (N_8869,N_8799,N_8778);
nor U8870 (N_8870,N_8791,N_8753);
or U8871 (N_8871,N_8748,N_8764);
or U8872 (N_8872,N_8767,N_8708);
nand U8873 (N_8873,N_8796,N_8732);
and U8874 (N_8874,N_8724,N_8712);
nand U8875 (N_8875,N_8713,N_8766);
xnor U8876 (N_8876,N_8713,N_8757);
nand U8877 (N_8877,N_8743,N_8739);
or U8878 (N_8878,N_8759,N_8780);
or U8879 (N_8879,N_8712,N_8713);
xor U8880 (N_8880,N_8751,N_8744);
nor U8881 (N_8881,N_8757,N_8704);
or U8882 (N_8882,N_8703,N_8775);
and U8883 (N_8883,N_8799,N_8758);
nand U8884 (N_8884,N_8775,N_8769);
xor U8885 (N_8885,N_8782,N_8712);
or U8886 (N_8886,N_8773,N_8777);
and U8887 (N_8887,N_8740,N_8723);
xnor U8888 (N_8888,N_8700,N_8771);
xor U8889 (N_8889,N_8740,N_8773);
nand U8890 (N_8890,N_8715,N_8747);
nand U8891 (N_8891,N_8737,N_8770);
nor U8892 (N_8892,N_8756,N_8705);
xor U8893 (N_8893,N_8775,N_8763);
nor U8894 (N_8894,N_8788,N_8735);
nand U8895 (N_8895,N_8772,N_8719);
or U8896 (N_8896,N_8735,N_8766);
or U8897 (N_8897,N_8795,N_8701);
and U8898 (N_8898,N_8710,N_8707);
and U8899 (N_8899,N_8774,N_8778);
or U8900 (N_8900,N_8892,N_8869);
xor U8901 (N_8901,N_8839,N_8825);
nand U8902 (N_8902,N_8840,N_8899);
xor U8903 (N_8903,N_8831,N_8894);
and U8904 (N_8904,N_8812,N_8821);
xnor U8905 (N_8905,N_8868,N_8804);
and U8906 (N_8906,N_8806,N_8852);
nand U8907 (N_8907,N_8860,N_8856);
nor U8908 (N_8908,N_8876,N_8830);
nand U8909 (N_8909,N_8887,N_8819);
and U8910 (N_8910,N_8855,N_8858);
nor U8911 (N_8911,N_8810,N_8870);
and U8912 (N_8912,N_8820,N_8891);
nand U8913 (N_8913,N_8882,N_8878);
and U8914 (N_8914,N_8871,N_8866);
nor U8915 (N_8915,N_8881,N_8875);
nand U8916 (N_8916,N_8802,N_8800);
or U8917 (N_8917,N_8807,N_8814);
and U8918 (N_8918,N_8826,N_8811);
or U8919 (N_8919,N_8862,N_8801);
nor U8920 (N_8920,N_8889,N_8824);
nand U8921 (N_8921,N_8850,N_8895);
and U8922 (N_8922,N_8816,N_8897);
xnor U8923 (N_8923,N_8827,N_8835);
and U8924 (N_8924,N_8846,N_8844);
nand U8925 (N_8925,N_8865,N_8867);
or U8926 (N_8926,N_8803,N_8815);
nor U8927 (N_8927,N_8833,N_8864);
nor U8928 (N_8928,N_8837,N_8813);
nand U8929 (N_8929,N_8809,N_8845);
nand U8930 (N_8930,N_8823,N_8890);
nand U8931 (N_8931,N_8888,N_8874);
nor U8932 (N_8932,N_8847,N_8854);
or U8933 (N_8933,N_8822,N_8849);
or U8934 (N_8934,N_8880,N_8883);
and U8935 (N_8935,N_8818,N_8838);
and U8936 (N_8936,N_8861,N_8836);
and U8937 (N_8937,N_8808,N_8829);
or U8938 (N_8938,N_8859,N_8841);
nand U8939 (N_8939,N_8877,N_8872);
and U8940 (N_8940,N_8834,N_8886);
and U8941 (N_8941,N_8884,N_8832);
nor U8942 (N_8942,N_8879,N_8885);
and U8943 (N_8943,N_8851,N_8896);
nand U8944 (N_8944,N_8898,N_8863);
nand U8945 (N_8945,N_8873,N_8848);
nand U8946 (N_8946,N_8817,N_8843);
xor U8947 (N_8947,N_8853,N_8857);
or U8948 (N_8948,N_8805,N_8828);
nor U8949 (N_8949,N_8893,N_8842);
nor U8950 (N_8950,N_8830,N_8821);
or U8951 (N_8951,N_8898,N_8865);
and U8952 (N_8952,N_8854,N_8826);
nor U8953 (N_8953,N_8852,N_8844);
or U8954 (N_8954,N_8896,N_8842);
and U8955 (N_8955,N_8803,N_8870);
or U8956 (N_8956,N_8836,N_8849);
nor U8957 (N_8957,N_8810,N_8833);
nor U8958 (N_8958,N_8894,N_8897);
nor U8959 (N_8959,N_8842,N_8834);
xnor U8960 (N_8960,N_8824,N_8842);
nand U8961 (N_8961,N_8822,N_8858);
nor U8962 (N_8962,N_8823,N_8893);
nor U8963 (N_8963,N_8814,N_8861);
nand U8964 (N_8964,N_8849,N_8815);
nor U8965 (N_8965,N_8873,N_8863);
or U8966 (N_8966,N_8829,N_8873);
or U8967 (N_8967,N_8832,N_8846);
nand U8968 (N_8968,N_8884,N_8852);
and U8969 (N_8969,N_8877,N_8841);
or U8970 (N_8970,N_8824,N_8814);
or U8971 (N_8971,N_8803,N_8816);
or U8972 (N_8972,N_8873,N_8847);
nor U8973 (N_8973,N_8816,N_8827);
nor U8974 (N_8974,N_8808,N_8816);
nor U8975 (N_8975,N_8816,N_8859);
and U8976 (N_8976,N_8805,N_8892);
nand U8977 (N_8977,N_8814,N_8820);
or U8978 (N_8978,N_8801,N_8839);
xnor U8979 (N_8979,N_8866,N_8813);
and U8980 (N_8980,N_8871,N_8831);
and U8981 (N_8981,N_8873,N_8804);
nor U8982 (N_8982,N_8899,N_8843);
and U8983 (N_8983,N_8868,N_8897);
nand U8984 (N_8984,N_8858,N_8837);
and U8985 (N_8985,N_8823,N_8895);
or U8986 (N_8986,N_8854,N_8887);
nor U8987 (N_8987,N_8802,N_8843);
and U8988 (N_8988,N_8828,N_8889);
xor U8989 (N_8989,N_8872,N_8832);
nand U8990 (N_8990,N_8879,N_8845);
and U8991 (N_8991,N_8888,N_8858);
xor U8992 (N_8992,N_8839,N_8871);
nand U8993 (N_8993,N_8858,N_8818);
or U8994 (N_8994,N_8806,N_8880);
nor U8995 (N_8995,N_8819,N_8820);
and U8996 (N_8996,N_8860,N_8852);
and U8997 (N_8997,N_8823,N_8806);
nand U8998 (N_8998,N_8855,N_8831);
and U8999 (N_8999,N_8895,N_8880);
nor U9000 (N_9000,N_8999,N_8937);
xor U9001 (N_9001,N_8951,N_8962);
nand U9002 (N_9002,N_8958,N_8927);
nor U9003 (N_9003,N_8947,N_8995);
xor U9004 (N_9004,N_8981,N_8975);
nor U9005 (N_9005,N_8938,N_8993);
or U9006 (N_9006,N_8916,N_8914);
or U9007 (N_9007,N_8992,N_8952);
nor U9008 (N_9008,N_8919,N_8930);
and U9009 (N_9009,N_8922,N_8908);
xnor U9010 (N_9010,N_8997,N_8905);
and U9011 (N_9011,N_8990,N_8907);
nand U9012 (N_9012,N_8988,N_8924);
xor U9013 (N_9013,N_8915,N_8954);
nor U9014 (N_9014,N_8972,N_8902);
or U9015 (N_9015,N_8998,N_8994);
xor U9016 (N_9016,N_8932,N_8904);
nor U9017 (N_9017,N_8973,N_8960);
xor U9018 (N_9018,N_8964,N_8943);
nor U9019 (N_9019,N_8959,N_8909);
nand U9020 (N_9020,N_8968,N_8911);
and U9021 (N_9021,N_8950,N_8940);
or U9022 (N_9022,N_8953,N_8939);
xor U9023 (N_9023,N_8957,N_8921);
nor U9024 (N_9024,N_8949,N_8946);
and U9025 (N_9025,N_8970,N_8918);
nand U9026 (N_9026,N_8903,N_8917);
or U9027 (N_9027,N_8933,N_8925);
nand U9028 (N_9028,N_8928,N_8945);
and U9029 (N_9029,N_8976,N_8906);
and U9030 (N_9030,N_8966,N_8987);
and U9031 (N_9031,N_8982,N_8955);
nor U9032 (N_9032,N_8984,N_8910);
nor U9033 (N_9033,N_8991,N_8920);
or U9034 (N_9034,N_8935,N_8929);
or U9035 (N_9035,N_8956,N_8989);
nor U9036 (N_9036,N_8971,N_8977);
nand U9037 (N_9037,N_8969,N_8961);
nand U9038 (N_9038,N_8985,N_8979);
and U9039 (N_9039,N_8948,N_8936);
nand U9040 (N_9040,N_8967,N_8996);
and U9041 (N_9041,N_8913,N_8983);
xnor U9042 (N_9042,N_8963,N_8934);
nand U9043 (N_9043,N_8942,N_8980);
nand U9044 (N_9044,N_8912,N_8923);
nor U9045 (N_9045,N_8926,N_8974);
nor U9046 (N_9046,N_8931,N_8978);
and U9047 (N_9047,N_8900,N_8986);
nand U9048 (N_9048,N_8901,N_8944);
and U9049 (N_9049,N_8965,N_8941);
xor U9050 (N_9050,N_8949,N_8932);
or U9051 (N_9051,N_8998,N_8946);
nand U9052 (N_9052,N_8999,N_8940);
or U9053 (N_9053,N_8946,N_8915);
nand U9054 (N_9054,N_8941,N_8917);
and U9055 (N_9055,N_8977,N_8984);
nor U9056 (N_9056,N_8983,N_8975);
xnor U9057 (N_9057,N_8967,N_8906);
nand U9058 (N_9058,N_8918,N_8900);
and U9059 (N_9059,N_8963,N_8985);
nand U9060 (N_9060,N_8967,N_8909);
nor U9061 (N_9061,N_8912,N_8956);
and U9062 (N_9062,N_8973,N_8977);
or U9063 (N_9063,N_8944,N_8923);
nand U9064 (N_9064,N_8974,N_8973);
nand U9065 (N_9065,N_8920,N_8977);
xnor U9066 (N_9066,N_8948,N_8986);
nor U9067 (N_9067,N_8971,N_8948);
nor U9068 (N_9068,N_8952,N_8978);
nor U9069 (N_9069,N_8911,N_8948);
nor U9070 (N_9070,N_8982,N_8914);
or U9071 (N_9071,N_8937,N_8997);
and U9072 (N_9072,N_8936,N_8958);
and U9073 (N_9073,N_8961,N_8987);
nor U9074 (N_9074,N_8956,N_8926);
nand U9075 (N_9075,N_8947,N_8921);
nand U9076 (N_9076,N_8953,N_8919);
xor U9077 (N_9077,N_8901,N_8964);
nor U9078 (N_9078,N_8964,N_8976);
nor U9079 (N_9079,N_8994,N_8919);
or U9080 (N_9080,N_8960,N_8988);
and U9081 (N_9081,N_8958,N_8926);
nor U9082 (N_9082,N_8938,N_8940);
nor U9083 (N_9083,N_8956,N_8920);
and U9084 (N_9084,N_8999,N_8946);
and U9085 (N_9085,N_8940,N_8960);
nand U9086 (N_9086,N_8929,N_8918);
xnor U9087 (N_9087,N_8916,N_8961);
nand U9088 (N_9088,N_8958,N_8917);
nor U9089 (N_9089,N_8993,N_8996);
nor U9090 (N_9090,N_8900,N_8931);
xnor U9091 (N_9091,N_8901,N_8984);
nand U9092 (N_9092,N_8971,N_8917);
nand U9093 (N_9093,N_8941,N_8981);
nand U9094 (N_9094,N_8990,N_8962);
and U9095 (N_9095,N_8924,N_8980);
xnor U9096 (N_9096,N_8937,N_8993);
nor U9097 (N_9097,N_8938,N_8900);
xor U9098 (N_9098,N_8916,N_8978);
nand U9099 (N_9099,N_8941,N_8964);
nand U9100 (N_9100,N_9055,N_9031);
nand U9101 (N_9101,N_9015,N_9057);
or U9102 (N_9102,N_9086,N_9018);
and U9103 (N_9103,N_9069,N_9022);
or U9104 (N_9104,N_9003,N_9020);
and U9105 (N_9105,N_9095,N_9039);
or U9106 (N_9106,N_9044,N_9063);
or U9107 (N_9107,N_9075,N_9077);
and U9108 (N_9108,N_9000,N_9088);
and U9109 (N_9109,N_9034,N_9084);
nor U9110 (N_9110,N_9079,N_9094);
nand U9111 (N_9111,N_9089,N_9065);
and U9112 (N_9112,N_9053,N_9011);
or U9113 (N_9113,N_9099,N_9040);
or U9114 (N_9114,N_9027,N_9038);
or U9115 (N_9115,N_9082,N_9014);
or U9116 (N_9116,N_9002,N_9046);
nand U9117 (N_9117,N_9001,N_9073);
nand U9118 (N_9118,N_9090,N_9029);
nor U9119 (N_9119,N_9045,N_9081);
or U9120 (N_9120,N_9052,N_9051);
or U9121 (N_9121,N_9096,N_9025);
or U9122 (N_9122,N_9035,N_9071);
or U9123 (N_9123,N_9097,N_9013);
nor U9124 (N_9124,N_9030,N_9005);
or U9125 (N_9125,N_9093,N_9064);
nand U9126 (N_9126,N_9012,N_9058);
and U9127 (N_9127,N_9050,N_9048);
nor U9128 (N_9128,N_9083,N_9033);
and U9129 (N_9129,N_9042,N_9043);
nor U9130 (N_9130,N_9068,N_9007);
or U9131 (N_9131,N_9092,N_9047);
nor U9132 (N_9132,N_9019,N_9010);
nor U9133 (N_9133,N_9087,N_9056);
nand U9134 (N_9134,N_9009,N_9091);
nor U9135 (N_9135,N_9098,N_9078);
nand U9136 (N_9136,N_9067,N_9017);
and U9137 (N_9137,N_9036,N_9037);
or U9138 (N_9138,N_9004,N_9032);
nand U9139 (N_9139,N_9061,N_9026);
nor U9140 (N_9140,N_9028,N_9062);
nand U9141 (N_9141,N_9080,N_9085);
nor U9142 (N_9142,N_9024,N_9072);
nand U9143 (N_9143,N_9016,N_9041);
nor U9144 (N_9144,N_9076,N_9008);
xor U9145 (N_9145,N_9023,N_9060);
nand U9146 (N_9146,N_9066,N_9074);
or U9147 (N_9147,N_9021,N_9070);
nand U9148 (N_9148,N_9054,N_9049);
and U9149 (N_9149,N_9006,N_9059);
nor U9150 (N_9150,N_9073,N_9042);
or U9151 (N_9151,N_9020,N_9013);
or U9152 (N_9152,N_9017,N_9078);
and U9153 (N_9153,N_9068,N_9097);
and U9154 (N_9154,N_9006,N_9093);
nand U9155 (N_9155,N_9092,N_9079);
nor U9156 (N_9156,N_9072,N_9083);
nand U9157 (N_9157,N_9046,N_9045);
or U9158 (N_9158,N_9078,N_9041);
and U9159 (N_9159,N_9070,N_9097);
nor U9160 (N_9160,N_9023,N_9048);
nand U9161 (N_9161,N_9091,N_9013);
and U9162 (N_9162,N_9025,N_9008);
nor U9163 (N_9163,N_9035,N_9069);
or U9164 (N_9164,N_9085,N_9071);
nand U9165 (N_9165,N_9010,N_9038);
or U9166 (N_9166,N_9070,N_9036);
nor U9167 (N_9167,N_9063,N_9006);
xor U9168 (N_9168,N_9094,N_9065);
xnor U9169 (N_9169,N_9012,N_9032);
nand U9170 (N_9170,N_9072,N_9067);
and U9171 (N_9171,N_9039,N_9041);
and U9172 (N_9172,N_9058,N_9032);
nor U9173 (N_9173,N_9056,N_9022);
nor U9174 (N_9174,N_9076,N_9050);
or U9175 (N_9175,N_9036,N_9035);
nand U9176 (N_9176,N_9028,N_9020);
xnor U9177 (N_9177,N_9093,N_9083);
nor U9178 (N_9178,N_9059,N_9048);
and U9179 (N_9179,N_9081,N_9097);
or U9180 (N_9180,N_9049,N_9017);
or U9181 (N_9181,N_9046,N_9012);
or U9182 (N_9182,N_9038,N_9064);
or U9183 (N_9183,N_9041,N_9027);
nand U9184 (N_9184,N_9064,N_9069);
or U9185 (N_9185,N_9040,N_9094);
xor U9186 (N_9186,N_9000,N_9082);
nor U9187 (N_9187,N_9033,N_9052);
and U9188 (N_9188,N_9046,N_9031);
xnor U9189 (N_9189,N_9022,N_9027);
or U9190 (N_9190,N_9001,N_9056);
nand U9191 (N_9191,N_9038,N_9007);
nand U9192 (N_9192,N_9044,N_9009);
and U9193 (N_9193,N_9066,N_9044);
or U9194 (N_9194,N_9071,N_9043);
nor U9195 (N_9195,N_9079,N_9054);
nor U9196 (N_9196,N_9003,N_9037);
xor U9197 (N_9197,N_9079,N_9017);
xor U9198 (N_9198,N_9032,N_9063);
nand U9199 (N_9199,N_9075,N_9089);
nand U9200 (N_9200,N_9134,N_9171);
and U9201 (N_9201,N_9157,N_9195);
xnor U9202 (N_9202,N_9153,N_9118);
or U9203 (N_9203,N_9168,N_9121);
nand U9204 (N_9204,N_9187,N_9114);
nor U9205 (N_9205,N_9196,N_9159);
nor U9206 (N_9206,N_9193,N_9173);
or U9207 (N_9207,N_9108,N_9188);
and U9208 (N_9208,N_9139,N_9128);
or U9209 (N_9209,N_9154,N_9122);
nor U9210 (N_9210,N_9156,N_9152);
nor U9211 (N_9211,N_9123,N_9142);
nand U9212 (N_9212,N_9101,N_9164);
nand U9213 (N_9213,N_9127,N_9172);
nand U9214 (N_9214,N_9178,N_9111);
nor U9215 (N_9215,N_9138,N_9151);
and U9216 (N_9216,N_9105,N_9125);
or U9217 (N_9217,N_9145,N_9180);
nor U9218 (N_9218,N_9102,N_9147);
xor U9219 (N_9219,N_9186,N_9174);
or U9220 (N_9220,N_9148,N_9144);
xnor U9221 (N_9221,N_9185,N_9115);
nand U9222 (N_9222,N_9192,N_9119);
nor U9223 (N_9223,N_9120,N_9198);
or U9224 (N_9224,N_9162,N_9112);
xor U9225 (N_9225,N_9191,N_9166);
or U9226 (N_9226,N_9103,N_9129);
nor U9227 (N_9227,N_9176,N_9189);
xnor U9228 (N_9228,N_9124,N_9169);
nand U9229 (N_9229,N_9133,N_9109);
and U9230 (N_9230,N_9137,N_9146);
xor U9231 (N_9231,N_9106,N_9140);
and U9232 (N_9232,N_9143,N_9117);
nor U9233 (N_9233,N_9104,N_9135);
xor U9234 (N_9234,N_9141,N_9130);
and U9235 (N_9235,N_9160,N_9136);
nor U9236 (N_9236,N_9161,N_9165);
nand U9237 (N_9237,N_9107,N_9170);
or U9238 (N_9238,N_9167,N_9184);
xor U9239 (N_9239,N_9110,N_9163);
or U9240 (N_9240,N_9177,N_9158);
nor U9241 (N_9241,N_9132,N_9131);
nand U9242 (N_9242,N_9116,N_9175);
xnor U9243 (N_9243,N_9182,N_9197);
and U9244 (N_9244,N_9183,N_9126);
nand U9245 (N_9245,N_9113,N_9149);
and U9246 (N_9246,N_9155,N_9194);
and U9247 (N_9247,N_9181,N_9199);
nand U9248 (N_9248,N_9179,N_9190);
nor U9249 (N_9249,N_9150,N_9100);
nand U9250 (N_9250,N_9173,N_9127);
and U9251 (N_9251,N_9169,N_9162);
and U9252 (N_9252,N_9168,N_9131);
or U9253 (N_9253,N_9120,N_9121);
nand U9254 (N_9254,N_9147,N_9184);
nand U9255 (N_9255,N_9193,N_9131);
nand U9256 (N_9256,N_9180,N_9117);
nor U9257 (N_9257,N_9141,N_9170);
nand U9258 (N_9258,N_9118,N_9186);
xnor U9259 (N_9259,N_9142,N_9110);
nand U9260 (N_9260,N_9123,N_9146);
nand U9261 (N_9261,N_9139,N_9196);
or U9262 (N_9262,N_9190,N_9173);
nor U9263 (N_9263,N_9179,N_9124);
xor U9264 (N_9264,N_9179,N_9155);
nor U9265 (N_9265,N_9193,N_9123);
nand U9266 (N_9266,N_9129,N_9164);
nand U9267 (N_9267,N_9195,N_9141);
nor U9268 (N_9268,N_9117,N_9153);
and U9269 (N_9269,N_9117,N_9130);
or U9270 (N_9270,N_9137,N_9172);
nand U9271 (N_9271,N_9154,N_9107);
nand U9272 (N_9272,N_9168,N_9148);
nor U9273 (N_9273,N_9170,N_9108);
nor U9274 (N_9274,N_9156,N_9119);
nand U9275 (N_9275,N_9156,N_9163);
nand U9276 (N_9276,N_9117,N_9129);
or U9277 (N_9277,N_9112,N_9165);
or U9278 (N_9278,N_9182,N_9125);
nand U9279 (N_9279,N_9194,N_9118);
and U9280 (N_9280,N_9153,N_9176);
nand U9281 (N_9281,N_9199,N_9198);
xnor U9282 (N_9282,N_9195,N_9182);
and U9283 (N_9283,N_9176,N_9105);
nand U9284 (N_9284,N_9169,N_9131);
or U9285 (N_9285,N_9128,N_9159);
nand U9286 (N_9286,N_9113,N_9177);
nand U9287 (N_9287,N_9150,N_9193);
and U9288 (N_9288,N_9117,N_9162);
nand U9289 (N_9289,N_9141,N_9172);
nor U9290 (N_9290,N_9134,N_9178);
nor U9291 (N_9291,N_9127,N_9137);
xnor U9292 (N_9292,N_9179,N_9143);
nand U9293 (N_9293,N_9183,N_9189);
xor U9294 (N_9294,N_9179,N_9158);
or U9295 (N_9295,N_9129,N_9121);
nand U9296 (N_9296,N_9102,N_9108);
nand U9297 (N_9297,N_9100,N_9136);
or U9298 (N_9298,N_9188,N_9158);
nor U9299 (N_9299,N_9179,N_9135);
and U9300 (N_9300,N_9227,N_9214);
and U9301 (N_9301,N_9264,N_9204);
nor U9302 (N_9302,N_9269,N_9275);
nand U9303 (N_9303,N_9293,N_9257);
nand U9304 (N_9304,N_9265,N_9222);
and U9305 (N_9305,N_9219,N_9274);
or U9306 (N_9306,N_9278,N_9289);
nor U9307 (N_9307,N_9273,N_9205);
nor U9308 (N_9308,N_9242,N_9288);
nand U9309 (N_9309,N_9280,N_9236);
or U9310 (N_9310,N_9213,N_9263);
nor U9311 (N_9311,N_9281,N_9232);
nand U9312 (N_9312,N_9206,N_9259);
nand U9313 (N_9313,N_9233,N_9279);
or U9314 (N_9314,N_9209,N_9229);
nand U9315 (N_9315,N_9255,N_9210);
and U9316 (N_9316,N_9271,N_9287);
nor U9317 (N_9317,N_9215,N_9299);
or U9318 (N_9318,N_9211,N_9297);
nor U9319 (N_9319,N_9241,N_9260);
or U9320 (N_9320,N_9207,N_9261);
nor U9321 (N_9321,N_9248,N_9290);
nor U9322 (N_9322,N_9258,N_9235);
xnor U9323 (N_9323,N_9203,N_9249);
and U9324 (N_9324,N_9225,N_9208);
xnor U9325 (N_9325,N_9294,N_9262);
nor U9326 (N_9326,N_9251,N_9277);
or U9327 (N_9327,N_9224,N_9234);
or U9328 (N_9328,N_9237,N_9256);
nand U9329 (N_9329,N_9266,N_9267);
nor U9330 (N_9330,N_9268,N_9272);
or U9331 (N_9331,N_9230,N_9292);
and U9332 (N_9332,N_9220,N_9218);
or U9333 (N_9333,N_9252,N_9284);
or U9334 (N_9334,N_9212,N_9226);
nor U9335 (N_9335,N_9253,N_9291);
or U9336 (N_9336,N_9216,N_9231);
or U9337 (N_9337,N_9296,N_9295);
nor U9338 (N_9338,N_9250,N_9201);
nand U9339 (N_9339,N_9217,N_9298);
and U9340 (N_9340,N_9276,N_9238);
xor U9341 (N_9341,N_9245,N_9286);
nand U9342 (N_9342,N_9254,N_9270);
or U9343 (N_9343,N_9240,N_9200);
and U9344 (N_9344,N_9247,N_9282);
nand U9345 (N_9345,N_9243,N_9228);
or U9346 (N_9346,N_9244,N_9223);
nand U9347 (N_9347,N_9239,N_9283);
nand U9348 (N_9348,N_9221,N_9202);
or U9349 (N_9349,N_9246,N_9285);
nand U9350 (N_9350,N_9208,N_9265);
xnor U9351 (N_9351,N_9218,N_9213);
and U9352 (N_9352,N_9249,N_9229);
or U9353 (N_9353,N_9207,N_9222);
nand U9354 (N_9354,N_9259,N_9214);
and U9355 (N_9355,N_9226,N_9247);
nand U9356 (N_9356,N_9273,N_9235);
nand U9357 (N_9357,N_9251,N_9253);
nor U9358 (N_9358,N_9266,N_9206);
and U9359 (N_9359,N_9289,N_9292);
and U9360 (N_9360,N_9265,N_9210);
or U9361 (N_9361,N_9225,N_9235);
nand U9362 (N_9362,N_9266,N_9223);
or U9363 (N_9363,N_9201,N_9246);
nor U9364 (N_9364,N_9272,N_9285);
nand U9365 (N_9365,N_9204,N_9240);
nand U9366 (N_9366,N_9208,N_9277);
and U9367 (N_9367,N_9244,N_9288);
nor U9368 (N_9368,N_9238,N_9234);
nand U9369 (N_9369,N_9274,N_9215);
nand U9370 (N_9370,N_9214,N_9258);
nor U9371 (N_9371,N_9254,N_9256);
xnor U9372 (N_9372,N_9282,N_9293);
xor U9373 (N_9373,N_9246,N_9217);
nand U9374 (N_9374,N_9284,N_9245);
nor U9375 (N_9375,N_9271,N_9206);
xnor U9376 (N_9376,N_9210,N_9244);
nor U9377 (N_9377,N_9204,N_9224);
nand U9378 (N_9378,N_9252,N_9245);
xnor U9379 (N_9379,N_9208,N_9264);
or U9380 (N_9380,N_9231,N_9269);
nand U9381 (N_9381,N_9273,N_9262);
nand U9382 (N_9382,N_9238,N_9212);
nor U9383 (N_9383,N_9200,N_9268);
and U9384 (N_9384,N_9232,N_9265);
nand U9385 (N_9385,N_9265,N_9234);
and U9386 (N_9386,N_9289,N_9234);
nand U9387 (N_9387,N_9282,N_9260);
and U9388 (N_9388,N_9235,N_9222);
and U9389 (N_9389,N_9219,N_9241);
or U9390 (N_9390,N_9276,N_9212);
or U9391 (N_9391,N_9239,N_9297);
and U9392 (N_9392,N_9203,N_9206);
nand U9393 (N_9393,N_9214,N_9237);
nand U9394 (N_9394,N_9283,N_9269);
xor U9395 (N_9395,N_9244,N_9259);
and U9396 (N_9396,N_9239,N_9205);
and U9397 (N_9397,N_9280,N_9252);
nor U9398 (N_9398,N_9279,N_9285);
and U9399 (N_9399,N_9288,N_9298);
and U9400 (N_9400,N_9347,N_9352);
and U9401 (N_9401,N_9319,N_9308);
nand U9402 (N_9402,N_9353,N_9344);
and U9403 (N_9403,N_9372,N_9326);
and U9404 (N_9404,N_9395,N_9329);
nand U9405 (N_9405,N_9390,N_9374);
nor U9406 (N_9406,N_9322,N_9306);
or U9407 (N_9407,N_9399,N_9398);
nor U9408 (N_9408,N_9356,N_9392);
nand U9409 (N_9409,N_9314,N_9324);
nand U9410 (N_9410,N_9303,N_9311);
and U9411 (N_9411,N_9340,N_9341);
or U9412 (N_9412,N_9370,N_9369);
nand U9413 (N_9413,N_9387,N_9349);
xnor U9414 (N_9414,N_9373,N_9382);
and U9415 (N_9415,N_9328,N_9338);
nand U9416 (N_9416,N_9331,N_9342);
or U9417 (N_9417,N_9307,N_9301);
xor U9418 (N_9418,N_9381,N_9379);
and U9419 (N_9419,N_9332,N_9302);
nand U9420 (N_9420,N_9391,N_9355);
nand U9421 (N_9421,N_9304,N_9330);
and U9422 (N_9422,N_9380,N_9351);
nand U9423 (N_9423,N_9315,N_9394);
nand U9424 (N_9424,N_9318,N_9362);
and U9425 (N_9425,N_9383,N_9359);
and U9426 (N_9426,N_9397,N_9313);
nand U9427 (N_9427,N_9388,N_9350);
nor U9428 (N_9428,N_9361,N_9327);
nand U9429 (N_9429,N_9375,N_9305);
nand U9430 (N_9430,N_9385,N_9354);
nor U9431 (N_9431,N_9360,N_9384);
xnor U9432 (N_9432,N_9366,N_9323);
nor U9433 (N_9433,N_9300,N_9365);
and U9434 (N_9434,N_9333,N_9336);
xor U9435 (N_9435,N_9378,N_9348);
and U9436 (N_9436,N_9312,N_9364);
nand U9437 (N_9437,N_9346,N_9386);
or U9438 (N_9438,N_9376,N_9396);
and U9439 (N_9439,N_9309,N_9317);
nand U9440 (N_9440,N_9358,N_9316);
nor U9441 (N_9441,N_9334,N_9389);
and U9442 (N_9442,N_9321,N_9371);
nand U9443 (N_9443,N_9339,N_9377);
nor U9444 (N_9444,N_9337,N_9357);
nor U9445 (N_9445,N_9310,N_9345);
nand U9446 (N_9446,N_9335,N_9393);
or U9447 (N_9447,N_9343,N_9320);
xnor U9448 (N_9448,N_9325,N_9368);
or U9449 (N_9449,N_9363,N_9367);
nand U9450 (N_9450,N_9323,N_9305);
nor U9451 (N_9451,N_9383,N_9375);
or U9452 (N_9452,N_9353,N_9337);
nand U9453 (N_9453,N_9314,N_9335);
xnor U9454 (N_9454,N_9355,N_9352);
and U9455 (N_9455,N_9307,N_9323);
or U9456 (N_9456,N_9330,N_9337);
or U9457 (N_9457,N_9366,N_9357);
or U9458 (N_9458,N_9376,N_9383);
nand U9459 (N_9459,N_9328,N_9340);
nor U9460 (N_9460,N_9334,N_9332);
nor U9461 (N_9461,N_9380,N_9354);
nor U9462 (N_9462,N_9333,N_9352);
nand U9463 (N_9463,N_9301,N_9396);
nand U9464 (N_9464,N_9310,N_9338);
nor U9465 (N_9465,N_9386,N_9357);
or U9466 (N_9466,N_9315,N_9377);
or U9467 (N_9467,N_9352,N_9345);
xnor U9468 (N_9468,N_9320,N_9372);
and U9469 (N_9469,N_9363,N_9308);
and U9470 (N_9470,N_9339,N_9355);
and U9471 (N_9471,N_9384,N_9323);
and U9472 (N_9472,N_9322,N_9392);
and U9473 (N_9473,N_9391,N_9380);
and U9474 (N_9474,N_9385,N_9386);
nand U9475 (N_9475,N_9352,N_9327);
nand U9476 (N_9476,N_9312,N_9391);
nor U9477 (N_9477,N_9355,N_9346);
xnor U9478 (N_9478,N_9334,N_9336);
nand U9479 (N_9479,N_9366,N_9361);
nand U9480 (N_9480,N_9388,N_9344);
nor U9481 (N_9481,N_9340,N_9345);
nand U9482 (N_9482,N_9303,N_9305);
or U9483 (N_9483,N_9371,N_9357);
nand U9484 (N_9484,N_9336,N_9391);
nor U9485 (N_9485,N_9339,N_9338);
nand U9486 (N_9486,N_9333,N_9358);
nand U9487 (N_9487,N_9325,N_9378);
nand U9488 (N_9488,N_9355,N_9344);
or U9489 (N_9489,N_9398,N_9370);
xor U9490 (N_9490,N_9342,N_9350);
or U9491 (N_9491,N_9312,N_9331);
xnor U9492 (N_9492,N_9340,N_9300);
and U9493 (N_9493,N_9311,N_9317);
nor U9494 (N_9494,N_9339,N_9311);
and U9495 (N_9495,N_9329,N_9320);
nor U9496 (N_9496,N_9302,N_9354);
xor U9497 (N_9497,N_9318,N_9311);
xor U9498 (N_9498,N_9351,N_9337);
or U9499 (N_9499,N_9361,N_9304);
nor U9500 (N_9500,N_9456,N_9423);
nand U9501 (N_9501,N_9428,N_9433);
and U9502 (N_9502,N_9437,N_9499);
nor U9503 (N_9503,N_9409,N_9462);
nand U9504 (N_9504,N_9474,N_9401);
or U9505 (N_9505,N_9492,N_9411);
and U9506 (N_9506,N_9413,N_9436);
xnor U9507 (N_9507,N_9458,N_9479);
nor U9508 (N_9508,N_9419,N_9468);
xor U9509 (N_9509,N_9444,N_9426);
xor U9510 (N_9510,N_9450,N_9490);
or U9511 (N_9511,N_9480,N_9454);
or U9512 (N_9512,N_9459,N_9466);
nand U9513 (N_9513,N_9495,N_9445);
or U9514 (N_9514,N_9488,N_9469);
and U9515 (N_9515,N_9482,N_9489);
nand U9516 (N_9516,N_9431,N_9418);
or U9517 (N_9517,N_9406,N_9452);
nand U9518 (N_9518,N_9415,N_9476);
and U9519 (N_9519,N_9477,N_9439);
nand U9520 (N_9520,N_9457,N_9441);
nand U9521 (N_9521,N_9449,N_9494);
or U9522 (N_9522,N_9475,N_9414);
nand U9523 (N_9523,N_9461,N_9404);
or U9524 (N_9524,N_9487,N_9416);
or U9525 (N_9525,N_9408,N_9472);
and U9526 (N_9526,N_9402,N_9446);
or U9527 (N_9527,N_9493,N_9435);
nor U9528 (N_9528,N_9470,N_9432);
xnor U9529 (N_9529,N_9484,N_9498);
nor U9530 (N_9530,N_9427,N_9429);
or U9531 (N_9531,N_9420,N_9410);
nand U9532 (N_9532,N_9438,N_9453);
nand U9533 (N_9533,N_9407,N_9486);
nand U9534 (N_9534,N_9463,N_9497);
and U9535 (N_9535,N_9425,N_9478);
nand U9536 (N_9536,N_9424,N_9434);
nor U9537 (N_9537,N_9447,N_9460);
nor U9538 (N_9538,N_9417,N_9481);
or U9539 (N_9539,N_9442,N_9455);
and U9540 (N_9540,N_9443,N_9465);
nor U9541 (N_9541,N_9403,N_9496);
nand U9542 (N_9542,N_9405,N_9491);
nand U9543 (N_9543,N_9422,N_9400);
nand U9544 (N_9544,N_9485,N_9467);
and U9545 (N_9545,N_9440,N_9430);
or U9546 (N_9546,N_9421,N_9412);
or U9547 (N_9547,N_9471,N_9448);
nor U9548 (N_9548,N_9464,N_9451);
and U9549 (N_9549,N_9473,N_9483);
or U9550 (N_9550,N_9442,N_9441);
or U9551 (N_9551,N_9475,N_9499);
or U9552 (N_9552,N_9436,N_9446);
and U9553 (N_9553,N_9465,N_9449);
and U9554 (N_9554,N_9482,N_9476);
nand U9555 (N_9555,N_9467,N_9418);
nand U9556 (N_9556,N_9466,N_9492);
nor U9557 (N_9557,N_9403,N_9487);
nor U9558 (N_9558,N_9452,N_9442);
nand U9559 (N_9559,N_9496,N_9430);
nor U9560 (N_9560,N_9474,N_9464);
nor U9561 (N_9561,N_9417,N_9427);
xor U9562 (N_9562,N_9458,N_9410);
or U9563 (N_9563,N_9493,N_9418);
or U9564 (N_9564,N_9452,N_9407);
or U9565 (N_9565,N_9478,N_9410);
nor U9566 (N_9566,N_9455,N_9427);
nand U9567 (N_9567,N_9434,N_9469);
nor U9568 (N_9568,N_9409,N_9425);
and U9569 (N_9569,N_9430,N_9475);
nor U9570 (N_9570,N_9406,N_9454);
nand U9571 (N_9571,N_9478,N_9430);
or U9572 (N_9572,N_9421,N_9411);
nand U9573 (N_9573,N_9475,N_9408);
or U9574 (N_9574,N_9417,N_9453);
or U9575 (N_9575,N_9405,N_9486);
or U9576 (N_9576,N_9416,N_9481);
nor U9577 (N_9577,N_9444,N_9463);
nand U9578 (N_9578,N_9478,N_9416);
nor U9579 (N_9579,N_9443,N_9454);
nor U9580 (N_9580,N_9470,N_9471);
or U9581 (N_9581,N_9415,N_9468);
nand U9582 (N_9582,N_9499,N_9452);
or U9583 (N_9583,N_9496,N_9491);
or U9584 (N_9584,N_9470,N_9493);
nor U9585 (N_9585,N_9452,N_9455);
or U9586 (N_9586,N_9442,N_9437);
nand U9587 (N_9587,N_9409,N_9494);
or U9588 (N_9588,N_9433,N_9447);
nor U9589 (N_9589,N_9447,N_9451);
nor U9590 (N_9590,N_9440,N_9449);
xnor U9591 (N_9591,N_9459,N_9463);
xnor U9592 (N_9592,N_9495,N_9412);
and U9593 (N_9593,N_9479,N_9495);
nand U9594 (N_9594,N_9492,N_9432);
and U9595 (N_9595,N_9425,N_9454);
nand U9596 (N_9596,N_9421,N_9473);
and U9597 (N_9597,N_9498,N_9419);
xor U9598 (N_9598,N_9417,N_9462);
or U9599 (N_9599,N_9400,N_9469);
or U9600 (N_9600,N_9535,N_9594);
nor U9601 (N_9601,N_9595,N_9509);
nand U9602 (N_9602,N_9562,N_9565);
and U9603 (N_9603,N_9530,N_9527);
nand U9604 (N_9604,N_9598,N_9597);
nand U9605 (N_9605,N_9502,N_9554);
nand U9606 (N_9606,N_9569,N_9556);
and U9607 (N_9607,N_9513,N_9573);
and U9608 (N_9608,N_9552,N_9593);
or U9609 (N_9609,N_9567,N_9533);
or U9610 (N_9610,N_9558,N_9540);
nor U9611 (N_9611,N_9521,N_9583);
xor U9612 (N_9612,N_9525,N_9577);
nand U9613 (N_9613,N_9505,N_9588);
nand U9614 (N_9614,N_9572,N_9579);
or U9615 (N_9615,N_9599,N_9589);
and U9616 (N_9616,N_9526,N_9529);
xor U9617 (N_9617,N_9538,N_9547);
nor U9618 (N_9618,N_9563,N_9517);
and U9619 (N_9619,N_9549,N_9534);
and U9620 (N_9620,N_9586,N_9542);
nand U9621 (N_9621,N_9512,N_9571);
or U9622 (N_9622,N_9543,N_9584);
nor U9623 (N_9623,N_9522,N_9566);
nand U9624 (N_9624,N_9585,N_9532);
or U9625 (N_9625,N_9500,N_9591);
nand U9626 (N_9626,N_9574,N_9555);
nand U9627 (N_9627,N_9548,N_9596);
nor U9628 (N_9628,N_9507,N_9559);
nor U9629 (N_9629,N_9557,N_9524);
nand U9630 (N_9630,N_9546,N_9516);
nand U9631 (N_9631,N_9581,N_9582);
and U9632 (N_9632,N_9523,N_9578);
nor U9633 (N_9633,N_9560,N_9515);
nand U9634 (N_9634,N_9576,N_9519);
xnor U9635 (N_9635,N_9541,N_9506);
nand U9636 (N_9636,N_9551,N_9510);
and U9637 (N_9637,N_9550,N_9501);
nand U9638 (N_9638,N_9537,N_9590);
nor U9639 (N_9639,N_9561,N_9514);
nand U9640 (N_9640,N_9570,N_9508);
nor U9641 (N_9641,N_9544,N_9518);
and U9642 (N_9642,N_9511,N_9520);
and U9643 (N_9643,N_9564,N_9587);
nor U9644 (N_9644,N_9536,N_9503);
or U9645 (N_9645,N_9553,N_9528);
and U9646 (N_9646,N_9575,N_9504);
xnor U9647 (N_9647,N_9568,N_9592);
or U9648 (N_9648,N_9539,N_9531);
and U9649 (N_9649,N_9545,N_9580);
nor U9650 (N_9650,N_9519,N_9595);
or U9651 (N_9651,N_9523,N_9581);
or U9652 (N_9652,N_9566,N_9555);
nor U9653 (N_9653,N_9564,N_9576);
or U9654 (N_9654,N_9531,N_9594);
nand U9655 (N_9655,N_9562,N_9512);
nor U9656 (N_9656,N_9540,N_9523);
and U9657 (N_9657,N_9587,N_9568);
nor U9658 (N_9658,N_9599,N_9562);
or U9659 (N_9659,N_9584,N_9560);
or U9660 (N_9660,N_9548,N_9507);
nor U9661 (N_9661,N_9582,N_9559);
nand U9662 (N_9662,N_9571,N_9575);
and U9663 (N_9663,N_9564,N_9586);
xor U9664 (N_9664,N_9552,N_9536);
xor U9665 (N_9665,N_9506,N_9559);
and U9666 (N_9666,N_9528,N_9511);
and U9667 (N_9667,N_9525,N_9570);
or U9668 (N_9668,N_9532,N_9569);
or U9669 (N_9669,N_9518,N_9576);
nor U9670 (N_9670,N_9515,N_9523);
or U9671 (N_9671,N_9502,N_9526);
nor U9672 (N_9672,N_9563,N_9574);
xor U9673 (N_9673,N_9554,N_9573);
or U9674 (N_9674,N_9527,N_9529);
and U9675 (N_9675,N_9508,N_9564);
nor U9676 (N_9676,N_9535,N_9584);
and U9677 (N_9677,N_9566,N_9514);
or U9678 (N_9678,N_9562,N_9506);
and U9679 (N_9679,N_9510,N_9518);
or U9680 (N_9680,N_9502,N_9524);
nor U9681 (N_9681,N_9523,N_9573);
or U9682 (N_9682,N_9554,N_9582);
or U9683 (N_9683,N_9570,N_9580);
and U9684 (N_9684,N_9549,N_9520);
or U9685 (N_9685,N_9543,N_9598);
nand U9686 (N_9686,N_9569,N_9592);
or U9687 (N_9687,N_9588,N_9564);
nand U9688 (N_9688,N_9519,N_9538);
nor U9689 (N_9689,N_9569,N_9591);
nor U9690 (N_9690,N_9593,N_9582);
nand U9691 (N_9691,N_9516,N_9596);
xor U9692 (N_9692,N_9594,N_9552);
or U9693 (N_9693,N_9595,N_9567);
and U9694 (N_9694,N_9571,N_9517);
nand U9695 (N_9695,N_9550,N_9514);
nand U9696 (N_9696,N_9560,N_9533);
and U9697 (N_9697,N_9596,N_9512);
or U9698 (N_9698,N_9507,N_9558);
nand U9699 (N_9699,N_9503,N_9508);
nand U9700 (N_9700,N_9627,N_9655);
or U9701 (N_9701,N_9622,N_9610);
nor U9702 (N_9702,N_9684,N_9617);
or U9703 (N_9703,N_9623,N_9687);
and U9704 (N_9704,N_9675,N_9681);
nand U9705 (N_9705,N_9647,N_9633);
nand U9706 (N_9706,N_9642,N_9648);
and U9707 (N_9707,N_9665,N_9603);
or U9708 (N_9708,N_9661,N_9654);
xnor U9709 (N_9709,N_9669,N_9663);
nand U9710 (N_9710,N_9635,N_9608);
nor U9711 (N_9711,N_9621,N_9676);
nand U9712 (N_9712,N_9695,N_9682);
or U9713 (N_9713,N_9628,N_9614);
xor U9714 (N_9714,N_9636,N_9692);
nor U9715 (N_9715,N_9656,N_9696);
nor U9716 (N_9716,N_9699,N_9658);
nor U9717 (N_9717,N_9697,N_9620);
nand U9718 (N_9718,N_9600,N_9650);
and U9719 (N_9719,N_9653,N_9688);
or U9720 (N_9720,N_9690,N_9686);
nor U9721 (N_9721,N_9689,N_9606);
and U9722 (N_9722,N_9629,N_9649);
nand U9723 (N_9723,N_9641,N_9601);
nand U9724 (N_9724,N_9612,N_9646);
nor U9725 (N_9725,N_9662,N_9677);
or U9726 (N_9726,N_9673,N_9643);
nand U9727 (N_9727,N_9667,N_9607);
and U9728 (N_9728,N_9664,N_9619);
nor U9729 (N_9729,N_9670,N_9634);
nor U9730 (N_9730,N_9605,N_9691);
and U9731 (N_9731,N_9657,N_9630);
nand U9732 (N_9732,N_9616,N_9685);
or U9733 (N_9733,N_9694,N_9625);
or U9734 (N_9734,N_9683,N_9698);
or U9735 (N_9735,N_9680,N_9674);
and U9736 (N_9736,N_9637,N_9604);
nand U9737 (N_9737,N_9659,N_9652);
nand U9738 (N_9738,N_9626,N_9624);
nand U9739 (N_9739,N_9631,N_9660);
xnor U9740 (N_9740,N_9609,N_9644);
nand U9741 (N_9741,N_9678,N_9618);
nor U9742 (N_9742,N_9651,N_9602);
xor U9743 (N_9743,N_9611,N_9672);
or U9744 (N_9744,N_9693,N_9615);
nor U9745 (N_9745,N_9639,N_9666);
and U9746 (N_9746,N_9640,N_9613);
nor U9747 (N_9747,N_9638,N_9645);
or U9748 (N_9748,N_9632,N_9668);
nand U9749 (N_9749,N_9671,N_9679);
and U9750 (N_9750,N_9610,N_9654);
nand U9751 (N_9751,N_9612,N_9608);
nor U9752 (N_9752,N_9670,N_9621);
and U9753 (N_9753,N_9697,N_9635);
and U9754 (N_9754,N_9639,N_9640);
nand U9755 (N_9755,N_9608,N_9621);
and U9756 (N_9756,N_9664,N_9656);
nor U9757 (N_9757,N_9699,N_9604);
nand U9758 (N_9758,N_9612,N_9633);
nor U9759 (N_9759,N_9602,N_9604);
and U9760 (N_9760,N_9640,N_9687);
and U9761 (N_9761,N_9656,N_9620);
or U9762 (N_9762,N_9689,N_9612);
xor U9763 (N_9763,N_9649,N_9684);
or U9764 (N_9764,N_9648,N_9661);
nand U9765 (N_9765,N_9622,N_9663);
and U9766 (N_9766,N_9617,N_9670);
or U9767 (N_9767,N_9663,N_9659);
nand U9768 (N_9768,N_9665,N_9645);
xor U9769 (N_9769,N_9650,N_9684);
xnor U9770 (N_9770,N_9693,N_9664);
nor U9771 (N_9771,N_9690,N_9672);
nor U9772 (N_9772,N_9682,N_9698);
and U9773 (N_9773,N_9617,N_9610);
nand U9774 (N_9774,N_9650,N_9620);
nand U9775 (N_9775,N_9688,N_9677);
or U9776 (N_9776,N_9664,N_9640);
or U9777 (N_9777,N_9613,N_9646);
nand U9778 (N_9778,N_9605,N_9685);
or U9779 (N_9779,N_9639,N_9677);
nor U9780 (N_9780,N_9642,N_9638);
nor U9781 (N_9781,N_9658,N_9635);
nor U9782 (N_9782,N_9675,N_9631);
nor U9783 (N_9783,N_9610,N_9614);
xor U9784 (N_9784,N_9615,N_9637);
and U9785 (N_9785,N_9696,N_9688);
nand U9786 (N_9786,N_9638,N_9653);
or U9787 (N_9787,N_9611,N_9630);
and U9788 (N_9788,N_9629,N_9661);
and U9789 (N_9789,N_9647,N_9622);
xor U9790 (N_9790,N_9629,N_9613);
nor U9791 (N_9791,N_9611,N_9673);
and U9792 (N_9792,N_9674,N_9604);
nor U9793 (N_9793,N_9617,N_9678);
nor U9794 (N_9794,N_9606,N_9651);
xor U9795 (N_9795,N_9621,N_9693);
nand U9796 (N_9796,N_9683,N_9629);
and U9797 (N_9797,N_9672,N_9643);
and U9798 (N_9798,N_9679,N_9696);
or U9799 (N_9799,N_9603,N_9644);
or U9800 (N_9800,N_9757,N_9713);
nand U9801 (N_9801,N_9733,N_9732);
or U9802 (N_9802,N_9779,N_9703);
nor U9803 (N_9803,N_9705,N_9785);
and U9804 (N_9804,N_9700,N_9775);
or U9805 (N_9805,N_9736,N_9794);
or U9806 (N_9806,N_9792,N_9774);
and U9807 (N_9807,N_9707,N_9750);
nand U9808 (N_9808,N_9742,N_9728);
or U9809 (N_9809,N_9796,N_9763);
nand U9810 (N_9810,N_9701,N_9778);
nor U9811 (N_9811,N_9767,N_9740);
xnor U9812 (N_9812,N_9752,N_9765);
or U9813 (N_9813,N_9766,N_9709);
nand U9814 (N_9814,N_9708,N_9731);
and U9815 (N_9815,N_9730,N_9738);
nor U9816 (N_9816,N_9754,N_9715);
nand U9817 (N_9817,N_9727,N_9726);
nor U9818 (N_9818,N_9753,N_9723);
or U9819 (N_9819,N_9748,N_9771);
nand U9820 (N_9820,N_9739,N_9702);
xor U9821 (N_9821,N_9725,N_9782);
or U9822 (N_9822,N_9716,N_9729);
and U9823 (N_9823,N_9737,N_9741);
and U9824 (N_9824,N_9790,N_9735);
and U9825 (N_9825,N_9777,N_9786);
nor U9826 (N_9826,N_9795,N_9798);
or U9827 (N_9827,N_9780,N_9706);
or U9828 (N_9828,N_9710,N_9764);
or U9829 (N_9829,N_9714,N_9747);
and U9830 (N_9830,N_9761,N_9745);
nor U9831 (N_9831,N_9720,N_9781);
and U9832 (N_9832,N_9721,N_9760);
nor U9833 (N_9833,N_9793,N_9719);
or U9834 (N_9834,N_9712,N_9784);
and U9835 (N_9835,N_9773,N_9724);
nand U9836 (N_9836,N_9743,N_9744);
or U9837 (N_9837,N_9722,N_9791);
nor U9838 (N_9838,N_9789,N_9769);
nor U9839 (N_9839,N_9776,N_9717);
xnor U9840 (N_9840,N_9751,N_9787);
xnor U9841 (N_9841,N_9749,N_9799);
nand U9842 (N_9842,N_9756,N_9718);
nand U9843 (N_9843,N_9762,N_9711);
and U9844 (N_9844,N_9783,N_9755);
nor U9845 (N_9845,N_9768,N_9770);
and U9846 (N_9846,N_9734,N_9759);
nand U9847 (N_9847,N_9788,N_9746);
and U9848 (N_9848,N_9758,N_9772);
or U9849 (N_9849,N_9797,N_9704);
or U9850 (N_9850,N_9773,N_9714);
xnor U9851 (N_9851,N_9705,N_9761);
and U9852 (N_9852,N_9708,N_9790);
nor U9853 (N_9853,N_9712,N_9730);
or U9854 (N_9854,N_9748,N_9793);
or U9855 (N_9855,N_9768,N_9730);
and U9856 (N_9856,N_9748,N_9795);
nor U9857 (N_9857,N_9702,N_9787);
nor U9858 (N_9858,N_9765,N_9700);
xor U9859 (N_9859,N_9742,N_9773);
xnor U9860 (N_9860,N_9724,N_9717);
nor U9861 (N_9861,N_9767,N_9748);
and U9862 (N_9862,N_9740,N_9741);
or U9863 (N_9863,N_9780,N_9715);
nand U9864 (N_9864,N_9784,N_9713);
or U9865 (N_9865,N_9776,N_9743);
nor U9866 (N_9866,N_9778,N_9741);
nand U9867 (N_9867,N_9700,N_9780);
nor U9868 (N_9868,N_9733,N_9754);
nand U9869 (N_9869,N_9734,N_9763);
or U9870 (N_9870,N_9777,N_9759);
and U9871 (N_9871,N_9709,N_9725);
or U9872 (N_9872,N_9746,N_9757);
or U9873 (N_9873,N_9729,N_9781);
or U9874 (N_9874,N_9797,N_9746);
nand U9875 (N_9875,N_9719,N_9791);
and U9876 (N_9876,N_9748,N_9772);
or U9877 (N_9877,N_9720,N_9719);
and U9878 (N_9878,N_9734,N_9789);
xnor U9879 (N_9879,N_9723,N_9783);
nor U9880 (N_9880,N_9700,N_9733);
or U9881 (N_9881,N_9737,N_9758);
and U9882 (N_9882,N_9715,N_9716);
and U9883 (N_9883,N_9759,N_9785);
or U9884 (N_9884,N_9721,N_9777);
and U9885 (N_9885,N_9729,N_9717);
nand U9886 (N_9886,N_9701,N_9772);
or U9887 (N_9887,N_9788,N_9714);
xor U9888 (N_9888,N_9728,N_9763);
and U9889 (N_9889,N_9788,N_9775);
and U9890 (N_9890,N_9728,N_9721);
nor U9891 (N_9891,N_9770,N_9727);
xor U9892 (N_9892,N_9713,N_9709);
and U9893 (N_9893,N_9770,N_9757);
nand U9894 (N_9894,N_9780,N_9793);
nand U9895 (N_9895,N_9728,N_9772);
or U9896 (N_9896,N_9769,N_9737);
and U9897 (N_9897,N_9726,N_9763);
nor U9898 (N_9898,N_9743,N_9786);
nor U9899 (N_9899,N_9786,N_9762);
nor U9900 (N_9900,N_9898,N_9801);
or U9901 (N_9901,N_9842,N_9810);
nor U9902 (N_9902,N_9815,N_9830);
nand U9903 (N_9903,N_9890,N_9897);
nand U9904 (N_9904,N_9826,N_9839);
or U9905 (N_9905,N_9888,N_9885);
and U9906 (N_9906,N_9873,N_9832);
nor U9907 (N_9907,N_9867,N_9875);
nor U9908 (N_9908,N_9825,N_9843);
nand U9909 (N_9909,N_9840,N_9824);
nand U9910 (N_9910,N_9865,N_9841);
nand U9911 (N_9911,N_9800,N_9848);
xor U9912 (N_9912,N_9846,N_9882);
and U9913 (N_9913,N_9861,N_9819);
or U9914 (N_9914,N_9817,N_9837);
or U9915 (N_9915,N_9828,N_9871);
nand U9916 (N_9916,N_9835,N_9881);
and U9917 (N_9917,N_9869,N_9862);
nor U9918 (N_9918,N_9812,N_9803);
and U9919 (N_9919,N_9821,N_9805);
or U9920 (N_9920,N_9886,N_9860);
nor U9921 (N_9921,N_9814,N_9852);
xnor U9922 (N_9922,N_9808,N_9836);
nor U9923 (N_9923,N_9856,N_9811);
nand U9924 (N_9924,N_9863,N_9877);
or U9925 (N_9925,N_9866,N_9878);
nand U9926 (N_9926,N_9807,N_9844);
nand U9927 (N_9927,N_9870,N_9818);
and U9928 (N_9928,N_9802,N_9879);
or U9929 (N_9929,N_9850,N_9851);
nor U9930 (N_9930,N_9816,N_9827);
or U9931 (N_9931,N_9847,N_9899);
and U9932 (N_9932,N_9822,N_9853);
nand U9933 (N_9933,N_9893,N_9833);
nand U9934 (N_9934,N_9838,N_9872);
and U9935 (N_9935,N_9809,N_9834);
or U9936 (N_9936,N_9829,N_9883);
nor U9937 (N_9937,N_9894,N_9855);
or U9938 (N_9938,N_9889,N_9891);
nand U9939 (N_9939,N_9813,N_9892);
or U9940 (N_9940,N_9806,N_9823);
nand U9941 (N_9941,N_9857,N_9804);
nor U9942 (N_9942,N_9859,N_9880);
nand U9943 (N_9943,N_9849,N_9831);
or U9944 (N_9944,N_9895,N_9874);
xor U9945 (N_9945,N_9896,N_9845);
or U9946 (N_9946,N_9887,N_9864);
nor U9947 (N_9947,N_9876,N_9884);
nor U9948 (N_9948,N_9854,N_9820);
and U9949 (N_9949,N_9858,N_9868);
or U9950 (N_9950,N_9862,N_9852);
nor U9951 (N_9951,N_9809,N_9847);
nor U9952 (N_9952,N_9806,N_9877);
nand U9953 (N_9953,N_9806,N_9841);
nand U9954 (N_9954,N_9804,N_9800);
and U9955 (N_9955,N_9825,N_9882);
nor U9956 (N_9956,N_9801,N_9887);
or U9957 (N_9957,N_9865,N_9833);
nand U9958 (N_9958,N_9882,N_9800);
nor U9959 (N_9959,N_9899,N_9828);
and U9960 (N_9960,N_9804,N_9802);
nand U9961 (N_9961,N_9866,N_9819);
and U9962 (N_9962,N_9873,N_9857);
xnor U9963 (N_9963,N_9867,N_9898);
or U9964 (N_9964,N_9843,N_9849);
and U9965 (N_9965,N_9827,N_9846);
nand U9966 (N_9966,N_9864,N_9871);
or U9967 (N_9967,N_9871,N_9821);
and U9968 (N_9968,N_9872,N_9824);
or U9969 (N_9969,N_9863,N_9855);
nand U9970 (N_9970,N_9871,N_9873);
or U9971 (N_9971,N_9886,N_9813);
nand U9972 (N_9972,N_9822,N_9825);
nand U9973 (N_9973,N_9887,N_9806);
and U9974 (N_9974,N_9836,N_9817);
and U9975 (N_9975,N_9812,N_9808);
nand U9976 (N_9976,N_9879,N_9892);
nor U9977 (N_9977,N_9803,N_9858);
nand U9978 (N_9978,N_9824,N_9887);
or U9979 (N_9979,N_9893,N_9825);
and U9980 (N_9980,N_9865,N_9897);
xnor U9981 (N_9981,N_9825,N_9894);
nor U9982 (N_9982,N_9877,N_9822);
nand U9983 (N_9983,N_9823,N_9898);
xnor U9984 (N_9984,N_9810,N_9817);
nand U9985 (N_9985,N_9860,N_9881);
xnor U9986 (N_9986,N_9853,N_9844);
xor U9987 (N_9987,N_9896,N_9805);
nand U9988 (N_9988,N_9874,N_9800);
or U9989 (N_9989,N_9809,N_9824);
nand U9990 (N_9990,N_9848,N_9830);
or U9991 (N_9991,N_9873,N_9895);
nand U9992 (N_9992,N_9883,N_9834);
xor U9993 (N_9993,N_9838,N_9814);
or U9994 (N_9994,N_9853,N_9807);
and U9995 (N_9995,N_9896,N_9811);
or U9996 (N_9996,N_9819,N_9820);
and U9997 (N_9997,N_9826,N_9899);
or U9998 (N_9998,N_9838,N_9817);
or U9999 (N_9999,N_9895,N_9812);
and UO_0 (O_0,N_9982,N_9967);
and UO_1 (O_1,N_9992,N_9917);
nand UO_2 (O_2,N_9990,N_9945);
xor UO_3 (O_3,N_9959,N_9946);
nor UO_4 (O_4,N_9952,N_9941);
and UO_5 (O_5,N_9902,N_9920);
and UO_6 (O_6,N_9977,N_9943);
and UO_7 (O_7,N_9984,N_9954);
or UO_8 (O_8,N_9947,N_9928);
nand UO_9 (O_9,N_9924,N_9932);
xnor UO_10 (O_10,N_9972,N_9933);
nand UO_11 (O_11,N_9939,N_9968);
nand UO_12 (O_12,N_9971,N_9937);
or UO_13 (O_13,N_9911,N_9938);
nand UO_14 (O_14,N_9970,N_9997);
xor UO_15 (O_15,N_9960,N_9916);
and UO_16 (O_16,N_9994,N_9965);
or UO_17 (O_17,N_9958,N_9998);
nand UO_18 (O_18,N_9995,N_9950);
and UO_19 (O_19,N_9964,N_9904);
or UO_20 (O_20,N_9999,N_9951);
and UO_21 (O_21,N_9957,N_9989);
xor UO_22 (O_22,N_9907,N_9987);
nand UO_23 (O_23,N_9979,N_9931);
or UO_24 (O_24,N_9918,N_9905);
and UO_25 (O_25,N_9978,N_9973);
nand UO_26 (O_26,N_9988,N_9961);
nor UO_27 (O_27,N_9929,N_9956);
xor UO_28 (O_28,N_9925,N_9903);
nor UO_29 (O_29,N_9901,N_9930);
xnor UO_30 (O_30,N_9909,N_9923);
xor UO_31 (O_31,N_9940,N_9926);
nand UO_32 (O_32,N_9906,N_9975);
and UO_33 (O_33,N_9966,N_9948);
or UO_34 (O_34,N_9914,N_9969);
nand UO_35 (O_35,N_9983,N_9963);
and UO_36 (O_36,N_9900,N_9953);
nor UO_37 (O_37,N_9934,N_9910);
and UO_38 (O_38,N_9996,N_9936);
nand UO_39 (O_39,N_9974,N_9919);
nand UO_40 (O_40,N_9976,N_9955);
and UO_41 (O_41,N_9922,N_9962);
nand UO_42 (O_42,N_9993,N_9944);
nor UO_43 (O_43,N_9908,N_9991);
nor UO_44 (O_44,N_9949,N_9913);
nor UO_45 (O_45,N_9921,N_9912);
xnor UO_46 (O_46,N_9980,N_9942);
nor UO_47 (O_47,N_9927,N_9985);
or UO_48 (O_48,N_9935,N_9986);
and UO_49 (O_49,N_9915,N_9981);
or UO_50 (O_50,N_9985,N_9909);
xnor UO_51 (O_51,N_9980,N_9934);
and UO_52 (O_52,N_9918,N_9952);
or UO_53 (O_53,N_9957,N_9940);
and UO_54 (O_54,N_9946,N_9999);
or UO_55 (O_55,N_9951,N_9982);
and UO_56 (O_56,N_9901,N_9918);
nor UO_57 (O_57,N_9971,N_9918);
nand UO_58 (O_58,N_9969,N_9967);
or UO_59 (O_59,N_9972,N_9970);
xor UO_60 (O_60,N_9944,N_9916);
nor UO_61 (O_61,N_9919,N_9972);
xnor UO_62 (O_62,N_9938,N_9996);
nor UO_63 (O_63,N_9918,N_9972);
nor UO_64 (O_64,N_9999,N_9957);
or UO_65 (O_65,N_9969,N_9903);
or UO_66 (O_66,N_9978,N_9991);
and UO_67 (O_67,N_9952,N_9966);
nor UO_68 (O_68,N_9943,N_9976);
or UO_69 (O_69,N_9920,N_9927);
and UO_70 (O_70,N_9900,N_9949);
xnor UO_71 (O_71,N_9999,N_9971);
nor UO_72 (O_72,N_9914,N_9929);
xor UO_73 (O_73,N_9916,N_9990);
nand UO_74 (O_74,N_9920,N_9910);
or UO_75 (O_75,N_9994,N_9904);
nand UO_76 (O_76,N_9978,N_9977);
or UO_77 (O_77,N_9915,N_9908);
nand UO_78 (O_78,N_9960,N_9959);
or UO_79 (O_79,N_9976,N_9998);
or UO_80 (O_80,N_9963,N_9965);
nand UO_81 (O_81,N_9977,N_9976);
and UO_82 (O_82,N_9986,N_9978);
nor UO_83 (O_83,N_9979,N_9941);
nand UO_84 (O_84,N_9931,N_9919);
or UO_85 (O_85,N_9947,N_9932);
nor UO_86 (O_86,N_9933,N_9980);
nand UO_87 (O_87,N_9945,N_9904);
nand UO_88 (O_88,N_9911,N_9965);
nor UO_89 (O_89,N_9925,N_9928);
nor UO_90 (O_90,N_9915,N_9975);
and UO_91 (O_91,N_9905,N_9961);
xor UO_92 (O_92,N_9928,N_9924);
and UO_93 (O_93,N_9935,N_9980);
and UO_94 (O_94,N_9928,N_9993);
nand UO_95 (O_95,N_9930,N_9910);
nor UO_96 (O_96,N_9962,N_9981);
and UO_97 (O_97,N_9988,N_9918);
and UO_98 (O_98,N_9990,N_9969);
nor UO_99 (O_99,N_9928,N_9955);
nand UO_100 (O_100,N_9974,N_9985);
nor UO_101 (O_101,N_9986,N_9941);
or UO_102 (O_102,N_9950,N_9927);
nor UO_103 (O_103,N_9917,N_9982);
nor UO_104 (O_104,N_9982,N_9966);
nand UO_105 (O_105,N_9968,N_9974);
and UO_106 (O_106,N_9992,N_9934);
nor UO_107 (O_107,N_9993,N_9931);
nor UO_108 (O_108,N_9985,N_9970);
nand UO_109 (O_109,N_9989,N_9911);
and UO_110 (O_110,N_9936,N_9919);
nand UO_111 (O_111,N_9996,N_9994);
or UO_112 (O_112,N_9975,N_9945);
or UO_113 (O_113,N_9976,N_9944);
nand UO_114 (O_114,N_9924,N_9926);
nand UO_115 (O_115,N_9962,N_9943);
or UO_116 (O_116,N_9958,N_9927);
nor UO_117 (O_117,N_9914,N_9913);
nor UO_118 (O_118,N_9916,N_9933);
and UO_119 (O_119,N_9922,N_9906);
and UO_120 (O_120,N_9950,N_9961);
and UO_121 (O_121,N_9945,N_9993);
nor UO_122 (O_122,N_9966,N_9953);
or UO_123 (O_123,N_9937,N_9980);
and UO_124 (O_124,N_9975,N_9959);
and UO_125 (O_125,N_9931,N_9966);
xnor UO_126 (O_126,N_9909,N_9918);
nand UO_127 (O_127,N_9997,N_9948);
and UO_128 (O_128,N_9960,N_9996);
xor UO_129 (O_129,N_9963,N_9975);
or UO_130 (O_130,N_9915,N_9986);
nor UO_131 (O_131,N_9961,N_9924);
nand UO_132 (O_132,N_9996,N_9978);
and UO_133 (O_133,N_9984,N_9993);
and UO_134 (O_134,N_9915,N_9905);
and UO_135 (O_135,N_9948,N_9933);
or UO_136 (O_136,N_9981,N_9973);
or UO_137 (O_137,N_9977,N_9942);
and UO_138 (O_138,N_9903,N_9926);
nand UO_139 (O_139,N_9912,N_9985);
nor UO_140 (O_140,N_9911,N_9942);
or UO_141 (O_141,N_9948,N_9951);
or UO_142 (O_142,N_9948,N_9959);
nand UO_143 (O_143,N_9960,N_9922);
and UO_144 (O_144,N_9900,N_9973);
or UO_145 (O_145,N_9998,N_9985);
nor UO_146 (O_146,N_9915,N_9954);
or UO_147 (O_147,N_9903,N_9928);
nand UO_148 (O_148,N_9959,N_9992);
nand UO_149 (O_149,N_9946,N_9909);
and UO_150 (O_150,N_9969,N_9926);
xnor UO_151 (O_151,N_9963,N_9921);
nand UO_152 (O_152,N_9952,N_9982);
or UO_153 (O_153,N_9957,N_9971);
or UO_154 (O_154,N_9962,N_9902);
nand UO_155 (O_155,N_9913,N_9916);
nand UO_156 (O_156,N_9948,N_9931);
nand UO_157 (O_157,N_9912,N_9970);
and UO_158 (O_158,N_9982,N_9973);
nor UO_159 (O_159,N_9912,N_9933);
xnor UO_160 (O_160,N_9953,N_9994);
or UO_161 (O_161,N_9907,N_9944);
or UO_162 (O_162,N_9963,N_9973);
nand UO_163 (O_163,N_9939,N_9914);
nand UO_164 (O_164,N_9974,N_9918);
or UO_165 (O_165,N_9903,N_9937);
nor UO_166 (O_166,N_9990,N_9942);
and UO_167 (O_167,N_9970,N_9968);
nor UO_168 (O_168,N_9917,N_9908);
nor UO_169 (O_169,N_9969,N_9930);
xor UO_170 (O_170,N_9943,N_9931);
and UO_171 (O_171,N_9991,N_9926);
nor UO_172 (O_172,N_9944,N_9925);
and UO_173 (O_173,N_9976,N_9931);
or UO_174 (O_174,N_9923,N_9912);
or UO_175 (O_175,N_9954,N_9916);
nor UO_176 (O_176,N_9992,N_9952);
xnor UO_177 (O_177,N_9933,N_9915);
xor UO_178 (O_178,N_9928,N_9929);
nor UO_179 (O_179,N_9967,N_9935);
nor UO_180 (O_180,N_9946,N_9966);
and UO_181 (O_181,N_9982,N_9974);
or UO_182 (O_182,N_9906,N_9950);
or UO_183 (O_183,N_9918,N_9984);
nand UO_184 (O_184,N_9931,N_9906);
nor UO_185 (O_185,N_9921,N_9950);
or UO_186 (O_186,N_9964,N_9927);
nor UO_187 (O_187,N_9907,N_9905);
nand UO_188 (O_188,N_9936,N_9912);
or UO_189 (O_189,N_9958,N_9975);
nand UO_190 (O_190,N_9993,N_9902);
xor UO_191 (O_191,N_9904,N_9947);
or UO_192 (O_192,N_9919,N_9902);
or UO_193 (O_193,N_9978,N_9931);
or UO_194 (O_194,N_9908,N_9944);
or UO_195 (O_195,N_9961,N_9973);
nand UO_196 (O_196,N_9912,N_9934);
or UO_197 (O_197,N_9937,N_9973);
xor UO_198 (O_198,N_9900,N_9944);
nor UO_199 (O_199,N_9943,N_9981);
and UO_200 (O_200,N_9949,N_9946);
or UO_201 (O_201,N_9978,N_9950);
nor UO_202 (O_202,N_9913,N_9964);
nand UO_203 (O_203,N_9945,N_9925);
nand UO_204 (O_204,N_9972,N_9983);
or UO_205 (O_205,N_9989,N_9941);
nor UO_206 (O_206,N_9928,N_9941);
nor UO_207 (O_207,N_9997,N_9900);
and UO_208 (O_208,N_9997,N_9911);
xor UO_209 (O_209,N_9903,N_9944);
or UO_210 (O_210,N_9984,N_9904);
nor UO_211 (O_211,N_9958,N_9995);
nor UO_212 (O_212,N_9904,N_9911);
nor UO_213 (O_213,N_9921,N_9955);
nor UO_214 (O_214,N_9931,N_9934);
nor UO_215 (O_215,N_9983,N_9903);
nand UO_216 (O_216,N_9962,N_9908);
or UO_217 (O_217,N_9973,N_9908);
and UO_218 (O_218,N_9964,N_9915);
or UO_219 (O_219,N_9993,N_9913);
nor UO_220 (O_220,N_9986,N_9954);
nor UO_221 (O_221,N_9973,N_9906);
and UO_222 (O_222,N_9934,N_9998);
nand UO_223 (O_223,N_9923,N_9949);
or UO_224 (O_224,N_9900,N_9931);
xor UO_225 (O_225,N_9972,N_9930);
nor UO_226 (O_226,N_9957,N_9992);
or UO_227 (O_227,N_9922,N_9924);
nand UO_228 (O_228,N_9993,N_9991);
nand UO_229 (O_229,N_9919,N_9993);
or UO_230 (O_230,N_9977,N_9956);
nand UO_231 (O_231,N_9973,N_9948);
nand UO_232 (O_232,N_9998,N_9990);
and UO_233 (O_233,N_9941,N_9973);
xor UO_234 (O_234,N_9925,N_9974);
and UO_235 (O_235,N_9954,N_9979);
or UO_236 (O_236,N_9935,N_9902);
nand UO_237 (O_237,N_9903,N_9921);
nor UO_238 (O_238,N_9943,N_9988);
nand UO_239 (O_239,N_9979,N_9972);
nand UO_240 (O_240,N_9932,N_9944);
and UO_241 (O_241,N_9927,N_9901);
nand UO_242 (O_242,N_9992,N_9923);
nor UO_243 (O_243,N_9950,N_9977);
nor UO_244 (O_244,N_9916,N_9966);
xor UO_245 (O_245,N_9912,N_9919);
nor UO_246 (O_246,N_9945,N_9901);
or UO_247 (O_247,N_9967,N_9993);
and UO_248 (O_248,N_9909,N_9955);
nand UO_249 (O_249,N_9984,N_9975);
and UO_250 (O_250,N_9977,N_9923);
nand UO_251 (O_251,N_9980,N_9964);
and UO_252 (O_252,N_9975,N_9952);
nor UO_253 (O_253,N_9909,N_9949);
nor UO_254 (O_254,N_9929,N_9940);
nor UO_255 (O_255,N_9967,N_9949);
and UO_256 (O_256,N_9978,N_9939);
and UO_257 (O_257,N_9997,N_9989);
or UO_258 (O_258,N_9944,N_9905);
nand UO_259 (O_259,N_9976,N_9988);
nor UO_260 (O_260,N_9989,N_9991);
nand UO_261 (O_261,N_9967,N_9939);
nand UO_262 (O_262,N_9976,N_9952);
or UO_263 (O_263,N_9907,N_9947);
nand UO_264 (O_264,N_9988,N_9936);
xnor UO_265 (O_265,N_9912,N_9953);
xor UO_266 (O_266,N_9997,N_9976);
nor UO_267 (O_267,N_9999,N_9963);
nor UO_268 (O_268,N_9908,N_9986);
nor UO_269 (O_269,N_9997,N_9999);
or UO_270 (O_270,N_9983,N_9916);
nand UO_271 (O_271,N_9984,N_9934);
nor UO_272 (O_272,N_9939,N_9956);
nand UO_273 (O_273,N_9906,N_9988);
or UO_274 (O_274,N_9945,N_9955);
or UO_275 (O_275,N_9990,N_9947);
nand UO_276 (O_276,N_9989,N_9995);
nand UO_277 (O_277,N_9998,N_9922);
xnor UO_278 (O_278,N_9984,N_9933);
or UO_279 (O_279,N_9979,N_9920);
and UO_280 (O_280,N_9923,N_9921);
nor UO_281 (O_281,N_9953,N_9997);
and UO_282 (O_282,N_9973,N_9949);
or UO_283 (O_283,N_9958,N_9930);
xor UO_284 (O_284,N_9930,N_9944);
nor UO_285 (O_285,N_9940,N_9937);
nor UO_286 (O_286,N_9920,N_9931);
and UO_287 (O_287,N_9986,N_9961);
and UO_288 (O_288,N_9945,N_9916);
nor UO_289 (O_289,N_9989,N_9925);
or UO_290 (O_290,N_9927,N_9938);
or UO_291 (O_291,N_9961,N_9957);
nand UO_292 (O_292,N_9976,N_9907);
and UO_293 (O_293,N_9975,N_9914);
xnor UO_294 (O_294,N_9923,N_9929);
and UO_295 (O_295,N_9972,N_9996);
and UO_296 (O_296,N_9964,N_9962);
nand UO_297 (O_297,N_9918,N_9998);
and UO_298 (O_298,N_9927,N_9942);
nor UO_299 (O_299,N_9946,N_9923);
or UO_300 (O_300,N_9967,N_9917);
or UO_301 (O_301,N_9925,N_9955);
xnor UO_302 (O_302,N_9986,N_9952);
and UO_303 (O_303,N_9982,N_9984);
and UO_304 (O_304,N_9967,N_9958);
and UO_305 (O_305,N_9913,N_9983);
and UO_306 (O_306,N_9966,N_9935);
or UO_307 (O_307,N_9917,N_9932);
or UO_308 (O_308,N_9970,N_9978);
or UO_309 (O_309,N_9972,N_9990);
or UO_310 (O_310,N_9932,N_9954);
and UO_311 (O_311,N_9970,N_9960);
nand UO_312 (O_312,N_9988,N_9941);
or UO_313 (O_313,N_9943,N_9928);
and UO_314 (O_314,N_9961,N_9991);
nand UO_315 (O_315,N_9972,N_9939);
nor UO_316 (O_316,N_9944,N_9961);
nand UO_317 (O_317,N_9950,N_9925);
nor UO_318 (O_318,N_9903,N_9967);
and UO_319 (O_319,N_9969,N_9982);
nand UO_320 (O_320,N_9950,N_9979);
nor UO_321 (O_321,N_9946,N_9969);
or UO_322 (O_322,N_9913,N_9917);
nand UO_323 (O_323,N_9905,N_9929);
nor UO_324 (O_324,N_9906,N_9911);
nor UO_325 (O_325,N_9934,N_9920);
or UO_326 (O_326,N_9919,N_9982);
nor UO_327 (O_327,N_9936,N_9971);
or UO_328 (O_328,N_9980,N_9953);
nor UO_329 (O_329,N_9930,N_9934);
nand UO_330 (O_330,N_9925,N_9946);
and UO_331 (O_331,N_9977,N_9925);
and UO_332 (O_332,N_9957,N_9944);
nor UO_333 (O_333,N_9966,N_9940);
and UO_334 (O_334,N_9900,N_9906);
xnor UO_335 (O_335,N_9900,N_9959);
nor UO_336 (O_336,N_9911,N_9988);
nand UO_337 (O_337,N_9981,N_9929);
nor UO_338 (O_338,N_9919,N_9960);
nand UO_339 (O_339,N_9963,N_9998);
and UO_340 (O_340,N_9927,N_9956);
and UO_341 (O_341,N_9992,N_9930);
and UO_342 (O_342,N_9910,N_9968);
xnor UO_343 (O_343,N_9987,N_9961);
or UO_344 (O_344,N_9937,N_9936);
or UO_345 (O_345,N_9915,N_9938);
or UO_346 (O_346,N_9964,N_9939);
or UO_347 (O_347,N_9912,N_9938);
nor UO_348 (O_348,N_9965,N_9993);
or UO_349 (O_349,N_9960,N_9975);
or UO_350 (O_350,N_9919,N_9932);
and UO_351 (O_351,N_9918,N_9907);
or UO_352 (O_352,N_9943,N_9978);
and UO_353 (O_353,N_9944,N_9962);
and UO_354 (O_354,N_9996,N_9981);
nand UO_355 (O_355,N_9916,N_9971);
xnor UO_356 (O_356,N_9931,N_9956);
nor UO_357 (O_357,N_9976,N_9947);
or UO_358 (O_358,N_9997,N_9928);
nand UO_359 (O_359,N_9997,N_9924);
or UO_360 (O_360,N_9983,N_9909);
xor UO_361 (O_361,N_9930,N_9947);
nand UO_362 (O_362,N_9935,N_9997);
or UO_363 (O_363,N_9936,N_9982);
and UO_364 (O_364,N_9926,N_9933);
and UO_365 (O_365,N_9996,N_9989);
nor UO_366 (O_366,N_9929,N_9906);
and UO_367 (O_367,N_9930,N_9980);
xnor UO_368 (O_368,N_9990,N_9971);
nor UO_369 (O_369,N_9948,N_9993);
and UO_370 (O_370,N_9979,N_9917);
nand UO_371 (O_371,N_9988,N_9946);
or UO_372 (O_372,N_9915,N_9952);
and UO_373 (O_373,N_9934,N_9950);
or UO_374 (O_374,N_9953,N_9969);
and UO_375 (O_375,N_9948,N_9923);
or UO_376 (O_376,N_9982,N_9944);
nor UO_377 (O_377,N_9919,N_9929);
nor UO_378 (O_378,N_9913,N_9982);
nand UO_379 (O_379,N_9942,N_9906);
or UO_380 (O_380,N_9960,N_9976);
or UO_381 (O_381,N_9907,N_9957);
nand UO_382 (O_382,N_9946,N_9977);
nand UO_383 (O_383,N_9956,N_9992);
or UO_384 (O_384,N_9954,N_9960);
and UO_385 (O_385,N_9954,N_9944);
nor UO_386 (O_386,N_9951,N_9909);
and UO_387 (O_387,N_9920,N_9933);
or UO_388 (O_388,N_9970,N_9922);
xor UO_389 (O_389,N_9974,N_9955);
xnor UO_390 (O_390,N_9980,N_9939);
or UO_391 (O_391,N_9983,N_9937);
or UO_392 (O_392,N_9930,N_9929);
and UO_393 (O_393,N_9934,N_9990);
xnor UO_394 (O_394,N_9920,N_9963);
xnor UO_395 (O_395,N_9969,N_9950);
or UO_396 (O_396,N_9987,N_9904);
or UO_397 (O_397,N_9957,N_9938);
nand UO_398 (O_398,N_9952,N_9925);
nand UO_399 (O_399,N_9918,N_9944);
nor UO_400 (O_400,N_9975,N_9930);
nand UO_401 (O_401,N_9936,N_9952);
and UO_402 (O_402,N_9924,N_9984);
nor UO_403 (O_403,N_9914,N_9982);
or UO_404 (O_404,N_9943,N_9975);
nand UO_405 (O_405,N_9918,N_9910);
nor UO_406 (O_406,N_9914,N_9956);
nor UO_407 (O_407,N_9960,N_9998);
nor UO_408 (O_408,N_9904,N_9992);
or UO_409 (O_409,N_9906,N_9985);
xnor UO_410 (O_410,N_9981,N_9940);
nor UO_411 (O_411,N_9947,N_9934);
nor UO_412 (O_412,N_9964,N_9950);
and UO_413 (O_413,N_9943,N_9923);
nor UO_414 (O_414,N_9999,N_9953);
nand UO_415 (O_415,N_9937,N_9970);
nand UO_416 (O_416,N_9986,N_9955);
nand UO_417 (O_417,N_9962,N_9984);
or UO_418 (O_418,N_9942,N_9972);
nand UO_419 (O_419,N_9982,N_9907);
and UO_420 (O_420,N_9969,N_9959);
or UO_421 (O_421,N_9994,N_9941);
xnor UO_422 (O_422,N_9974,N_9931);
or UO_423 (O_423,N_9981,N_9917);
nand UO_424 (O_424,N_9949,N_9937);
nand UO_425 (O_425,N_9978,N_9904);
nand UO_426 (O_426,N_9939,N_9991);
nand UO_427 (O_427,N_9938,N_9921);
and UO_428 (O_428,N_9981,N_9916);
or UO_429 (O_429,N_9951,N_9922);
and UO_430 (O_430,N_9935,N_9993);
xnor UO_431 (O_431,N_9984,N_9927);
nand UO_432 (O_432,N_9907,N_9916);
nor UO_433 (O_433,N_9907,N_9941);
nand UO_434 (O_434,N_9938,N_9942);
nand UO_435 (O_435,N_9919,N_9986);
nand UO_436 (O_436,N_9938,N_9940);
and UO_437 (O_437,N_9915,N_9960);
nand UO_438 (O_438,N_9909,N_9973);
or UO_439 (O_439,N_9918,N_9996);
or UO_440 (O_440,N_9906,N_9940);
nand UO_441 (O_441,N_9947,N_9922);
and UO_442 (O_442,N_9927,N_9925);
and UO_443 (O_443,N_9948,N_9928);
nand UO_444 (O_444,N_9963,N_9969);
nor UO_445 (O_445,N_9917,N_9914);
or UO_446 (O_446,N_9953,N_9996);
and UO_447 (O_447,N_9993,N_9974);
or UO_448 (O_448,N_9960,N_9943);
nand UO_449 (O_449,N_9981,N_9970);
nor UO_450 (O_450,N_9956,N_9923);
xor UO_451 (O_451,N_9915,N_9945);
or UO_452 (O_452,N_9955,N_9953);
and UO_453 (O_453,N_9948,N_9922);
and UO_454 (O_454,N_9933,N_9981);
or UO_455 (O_455,N_9968,N_9994);
nor UO_456 (O_456,N_9991,N_9960);
and UO_457 (O_457,N_9938,N_9901);
nand UO_458 (O_458,N_9910,N_9921);
nand UO_459 (O_459,N_9928,N_9915);
and UO_460 (O_460,N_9944,N_9933);
nand UO_461 (O_461,N_9975,N_9933);
and UO_462 (O_462,N_9977,N_9964);
nand UO_463 (O_463,N_9958,N_9956);
xor UO_464 (O_464,N_9934,N_9906);
nor UO_465 (O_465,N_9917,N_9926);
nand UO_466 (O_466,N_9934,N_9985);
nand UO_467 (O_467,N_9948,N_9968);
nor UO_468 (O_468,N_9966,N_9908);
and UO_469 (O_469,N_9971,N_9923);
or UO_470 (O_470,N_9961,N_9910);
xnor UO_471 (O_471,N_9974,N_9983);
nand UO_472 (O_472,N_9987,N_9947);
nor UO_473 (O_473,N_9906,N_9926);
nand UO_474 (O_474,N_9978,N_9920);
and UO_475 (O_475,N_9950,N_9919);
nand UO_476 (O_476,N_9952,N_9932);
nand UO_477 (O_477,N_9993,N_9986);
nand UO_478 (O_478,N_9937,N_9911);
nand UO_479 (O_479,N_9991,N_9932);
nand UO_480 (O_480,N_9987,N_9909);
nand UO_481 (O_481,N_9902,N_9971);
or UO_482 (O_482,N_9953,N_9904);
nor UO_483 (O_483,N_9978,N_9952);
and UO_484 (O_484,N_9946,N_9950);
nor UO_485 (O_485,N_9917,N_9969);
and UO_486 (O_486,N_9913,N_9937);
or UO_487 (O_487,N_9933,N_9939);
or UO_488 (O_488,N_9905,N_9964);
nor UO_489 (O_489,N_9975,N_9938);
and UO_490 (O_490,N_9951,N_9913);
nor UO_491 (O_491,N_9947,N_9965);
xor UO_492 (O_492,N_9962,N_9976);
or UO_493 (O_493,N_9966,N_9936);
and UO_494 (O_494,N_9977,N_9958);
nor UO_495 (O_495,N_9960,N_9949);
nor UO_496 (O_496,N_9906,N_9943);
nor UO_497 (O_497,N_9998,N_9904);
and UO_498 (O_498,N_9936,N_9908);
xnor UO_499 (O_499,N_9955,N_9908);
xor UO_500 (O_500,N_9940,N_9922);
and UO_501 (O_501,N_9950,N_9985);
and UO_502 (O_502,N_9941,N_9980);
nand UO_503 (O_503,N_9974,N_9920);
nand UO_504 (O_504,N_9931,N_9947);
or UO_505 (O_505,N_9971,N_9987);
or UO_506 (O_506,N_9976,N_9911);
xor UO_507 (O_507,N_9953,N_9975);
or UO_508 (O_508,N_9973,N_9983);
nor UO_509 (O_509,N_9969,N_9913);
or UO_510 (O_510,N_9925,N_9931);
nand UO_511 (O_511,N_9987,N_9985);
nor UO_512 (O_512,N_9927,N_9910);
or UO_513 (O_513,N_9963,N_9929);
and UO_514 (O_514,N_9952,N_9906);
nor UO_515 (O_515,N_9930,N_9988);
or UO_516 (O_516,N_9913,N_9959);
or UO_517 (O_517,N_9908,N_9951);
nor UO_518 (O_518,N_9960,N_9931);
or UO_519 (O_519,N_9938,N_9987);
nor UO_520 (O_520,N_9950,N_9928);
nand UO_521 (O_521,N_9956,N_9959);
or UO_522 (O_522,N_9908,N_9970);
or UO_523 (O_523,N_9923,N_9987);
and UO_524 (O_524,N_9955,N_9939);
nand UO_525 (O_525,N_9969,N_9975);
nor UO_526 (O_526,N_9941,N_9963);
nand UO_527 (O_527,N_9902,N_9943);
or UO_528 (O_528,N_9989,N_9910);
xnor UO_529 (O_529,N_9974,N_9997);
or UO_530 (O_530,N_9969,N_9974);
and UO_531 (O_531,N_9928,N_9931);
and UO_532 (O_532,N_9988,N_9905);
or UO_533 (O_533,N_9915,N_9935);
nor UO_534 (O_534,N_9986,N_9921);
nand UO_535 (O_535,N_9957,N_9972);
nand UO_536 (O_536,N_9974,N_9901);
or UO_537 (O_537,N_9962,N_9967);
xnor UO_538 (O_538,N_9988,N_9989);
nand UO_539 (O_539,N_9991,N_9970);
nand UO_540 (O_540,N_9988,N_9919);
and UO_541 (O_541,N_9921,N_9919);
or UO_542 (O_542,N_9904,N_9968);
and UO_543 (O_543,N_9964,N_9948);
nor UO_544 (O_544,N_9934,N_9921);
nor UO_545 (O_545,N_9946,N_9975);
nand UO_546 (O_546,N_9958,N_9939);
and UO_547 (O_547,N_9949,N_9943);
or UO_548 (O_548,N_9940,N_9980);
nand UO_549 (O_549,N_9933,N_9959);
or UO_550 (O_550,N_9977,N_9984);
nand UO_551 (O_551,N_9971,N_9939);
or UO_552 (O_552,N_9915,N_9969);
nor UO_553 (O_553,N_9968,N_9944);
and UO_554 (O_554,N_9911,N_9925);
nor UO_555 (O_555,N_9911,N_9959);
and UO_556 (O_556,N_9905,N_9937);
nand UO_557 (O_557,N_9988,N_9904);
and UO_558 (O_558,N_9967,N_9920);
or UO_559 (O_559,N_9900,N_9912);
nor UO_560 (O_560,N_9989,N_9931);
nor UO_561 (O_561,N_9911,N_9971);
or UO_562 (O_562,N_9913,N_9903);
xnor UO_563 (O_563,N_9923,N_9933);
or UO_564 (O_564,N_9989,N_9958);
nand UO_565 (O_565,N_9953,N_9961);
nand UO_566 (O_566,N_9994,N_9910);
or UO_567 (O_567,N_9989,N_9915);
or UO_568 (O_568,N_9987,N_9905);
nor UO_569 (O_569,N_9993,N_9912);
nand UO_570 (O_570,N_9922,N_9993);
or UO_571 (O_571,N_9940,N_9925);
or UO_572 (O_572,N_9942,N_9922);
and UO_573 (O_573,N_9980,N_9994);
nand UO_574 (O_574,N_9971,N_9984);
and UO_575 (O_575,N_9929,N_9954);
nand UO_576 (O_576,N_9931,N_9942);
xor UO_577 (O_577,N_9945,N_9976);
nand UO_578 (O_578,N_9952,N_9944);
nor UO_579 (O_579,N_9987,N_9978);
xnor UO_580 (O_580,N_9973,N_9956);
or UO_581 (O_581,N_9916,N_9965);
nand UO_582 (O_582,N_9972,N_9902);
or UO_583 (O_583,N_9970,N_9924);
nor UO_584 (O_584,N_9983,N_9956);
and UO_585 (O_585,N_9916,N_9900);
nand UO_586 (O_586,N_9987,N_9921);
nand UO_587 (O_587,N_9923,N_9963);
and UO_588 (O_588,N_9942,N_9998);
and UO_589 (O_589,N_9936,N_9923);
nand UO_590 (O_590,N_9914,N_9996);
nor UO_591 (O_591,N_9902,N_9966);
nand UO_592 (O_592,N_9941,N_9915);
nand UO_593 (O_593,N_9940,N_9961);
nor UO_594 (O_594,N_9900,N_9919);
and UO_595 (O_595,N_9986,N_9959);
and UO_596 (O_596,N_9958,N_9993);
nor UO_597 (O_597,N_9995,N_9931);
or UO_598 (O_598,N_9923,N_9917);
nor UO_599 (O_599,N_9923,N_9960);
nand UO_600 (O_600,N_9966,N_9930);
nand UO_601 (O_601,N_9966,N_9947);
nor UO_602 (O_602,N_9941,N_9987);
nor UO_603 (O_603,N_9904,N_9993);
and UO_604 (O_604,N_9999,N_9989);
nand UO_605 (O_605,N_9903,N_9966);
and UO_606 (O_606,N_9935,N_9918);
or UO_607 (O_607,N_9907,N_9930);
xnor UO_608 (O_608,N_9979,N_9923);
or UO_609 (O_609,N_9949,N_9982);
xor UO_610 (O_610,N_9914,N_9902);
xor UO_611 (O_611,N_9913,N_9973);
nor UO_612 (O_612,N_9968,N_9936);
nor UO_613 (O_613,N_9927,N_9931);
xor UO_614 (O_614,N_9905,N_9930);
or UO_615 (O_615,N_9902,N_9936);
or UO_616 (O_616,N_9986,N_9937);
xor UO_617 (O_617,N_9984,N_9963);
nor UO_618 (O_618,N_9928,N_9901);
and UO_619 (O_619,N_9976,N_9966);
and UO_620 (O_620,N_9943,N_9922);
or UO_621 (O_621,N_9900,N_9902);
nor UO_622 (O_622,N_9965,N_9904);
nor UO_623 (O_623,N_9947,N_9901);
and UO_624 (O_624,N_9973,N_9952);
nor UO_625 (O_625,N_9905,N_9983);
nand UO_626 (O_626,N_9994,N_9985);
and UO_627 (O_627,N_9969,N_9907);
and UO_628 (O_628,N_9989,N_9927);
nand UO_629 (O_629,N_9925,N_9951);
xor UO_630 (O_630,N_9995,N_9986);
and UO_631 (O_631,N_9910,N_9948);
and UO_632 (O_632,N_9962,N_9928);
nand UO_633 (O_633,N_9921,N_9909);
and UO_634 (O_634,N_9993,N_9961);
or UO_635 (O_635,N_9957,N_9959);
or UO_636 (O_636,N_9983,N_9976);
and UO_637 (O_637,N_9914,N_9945);
xnor UO_638 (O_638,N_9975,N_9993);
nor UO_639 (O_639,N_9914,N_9957);
nand UO_640 (O_640,N_9927,N_9988);
xor UO_641 (O_641,N_9914,N_9989);
xor UO_642 (O_642,N_9937,N_9984);
nand UO_643 (O_643,N_9976,N_9927);
and UO_644 (O_644,N_9914,N_9941);
nor UO_645 (O_645,N_9982,N_9989);
or UO_646 (O_646,N_9989,N_9922);
or UO_647 (O_647,N_9958,N_9914);
nand UO_648 (O_648,N_9910,N_9960);
nand UO_649 (O_649,N_9930,N_9902);
and UO_650 (O_650,N_9979,N_9904);
nor UO_651 (O_651,N_9993,N_9988);
nor UO_652 (O_652,N_9989,N_9990);
xor UO_653 (O_653,N_9979,N_9927);
nor UO_654 (O_654,N_9914,N_9998);
or UO_655 (O_655,N_9926,N_9970);
and UO_656 (O_656,N_9938,N_9982);
nand UO_657 (O_657,N_9995,N_9926);
and UO_658 (O_658,N_9975,N_9954);
or UO_659 (O_659,N_9943,N_9979);
and UO_660 (O_660,N_9981,N_9952);
nand UO_661 (O_661,N_9928,N_9912);
nand UO_662 (O_662,N_9961,N_9965);
and UO_663 (O_663,N_9997,N_9950);
xnor UO_664 (O_664,N_9963,N_9914);
xor UO_665 (O_665,N_9936,N_9934);
and UO_666 (O_666,N_9916,N_9973);
nor UO_667 (O_667,N_9963,N_9926);
nor UO_668 (O_668,N_9934,N_9904);
or UO_669 (O_669,N_9914,N_9930);
and UO_670 (O_670,N_9901,N_9983);
nor UO_671 (O_671,N_9934,N_9949);
and UO_672 (O_672,N_9979,N_9929);
or UO_673 (O_673,N_9936,N_9994);
nand UO_674 (O_674,N_9989,N_9965);
and UO_675 (O_675,N_9940,N_9975);
xnor UO_676 (O_676,N_9924,N_9909);
or UO_677 (O_677,N_9926,N_9986);
xnor UO_678 (O_678,N_9917,N_9938);
and UO_679 (O_679,N_9935,N_9946);
and UO_680 (O_680,N_9938,N_9922);
nor UO_681 (O_681,N_9993,N_9956);
nand UO_682 (O_682,N_9902,N_9978);
or UO_683 (O_683,N_9972,N_9964);
nor UO_684 (O_684,N_9943,N_9911);
or UO_685 (O_685,N_9998,N_9973);
nand UO_686 (O_686,N_9963,N_9925);
or UO_687 (O_687,N_9947,N_9926);
nand UO_688 (O_688,N_9990,N_9986);
nand UO_689 (O_689,N_9922,N_9917);
nand UO_690 (O_690,N_9981,N_9982);
or UO_691 (O_691,N_9915,N_9903);
nor UO_692 (O_692,N_9930,N_9951);
nor UO_693 (O_693,N_9985,N_9938);
and UO_694 (O_694,N_9972,N_9952);
nor UO_695 (O_695,N_9908,N_9928);
nand UO_696 (O_696,N_9977,N_9952);
nor UO_697 (O_697,N_9940,N_9928);
nand UO_698 (O_698,N_9985,N_9908);
nand UO_699 (O_699,N_9965,N_9906);
or UO_700 (O_700,N_9984,N_9987);
and UO_701 (O_701,N_9942,N_9941);
nand UO_702 (O_702,N_9926,N_9942);
xnor UO_703 (O_703,N_9949,N_9952);
xor UO_704 (O_704,N_9967,N_9979);
nand UO_705 (O_705,N_9939,N_9910);
and UO_706 (O_706,N_9953,N_9910);
nand UO_707 (O_707,N_9936,N_9978);
nand UO_708 (O_708,N_9992,N_9908);
nor UO_709 (O_709,N_9975,N_9991);
nand UO_710 (O_710,N_9939,N_9919);
nand UO_711 (O_711,N_9924,N_9966);
nor UO_712 (O_712,N_9932,N_9972);
nor UO_713 (O_713,N_9984,N_9961);
or UO_714 (O_714,N_9909,N_9957);
nor UO_715 (O_715,N_9937,N_9944);
nand UO_716 (O_716,N_9948,N_9919);
nor UO_717 (O_717,N_9981,N_9999);
and UO_718 (O_718,N_9983,N_9944);
or UO_719 (O_719,N_9974,N_9991);
and UO_720 (O_720,N_9900,N_9961);
nor UO_721 (O_721,N_9916,N_9905);
nor UO_722 (O_722,N_9998,N_9936);
nand UO_723 (O_723,N_9915,N_9940);
and UO_724 (O_724,N_9951,N_9967);
nand UO_725 (O_725,N_9935,N_9933);
nor UO_726 (O_726,N_9912,N_9998);
nand UO_727 (O_727,N_9954,N_9969);
or UO_728 (O_728,N_9908,N_9958);
and UO_729 (O_729,N_9930,N_9953);
or UO_730 (O_730,N_9934,N_9999);
or UO_731 (O_731,N_9972,N_9969);
or UO_732 (O_732,N_9990,N_9912);
xnor UO_733 (O_733,N_9934,N_9964);
xor UO_734 (O_734,N_9941,N_9910);
nand UO_735 (O_735,N_9931,N_9913);
nor UO_736 (O_736,N_9937,N_9958);
nor UO_737 (O_737,N_9953,N_9937);
or UO_738 (O_738,N_9943,N_9947);
nand UO_739 (O_739,N_9915,N_9943);
nor UO_740 (O_740,N_9940,N_9901);
nand UO_741 (O_741,N_9970,N_9983);
xor UO_742 (O_742,N_9992,N_9999);
nor UO_743 (O_743,N_9928,N_9918);
nand UO_744 (O_744,N_9990,N_9961);
and UO_745 (O_745,N_9938,N_9959);
and UO_746 (O_746,N_9969,N_9966);
nand UO_747 (O_747,N_9969,N_9916);
and UO_748 (O_748,N_9965,N_9957);
or UO_749 (O_749,N_9901,N_9997);
and UO_750 (O_750,N_9982,N_9965);
and UO_751 (O_751,N_9974,N_9937);
nor UO_752 (O_752,N_9923,N_9991);
xnor UO_753 (O_753,N_9990,N_9997);
nor UO_754 (O_754,N_9951,N_9968);
or UO_755 (O_755,N_9951,N_9935);
or UO_756 (O_756,N_9965,N_9962);
or UO_757 (O_757,N_9908,N_9945);
nor UO_758 (O_758,N_9968,N_9964);
nand UO_759 (O_759,N_9942,N_9946);
and UO_760 (O_760,N_9929,N_9913);
or UO_761 (O_761,N_9933,N_9921);
or UO_762 (O_762,N_9906,N_9972);
or UO_763 (O_763,N_9969,N_9978);
nor UO_764 (O_764,N_9910,N_9979);
xor UO_765 (O_765,N_9965,N_9903);
and UO_766 (O_766,N_9979,N_9928);
nand UO_767 (O_767,N_9950,N_9902);
xor UO_768 (O_768,N_9913,N_9955);
or UO_769 (O_769,N_9983,N_9946);
and UO_770 (O_770,N_9946,N_9912);
or UO_771 (O_771,N_9971,N_9955);
nand UO_772 (O_772,N_9935,N_9970);
nor UO_773 (O_773,N_9955,N_9964);
and UO_774 (O_774,N_9931,N_9982);
or UO_775 (O_775,N_9968,N_9982);
and UO_776 (O_776,N_9942,N_9912);
nand UO_777 (O_777,N_9968,N_9992);
nand UO_778 (O_778,N_9992,N_9919);
nor UO_779 (O_779,N_9990,N_9907);
or UO_780 (O_780,N_9999,N_9925);
nor UO_781 (O_781,N_9914,N_9901);
or UO_782 (O_782,N_9949,N_9917);
and UO_783 (O_783,N_9989,N_9956);
or UO_784 (O_784,N_9940,N_9993);
nor UO_785 (O_785,N_9907,N_9983);
nor UO_786 (O_786,N_9978,N_9971);
or UO_787 (O_787,N_9942,N_9987);
or UO_788 (O_788,N_9925,N_9932);
or UO_789 (O_789,N_9947,N_9986);
or UO_790 (O_790,N_9992,N_9966);
nor UO_791 (O_791,N_9906,N_9982);
and UO_792 (O_792,N_9942,N_9964);
xnor UO_793 (O_793,N_9963,N_9907);
nand UO_794 (O_794,N_9905,N_9966);
nor UO_795 (O_795,N_9923,N_9904);
xor UO_796 (O_796,N_9962,N_9992);
nor UO_797 (O_797,N_9974,N_9970);
xor UO_798 (O_798,N_9972,N_9937);
xnor UO_799 (O_799,N_9915,N_9910);
xnor UO_800 (O_800,N_9944,N_9902);
nand UO_801 (O_801,N_9912,N_9916);
and UO_802 (O_802,N_9953,N_9947);
or UO_803 (O_803,N_9914,N_9908);
nor UO_804 (O_804,N_9935,N_9921);
xnor UO_805 (O_805,N_9963,N_9942);
and UO_806 (O_806,N_9938,N_9952);
nor UO_807 (O_807,N_9915,N_9924);
or UO_808 (O_808,N_9946,N_9931);
and UO_809 (O_809,N_9989,N_9921);
xor UO_810 (O_810,N_9919,N_9958);
or UO_811 (O_811,N_9981,N_9961);
nand UO_812 (O_812,N_9984,N_9922);
nor UO_813 (O_813,N_9928,N_9944);
nand UO_814 (O_814,N_9959,N_9994);
or UO_815 (O_815,N_9991,N_9979);
nand UO_816 (O_816,N_9918,N_9919);
nor UO_817 (O_817,N_9945,N_9982);
or UO_818 (O_818,N_9987,N_9946);
nand UO_819 (O_819,N_9975,N_9917);
nand UO_820 (O_820,N_9935,N_9942);
nor UO_821 (O_821,N_9930,N_9917);
and UO_822 (O_822,N_9937,N_9962);
and UO_823 (O_823,N_9968,N_9999);
or UO_824 (O_824,N_9979,N_9976);
and UO_825 (O_825,N_9993,N_9973);
or UO_826 (O_826,N_9919,N_9963);
xnor UO_827 (O_827,N_9932,N_9913);
xor UO_828 (O_828,N_9959,N_9963);
and UO_829 (O_829,N_9940,N_9988);
nand UO_830 (O_830,N_9961,N_9964);
xor UO_831 (O_831,N_9905,N_9957);
xor UO_832 (O_832,N_9908,N_9998);
nor UO_833 (O_833,N_9960,N_9990);
or UO_834 (O_834,N_9997,N_9977);
and UO_835 (O_835,N_9957,N_9995);
or UO_836 (O_836,N_9969,N_9976);
nor UO_837 (O_837,N_9939,N_9931);
xor UO_838 (O_838,N_9914,N_9947);
xnor UO_839 (O_839,N_9995,N_9945);
nand UO_840 (O_840,N_9959,N_9947);
and UO_841 (O_841,N_9964,N_9921);
xnor UO_842 (O_842,N_9927,N_9951);
and UO_843 (O_843,N_9915,N_9968);
and UO_844 (O_844,N_9909,N_9901);
or UO_845 (O_845,N_9950,N_9962);
xnor UO_846 (O_846,N_9990,N_9999);
nor UO_847 (O_847,N_9938,N_9960);
and UO_848 (O_848,N_9931,N_9938);
nor UO_849 (O_849,N_9986,N_9992);
nor UO_850 (O_850,N_9930,N_9932);
or UO_851 (O_851,N_9969,N_9927);
nor UO_852 (O_852,N_9941,N_9956);
nand UO_853 (O_853,N_9961,N_9979);
and UO_854 (O_854,N_9975,N_9948);
nor UO_855 (O_855,N_9900,N_9913);
nand UO_856 (O_856,N_9926,N_9916);
nor UO_857 (O_857,N_9914,N_9986);
nand UO_858 (O_858,N_9952,N_9907);
or UO_859 (O_859,N_9907,N_9946);
nand UO_860 (O_860,N_9947,N_9929);
or UO_861 (O_861,N_9976,N_9926);
and UO_862 (O_862,N_9983,N_9960);
nor UO_863 (O_863,N_9918,N_9989);
or UO_864 (O_864,N_9989,N_9980);
or UO_865 (O_865,N_9929,N_9909);
and UO_866 (O_866,N_9901,N_9908);
xnor UO_867 (O_867,N_9922,N_9918);
or UO_868 (O_868,N_9955,N_9918);
xor UO_869 (O_869,N_9912,N_9927);
nor UO_870 (O_870,N_9967,N_9919);
nor UO_871 (O_871,N_9957,N_9925);
nor UO_872 (O_872,N_9905,N_9986);
nand UO_873 (O_873,N_9945,N_9992);
or UO_874 (O_874,N_9992,N_9915);
nor UO_875 (O_875,N_9908,N_9939);
and UO_876 (O_876,N_9928,N_9951);
nor UO_877 (O_877,N_9989,N_9979);
nand UO_878 (O_878,N_9954,N_9938);
nor UO_879 (O_879,N_9961,N_9983);
nor UO_880 (O_880,N_9955,N_9949);
and UO_881 (O_881,N_9915,N_9976);
or UO_882 (O_882,N_9962,N_9989);
nand UO_883 (O_883,N_9951,N_9969);
and UO_884 (O_884,N_9973,N_9925);
nand UO_885 (O_885,N_9931,N_9967);
xor UO_886 (O_886,N_9929,N_9942);
and UO_887 (O_887,N_9923,N_9914);
nand UO_888 (O_888,N_9924,N_9993);
or UO_889 (O_889,N_9916,N_9923);
nand UO_890 (O_890,N_9991,N_9921);
or UO_891 (O_891,N_9998,N_9926);
nor UO_892 (O_892,N_9912,N_9944);
and UO_893 (O_893,N_9956,N_9930);
or UO_894 (O_894,N_9926,N_9945);
and UO_895 (O_895,N_9930,N_9909);
nor UO_896 (O_896,N_9919,N_9983);
or UO_897 (O_897,N_9928,N_9973);
xor UO_898 (O_898,N_9903,N_9941);
xnor UO_899 (O_899,N_9956,N_9922);
or UO_900 (O_900,N_9917,N_9928);
nand UO_901 (O_901,N_9998,N_9978);
and UO_902 (O_902,N_9922,N_9927);
nor UO_903 (O_903,N_9940,N_9943);
nand UO_904 (O_904,N_9940,N_9909);
and UO_905 (O_905,N_9933,N_9936);
or UO_906 (O_906,N_9936,N_9926);
and UO_907 (O_907,N_9991,N_9919);
nand UO_908 (O_908,N_9910,N_9984);
and UO_909 (O_909,N_9910,N_9903);
nand UO_910 (O_910,N_9968,N_9928);
nand UO_911 (O_911,N_9986,N_9907);
or UO_912 (O_912,N_9942,N_9959);
xnor UO_913 (O_913,N_9968,N_9953);
nand UO_914 (O_914,N_9992,N_9921);
nor UO_915 (O_915,N_9940,N_9954);
nor UO_916 (O_916,N_9984,N_9994);
and UO_917 (O_917,N_9953,N_9903);
and UO_918 (O_918,N_9941,N_9975);
and UO_919 (O_919,N_9940,N_9955);
xnor UO_920 (O_920,N_9924,N_9988);
nor UO_921 (O_921,N_9996,N_9916);
nor UO_922 (O_922,N_9904,N_9913);
nor UO_923 (O_923,N_9927,N_9929);
or UO_924 (O_924,N_9982,N_9933);
and UO_925 (O_925,N_9904,N_9963);
and UO_926 (O_926,N_9952,N_9924);
and UO_927 (O_927,N_9991,N_9913);
nor UO_928 (O_928,N_9977,N_9915);
or UO_929 (O_929,N_9944,N_9977);
and UO_930 (O_930,N_9908,N_9996);
and UO_931 (O_931,N_9986,N_9975);
nand UO_932 (O_932,N_9910,N_9986);
nand UO_933 (O_933,N_9964,N_9975);
or UO_934 (O_934,N_9964,N_9982);
nand UO_935 (O_935,N_9911,N_9903);
nor UO_936 (O_936,N_9995,N_9936);
nand UO_937 (O_937,N_9983,N_9985);
nor UO_938 (O_938,N_9931,N_9958);
and UO_939 (O_939,N_9905,N_9994);
nor UO_940 (O_940,N_9934,N_9908);
or UO_941 (O_941,N_9913,N_9960);
or UO_942 (O_942,N_9961,N_9938);
or UO_943 (O_943,N_9927,N_9940);
nand UO_944 (O_944,N_9931,N_9954);
xnor UO_945 (O_945,N_9954,N_9934);
and UO_946 (O_946,N_9937,N_9982);
or UO_947 (O_947,N_9901,N_9985);
nand UO_948 (O_948,N_9999,N_9924);
nand UO_949 (O_949,N_9995,N_9955);
or UO_950 (O_950,N_9979,N_9934);
and UO_951 (O_951,N_9992,N_9984);
or UO_952 (O_952,N_9989,N_9908);
or UO_953 (O_953,N_9956,N_9974);
nor UO_954 (O_954,N_9963,N_9924);
or UO_955 (O_955,N_9934,N_9933);
nand UO_956 (O_956,N_9928,N_9991);
and UO_957 (O_957,N_9943,N_9992);
nand UO_958 (O_958,N_9912,N_9996);
nor UO_959 (O_959,N_9925,N_9993);
nand UO_960 (O_960,N_9956,N_9943);
and UO_961 (O_961,N_9987,N_9916);
and UO_962 (O_962,N_9965,N_9941);
or UO_963 (O_963,N_9946,N_9964);
and UO_964 (O_964,N_9911,N_9999);
and UO_965 (O_965,N_9937,N_9912);
and UO_966 (O_966,N_9941,N_9925);
or UO_967 (O_967,N_9955,N_9997);
or UO_968 (O_968,N_9977,N_9917);
xor UO_969 (O_969,N_9950,N_9901);
or UO_970 (O_970,N_9996,N_9901);
or UO_971 (O_971,N_9960,N_9993);
xnor UO_972 (O_972,N_9938,N_9953);
nand UO_973 (O_973,N_9946,N_9914);
and UO_974 (O_974,N_9973,N_9945);
nor UO_975 (O_975,N_9935,N_9911);
or UO_976 (O_976,N_9959,N_9936);
and UO_977 (O_977,N_9926,N_9931);
or UO_978 (O_978,N_9968,N_9963);
or UO_979 (O_979,N_9957,N_9922);
xor UO_980 (O_980,N_9943,N_9920);
nand UO_981 (O_981,N_9907,N_9927);
and UO_982 (O_982,N_9988,N_9981);
nor UO_983 (O_983,N_9992,N_9989);
nor UO_984 (O_984,N_9932,N_9955);
nand UO_985 (O_985,N_9990,N_9957);
nand UO_986 (O_986,N_9948,N_9958);
nor UO_987 (O_987,N_9965,N_9952);
nor UO_988 (O_988,N_9958,N_9980);
or UO_989 (O_989,N_9924,N_9901);
or UO_990 (O_990,N_9926,N_9901);
nor UO_991 (O_991,N_9946,N_9976);
and UO_992 (O_992,N_9966,N_9938);
and UO_993 (O_993,N_9933,N_9999);
xnor UO_994 (O_994,N_9956,N_9998);
nor UO_995 (O_995,N_9911,N_9928);
nand UO_996 (O_996,N_9912,N_9969);
xnor UO_997 (O_997,N_9932,N_9988);
and UO_998 (O_998,N_9927,N_9911);
xnor UO_999 (O_999,N_9949,N_9904);
or UO_1000 (O_1000,N_9979,N_9918);
nand UO_1001 (O_1001,N_9904,N_9909);
or UO_1002 (O_1002,N_9962,N_9987);
and UO_1003 (O_1003,N_9919,N_9914);
and UO_1004 (O_1004,N_9973,N_9921);
and UO_1005 (O_1005,N_9910,N_9914);
and UO_1006 (O_1006,N_9936,N_9925);
and UO_1007 (O_1007,N_9944,N_9956);
nor UO_1008 (O_1008,N_9924,N_9985);
nor UO_1009 (O_1009,N_9911,N_9978);
or UO_1010 (O_1010,N_9943,N_9991);
nor UO_1011 (O_1011,N_9978,N_9921);
nand UO_1012 (O_1012,N_9971,N_9982);
nor UO_1013 (O_1013,N_9997,N_9905);
nand UO_1014 (O_1014,N_9994,N_9971);
or UO_1015 (O_1015,N_9927,N_9986);
nor UO_1016 (O_1016,N_9983,N_9928);
xor UO_1017 (O_1017,N_9936,N_9975);
nand UO_1018 (O_1018,N_9986,N_9943);
nand UO_1019 (O_1019,N_9947,N_9982);
xor UO_1020 (O_1020,N_9924,N_9931);
nor UO_1021 (O_1021,N_9933,N_9922);
nand UO_1022 (O_1022,N_9908,N_9969);
or UO_1023 (O_1023,N_9901,N_9964);
nor UO_1024 (O_1024,N_9931,N_9937);
or UO_1025 (O_1025,N_9941,N_9947);
nand UO_1026 (O_1026,N_9937,N_9902);
nor UO_1027 (O_1027,N_9938,N_9919);
nand UO_1028 (O_1028,N_9961,N_9975);
nand UO_1029 (O_1029,N_9956,N_9980);
or UO_1030 (O_1030,N_9963,N_9939);
nand UO_1031 (O_1031,N_9992,N_9922);
xnor UO_1032 (O_1032,N_9975,N_9947);
nor UO_1033 (O_1033,N_9935,N_9999);
nand UO_1034 (O_1034,N_9962,N_9936);
or UO_1035 (O_1035,N_9971,N_9991);
nor UO_1036 (O_1036,N_9985,N_9996);
nand UO_1037 (O_1037,N_9960,N_9940);
nor UO_1038 (O_1038,N_9985,N_9956);
xnor UO_1039 (O_1039,N_9960,N_9906);
or UO_1040 (O_1040,N_9926,N_9966);
nor UO_1041 (O_1041,N_9991,N_9986);
or UO_1042 (O_1042,N_9987,N_9968);
and UO_1043 (O_1043,N_9949,N_9997);
and UO_1044 (O_1044,N_9946,N_9910);
xor UO_1045 (O_1045,N_9929,N_9917);
or UO_1046 (O_1046,N_9907,N_9950);
and UO_1047 (O_1047,N_9964,N_9936);
and UO_1048 (O_1048,N_9975,N_9919);
nand UO_1049 (O_1049,N_9969,N_9918);
nor UO_1050 (O_1050,N_9922,N_9900);
and UO_1051 (O_1051,N_9978,N_9912);
xor UO_1052 (O_1052,N_9929,N_9957);
or UO_1053 (O_1053,N_9989,N_9947);
and UO_1054 (O_1054,N_9958,N_9966);
nand UO_1055 (O_1055,N_9999,N_9909);
xor UO_1056 (O_1056,N_9907,N_9937);
and UO_1057 (O_1057,N_9953,N_9907);
xnor UO_1058 (O_1058,N_9902,N_9956);
nand UO_1059 (O_1059,N_9976,N_9965);
nand UO_1060 (O_1060,N_9980,N_9992);
and UO_1061 (O_1061,N_9978,N_9963);
nand UO_1062 (O_1062,N_9941,N_9900);
and UO_1063 (O_1063,N_9950,N_9984);
or UO_1064 (O_1064,N_9948,N_9917);
or UO_1065 (O_1065,N_9921,N_9904);
nor UO_1066 (O_1066,N_9964,N_9933);
nor UO_1067 (O_1067,N_9952,N_9957);
nand UO_1068 (O_1068,N_9905,N_9979);
or UO_1069 (O_1069,N_9902,N_9955);
nand UO_1070 (O_1070,N_9959,N_9904);
and UO_1071 (O_1071,N_9995,N_9934);
and UO_1072 (O_1072,N_9987,N_9911);
nand UO_1073 (O_1073,N_9964,N_9976);
xnor UO_1074 (O_1074,N_9996,N_9976);
nor UO_1075 (O_1075,N_9927,N_9987);
and UO_1076 (O_1076,N_9964,N_9981);
xnor UO_1077 (O_1077,N_9983,N_9953);
or UO_1078 (O_1078,N_9977,N_9938);
nor UO_1079 (O_1079,N_9960,N_9903);
nand UO_1080 (O_1080,N_9978,N_9929);
or UO_1081 (O_1081,N_9917,N_9911);
nor UO_1082 (O_1082,N_9987,N_9928);
xnor UO_1083 (O_1083,N_9999,N_9949);
or UO_1084 (O_1084,N_9967,N_9934);
and UO_1085 (O_1085,N_9952,N_9911);
and UO_1086 (O_1086,N_9940,N_9913);
nand UO_1087 (O_1087,N_9991,N_9927);
nor UO_1088 (O_1088,N_9934,N_9907);
nor UO_1089 (O_1089,N_9952,N_9913);
or UO_1090 (O_1090,N_9969,N_9983);
nand UO_1091 (O_1091,N_9921,N_9932);
or UO_1092 (O_1092,N_9919,N_9987);
xnor UO_1093 (O_1093,N_9920,N_9924);
nand UO_1094 (O_1094,N_9997,N_9951);
or UO_1095 (O_1095,N_9946,N_9919);
nor UO_1096 (O_1096,N_9988,N_9973);
xor UO_1097 (O_1097,N_9975,N_9934);
xnor UO_1098 (O_1098,N_9947,N_9991);
and UO_1099 (O_1099,N_9934,N_9937);
or UO_1100 (O_1100,N_9957,N_9993);
and UO_1101 (O_1101,N_9913,N_9954);
nand UO_1102 (O_1102,N_9936,N_9997);
or UO_1103 (O_1103,N_9969,N_9909);
nor UO_1104 (O_1104,N_9947,N_9908);
or UO_1105 (O_1105,N_9997,N_9913);
or UO_1106 (O_1106,N_9943,N_9914);
or UO_1107 (O_1107,N_9981,N_9990);
or UO_1108 (O_1108,N_9918,N_9995);
nor UO_1109 (O_1109,N_9967,N_9968);
nor UO_1110 (O_1110,N_9938,N_9926);
and UO_1111 (O_1111,N_9946,N_9991);
nor UO_1112 (O_1112,N_9976,N_9967);
nand UO_1113 (O_1113,N_9918,N_9946);
or UO_1114 (O_1114,N_9953,N_9958);
nand UO_1115 (O_1115,N_9936,N_9960);
nor UO_1116 (O_1116,N_9910,N_9964);
or UO_1117 (O_1117,N_9976,N_9939);
and UO_1118 (O_1118,N_9917,N_9990);
and UO_1119 (O_1119,N_9940,N_9912);
nor UO_1120 (O_1120,N_9924,N_9979);
nand UO_1121 (O_1121,N_9953,N_9979);
nor UO_1122 (O_1122,N_9981,N_9902);
or UO_1123 (O_1123,N_9956,N_9978);
nand UO_1124 (O_1124,N_9946,N_9924);
nand UO_1125 (O_1125,N_9953,N_9959);
nor UO_1126 (O_1126,N_9993,N_9953);
and UO_1127 (O_1127,N_9945,N_9936);
nand UO_1128 (O_1128,N_9980,N_9918);
nand UO_1129 (O_1129,N_9961,N_9930);
or UO_1130 (O_1130,N_9972,N_9946);
or UO_1131 (O_1131,N_9928,N_9981);
nor UO_1132 (O_1132,N_9979,N_9902);
or UO_1133 (O_1133,N_9963,N_9917);
or UO_1134 (O_1134,N_9979,N_9971);
xnor UO_1135 (O_1135,N_9983,N_9908);
or UO_1136 (O_1136,N_9914,N_9948);
xnor UO_1137 (O_1137,N_9965,N_9974);
nand UO_1138 (O_1138,N_9951,N_9986);
and UO_1139 (O_1139,N_9968,N_9912);
or UO_1140 (O_1140,N_9948,N_9926);
and UO_1141 (O_1141,N_9920,N_9917);
nand UO_1142 (O_1142,N_9903,N_9962);
xor UO_1143 (O_1143,N_9942,N_9944);
xnor UO_1144 (O_1144,N_9934,N_9983);
or UO_1145 (O_1145,N_9969,N_9984);
or UO_1146 (O_1146,N_9909,N_9906);
or UO_1147 (O_1147,N_9995,N_9901);
and UO_1148 (O_1148,N_9998,N_9911);
and UO_1149 (O_1149,N_9908,N_9927);
and UO_1150 (O_1150,N_9942,N_9992);
nand UO_1151 (O_1151,N_9913,N_9994);
nor UO_1152 (O_1152,N_9971,N_9997);
nand UO_1153 (O_1153,N_9944,N_9999);
nor UO_1154 (O_1154,N_9919,N_9907);
and UO_1155 (O_1155,N_9946,N_9930);
xnor UO_1156 (O_1156,N_9962,N_9998);
or UO_1157 (O_1157,N_9923,N_9945);
xnor UO_1158 (O_1158,N_9998,N_9964);
xnor UO_1159 (O_1159,N_9973,N_9999);
xor UO_1160 (O_1160,N_9922,N_9964);
and UO_1161 (O_1161,N_9968,N_9981);
xor UO_1162 (O_1162,N_9946,N_9936);
nand UO_1163 (O_1163,N_9916,N_9948);
nor UO_1164 (O_1164,N_9951,N_9959);
or UO_1165 (O_1165,N_9945,N_9900);
nand UO_1166 (O_1166,N_9948,N_9980);
nor UO_1167 (O_1167,N_9929,N_9960);
nor UO_1168 (O_1168,N_9981,N_9944);
and UO_1169 (O_1169,N_9962,N_9946);
nand UO_1170 (O_1170,N_9906,N_9980);
nand UO_1171 (O_1171,N_9935,N_9948);
nand UO_1172 (O_1172,N_9999,N_9915);
or UO_1173 (O_1173,N_9986,N_9957);
or UO_1174 (O_1174,N_9967,N_9978);
nor UO_1175 (O_1175,N_9948,N_9929);
and UO_1176 (O_1176,N_9949,N_9950);
nand UO_1177 (O_1177,N_9979,N_9945);
and UO_1178 (O_1178,N_9909,N_9981);
and UO_1179 (O_1179,N_9971,N_9969);
nand UO_1180 (O_1180,N_9923,N_9901);
or UO_1181 (O_1181,N_9914,N_9934);
xor UO_1182 (O_1182,N_9966,N_9929);
or UO_1183 (O_1183,N_9909,N_9980);
nor UO_1184 (O_1184,N_9992,N_9939);
nand UO_1185 (O_1185,N_9984,N_9953);
or UO_1186 (O_1186,N_9916,N_9992);
or UO_1187 (O_1187,N_9926,N_9908);
and UO_1188 (O_1188,N_9976,N_9906);
and UO_1189 (O_1189,N_9935,N_9931);
or UO_1190 (O_1190,N_9930,N_9933);
and UO_1191 (O_1191,N_9943,N_9924);
xnor UO_1192 (O_1192,N_9908,N_9943);
nand UO_1193 (O_1193,N_9949,N_9922);
or UO_1194 (O_1194,N_9994,N_9946);
and UO_1195 (O_1195,N_9956,N_9971);
or UO_1196 (O_1196,N_9998,N_9909);
xor UO_1197 (O_1197,N_9903,N_9939);
nand UO_1198 (O_1198,N_9911,N_9913);
or UO_1199 (O_1199,N_9915,N_9939);
and UO_1200 (O_1200,N_9985,N_9952);
xnor UO_1201 (O_1201,N_9927,N_9903);
nor UO_1202 (O_1202,N_9936,N_9993);
nand UO_1203 (O_1203,N_9911,N_9981);
nand UO_1204 (O_1204,N_9997,N_9966);
or UO_1205 (O_1205,N_9935,N_9995);
and UO_1206 (O_1206,N_9906,N_9964);
nor UO_1207 (O_1207,N_9912,N_9907);
nand UO_1208 (O_1208,N_9942,N_9934);
and UO_1209 (O_1209,N_9994,N_9903);
or UO_1210 (O_1210,N_9952,N_9962);
xor UO_1211 (O_1211,N_9960,N_9987);
xor UO_1212 (O_1212,N_9973,N_9907);
and UO_1213 (O_1213,N_9925,N_9934);
nor UO_1214 (O_1214,N_9935,N_9957);
nor UO_1215 (O_1215,N_9987,N_9949);
nor UO_1216 (O_1216,N_9982,N_9918);
nand UO_1217 (O_1217,N_9911,N_9964);
nand UO_1218 (O_1218,N_9933,N_9973);
nor UO_1219 (O_1219,N_9911,N_9946);
nor UO_1220 (O_1220,N_9984,N_9945);
nand UO_1221 (O_1221,N_9990,N_9935);
nand UO_1222 (O_1222,N_9993,N_9905);
nand UO_1223 (O_1223,N_9933,N_9947);
and UO_1224 (O_1224,N_9949,N_9929);
or UO_1225 (O_1225,N_9990,N_9965);
nand UO_1226 (O_1226,N_9992,N_9997);
and UO_1227 (O_1227,N_9933,N_9914);
and UO_1228 (O_1228,N_9934,N_9958);
and UO_1229 (O_1229,N_9928,N_9922);
nor UO_1230 (O_1230,N_9996,N_9952);
nor UO_1231 (O_1231,N_9929,N_9915);
and UO_1232 (O_1232,N_9982,N_9955);
and UO_1233 (O_1233,N_9986,N_9929);
nor UO_1234 (O_1234,N_9972,N_9907);
nor UO_1235 (O_1235,N_9949,N_9978);
and UO_1236 (O_1236,N_9916,N_9937);
nor UO_1237 (O_1237,N_9923,N_9935);
or UO_1238 (O_1238,N_9923,N_9996);
or UO_1239 (O_1239,N_9914,N_9964);
nor UO_1240 (O_1240,N_9968,N_9917);
and UO_1241 (O_1241,N_9923,N_9997);
nand UO_1242 (O_1242,N_9988,N_9908);
nand UO_1243 (O_1243,N_9994,N_9902);
nand UO_1244 (O_1244,N_9923,N_9930);
nor UO_1245 (O_1245,N_9973,N_9987);
xor UO_1246 (O_1246,N_9905,N_9926);
or UO_1247 (O_1247,N_9920,N_9938);
and UO_1248 (O_1248,N_9936,N_9965);
nand UO_1249 (O_1249,N_9975,N_9982);
or UO_1250 (O_1250,N_9933,N_9906);
nand UO_1251 (O_1251,N_9995,N_9956);
and UO_1252 (O_1252,N_9936,N_9991);
nor UO_1253 (O_1253,N_9951,N_9962);
xor UO_1254 (O_1254,N_9994,N_9954);
xor UO_1255 (O_1255,N_9958,N_9917);
and UO_1256 (O_1256,N_9987,N_9992);
nand UO_1257 (O_1257,N_9900,N_9901);
or UO_1258 (O_1258,N_9953,N_9964);
and UO_1259 (O_1259,N_9935,N_9929);
nor UO_1260 (O_1260,N_9957,N_9987);
nand UO_1261 (O_1261,N_9953,N_9998);
xnor UO_1262 (O_1262,N_9994,N_9909);
or UO_1263 (O_1263,N_9947,N_9921);
or UO_1264 (O_1264,N_9948,N_9908);
nor UO_1265 (O_1265,N_9949,N_9935);
nor UO_1266 (O_1266,N_9914,N_9961);
and UO_1267 (O_1267,N_9968,N_9965);
and UO_1268 (O_1268,N_9914,N_9960);
nor UO_1269 (O_1269,N_9986,N_9930);
and UO_1270 (O_1270,N_9913,N_9925);
xnor UO_1271 (O_1271,N_9940,N_9946);
nor UO_1272 (O_1272,N_9965,N_9942);
or UO_1273 (O_1273,N_9990,N_9968);
or UO_1274 (O_1274,N_9935,N_9944);
nand UO_1275 (O_1275,N_9942,N_9984);
nor UO_1276 (O_1276,N_9921,N_9907);
or UO_1277 (O_1277,N_9917,N_9986);
nor UO_1278 (O_1278,N_9996,N_9924);
nor UO_1279 (O_1279,N_9920,N_9953);
xnor UO_1280 (O_1280,N_9919,N_9920);
and UO_1281 (O_1281,N_9998,N_9939);
and UO_1282 (O_1282,N_9900,N_9979);
or UO_1283 (O_1283,N_9992,N_9978);
nand UO_1284 (O_1284,N_9942,N_9981);
nand UO_1285 (O_1285,N_9980,N_9990);
and UO_1286 (O_1286,N_9987,N_9902);
and UO_1287 (O_1287,N_9978,N_9926);
and UO_1288 (O_1288,N_9944,N_9929);
nand UO_1289 (O_1289,N_9979,N_9983);
xnor UO_1290 (O_1290,N_9971,N_9967);
and UO_1291 (O_1291,N_9963,N_9909);
nand UO_1292 (O_1292,N_9941,N_9967);
nor UO_1293 (O_1293,N_9977,N_9998);
or UO_1294 (O_1294,N_9940,N_9974);
nor UO_1295 (O_1295,N_9966,N_9999);
nand UO_1296 (O_1296,N_9927,N_9932);
nand UO_1297 (O_1297,N_9910,N_9972);
and UO_1298 (O_1298,N_9910,N_9963);
nand UO_1299 (O_1299,N_9952,N_9970);
nor UO_1300 (O_1300,N_9918,N_9959);
nor UO_1301 (O_1301,N_9918,N_9942);
or UO_1302 (O_1302,N_9989,N_9923);
or UO_1303 (O_1303,N_9934,N_9911);
xor UO_1304 (O_1304,N_9941,N_9908);
nand UO_1305 (O_1305,N_9998,N_9981);
or UO_1306 (O_1306,N_9961,N_9997);
nor UO_1307 (O_1307,N_9946,N_9928);
or UO_1308 (O_1308,N_9952,N_9988);
nand UO_1309 (O_1309,N_9990,N_9906);
and UO_1310 (O_1310,N_9956,N_9991);
nor UO_1311 (O_1311,N_9994,N_9992);
and UO_1312 (O_1312,N_9947,N_9956);
nor UO_1313 (O_1313,N_9940,N_9908);
nor UO_1314 (O_1314,N_9981,N_9995);
and UO_1315 (O_1315,N_9904,N_9920);
nand UO_1316 (O_1316,N_9912,N_9941);
nor UO_1317 (O_1317,N_9996,N_9956);
or UO_1318 (O_1318,N_9979,N_9965);
nor UO_1319 (O_1319,N_9933,N_9991);
and UO_1320 (O_1320,N_9979,N_9993);
and UO_1321 (O_1321,N_9957,N_9910);
or UO_1322 (O_1322,N_9916,N_9911);
and UO_1323 (O_1323,N_9921,N_9976);
or UO_1324 (O_1324,N_9935,N_9964);
and UO_1325 (O_1325,N_9992,N_9955);
nor UO_1326 (O_1326,N_9978,N_9942);
nand UO_1327 (O_1327,N_9987,N_9906);
xnor UO_1328 (O_1328,N_9978,N_9903);
nand UO_1329 (O_1329,N_9903,N_9970);
and UO_1330 (O_1330,N_9984,N_9923);
and UO_1331 (O_1331,N_9942,N_9908);
and UO_1332 (O_1332,N_9916,N_9964);
or UO_1333 (O_1333,N_9910,N_9958);
nand UO_1334 (O_1334,N_9904,N_9955);
xor UO_1335 (O_1335,N_9958,N_9962);
xnor UO_1336 (O_1336,N_9952,N_9935);
xnor UO_1337 (O_1337,N_9974,N_9911);
nand UO_1338 (O_1338,N_9937,N_9924);
and UO_1339 (O_1339,N_9979,N_9966);
nand UO_1340 (O_1340,N_9920,N_9954);
nor UO_1341 (O_1341,N_9982,N_9909);
or UO_1342 (O_1342,N_9955,N_9906);
or UO_1343 (O_1343,N_9920,N_9949);
nor UO_1344 (O_1344,N_9922,N_9971);
or UO_1345 (O_1345,N_9922,N_9978);
and UO_1346 (O_1346,N_9973,N_9932);
nor UO_1347 (O_1347,N_9972,N_9943);
nor UO_1348 (O_1348,N_9967,N_9905);
nand UO_1349 (O_1349,N_9937,N_9947);
nor UO_1350 (O_1350,N_9939,N_9993);
nand UO_1351 (O_1351,N_9918,N_9911);
and UO_1352 (O_1352,N_9931,N_9990);
nand UO_1353 (O_1353,N_9900,N_9935);
nand UO_1354 (O_1354,N_9911,N_9949);
nor UO_1355 (O_1355,N_9946,N_9982);
nand UO_1356 (O_1356,N_9903,N_9936);
or UO_1357 (O_1357,N_9933,N_9963);
or UO_1358 (O_1358,N_9964,N_9908);
nor UO_1359 (O_1359,N_9952,N_9927);
nor UO_1360 (O_1360,N_9931,N_9997);
or UO_1361 (O_1361,N_9964,N_9912);
xnor UO_1362 (O_1362,N_9942,N_9996);
xnor UO_1363 (O_1363,N_9989,N_9954);
nor UO_1364 (O_1364,N_9984,N_9959);
and UO_1365 (O_1365,N_9900,N_9917);
nor UO_1366 (O_1366,N_9972,N_9915);
nor UO_1367 (O_1367,N_9987,N_9952);
nand UO_1368 (O_1368,N_9932,N_9916);
nor UO_1369 (O_1369,N_9907,N_9906);
or UO_1370 (O_1370,N_9962,N_9918);
xnor UO_1371 (O_1371,N_9940,N_9942);
and UO_1372 (O_1372,N_9954,N_9962);
or UO_1373 (O_1373,N_9932,N_9926);
nor UO_1374 (O_1374,N_9931,N_9916);
nor UO_1375 (O_1375,N_9907,N_9917);
and UO_1376 (O_1376,N_9975,N_9989);
or UO_1377 (O_1377,N_9913,N_9927);
nand UO_1378 (O_1378,N_9935,N_9941);
nor UO_1379 (O_1379,N_9907,N_9981);
or UO_1380 (O_1380,N_9948,N_9983);
nor UO_1381 (O_1381,N_9920,N_9930);
or UO_1382 (O_1382,N_9976,N_9982);
nor UO_1383 (O_1383,N_9917,N_9960);
nor UO_1384 (O_1384,N_9983,N_9967);
and UO_1385 (O_1385,N_9990,N_9928);
and UO_1386 (O_1386,N_9983,N_9982);
nor UO_1387 (O_1387,N_9973,N_9904);
nor UO_1388 (O_1388,N_9961,N_9934);
nand UO_1389 (O_1389,N_9905,N_9973);
or UO_1390 (O_1390,N_9901,N_9992);
and UO_1391 (O_1391,N_9934,N_9969);
nor UO_1392 (O_1392,N_9973,N_9957);
nand UO_1393 (O_1393,N_9979,N_9995);
or UO_1394 (O_1394,N_9945,N_9964);
nand UO_1395 (O_1395,N_9920,N_9937);
nor UO_1396 (O_1396,N_9999,N_9967);
nor UO_1397 (O_1397,N_9990,N_9938);
nand UO_1398 (O_1398,N_9999,N_9947);
and UO_1399 (O_1399,N_9901,N_9919);
or UO_1400 (O_1400,N_9902,N_9908);
or UO_1401 (O_1401,N_9992,N_9937);
xnor UO_1402 (O_1402,N_9931,N_9992);
nor UO_1403 (O_1403,N_9941,N_9944);
nor UO_1404 (O_1404,N_9986,N_9903);
nand UO_1405 (O_1405,N_9971,N_9912);
xor UO_1406 (O_1406,N_9940,N_9914);
nor UO_1407 (O_1407,N_9905,N_9901);
nor UO_1408 (O_1408,N_9946,N_9900);
nor UO_1409 (O_1409,N_9921,N_9995);
nor UO_1410 (O_1410,N_9929,N_9953);
and UO_1411 (O_1411,N_9957,N_9924);
nor UO_1412 (O_1412,N_9977,N_9947);
or UO_1413 (O_1413,N_9978,N_9916);
or UO_1414 (O_1414,N_9920,N_9976);
nor UO_1415 (O_1415,N_9914,N_9970);
nand UO_1416 (O_1416,N_9976,N_9948);
nor UO_1417 (O_1417,N_9919,N_9984);
nor UO_1418 (O_1418,N_9969,N_9920);
nor UO_1419 (O_1419,N_9976,N_9954);
nor UO_1420 (O_1420,N_9984,N_9917);
nand UO_1421 (O_1421,N_9956,N_9951);
nor UO_1422 (O_1422,N_9917,N_9985);
nand UO_1423 (O_1423,N_9933,N_9911);
nor UO_1424 (O_1424,N_9987,N_9918);
or UO_1425 (O_1425,N_9959,N_9930);
nor UO_1426 (O_1426,N_9915,N_9951);
or UO_1427 (O_1427,N_9904,N_9906);
or UO_1428 (O_1428,N_9903,N_9912);
or UO_1429 (O_1429,N_9900,N_9954);
xor UO_1430 (O_1430,N_9968,N_9919);
and UO_1431 (O_1431,N_9947,N_9902);
xnor UO_1432 (O_1432,N_9943,N_9926);
or UO_1433 (O_1433,N_9989,N_9971);
nand UO_1434 (O_1434,N_9975,N_9939);
and UO_1435 (O_1435,N_9936,N_9920);
and UO_1436 (O_1436,N_9999,N_9941);
nand UO_1437 (O_1437,N_9915,N_9971);
and UO_1438 (O_1438,N_9916,N_9980);
and UO_1439 (O_1439,N_9996,N_9903);
nor UO_1440 (O_1440,N_9977,N_9909);
nand UO_1441 (O_1441,N_9946,N_9990);
nand UO_1442 (O_1442,N_9959,N_9977);
nor UO_1443 (O_1443,N_9990,N_9901);
and UO_1444 (O_1444,N_9980,N_9951);
nor UO_1445 (O_1445,N_9943,N_9965);
xor UO_1446 (O_1446,N_9974,N_9998);
or UO_1447 (O_1447,N_9915,N_9900);
or UO_1448 (O_1448,N_9981,N_9901);
xnor UO_1449 (O_1449,N_9967,N_9959);
or UO_1450 (O_1450,N_9949,N_9902);
nand UO_1451 (O_1451,N_9967,N_9900);
nor UO_1452 (O_1452,N_9973,N_9917);
and UO_1453 (O_1453,N_9986,N_9988);
and UO_1454 (O_1454,N_9972,N_9988);
or UO_1455 (O_1455,N_9996,N_9974);
and UO_1456 (O_1456,N_9970,N_9999);
and UO_1457 (O_1457,N_9944,N_9913);
nand UO_1458 (O_1458,N_9980,N_9944);
or UO_1459 (O_1459,N_9968,N_9980);
nand UO_1460 (O_1460,N_9918,N_9963);
nor UO_1461 (O_1461,N_9978,N_9960);
or UO_1462 (O_1462,N_9941,N_9997);
and UO_1463 (O_1463,N_9924,N_9947);
and UO_1464 (O_1464,N_9997,N_9995);
nand UO_1465 (O_1465,N_9995,N_9993);
or UO_1466 (O_1466,N_9935,N_9969);
and UO_1467 (O_1467,N_9935,N_9937);
or UO_1468 (O_1468,N_9956,N_9954);
and UO_1469 (O_1469,N_9923,N_9966);
or UO_1470 (O_1470,N_9997,N_9943);
or UO_1471 (O_1471,N_9934,N_9918);
and UO_1472 (O_1472,N_9941,N_9957);
nand UO_1473 (O_1473,N_9913,N_9941);
and UO_1474 (O_1474,N_9955,N_9956);
xnor UO_1475 (O_1475,N_9963,N_9986);
or UO_1476 (O_1476,N_9955,N_9900);
nand UO_1477 (O_1477,N_9956,N_9919);
nor UO_1478 (O_1478,N_9980,N_9975);
nand UO_1479 (O_1479,N_9932,N_9922);
and UO_1480 (O_1480,N_9924,N_9942);
nand UO_1481 (O_1481,N_9972,N_9991);
nand UO_1482 (O_1482,N_9999,N_9955);
nand UO_1483 (O_1483,N_9952,N_9979);
and UO_1484 (O_1484,N_9976,N_9963);
and UO_1485 (O_1485,N_9912,N_9959);
nand UO_1486 (O_1486,N_9943,N_9987);
nand UO_1487 (O_1487,N_9969,N_9924);
or UO_1488 (O_1488,N_9903,N_9999);
nand UO_1489 (O_1489,N_9922,N_9954);
nor UO_1490 (O_1490,N_9937,N_9942);
or UO_1491 (O_1491,N_9998,N_9975);
xnor UO_1492 (O_1492,N_9971,N_9964);
nand UO_1493 (O_1493,N_9905,N_9968);
nor UO_1494 (O_1494,N_9990,N_9915);
nand UO_1495 (O_1495,N_9993,N_9990);
or UO_1496 (O_1496,N_9973,N_9962);
nor UO_1497 (O_1497,N_9934,N_9957);
and UO_1498 (O_1498,N_9998,N_9935);
or UO_1499 (O_1499,N_9915,N_9913);
endmodule